module basic_1500_15000_2000_5_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_431,In_289);
nor U1 (N_1,In_1053,In_1286);
nor U2 (N_2,In_1197,In_1034);
or U3 (N_3,In_1374,In_843);
nand U4 (N_4,In_820,In_206);
nand U5 (N_5,In_36,In_1153);
and U6 (N_6,In_819,In_801);
nand U7 (N_7,In_31,In_974);
nor U8 (N_8,In_675,In_804);
nor U9 (N_9,In_1460,In_597);
nor U10 (N_10,In_960,In_962);
nand U11 (N_11,In_1031,In_645);
xnor U12 (N_12,In_1438,In_1100);
or U13 (N_13,In_1491,In_996);
nand U14 (N_14,In_827,In_307);
or U15 (N_15,In_761,In_368);
nor U16 (N_16,In_977,In_1224);
or U17 (N_17,In_1308,In_254);
or U18 (N_18,In_391,In_252);
and U19 (N_19,In_949,In_743);
nand U20 (N_20,In_253,In_470);
and U21 (N_21,In_1190,In_88);
or U22 (N_22,In_10,In_82);
and U23 (N_23,In_1146,In_1332);
or U24 (N_24,In_559,In_337);
nor U25 (N_25,In_377,In_747);
and U26 (N_26,In_237,In_961);
nand U27 (N_27,In_1135,In_746);
and U28 (N_28,In_256,In_1274);
and U29 (N_29,In_1305,In_44);
nor U30 (N_30,In_1273,In_1233);
and U31 (N_31,In_1411,In_1096);
and U32 (N_32,In_509,In_1284);
nor U33 (N_33,In_854,In_154);
nor U34 (N_34,In_13,In_224);
and U35 (N_35,In_434,In_401);
or U36 (N_36,In_934,In_896);
nand U37 (N_37,In_1128,In_528);
and U38 (N_38,In_441,In_808);
or U39 (N_39,In_1439,In_282);
nand U40 (N_40,In_1481,In_361);
nand U41 (N_41,In_793,In_1117);
and U42 (N_42,In_1014,In_553);
and U43 (N_43,In_92,In_416);
xnor U44 (N_44,In_1016,In_504);
xor U45 (N_45,In_152,In_158);
nand U46 (N_46,In_823,In_175);
and U47 (N_47,In_702,In_978);
nor U48 (N_48,In_1140,In_239);
nor U49 (N_49,In_1176,In_28);
and U50 (N_50,In_321,In_1363);
nand U51 (N_51,In_352,In_6);
and U52 (N_52,In_536,In_846);
and U53 (N_53,In_378,In_1183);
nor U54 (N_54,In_399,In_116);
nor U55 (N_55,In_1152,In_366);
and U56 (N_56,In_939,In_710);
and U57 (N_57,In_581,In_765);
xor U58 (N_58,In_1495,In_519);
and U59 (N_59,In_678,In_1384);
nor U60 (N_60,In_139,In_1242);
nand U61 (N_61,In_855,In_471);
nand U62 (N_62,In_570,In_350);
or U63 (N_63,In_1063,In_622);
and U64 (N_64,In_880,In_1292);
nor U65 (N_65,In_807,In_1487);
nor U66 (N_66,In_1383,In_999);
nor U67 (N_67,In_1321,In_40);
nor U68 (N_68,In_341,In_1032);
and U69 (N_69,In_692,In_875);
and U70 (N_70,In_969,In_24);
or U71 (N_71,In_261,In_660);
or U72 (N_72,In_1248,In_490);
or U73 (N_73,In_1236,In_555);
nor U74 (N_74,In_631,In_1436);
or U75 (N_75,In_693,In_1098);
xnor U76 (N_76,In_1237,In_125);
and U77 (N_77,In_1205,In_748);
or U78 (N_78,In_1073,In_179);
or U79 (N_79,In_111,In_964);
xnor U80 (N_80,In_283,In_310);
nor U81 (N_81,In_1262,In_810);
nor U82 (N_82,In_1023,In_1173);
or U83 (N_83,In_229,In_1093);
nor U84 (N_84,In_66,In_23);
nor U85 (N_85,In_184,In_639);
and U86 (N_86,In_1226,In_327);
and U87 (N_87,In_1428,In_1360);
nand U88 (N_88,In_772,In_1334);
or U89 (N_89,In_561,In_1157);
xor U90 (N_90,In_565,In_756);
or U91 (N_91,In_988,In_971);
xnor U92 (N_92,In_1120,In_1486);
nand U93 (N_93,In_1036,In_19);
nand U94 (N_94,In_435,In_1364);
and U95 (N_95,In_1365,In_1108);
xor U96 (N_96,In_607,In_144);
xnor U97 (N_97,In_1437,In_1201);
or U98 (N_98,In_1109,In_1377);
and U99 (N_99,In_458,In_143);
nor U100 (N_100,In_81,In_22);
and U101 (N_101,In_1241,In_757);
or U102 (N_102,In_665,In_402);
or U103 (N_103,In_113,In_1294);
and U104 (N_104,In_1368,In_1299);
xor U105 (N_105,In_518,In_1);
or U106 (N_106,In_1263,In_1429);
nor U107 (N_107,In_674,In_345);
nor U108 (N_108,In_835,In_1257);
nor U109 (N_109,In_510,In_572);
and U110 (N_110,In_172,In_1345);
nor U111 (N_111,In_1103,In_850);
nor U112 (N_112,In_904,In_697);
or U113 (N_113,In_1177,In_718);
nor U114 (N_114,In_67,In_929);
nor U115 (N_115,In_822,In_840);
and U116 (N_116,In_1245,In_178);
and U117 (N_117,In_1085,In_48);
xor U118 (N_118,In_837,In_842);
nand U119 (N_119,In_566,In_611);
and U120 (N_120,In_1361,In_594);
or U121 (N_121,In_844,In_147);
nor U122 (N_122,In_1024,In_780);
nor U123 (N_123,In_186,In_429);
nand U124 (N_124,In_538,In_1194);
and U125 (N_125,In_277,In_1039);
nor U126 (N_126,In_942,In_1217);
nand U127 (N_127,In_647,In_853);
xnor U128 (N_128,In_549,In_1225);
nor U129 (N_129,In_486,In_918);
nand U130 (N_130,In_478,In_1001);
xnor U131 (N_131,In_1403,In_372);
nor U132 (N_132,In_201,In_750);
and U133 (N_133,In_1319,In_308);
and U134 (N_134,In_1249,In_1206);
nor U135 (N_135,In_395,In_1422);
nand U136 (N_136,In_602,In_417);
nor U137 (N_137,In_1326,In_1078);
nor U138 (N_138,In_655,In_16);
or U139 (N_139,In_1269,In_209);
and U140 (N_140,In_963,In_595);
nor U141 (N_141,In_1306,In_573);
nor U142 (N_142,In_1082,In_706);
nor U143 (N_143,In_1070,In_1317);
nor U144 (N_144,In_290,In_159);
xnor U145 (N_145,In_879,In_1449);
and U146 (N_146,In_1134,In_1404);
and U147 (N_147,In_1490,In_601);
or U148 (N_148,In_1347,In_1342);
and U149 (N_149,In_1051,In_856);
or U150 (N_150,In_1366,In_295);
or U151 (N_151,In_1265,In_907);
or U152 (N_152,In_604,In_250);
and U153 (N_153,In_590,In_792);
and U154 (N_154,In_318,In_861);
nor U155 (N_155,In_344,In_35);
nand U156 (N_156,In_332,In_865);
nor U157 (N_157,In_728,In_1255);
nand U158 (N_158,In_1025,In_210);
nor U159 (N_159,In_118,In_475);
xnor U160 (N_160,In_1189,In_188);
or U161 (N_161,In_739,In_218);
nand U162 (N_162,In_195,In_859);
nor U163 (N_163,In_1182,In_292);
nand U164 (N_164,In_1095,In_523);
or U165 (N_165,In_1401,In_207);
and U166 (N_166,In_1488,In_1198);
nand U167 (N_167,In_374,In_931);
and U168 (N_168,In_1111,In_1002);
nand U169 (N_169,In_1026,In_1112);
xor U170 (N_170,In_1489,In_280);
nand U171 (N_171,In_670,In_740);
or U172 (N_172,In_713,In_894);
nor U173 (N_173,In_240,In_498);
nor U174 (N_174,In_500,In_893);
nor U175 (N_175,In_546,In_909);
nor U176 (N_176,In_293,In_432);
or U177 (N_177,In_719,In_970);
xor U178 (N_178,In_131,In_356);
nand U179 (N_179,In_579,In_571);
or U180 (N_180,In_142,In_862);
xnor U181 (N_181,In_369,In_889);
and U182 (N_182,In_110,In_609);
nor U183 (N_183,In_383,In_1370);
and U184 (N_184,In_335,In_552);
nand U185 (N_185,In_531,In_1030);
or U186 (N_186,In_442,In_491);
or U187 (N_187,In_365,In_811);
nor U188 (N_188,In_1106,In_1296);
nor U189 (N_189,In_932,In_348);
and U190 (N_190,In_683,In_1188);
or U191 (N_191,In_1028,In_77);
xnor U192 (N_192,In_45,In_895);
and U193 (N_193,In_1270,In_430);
nand U194 (N_194,In_1258,In_1171);
nor U195 (N_195,In_137,In_1426);
nand U196 (N_196,In_1327,In_1075);
and U197 (N_197,In_1048,In_657);
nand U198 (N_198,In_1208,In_754);
and U199 (N_199,In_868,In_599);
nor U200 (N_200,In_1144,In_664);
nor U201 (N_201,In_1022,In_1393);
and U202 (N_202,In_454,In_1318);
nand U203 (N_203,In_241,In_1083);
xnor U204 (N_204,In_717,In_900);
and U205 (N_205,In_829,In_938);
nor U206 (N_206,In_480,In_625);
nor U207 (N_207,In_149,In_349);
or U208 (N_208,In_917,In_589);
nor U209 (N_209,In_324,In_364);
and U210 (N_210,In_1250,In_476);
and U211 (N_211,In_232,In_1254);
and U212 (N_212,In_262,In_1040);
or U213 (N_213,In_1044,In_550);
xor U214 (N_214,In_408,In_641);
and U215 (N_215,In_216,In_18);
nor U216 (N_216,In_684,In_1155);
nand U217 (N_217,In_857,In_951);
nor U218 (N_218,In_1038,In_914);
nor U219 (N_219,In_708,In_314);
and U220 (N_220,In_543,In_731);
nand U221 (N_221,In_1339,In_1215);
nand U222 (N_222,In_150,In_1165);
nor U223 (N_223,In_1298,In_1042);
and U224 (N_224,In_502,In_634);
and U225 (N_225,In_1389,In_891);
or U226 (N_226,In_669,In_965);
nor U227 (N_227,In_233,In_326);
or U228 (N_228,In_1251,In_1397);
nor U229 (N_229,In_306,In_809);
or U230 (N_230,In_636,In_71);
nor U231 (N_231,In_1267,In_762);
or U232 (N_232,In_439,In_1291);
or U233 (N_233,In_212,In_1323);
nor U234 (N_234,In_1315,In_577);
xnor U235 (N_235,In_632,In_1094);
or U236 (N_236,In_214,In_1220);
nand U237 (N_237,In_1057,In_956);
nand U238 (N_238,In_987,In_1187);
or U239 (N_239,In_427,In_340);
nor U240 (N_240,In_452,In_1172);
or U241 (N_241,In_259,In_919);
nand U242 (N_242,In_1033,In_1047);
or U243 (N_243,In_80,In_1340);
nand U244 (N_244,In_913,In_438);
and U245 (N_245,In_723,In_517);
nand U246 (N_246,In_920,In_246);
nand U247 (N_247,In_460,In_802);
and U248 (N_248,In_336,In_638);
nor U249 (N_249,In_1065,In_1282);
xnor U250 (N_250,In_343,In_169);
nand U251 (N_251,In_1473,In_123);
nand U252 (N_252,In_911,In_580);
nor U253 (N_253,In_469,In_1137);
xor U254 (N_254,In_230,In_1402);
and U255 (N_255,In_1229,In_952);
or U256 (N_256,In_927,In_61);
xor U257 (N_257,In_881,In_1150);
nor U258 (N_258,In_1337,In_1092);
or U259 (N_259,In_182,In_433);
and U260 (N_260,In_34,In_27);
or U261 (N_261,In_1055,In_1376);
or U262 (N_262,In_784,In_1464);
or U263 (N_263,In_462,In_1214);
nor U264 (N_264,In_473,In_1018);
or U265 (N_265,In_245,In_925);
and U266 (N_266,In_915,In_271);
nand U267 (N_267,In_309,In_1129);
nor U268 (N_268,In_858,In_775);
xor U269 (N_269,In_1107,In_520);
xnor U270 (N_270,In_342,In_347);
nor U271 (N_271,In_773,In_1420);
or U272 (N_272,In_983,In_1329);
nor U273 (N_273,In_1043,In_260);
and U274 (N_274,In_1453,In_1114);
nand U275 (N_275,In_75,In_696);
or U276 (N_276,In_141,In_884);
xnor U277 (N_277,In_511,In_69);
and U278 (N_278,In_1061,In_1223);
and U279 (N_279,In_1170,In_560);
xnor U280 (N_280,In_874,In_1355);
nor U281 (N_281,In_541,In_1253);
and U282 (N_282,In_616,In_5);
or U283 (N_283,In_1432,In_217);
nor U284 (N_284,In_215,In_643);
or U285 (N_285,In_426,In_73);
nor U286 (N_286,In_185,In_1406);
nand U287 (N_287,In_495,In_1132);
or U288 (N_288,In_720,In_140);
or U289 (N_289,In_56,In_989);
and U290 (N_290,In_474,In_1445);
nor U291 (N_291,In_556,In_672);
nand U292 (N_292,In_958,In_1207);
and U293 (N_293,In_398,In_1278);
and U294 (N_294,In_46,In_738);
and U295 (N_295,In_109,In_812);
or U296 (N_296,In_791,In_1167);
nand U297 (N_297,In_1232,In_629);
nor U298 (N_298,In_1231,In_409);
xnor U299 (N_299,In_902,In_973);
xnor U300 (N_300,In_845,In_753);
or U301 (N_301,In_749,In_992);
nand U302 (N_302,In_187,In_193);
and U303 (N_303,In_596,In_1290);
nor U304 (N_304,In_1102,In_330);
nand U305 (N_305,In_1302,In_359);
nand U306 (N_306,In_393,In_626);
nand U307 (N_307,In_1392,In_134);
nor U308 (N_308,In_1396,In_725);
nor U309 (N_309,In_1276,In_381);
xor U310 (N_310,In_196,In_910);
and U311 (N_311,In_74,In_933);
nand U312 (N_312,In_976,In_1193);
or U313 (N_313,In_311,In_1476);
nand U314 (N_314,In_637,In_315);
or U315 (N_315,In_703,In_709);
nor U316 (N_316,In_617,In_1169);
and U317 (N_317,In_1184,In_821);
or U318 (N_318,In_1121,In_1322);
or U319 (N_319,In_1477,In_79);
nor U320 (N_320,In_985,In_943);
nand U321 (N_321,In_1003,In_136);
nor U322 (N_322,In_582,In_62);
nand U323 (N_323,In_472,In_457);
nand U324 (N_324,In_461,In_1472);
nor U325 (N_325,In_781,In_1373);
or U326 (N_326,In_382,In_785);
xnor U327 (N_327,In_1164,In_662);
and U328 (N_328,In_1281,In_1465);
nand U329 (N_329,In_211,In_1338);
nor U330 (N_330,In_489,In_576);
nor U331 (N_331,In_1483,In_997);
xnor U332 (N_332,In_97,In_11);
nor U333 (N_333,In_1077,In_524);
and U334 (N_334,In_183,In_387);
and U335 (N_335,In_1418,In_1049);
nand U336 (N_336,In_453,In_885);
nor U337 (N_337,In_1394,In_1099);
nand U338 (N_338,In_621,In_33);
or U339 (N_339,In_379,In_870);
nor U340 (N_340,In_1133,In_1463);
and U341 (N_341,In_598,In_763);
nor U342 (N_342,In_1086,In_117);
or U343 (N_343,In_4,In_1341);
or U344 (N_344,In_529,In_1415);
nor U345 (N_345,In_1256,In_569);
xnor U346 (N_346,In_1325,In_112);
nand U347 (N_347,In_514,In_1412);
nand U348 (N_348,In_776,In_1320);
nor U349 (N_349,In_800,In_1441);
or U350 (N_350,In_121,In_796);
nand U351 (N_351,In_1213,In_1056);
and U352 (N_352,In_707,In_21);
xor U353 (N_353,In_1468,In_355);
or U354 (N_354,In_1378,In_482);
or U355 (N_355,In_1433,In_1260);
nand U356 (N_356,In_1119,In_816);
nand U357 (N_357,In_711,In_492);
and U358 (N_358,In_1211,In_194);
nor U359 (N_359,In_122,In_1154);
nor U360 (N_360,In_1498,In_1440);
nor U361 (N_361,In_1280,In_652);
nor U362 (N_362,In_1369,In_608);
xnor U363 (N_363,In_353,In_779);
and U364 (N_364,In_724,In_1357);
nand U365 (N_365,In_317,In_659);
and U366 (N_366,In_181,In_1382);
nand U367 (N_367,In_1052,In_132);
nand U368 (N_368,In_269,In_107);
and U369 (N_369,In_866,In_394);
or U370 (N_370,In_276,In_535);
nor U371 (N_371,In_274,In_114);
or U372 (N_372,In_0,In_300);
or U373 (N_373,In_764,In_1354);
or U374 (N_374,In_727,In_1466);
xnor U375 (N_375,In_410,In_1407);
and U376 (N_376,In_1029,In_1162);
nand U377 (N_377,In_405,In_1410);
xor U378 (N_378,In_59,In_226);
and U379 (N_379,In_464,In_1434);
nor U380 (N_380,In_1451,In_1259);
or U381 (N_381,In_89,In_487);
and U382 (N_382,In_968,In_168);
nand U383 (N_383,In_287,In_745);
and U384 (N_384,In_1311,In_244);
and U385 (N_385,In_396,In_1239);
nand U386 (N_386,In_1244,In_568);
or U387 (N_387,In_799,In_1212);
xor U388 (N_388,In_1045,In_852);
nand U389 (N_389,In_463,In_1386);
nor U390 (N_390,In_57,In_1158);
or U391 (N_391,In_466,In_305);
nand U392 (N_392,In_1425,In_20);
or U393 (N_393,In_54,In_774);
nor U394 (N_394,In_1230,In_867);
or U395 (N_395,In_257,In_95);
nor U396 (N_396,In_712,In_331);
and U397 (N_397,In_477,In_1417);
nand U398 (N_398,In_248,In_1362);
nand U399 (N_399,In_924,In_755);
nand U400 (N_400,In_1068,In_790);
nor U401 (N_401,In_751,In_1174);
xor U402 (N_402,In_1470,In_921);
nand U403 (N_403,In_787,In_1159);
nand U404 (N_404,In_928,In_138);
nor U405 (N_405,In_213,In_86);
nand U406 (N_406,In_263,In_1191);
nand U407 (N_407,In_444,In_291);
nand U408 (N_408,In_741,In_685);
nor U409 (N_409,In_400,In_322);
nor U410 (N_410,In_1139,In_554);
nand U411 (N_411,In_898,In_588);
xor U412 (N_412,In_567,In_771);
nand U413 (N_413,In_1240,In_78);
or U414 (N_414,In_610,In_231);
and U415 (N_415,In_161,In_547);
or U416 (N_416,In_847,In_281);
and U417 (N_417,In_198,In_205);
nand U418 (N_418,In_85,In_1398);
xor U419 (N_419,In_687,In_1351);
or U420 (N_420,In_767,In_1041);
nand U421 (N_421,In_297,In_975);
nor U422 (N_422,In_623,In_1293);
or U423 (N_423,In_940,In_817);
xor U424 (N_424,In_423,In_864);
and U425 (N_425,In_127,In_945);
nor U426 (N_426,In_966,In_649);
xnor U427 (N_427,In_171,In_777);
xnor U428 (N_428,In_413,In_238);
or U429 (N_429,In_468,In_1492);
xor U430 (N_430,In_813,In_586);
nand U431 (N_431,In_1330,In_1252);
nor U432 (N_432,In_493,In_51);
nor U433 (N_433,In_690,In_102);
or U434 (N_434,In_783,In_1275);
nand U435 (N_435,In_329,In_640);
nand U436 (N_436,In_1125,In_304);
nand U437 (N_437,In_1448,In_285);
xnor U438 (N_438,In_1064,In_1127);
nor U439 (N_439,In_53,In_485);
and U440 (N_440,In_1216,In_1399);
nand U441 (N_441,In_600,In_686);
nand U442 (N_442,In_72,In_627);
or U443 (N_443,In_167,In_1080);
nand U444 (N_444,In_668,In_908);
nor U445 (N_445,In_160,In_794);
or U446 (N_446,In_101,In_1161);
or U447 (N_447,In_612,In_564);
nand U448 (N_448,In_84,In_1391);
nand U449 (N_449,In_47,In_730);
and U450 (N_450,In_545,In_49);
nand U451 (N_451,In_94,In_1494);
or U452 (N_452,In_362,In_1452);
and U453 (N_453,In_220,In_299);
nor U454 (N_454,In_1136,In_937);
and U455 (N_455,In_303,In_782);
nand U456 (N_456,In_1021,In_499);
or U457 (N_457,In_1246,In_912);
and U458 (N_458,In_76,In_180);
and U459 (N_459,In_1124,In_1079);
nor U460 (N_460,In_43,In_126);
and U461 (N_461,In_1020,In_176);
nor U462 (N_462,In_106,In_1419);
or U463 (N_463,In_390,In_1356);
nand U464 (N_464,In_451,In_145);
xnor U465 (N_465,In_1059,In_32);
nand U466 (N_466,In_412,In_505);
or U467 (N_467,In_1149,In_644);
or U468 (N_468,In_680,In_848);
or U469 (N_469,In_41,In_133);
xnor U470 (N_470,In_766,In_941);
and U471 (N_471,In_1335,In_1331);
nor U472 (N_472,In_334,In_1088);
or U473 (N_473,In_1381,In_704);
nand U474 (N_474,In_1455,In_620);
nand U475 (N_475,In_418,In_3);
and U476 (N_476,In_333,In_883);
and U477 (N_477,In_68,In_124);
nor U478 (N_478,In_251,In_967);
nand U479 (N_479,In_1228,In_614);
nand U480 (N_480,In_407,In_64);
nor U481 (N_481,In_994,In_1405);
nand U482 (N_482,In_1300,In_878);
nor U483 (N_483,In_103,In_8);
nand U484 (N_484,In_1178,In_449);
nand U485 (N_485,In_633,In_1131);
or U486 (N_486,In_681,In_1066);
or U487 (N_487,In_721,In_1105);
nor U488 (N_488,In_795,In_1336);
or U489 (N_489,In_1314,In_1074);
nand U490 (N_490,In_1408,In_1062);
nor U491 (N_491,In_380,In_1235);
or U492 (N_492,In_876,In_1409);
or U493 (N_493,In_591,In_1054);
or U494 (N_494,In_1202,In_752);
nand U495 (N_495,In_397,In_944);
or U496 (N_496,In_1288,In_1199);
or U497 (N_497,In_354,In_284);
xnor U498 (N_498,In_279,In_1268);
nand U499 (N_499,In_1015,In_742);
and U500 (N_500,In_1421,In_786);
nand U501 (N_501,In_592,In_1175);
and U502 (N_502,In_406,In_105);
or U503 (N_503,In_758,In_1122);
or U504 (N_504,In_798,In_249);
nand U505 (N_505,In_1423,In_676);
and U506 (N_506,In_243,In_860);
nand U507 (N_507,In_1143,In_722);
nor U508 (N_508,In_532,In_1349);
and U509 (N_509,In_128,In_991);
and U510 (N_510,In_955,In_1141);
and U511 (N_511,In_759,In_982);
nor U512 (N_512,In_42,In_446);
and U513 (N_513,In_302,In_456);
and U514 (N_514,In_90,In_1431);
and U515 (N_515,In_437,In_551);
or U516 (N_516,In_1243,In_1081);
xnor U517 (N_517,In_129,In_1304);
nor U518 (N_518,In_421,In_104);
and U519 (N_519,In_266,In_658);
and U520 (N_520,In_654,In_642);
or U521 (N_521,In_513,In_1350);
nor U522 (N_522,In_219,In_25);
or U523 (N_523,In_312,In_1289);
or U524 (N_524,In_1482,In_443);
nor U525 (N_525,In_849,In_414);
nor U526 (N_526,In_990,In_420);
and U527 (N_527,In_1097,In_923);
and U528 (N_528,In_1104,In_1209);
or U529 (N_529,In_770,In_419);
and U530 (N_530,In_521,In_841);
nand U531 (N_531,In_91,In_558);
nor U532 (N_532,In_899,In_897);
or U533 (N_533,In_1192,In_877);
nand U534 (N_534,In_268,In_1348);
and U535 (N_535,In_1462,In_1087);
and U536 (N_536,In_1456,In_673);
and U537 (N_537,In_389,In_119);
and U538 (N_538,In_744,In_26);
or U539 (N_539,In_1007,In_1479);
xnor U540 (N_540,In_769,In_508);
nor U541 (N_541,In_788,In_1484);
and U542 (N_542,In_1450,In_1035);
nand U543 (N_543,In_151,In_530);
or U544 (N_544,In_455,In_189);
and U545 (N_545,In_1221,In_415);
nor U546 (N_546,In_202,In_733);
and U547 (N_547,In_1156,In_1388);
nand U548 (N_548,In_584,In_888);
or U549 (N_549,In_948,In_15);
nor U550 (N_550,In_656,In_688);
nand U551 (N_551,In_96,In_507);
or U552 (N_552,In_527,In_922);
or U553 (N_553,In_1179,In_494);
xnor U554 (N_554,In_385,In_200);
and U555 (N_555,In_563,In_296);
nor U556 (N_556,In_1147,In_1266);
nand U557 (N_557,In_1310,In_1316);
nand U558 (N_558,In_428,In_1130);
nor U559 (N_559,In_905,In_234);
xnor U560 (N_560,In_578,In_1017);
nand U561 (N_561,In_425,In_946);
and U562 (N_562,In_323,In_1475);
nand U563 (N_563,In_488,In_574);
nand U564 (N_564,In_1312,In_650);
or U565 (N_565,In_1346,In_1277);
nor U566 (N_566,In_663,In_926);
nor U567 (N_567,In_1400,In_824);
xor U568 (N_568,In_203,In_1203);
nor U569 (N_569,In_1247,In_814);
nor U570 (N_570,In_1480,In_1037);
or U571 (N_571,In_603,In_995);
or U572 (N_572,In_1148,In_695);
nor U573 (N_573,In_12,In_17);
or U574 (N_574,In_346,In_328);
and U575 (N_575,In_484,In_1185);
nand U576 (N_576,In_339,In_1430);
and U577 (N_577,In_562,In_768);
and U578 (N_578,In_1219,In_830);
and U579 (N_579,In_1181,In_481);
nand U580 (N_580,In_371,In_1307);
xnor U581 (N_581,In_170,In_630);
and U582 (N_582,In_316,In_522);
and U583 (N_583,In_980,In_1469);
or U584 (N_584,In_190,In_863);
and U585 (N_585,In_165,In_236);
nand U586 (N_586,In_1072,In_515);
xor U587 (N_587,In_87,In_901);
nor U588 (N_588,In_63,In_1116);
or U589 (N_589,In_1180,In_839);
xnor U590 (N_590,In_1271,In_916);
or U591 (N_591,In_275,In_615);
and U592 (N_592,In_99,In_691);
nor U593 (N_593,In_286,In_37);
nor U594 (N_594,In_736,In_828);
nand U595 (N_595,In_1496,In_1309);
and U596 (N_596,In_29,In_1006);
xnor U597 (N_597,In_83,In_1261);
nand U598 (N_598,In_832,In_729);
or U599 (N_599,In_1324,In_376);
nand U600 (N_600,In_1058,In_1084);
nand U601 (N_601,In_957,In_1113);
and U602 (N_602,In_148,In_1123);
or U603 (N_603,In_1000,In_1371);
or U604 (N_604,In_360,In_715);
nand U605 (N_605,In_270,In_557);
and U606 (N_606,In_386,In_108);
nor U607 (N_607,In_993,In_1089);
nand U608 (N_608,In_1027,In_52);
or U609 (N_609,In_267,In_1091);
or U610 (N_610,In_525,In_14);
nor U611 (N_611,In_694,In_447);
nand U612 (N_612,In_585,In_1444);
nand U613 (N_613,In_1390,In_1485);
nor U614 (N_614,In_805,In_358);
nor U615 (N_615,In_265,In_363);
and U616 (N_616,In_1352,In_1493);
and U617 (N_617,In_903,In_392);
xor U618 (N_618,In_135,In_459);
nor U619 (N_619,In_872,In_1283);
nor U620 (N_620,In_661,In_886);
nand U621 (N_621,In_890,In_1285);
nor U622 (N_622,In_1234,In_1478);
and U623 (N_623,In_869,In_479);
or U624 (N_624,In_228,In_1295);
nor U625 (N_625,In_1011,In_981);
xnor U626 (N_626,In_157,In_93);
or U627 (N_627,In_1005,In_483);
nor U628 (N_628,In_235,In_384);
nand U629 (N_629,In_998,In_1013);
and U630 (N_630,In_533,In_1218);
nor U631 (N_631,In_1442,In_325);
nor U632 (N_632,In_1343,In_732);
and U633 (N_633,In_714,In_1367);
and U634 (N_634,In_367,In_370);
and U635 (N_635,In_1467,In_984);
nand U636 (N_636,In_1200,In_319);
nor U637 (N_637,In_539,In_534);
or U638 (N_638,In_1101,In_375);
and U639 (N_639,In_1328,In_698);
nor U640 (N_640,In_496,In_1497);
nor U641 (N_641,In_1004,In_9);
nor U642 (N_642,In_1359,In_177);
or U643 (N_643,In_403,In_1447);
nor U644 (N_644,In_272,In_947);
nand U645 (N_645,In_278,In_815);
nor U646 (N_646,In_677,In_806);
xnor U647 (N_647,In_465,In_162);
nand U648 (N_648,In_338,In_448);
nor U649 (N_649,In_227,In_258);
nand U650 (N_650,In_38,In_440);
nand U651 (N_651,In_1424,In_953);
nor U652 (N_652,In_760,In_255);
nor U653 (N_653,In_797,In_526);
or U654 (N_654,In_1458,In_1071);
or U655 (N_655,In_1186,In_404);
and U656 (N_656,In_930,In_411);
or U657 (N_657,In_834,In_651);
and U658 (N_658,In_666,In_373);
or U659 (N_659,In_146,In_320);
and U660 (N_660,In_1375,In_166);
and U661 (N_661,In_301,In_1353);
or U662 (N_662,In_1264,In_60);
and U663 (N_663,In_605,In_1499);
nor U664 (N_664,In_871,In_223);
and U665 (N_665,In_155,In_100);
nand U666 (N_666,In_1009,In_735);
or U667 (N_667,In_115,In_1333);
xor U668 (N_668,In_1196,In_1459);
and U669 (N_669,In_1435,In_1461);
or U670 (N_670,In_1303,In_972);
and U671 (N_671,In_351,In_1126);
xor U672 (N_672,In_1427,In_1227);
and U673 (N_673,In_1387,In_1163);
or U674 (N_674,In_1142,In_1019);
and U675 (N_675,In_648,In_1385);
nand U676 (N_676,In_436,In_516);
xnor U677 (N_677,In_445,In_1138);
or U678 (N_678,In_1060,In_1151);
nand U679 (N_679,In_197,In_1380);
xor U680 (N_680,In_906,In_700);
nor U681 (N_681,In_1413,In_699);
or U682 (N_682,In_667,In_153);
and U683 (N_683,In_1416,In_65);
or U684 (N_684,In_778,In_593);
xor U685 (N_685,In_242,In_986);
or U686 (N_686,In_173,In_705);
and U687 (N_687,In_221,In_1010);
nand U688 (N_688,In_512,In_1301);
and U689 (N_689,In_548,In_689);
nand U690 (N_690,In_619,In_174);
or U691 (N_691,In_838,In_1446);
or U692 (N_692,In_450,In_624);
or U693 (N_693,In_2,In_1168);
or U694 (N_694,In_1474,In_950);
or U695 (N_695,In_1195,In_935);
or U696 (N_696,In_825,In_1287);
and U697 (N_697,In_288,In_701);
and U698 (N_698,In_70,In_716);
nor U699 (N_699,In_737,In_979);
nand U700 (N_700,In_1115,In_156);
or U701 (N_701,In_613,In_39);
nor U702 (N_702,In_789,In_726);
or U703 (N_703,In_1297,In_30);
or U704 (N_704,In_50,In_247);
nor U705 (N_705,In_542,In_1344);
nand U706 (N_706,In_1372,In_1166);
or U707 (N_707,In_1008,In_682);
nor U708 (N_708,In_199,In_424);
or U709 (N_709,In_606,In_1046);
and U710 (N_710,In_959,In_501);
nor U711 (N_711,In_836,In_1160);
and U712 (N_712,In_1358,In_1414);
nor U713 (N_713,In_1069,In_882);
nand U714 (N_714,In_628,In_298);
nand U715 (N_715,In_98,In_1118);
or U716 (N_716,In_679,In_851);
and U717 (N_717,In_163,In_422);
and U718 (N_718,In_803,In_313);
or U719 (N_719,In_388,In_58);
or U720 (N_720,In_653,In_833);
nor U721 (N_721,In_734,In_646);
or U722 (N_722,In_1471,In_164);
and U723 (N_723,In_204,In_1067);
or U724 (N_724,In_583,In_191);
and U725 (N_725,In_1379,In_55);
nand U726 (N_726,In_587,In_225);
nand U727 (N_727,In_192,In_887);
or U728 (N_728,In_1238,In_1279);
or U729 (N_729,In_1454,In_1443);
nand U730 (N_730,In_506,In_826);
or U731 (N_731,In_818,In_1395);
xnor U732 (N_732,In_1272,In_575);
and U733 (N_733,In_503,In_1313);
and U734 (N_734,In_1457,In_540);
nor U735 (N_735,In_7,In_467);
or U736 (N_736,In_635,In_537);
nor U737 (N_737,In_1110,In_1012);
nor U738 (N_738,In_273,In_1210);
or U739 (N_739,In_222,In_954);
nand U740 (N_740,In_264,In_544);
nor U741 (N_741,In_497,In_208);
and U742 (N_742,In_1145,In_831);
and U743 (N_743,In_1050,In_120);
nand U744 (N_744,In_1204,In_294);
nand U745 (N_745,In_618,In_130);
and U746 (N_746,In_892,In_936);
nor U747 (N_747,In_873,In_671);
or U748 (N_748,In_1222,In_1090);
xnor U749 (N_749,In_1076,In_357);
and U750 (N_750,In_992,In_604);
and U751 (N_751,In_187,In_1301);
xnor U752 (N_752,In_1109,In_6);
nor U753 (N_753,In_1448,In_177);
and U754 (N_754,In_386,In_737);
nand U755 (N_755,In_512,In_208);
nand U756 (N_756,In_1152,In_880);
or U757 (N_757,In_1184,In_329);
nor U758 (N_758,In_1158,In_1125);
nand U759 (N_759,In_594,In_1186);
or U760 (N_760,In_528,In_765);
and U761 (N_761,In_1228,In_231);
or U762 (N_762,In_1025,In_283);
nor U763 (N_763,In_512,In_995);
nand U764 (N_764,In_573,In_46);
or U765 (N_765,In_171,In_1414);
and U766 (N_766,In_1032,In_706);
and U767 (N_767,In_469,In_220);
nand U768 (N_768,In_1116,In_718);
nor U769 (N_769,In_454,In_941);
and U770 (N_770,In_919,In_561);
nand U771 (N_771,In_414,In_1149);
or U772 (N_772,In_661,In_693);
or U773 (N_773,In_861,In_954);
or U774 (N_774,In_909,In_64);
or U775 (N_775,In_1283,In_121);
nand U776 (N_776,In_907,In_1125);
xor U777 (N_777,In_457,In_913);
xnor U778 (N_778,In_602,In_519);
and U779 (N_779,In_101,In_1251);
xor U780 (N_780,In_511,In_77);
nor U781 (N_781,In_1306,In_798);
and U782 (N_782,In_901,In_86);
and U783 (N_783,In_682,In_595);
nand U784 (N_784,In_1404,In_1228);
or U785 (N_785,In_476,In_658);
and U786 (N_786,In_1118,In_739);
nand U787 (N_787,In_1308,In_917);
or U788 (N_788,In_1106,In_897);
or U789 (N_789,In_1346,In_1021);
nor U790 (N_790,In_456,In_1065);
and U791 (N_791,In_840,In_954);
nor U792 (N_792,In_1051,In_426);
or U793 (N_793,In_990,In_909);
nor U794 (N_794,In_866,In_543);
or U795 (N_795,In_88,In_758);
or U796 (N_796,In_782,In_1220);
xnor U797 (N_797,In_1040,In_1082);
or U798 (N_798,In_1178,In_1044);
nor U799 (N_799,In_341,In_1114);
nand U800 (N_800,In_470,In_823);
nand U801 (N_801,In_560,In_1009);
nor U802 (N_802,In_30,In_222);
xor U803 (N_803,In_366,In_1457);
xnor U804 (N_804,In_1048,In_38);
nand U805 (N_805,In_1176,In_327);
nor U806 (N_806,In_1037,In_1107);
or U807 (N_807,In_693,In_706);
nand U808 (N_808,In_1059,In_1301);
and U809 (N_809,In_1124,In_1044);
or U810 (N_810,In_1368,In_471);
nor U811 (N_811,In_60,In_1430);
or U812 (N_812,In_213,In_1412);
or U813 (N_813,In_367,In_616);
or U814 (N_814,In_202,In_32);
and U815 (N_815,In_688,In_1280);
nand U816 (N_816,In_670,In_1186);
nor U817 (N_817,In_1166,In_788);
nor U818 (N_818,In_228,In_520);
or U819 (N_819,In_683,In_1005);
xor U820 (N_820,In_291,In_1082);
or U821 (N_821,In_571,In_661);
nand U822 (N_822,In_437,In_378);
or U823 (N_823,In_582,In_1139);
nand U824 (N_824,In_1430,In_859);
nor U825 (N_825,In_79,In_1174);
nand U826 (N_826,In_1323,In_910);
nor U827 (N_827,In_477,In_801);
and U828 (N_828,In_918,In_426);
or U829 (N_829,In_493,In_155);
and U830 (N_830,In_495,In_394);
and U831 (N_831,In_1122,In_659);
and U832 (N_832,In_161,In_1238);
nor U833 (N_833,In_1274,In_1142);
xor U834 (N_834,In_1101,In_367);
and U835 (N_835,In_1367,In_1322);
nand U836 (N_836,In_953,In_239);
and U837 (N_837,In_1337,In_255);
or U838 (N_838,In_531,In_97);
nor U839 (N_839,In_991,In_1033);
or U840 (N_840,In_253,In_583);
and U841 (N_841,In_135,In_906);
and U842 (N_842,In_1006,In_1463);
or U843 (N_843,In_1256,In_408);
xor U844 (N_844,In_1062,In_101);
and U845 (N_845,In_225,In_611);
nor U846 (N_846,In_887,In_789);
or U847 (N_847,In_990,In_416);
and U848 (N_848,In_566,In_1450);
nor U849 (N_849,In_538,In_404);
and U850 (N_850,In_734,In_1290);
nor U851 (N_851,In_947,In_864);
xor U852 (N_852,In_303,In_366);
nand U853 (N_853,In_742,In_976);
xnor U854 (N_854,In_24,In_752);
nor U855 (N_855,In_713,In_578);
or U856 (N_856,In_1166,In_647);
nor U857 (N_857,In_1048,In_120);
nor U858 (N_858,In_593,In_808);
nor U859 (N_859,In_483,In_569);
nand U860 (N_860,In_1295,In_1101);
and U861 (N_861,In_685,In_738);
or U862 (N_862,In_593,In_109);
or U863 (N_863,In_532,In_262);
nand U864 (N_864,In_84,In_99);
nand U865 (N_865,In_289,In_1415);
nand U866 (N_866,In_718,In_90);
nand U867 (N_867,In_640,In_800);
nor U868 (N_868,In_1401,In_457);
or U869 (N_869,In_1063,In_333);
and U870 (N_870,In_1342,In_54);
or U871 (N_871,In_369,In_1262);
and U872 (N_872,In_453,In_1361);
nor U873 (N_873,In_1393,In_215);
or U874 (N_874,In_392,In_1430);
nand U875 (N_875,In_108,In_516);
nor U876 (N_876,In_488,In_812);
nand U877 (N_877,In_1227,In_875);
nor U878 (N_878,In_427,In_681);
xnor U879 (N_879,In_254,In_1073);
and U880 (N_880,In_43,In_309);
and U881 (N_881,In_420,In_480);
nand U882 (N_882,In_929,In_11);
and U883 (N_883,In_804,In_275);
or U884 (N_884,In_1331,In_1263);
nor U885 (N_885,In_494,In_1242);
or U886 (N_886,In_792,In_1283);
or U887 (N_887,In_1164,In_590);
or U888 (N_888,In_271,In_443);
or U889 (N_889,In_1119,In_551);
xor U890 (N_890,In_689,In_981);
and U891 (N_891,In_612,In_473);
nand U892 (N_892,In_598,In_1367);
or U893 (N_893,In_434,In_1248);
or U894 (N_894,In_873,In_175);
nand U895 (N_895,In_592,In_204);
and U896 (N_896,In_700,In_863);
nand U897 (N_897,In_380,In_601);
and U898 (N_898,In_798,In_636);
nor U899 (N_899,In_1377,In_1208);
nand U900 (N_900,In_1037,In_820);
or U901 (N_901,In_448,In_382);
nor U902 (N_902,In_400,In_1269);
nand U903 (N_903,In_592,In_1392);
or U904 (N_904,In_693,In_287);
nor U905 (N_905,In_800,In_1370);
nand U906 (N_906,In_1263,In_439);
nand U907 (N_907,In_367,In_18);
nor U908 (N_908,In_1082,In_829);
nand U909 (N_909,In_1023,In_853);
nor U910 (N_910,In_212,In_645);
nor U911 (N_911,In_1450,In_66);
or U912 (N_912,In_868,In_229);
nand U913 (N_913,In_1123,In_259);
nand U914 (N_914,In_1184,In_966);
xnor U915 (N_915,In_868,In_1315);
and U916 (N_916,In_271,In_193);
nand U917 (N_917,In_122,In_1383);
or U918 (N_918,In_765,In_185);
or U919 (N_919,In_52,In_1064);
or U920 (N_920,In_617,In_1383);
or U921 (N_921,In_1060,In_1016);
nand U922 (N_922,In_564,In_1480);
nor U923 (N_923,In_102,In_1453);
or U924 (N_924,In_182,In_1073);
xor U925 (N_925,In_1066,In_1160);
or U926 (N_926,In_1188,In_145);
xor U927 (N_927,In_586,In_551);
or U928 (N_928,In_70,In_83);
and U929 (N_929,In_917,In_1406);
nor U930 (N_930,In_518,In_442);
nand U931 (N_931,In_1376,In_248);
nor U932 (N_932,In_479,In_822);
nand U933 (N_933,In_1300,In_398);
and U934 (N_934,In_1295,In_214);
or U935 (N_935,In_620,In_1174);
or U936 (N_936,In_445,In_691);
and U937 (N_937,In_922,In_148);
nor U938 (N_938,In_1062,In_1349);
nor U939 (N_939,In_1266,In_902);
xor U940 (N_940,In_402,In_307);
nor U941 (N_941,In_447,In_726);
or U942 (N_942,In_1495,In_602);
nor U943 (N_943,In_78,In_567);
and U944 (N_944,In_52,In_224);
or U945 (N_945,In_28,In_699);
and U946 (N_946,In_531,In_1394);
or U947 (N_947,In_497,In_242);
nor U948 (N_948,In_1420,In_414);
nor U949 (N_949,In_1449,In_162);
nand U950 (N_950,In_412,In_943);
nor U951 (N_951,In_1199,In_32);
xnor U952 (N_952,In_1489,In_553);
nand U953 (N_953,In_822,In_1449);
nor U954 (N_954,In_166,In_725);
nand U955 (N_955,In_725,In_1488);
and U956 (N_956,In_330,In_950);
nor U957 (N_957,In_1454,In_822);
xnor U958 (N_958,In_1407,In_1081);
xnor U959 (N_959,In_686,In_943);
or U960 (N_960,In_1121,In_11);
and U961 (N_961,In_897,In_854);
xnor U962 (N_962,In_281,In_156);
or U963 (N_963,In_967,In_48);
nor U964 (N_964,In_458,In_651);
and U965 (N_965,In_575,In_1090);
nor U966 (N_966,In_344,In_1282);
xor U967 (N_967,In_1076,In_709);
xor U968 (N_968,In_944,In_870);
nand U969 (N_969,In_767,In_55);
or U970 (N_970,In_1296,In_867);
nor U971 (N_971,In_1128,In_185);
or U972 (N_972,In_70,In_1447);
nor U973 (N_973,In_1157,In_392);
or U974 (N_974,In_577,In_143);
or U975 (N_975,In_989,In_111);
and U976 (N_976,In_6,In_1234);
nor U977 (N_977,In_300,In_1133);
or U978 (N_978,In_1457,In_1182);
xor U979 (N_979,In_887,In_682);
nor U980 (N_980,In_1166,In_887);
or U981 (N_981,In_1098,In_1325);
nor U982 (N_982,In_1321,In_586);
nand U983 (N_983,In_764,In_752);
or U984 (N_984,In_1252,In_1196);
nor U985 (N_985,In_913,In_1230);
xor U986 (N_986,In_1162,In_984);
or U987 (N_987,In_724,In_989);
nand U988 (N_988,In_548,In_227);
and U989 (N_989,In_1057,In_88);
and U990 (N_990,In_1324,In_884);
or U991 (N_991,In_344,In_1445);
and U992 (N_992,In_1313,In_595);
or U993 (N_993,In_825,In_595);
and U994 (N_994,In_1487,In_1094);
or U995 (N_995,In_671,In_1425);
xnor U996 (N_996,In_582,In_513);
xor U997 (N_997,In_95,In_660);
and U998 (N_998,In_926,In_1400);
and U999 (N_999,In_1211,In_1311);
and U1000 (N_1000,In_979,In_199);
or U1001 (N_1001,In_1091,In_880);
or U1002 (N_1002,In_941,In_662);
or U1003 (N_1003,In_706,In_849);
or U1004 (N_1004,In_641,In_850);
xor U1005 (N_1005,In_1068,In_1137);
and U1006 (N_1006,In_959,In_573);
and U1007 (N_1007,In_135,In_479);
nand U1008 (N_1008,In_450,In_809);
nand U1009 (N_1009,In_407,In_1449);
nor U1010 (N_1010,In_557,In_631);
and U1011 (N_1011,In_1070,In_734);
or U1012 (N_1012,In_558,In_1168);
nand U1013 (N_1013,In_392,In_97);
nand U1014 (N_1014,In_1018,In_288);
and U1015 (N_1015,In_1177,In_701);
xor U1016 (N_1016,In_1269,In_389);
or U1017 (N_1017,In_688,In_965);
xor U1018 (N_1018,In_1442,In_7);
or U1019 (N_1019,In_776,In_1469);
nand U1020 (N_1020,In_307,In_830);
and U1021 (N_1021,In_616,In_1266);
nand U1022 (N_1022,In_1359,In_249);
nor U1023 (N_1023,In_677,In_542);
or U1024 (N_1024,In_671,In_395);
nand U1025 (N_1025,In_298,In_1474);
nor U1026 (N_1026,In_17,In_797);
xnor U1027 (N_1027,In_597,In_1120);
nor U1028 (N_1028,In_1274,In_955);
or U1029 (N_1029,In_1215,In_614);
xnor U1030 (N_1030,In_687,In_699);
and U1031 (N_1031,In_1328,In_1448);
or U1032 (N_1032,In_16,In_612);
and U1033 (N_1033,In_425,In_978);
nand U1034 (N_1034,In_1118,In_1389);
xnor U1035 (N_1035,In_364,In_272);
nand U1036 (N_1036,In_1052,In_372);
and U1037 (N_1037,In_387,In_1267);
xor U1038 (N_1038,In_1305,In_709);
xor U1039 (N_1039,In_822,In_301);
and U1040 (N_1040,In_860,In_1295);
and U1041 (N_1041,In_395,In_567);
nand U1042 (N_1042,In_514,In_524);
nand U1043 (N_1043,In_386,In_73);
and U1044 (N_1044,In_872,In_13);
nand U1045 (N_1045,In_1013,In_338);
nor U1046 (N_1046,In_1307,In_358);
nand U1047 (N_1047,In_722,In_97);
nor U1048 (N_1048,In_539,In_474);
nor U1049 (N_1049,In_1413,In_1022);
nor U1050 (N_1050,In_1211,In_1333);
and U1051 (N_1051,In_184,In_214);
xor U1052 (N_1052,In_549,In_1459);
or U1053 (N_1053,In_943,In_1140);
nor U1054 (N_1054,In_219,In_1270);
xor U1055 (N_1055,In_913,In_1442);
xnor U1056 (N_1056,In_982,In_757);
and U1057 (N_1057,In_593,In_749);
and U1058 (N_1058,In_349,In_541);
and U1059 (N_1059,In_773,In_239);
nor U1060 (N_1060,In_422,In_190);
or U1061 (N_1061,In_929,In_1414);
nand U1062 (N_1062,In_861,In_533);
or U1063 (N_1063,In_1378,In_441);
or U1064 (N_1064,In_276,In_861);
or U1065 (N_1065,In_1161,In_119);
and U1066 (N_1066,In_1460,In_399);
nor U1067 (N_1067,In_1491,In_538);
xor U1068 (N_1068,In_276,In_926);
nand U1069 (N_1069,In_500,In_892);
or U1070 (N_1070,In_146,In_784);
or U1071 (N_1071,In_1155,In_896);
or U1072 (N_1072,In_1291,In_79);
and U1073 (N_1073,In_970,In_784);
and U1074 (N_1074,In_1315,In_788);
and U1075 (N_1075,In_696,In_393);
xnor U1076 (N_1076,In_776,In_1353);
nand U1077 (N_1077,In_561,In_503);
and U1078 (N_1078,In_256,In_415);
nor U1079 (N_1079,In_1406,In_162);
nand U1080 (N_1080,In_804,In_1016);
xnor U1081 (N_1081,In_529,In_344);
and U1082 (N_1082,In_214,In_909);
and U1083 (N_1083,In_736,In_680);
or U1084 (N_1084,In_736,In_427);
xor U1085 (N_1085,In_981,In_1334);
xnor U1086 (N_1086,In_1258,In_229);
nor U1087 (N_1087,In_143,In_798);
nor U1088 (N_1088,In_489,In_48);
nor U1089 (N_1089,In_1395,In_1471);
nor U1090 (N_1090,In_386,In_1397);
and U1091 (N_1091,In_86,In_479);
or U1092 (N_1092,In_166,In_432);
nor U1093 (N_1093,In_686,In_1318);
nand U1094 (N_1094,In_1045,In_833);
and U1095 (N_1095,In_87,In_956);
nor U1096 (N_1096,In_1153,In_385);
nand U1097 (N_1097,In_938,In_1229);
or U1098 (N_1098,In_403,In_450);
or U1099 (N_1099,In_165,In_989);
or U1100 (N_1100,In_709,In_394);
or U1101 (N_1101,In_851,In_53);
nand U1102 (N_1102,In_758,In_710);
and U1103 (N_1103,In_844,In_356);
and U1104 (N_1104,In_1073,In_1365);
and U1105 (N_1105,In_496,In_393);
nand U1106 (N_1106,In_984,In_1373);
nor U1107 (N_1107,In_1468,In_1064);
or U1108 (N_1108,In_1215,In_460);
nand U1109 (N_1109,In_650,In_644);
nor U1110 (N_1110,In_1171,In_162);
or U1111 (N_1111,In_122,In_35);
nand U1112 (N_1112,In_135,In_1018);
and U1113 (N_1113,In_690,In_1327);
and U1114 (N_1114,In_490,In_960);
nand U1115 (N_1115,In_1406,In_425);
nand U1116 (N_1116,In_1283,In_71);
or U1117 (N_1117,In_680,In_1470);
nand U1118 (N_1118,In_775,In_339);
or U1119 (N_1119,In_871,In_348);
and U1120 (N_1120,In_1273,In_832);
nand U1121 (N_1121,In_1219,In_1098);
and U1122 (N_1122,In_883,In_544);
or U1123 (N_1123,In_700,In_986);
nand U1124 (N_1124,In_650,In_1119);
and U1125 (N_1125,In_803,In_267);
and U1126 (N_1126,In_1324,In_741);
or U1127 (N_1127,In_869,In_1271);
and U1128 (N_1128,In_1442,In_974);
or U1129 (N_1129,In_1145,In_383);
and U1130 (N_1130,In_926,In_137);
or U1131 (N_1131,In_1294,In_205);
nor U1132 (N_1132,In_630,In_825);
and U1133 (N_1133,In_1362,In_1449);
nor U1134 (N_1134,In_694,In_63);
or U1135 (N_1135,In_1004,In_403);
and U1136 (N_1136,In_1028,In_1111);
xnor U1137 (N_1137,In_209,In_799);
and U1138 (N_1138,In_1215,In_36);
or U1139 (N_1139,In_1486,In_1033);
and U1140 (N_1140,In_876,In_618);
and U1141 (N_1141,In_1284,In_149);
nand U1142 (N_1142,In_491,In_540);
xor U1143 (N_1143,In_218,In_846);
nor U1144 (N_1144,In_410,In_1173);
nor U1145 (N_1145,In_1175,In_293);
and U1146 (N_1146,In_638,In_210);
or U1147 (N_1147,In_1432,In_1302);
or U1148 (N_1148,In_303,In_496);
and U1149 (N_1149,In_286,In_34);
nor U1150 (N_1150,In_896,In_1422);
or U1151 (N_1151,In_671,In_1240);
nor U1152 (N_1152,In_464,In_1182);
nand U1153 (N_1153,In_330,In_1083);
or U1154 (N_1154,In_837,In_928);
xor U1155 (N_1155,In_1145,In_392);
nand U1156 (N_1156,In_675,In_158);
nor U1157 (N_1157,In_784,In_1210);
nand U1158 (N_1158,In_896,In_1002);
or U1159 (N_1159,In_161,In_1463);
nor U1160 (N_1160,In_646,In_958);
or U1161 (N_1161,In_575,In_1023);
or U1162 (N_1162,In_129,In_407);
nand U1163 (N_1163,In_696,In_1324);
or U1164 (N_1164,In_903,In_250);
nand U1165 (N_1165,In_896,In_494);
and U1166 (N_1166,In_319,In_282);
or U1167 (N_1167,In_1117,In_1170);
and U1168 (N_1168,In_339,In_756);
or U1169 (N_1169,In_469,In_664);
and U1170 (N_1170,In_995,In_1299);
or U1171 (N_1171,In_1019,In_100);
nand U1172 (N_1172,In_1061,In_768);
and U1173 (N_1173,In_193,In_1201);
or U1174 (N_1174,In_885,In_163);
and U1175 (N_1175,In_1345,In_15);
and U1176 (N_1176,In_13,In_1027);
nand U1177 (N_1177,In_689,In_801);
or U1178 (N_1178,In_698,In_1309);
nor U1179 (N_1179,In_93,In_73);
nor U1180 (N_1180,In_1315,In_943);
xor U1181 (N_1181,In_478,In_428);
or U1182 (N_1182,In_795,In_1055);
or U1183 (N_1183,In_852,In_105);
or U1184 (N_1184,In_1169,In_997);
and U1185 (N_1185,In_702,In_1251);
xor U1186 (N_1186,In_563,In_1324);
nand U1187 (N_1187,In_810,In_1226);
nor U1188 (N_1188,In_291,In_66);
nor U1189 (N_1189,In_312,In_335);
or U1190 (N_1190,In_598,In_968);
or U1191 (N_1191,In_203,In_1063);
nand U1192 (N_1192,In_244,In_475);
and U1193 (N_1193,In_1313,In_1345);
nand U1194 (N_1194,In_1108,In_81);
and U1195 (N_1195,In_167,In_1444);
and U1196 (N_1196,In_1278,In_1129);
and U1197 (N_1197,In_1222,In_841);
or U1198 (N_1198,In_43,In_1380);
and U1199 (N_1199,In_198,In_117);
nand U1200 (N_1200,In_1240,In_387);
and U1201 (N_1201,In_600,In_1336);
and U1202 (N_1202,In_1159,In_453);
or U1203 (N_1203,In_406,In_1355);
and U1204 (N_1204,In_1138,In_1162);
xnor U1205 (N_1205,In_578,In_188);
or U1206 (N_1206,In_1021,In_1371);
nor U1207 (N_1207,In_942,In_1118);
and U1208 (N_1208,In_202,In_349);
or U1209 (N_1209,In_428,In_976);
xnor U1210 (N_1210,In_1182,In_46);
nor U1211 (N_1211,In_76,In_567);
nor U1212 (N_1212,In_1113,In_334);
xor U1213 (N_1213,In_860,In_1194);
nand U1214 (N_1214,In_92,In_265);
or U1215 (N_1215,In_1009,In_18);
or U1216 (N_1216,In_426,In_940);
nand U1217 (N_1217,In_129,In_244);
nand U1218 (N_1218,In_1022,In_448);
and U1219 (N_1219,In_111,In_252);
or U1220 (N_1220,In_852,In_1054);
nor U1221 (N_1221,In_1390,In_944);
nand U1222 (N_1222,In_1124,In_1177);
nand U1223 (N_1223,In_649,In_533);
nand U1224 (N_1224,In_726,In_1386);
nor U1225 (N_1225,In_1496,In_126);
nor U1226 (N_1226,In_819,In_1230);
xnor U1227 (N_1227,In_341,In_398);
nand U1228 (N_1228,In_756,In_412);
nor U1229 (N_1229,In_0,In_610);
nor U1230 (N_1230,In_1389,In_363);
or U1231 (N_1231,In_147,In_207);
nand U1232 (N_1232,In_1113,In_1372);
nor U1233 (N_1233,In_40,In_925);
nor U1234 (N_1234,In_1354,In_155);
xnor U1235 (N_1235,In_456,In_1024);
xor U1236 (N_1236,In_718,In_575);
or U1237 (N_1237,In_599,In_517);
or U1238 (N_1238,In_823,In_1386);
and U1239 (N_1239,In_1212,In_691);
nor U1240 (N_1240,In_723,In_487);
nand U1241 (N_1241,In_746,In_7);
and U1242 (N_1242,In_977,In_968);
and U1243 (N_1243,In_974,In_527);
xor U1244 (N_1244,In_1156,In_442);
and U1245 (N_1245,In_1118,In_433);
xnor U1246 (N_1246,In_498,In_172);
nor U1247 (N_1247,In_1096,In_183);
nor U1248 (N_1248,In_1077,In_150);
nand U1249 (N_1249,In_155,In_1306);
or U1250 (N_1250,In_649,In_775);
xor U1251 (N_1251,In_858,In_780);
or U1252 (N_1252,In_1099,In_922);
or U1253 (N_1253,In_1200,In_220);
and U1254 (N_1254,In_19,In_630);
nand U1255 (N_1255,In_107,In_1202);
xor U1256 (N_1256,In_853,In_1020);
nor U1257 (N_1257,In_139,In_1264);
nor U1258 (N_1258,In_442,In_704);
and U1259 (N_1259,In_1207,In_597);
nand U1260 (N_1260,In_711,In_1403);
nor U1261 (N_1261,In_888,In_164);
or U1262 (N_1262,In_720,In_46);
nand U1263 (N_1263,In_840,In_1150);
nand U1264 (N_1264,In_197,In_81);
and U1265 (N_1265,In_27,In_440);
or U1266 (N_1266,In_1421,In_1361);
nand U1267 (N_1267,In_1302,In_1350);
nand U1268 (N_1268,In_681,In_623);
and U1269 (N_1269,In_1452,In_302);
xnor U1270 (N_1270,In_1221,In_751);
nand U1271 (N_1271,In_550,In_1353);
or U1272 (N_1272,In_1152,In_596);
and U1273 (N_1273,In_753,In_515);
xnor U1274 (N_1274,In_1318,In_629);
nand U1275 (N_1275,In_227,In_83);
xor U1276 (N_1276,In_1428,In_591);
nor U1277 (N_1277,In_432,In_1315);
xor U1278 (N_1278,In_967,In_677);
and U1279 (N_1279,In_259,In_363);
xnor U1280 (N_1280,In_764,In_731);
or U1281 (N_1281,In_25,In_1080);
or U1282 (N_1282,In_180,In_243);
and U1283 (N_1283,In_497,In_448);
nand U1284 (N_1284,In_59,In_866);
xnor U1285 (N_1285,In_1477,In_1062);
nor U1286 (N_1286,In_1401,In_973);
nand U1287 (N_1287,In_1331,In_702);
nor U1288 (N_1288,In_418,In_1230);
nor U1289 (N_1289,In_1292,In_53);
and U1290 (N_1290,In_145,In_1085);
nor U1291 (N_1291,In_888,In_1234);
nor U1292 (N_1292,In_1434,In_1044);
xnor U1293 (N_1293,In_1432,In_388);
nor U1294 (N_1294,In_700,In_279);
xnor U1295 (N_1295,In_250,In_419);
xor U1296 (N_1296,In_776,In_870);
or U1297 (N_1297,In_912,In_528);
or U1298 (N_1298,In_1314,In_555);
or U1299 (N_1299,In_1005,In_1334);
nand U1300 (N_1300,In_246,In_777);
or U1301 (N_1301,In_934,In_564);
nor U1302 (N_1302,In_568,In_931);
and U1303 (N_1303,In_1189,In_1021);
nor U1304 (N_1304,In_811,In_396);
and U1305 (N_1305,In_142,In_1);
nand U1306 (N_1306,In_800,In_1173);
and U1307 (N_1307,In_9,In_827);
and U1308 (N_1308,In_175,In_1285);
nor U1309 (N_1309,In_386,In_1170);
or U1310 (N_1310,In_495,In_832);
nand U1311 (N_1311,In_794,In_1479);
or U1312 (N_1312,In_846,In_1273);
nor U1313 (N_1313,In_1495,In_466);
nand U1314 (N_1314,In_232,In_685);
nand U1315 (N_1315,In_752,In_602);
and U1316 (N_1316,In_1037,In_1410);
and U1317 (N_1317,In_792,In_709);
nand U1318 (N_1318,In_278,In_508);
nor U1319 (N_1319,In_1200,In_801);
and U1320 (N_1320,In_499,In_1269);
nor U1321 (N_1321,In_100,In_959);
nand U1322 (N_1322,In_599,In_1337);
or U1323 (N_1323,In_103,In_169);
or U1324 (N_1324,In_910,In_665);
or U1325 (N_1325,In_1090,In_921);
nor U1326 (N_1326,In_1436,In_861);
nand U1327 (N_1327,In_274,In_677);
nor U1328 (N_1328,In_753,In_583);
or U1329 (N_1329,In_535,In_473);
nor U1330 (N_1330,In_650,In_720);
nor U1331 (N_1331,In_927,In_584);
and U1332 (N_1332,In_971,In_520);
or U1333 (N_1333,In_434,In_1216);
nand U1334 (N_1334,In_479,In_1235);
or U1335 (N_1335,In_840,In_1461);
and U1336 (N_1336,In_1396,In_1157);
and U1337 (N_1337,In_1027,In_219);
and U1338 (N_1338,In_367,In_767);
and U1339 (N_1339,In_1359,In_1282);
xnor U1340 (N_1340,In_580,In_255);
nand U1341 (N_1341,In_1189,In_1044);
and U1342 (N_1342,In_377,In_179);
or U1343 (N_1343,In_366,In_777);
nand U1344 (N_1344,In_173,In_1031);
nor U1345 (N_1345,In_843,In_35);
or U1346 (N_1346,In_672,In_222);
and U1347 (N_1347,In_732,In_1338);
nand U1348 (N_1348,In_1129,In_217);
nor U1349 (N_1349,In_26,In_902);
xnor U1350 (N_1350,In_750,In_1009);
and U1351 (N_1351,In_398,In_1071);
or U1352 (N_1352,In_365,In_510);
nor U1353 (N_1353,In_1357,In_1155);
nand U1354 (N_1354,In_158,In_878);
nand U1355 (N_1355,In_104,In_38);
or U1356 (N_1356,In_1260,In_604);
nand U1357 (N_1357,In_252,In_378);
nor U1358 (N_1358,In_641,In_1067);
nand U1359 (N_1359,In_872,In_1341);
xnor U1360 (N_1360,In_751,In_928);
nor U1361 (N_1361,In_933,In_1142);
nor U1362 (N_1362,In_1257,In_657);
nor U1363 (N_1363,In_123,In_483);
and U1364 (N_1364,In_263,In_1162);
xor U1365 (N_1365,In_1246,In_318);
and U1366 (N_1366,In_635,In_346);
nor U1367 (N_1367,In_1361,In_763);
or U1368 (N_1368,In_35,In_1022);
or U1369 (N_1369,In_957,In_663);
nor U1370 (N_1370,In_1112,In_905);
and U1371 (N_1371,In_254,In_1443);
nor U1372 (N_1372,In_1138,In_1277);
or U1373 (N_1373,In_1317,In_858);
and U1374 (N_1374,In_377,In_463);
nor U1375 (N_1375,In_526,In_841);
or U1376 (N_1376,In_448,In_1000);
nor U1377 (N_1377,In_580,In_845);
or U1378 (N_1378,In_48,In_1192);
and U1379 (N_1379,In_1241,In_1427);
nor U1380 (N_1380,In_92,In_854);
and U1381 (N_1381,In_230,In_855);
and U1382 (N_1382,In_1315,In_1329);
nor U1383 (N_1383,In_1235,In_632);
nand U1384 (N_1384,In_342,In_643);
nand U1385 (N_1385,In_1493,In_582);
xnor U1386 (N_1386,In_1092,In_482);
nand U1387 (N_1387,In_105,In_1094);
or U1388 (N_1388,In_1335,In_910);
and U1389 (N_1389,In_864,In_532);
nand U1390 (N_1390,In_433,In_1222);
and U1391 (N_1391,In_871,In_1196);
nor U1392 (N_1392,In_153,In_1278);
or U1393 (N_1393,In_173,In_140);
nor U1394 (N_1394,In_923,In_1153);
or U1395 (N_1395,In_1272,In_1279);
nand U1396 (N_1396,In_687,In_459);
and U1397 (N_1397,In_5,In_1373);
or U1398 (N_1398,In_1349,In_714);
nand U1399 (N_1399,In_615,In_134);
xor U1400 (N_1400,In_994,In_1130);
nand U1401 (N_1401,In_858,In_1231);
or U1402 (N_1402,In_0,In_1304);
and U1403 (N_1403,In_716,In_118);
nand U1404 (N_1404,In_689,In_329);
nor U1405 (N_1405,In_38,In_103);
nor U1406 (N_1406,In_572,In_1006);
or U1407 (N_1407,In_1055,In_929);
and U1408 (N_1408,In_1429,In_1377);
nand U1409 (N_1409,In_157,In_579);
or U1410 (N_1410,In_687,In_669);
nor U1411 (N_1411,In_424,In_1138);
and U1412 (N_1412,In_621,In_337);
nor U1413 (N_1413,In_1005,In_1285);
nand U1414 (N_1414,In_1171,In_482);
or U1415 (N_1415,In_1269,In_1443);
nor U1416 (N_1416,In_917,In_1443);
nor U1417 (N_1417,In_1140,In_975);
xor U1418 (N_1418,In_1166,In_843);
nand U1419 (N_1419,In_1026,In_1358);
nand U1420 (N_1420,In_887,In_1139);
or U1421 (N_1421,In_35,In_456);
nor U1422 (N_1422,In_194,In_687);
nand U1423 (N_1423,In_1241,In_1485);
or U1424 (N_1424,In_489,In_54);
nand U1425 (N_1425,In_71,In_1299);
or U1426 (N_1426,In_183,In_914);
or U1427 (N_1427,In_834,In_93);
or U1428 (N_1428,In_627,In_391);
nor U1429 (N_1429,In_1145,In_410);
or U1430 (N_1430,In_1248,In_481);
nand U1431 (N_1431,In_1017,In_320);
nand U1432 (N_1432,In_1431,In_620);
or U1433 (N_1433,In_645,In_1017);
nand U1434 (N_1434,In_583,In_367);
nand U1435 (N_1435,In_972,In_233);
and U1436 (N_1436,In_479,In_1493);
nand U1437 (N_1437,In_1467,In_1189);
xnor U1438 (N_1438,In_186,In_881);
nand U1439 (N_1439,In_1444,In_552);
nand U1440 (N_1440,In_196,In_640);
and U1441 (N_1441,In_1255,In_1119);
or U1442 (N_1442,In_559,In_99);
nor U1443 (N_1443,In_1494,In_1034);
nor U1444 (N_1444,In_907,In_1301);
nor U1445 (N_1445,In_1246,In_234);
nand U1446 (N_1446,In_1042,In_337);
nand U1447 (N_1447,In_128,In_174);
nor U1448 (N_1448,In_128,In_712);
nand U1449 (N_1449,In_744,In_198);
nand U1450 (N_1450,In_896,In_3);
nor U1451 (N_1451,In_154,In_1256);
nor U1452 (N_1452,In_92,In_826);
and U1453 (N_1453,In_22,In_1314);
and U1454 (N_1454,In_1193,In_744);
and U1455 (N_1455,In_597,In_979);
and U1456 (N_1456,In_652,In_896);
nand U1457 (N_1457,In_1054,In_855);
and U1458 (N_1458,In_1378,In_923);
or U1459 (N_1459,In_1290,In_445);
and U1460 (N_1460,In_1420,In_626);
and U1461 (N_1461,In_1291,In_1081);
xor U1462 (N_1462,In_199,In_940);
and U1463 (N_1463,In_31,In_1167);
nor U1464 (N_1464,In_1380,In_1158);
and U1465 (N_1465,In_1498,In_1426);
and U1466 (N_1466,In_193,In_322);
nand U1467 (N_1467,In_1457,In_219);
or U1468 (N_1468,In_1038,In_1112);
nand U1469 (N_1469,In_81,In_890);
xnor U1470 (N_1470,In_826,In_173);
nor U1471 (N_1471,In_230,In_282);
nor U1472 (N_1472,In_1390,In_1364);
nor U1473 (N_1473,In_398,In_889);
and U1474 (N_1474,In_912,In_33);
nor U1475 (N_1475,In_1068,In_716);
nand U1476 (N_1476,In_1140,In_1353);
nand U1477 (N_1477,In_1126,In_324);
and U1478 (N_1478,In_1018,In_1367);
nand U1479 (N_1479,In_88,In_1222);
or U1480 (N_1480,In_315,In_533);
nand U1481 (N_1481,In_279,In_1180);
and U1482 (N_1482,In_9,In_943);
nor U1483 (N_1483,In_1441,In_604);
and U1484 (N_1484,In_1054,In_194);
nor U1485 (N_1485,In_1288,In_916);
nand U1486 (N_1486,In_785,In_839);
nand U1487 (N_1487,In_435,In_1349);
and U1488 (N_1488,In_1133,In_1276);
nand U1489 (N_1489,In_1073,In_1291);
nand U1490 (N_1490,In_1215,In_1231);
or U1491 (N_1491,In_1222,In_1304);
xor U1492 (N_1492,In_896,In_953);
xnor U1493 (N_1493,In_942,In_330);
nand U1494 (N_1494,In_653,In_171);
nor U1495 (N_1495,In_1034,In_821);
nand U1496 (N_1496,In_1310,In_1360);
nand U1497 (N_1497,In_252,In_55);
and U1498 (N_1498,In_354,In_597);
and U1499 (N_1499,In_67,In_816);
or U1500 (N_1500,In_515,In_265);
nor U1501 (N_1501,In_308,In_1344);
and U1502 (N_1502,In_1398,In_353);
nor U1503 (N_1503,In_1406,In_1124);
and U1504 (N_1504,In_446,In_1141);
nand U1505 (N_1505,In_648,In_148);
nor U1506 (N_1506,In_322,In_1410);
nand U1507 (N_1507,In_1141,In_1386);
nand U1508 (N_1508,In_20,In_435);
nor U1509 (N_1509,In_1387,In_164);
or U1510 (N_1510,In_1079,In_316);
and U1511 (N_1511,In_1039,In_841);
and U1512 (N_1512,In_96,In_354);
nor U1513 (N_1513,In_1412,In_883);
and U1514 (N_1514,In_1478,In_259);
nor U1515 (N_1515,In_1474,In_1445);
nand U1516 (N_1516,In_1077,In_1020);
or U1517 (N_1517,In_1292,In_993);
or U1518 (N_1518,In_407,In_1356);
nand U1519 (N_1519,In_1487,In_436);
or U1520 (N_1520,In_656,In_189);
nor U1521 (N_1521,In_436,In_829);
nor U1522 (N_1522,In_682,In_1105);
and U1523 (N_1523,In_336,In_593);
nor U1524 (N_1524,In_1473,In_764);
and U1525 (N_1525,In_782,In_332);
nand U1526 (N_1526,In_995,In_167);
and U1527 (N_1527,In_270,In_1313);
and U1528 (N_1528,In_1271,In_1383);
nand U1529 (N_1529,In_1196,In_429);
or U1530 (N_1530,In_1058,In_727);
and U1531 (N_1531,In_1064,In_357);
or U1532 (N_1532,In_1304,In_170);
nand U1533 (N_1533,In_1319,In_548);
xnor U1534 (N_1534,In_563,In_290);
xnor U1535 (N_1535,In_1401,In_1106);
xor U1536 (N_1536,In_1357,In_1004);
and U1537 (N_1537,In_1066,In_1127);
nor U1538 (N_1538,In_714,In_10);
nand U1539 (N_1539,In_647,In_863);
nand U1540 (N_1540,In_707,In_446);
nor U1541 (N_1541,In_1050,In_923);
xor U1542 (N_1542,In_921,In_1045);
nand U1543 (N_1543,In_130,In_1378);
nor U1544 (N_1544,In_1177,In_84);
or U1545 (N_1545,In_188,In_1331);
or U1546 (N_1546,In_692,In_761);
and U1547 (N_1547,In_767,In_681);
nand U1548 (N_1548,In_1118,In_1175);
or U1549 (N_1549,In_1189,In_1217);
xnor U1550 (N_1550,In_1018,In_625);
and U1551 (N_1551,In_364,In_107);
or U1552 (N_1552,In_1489,In_899);
nor U1553 (N_1553,In_186,In_571);
or U1554 (N_1554,In_1188,In_638);
and U1555 (N_1555,In_212,In_865);
or U1556 (N_1556,In_1079,In_623);
nand U1557 (N_1557,In_652,In_1369);
and U1558 (N_1558,In_710,In_910);
nand U1559 (N_1559,In_662,In_877);
xor U1560 (N_1560,In_242,In_1172);
and U1561 (N_1561,In_282,In_1254);
or U1562 (N_1562,In_1069,In_1016);
or U1563 (N_1563,In_417,In_568);
nand U1564 (N_1564,In_859,In_652);
nand U1565 (N_1565,In_1306,In_463);
nand U1566 (N_1566,In_335,In_1374);
xor U1567 (N_1567,In_1365,In_1352);
nor U1568 (N_1568,In_111,In_1226);
xnor U1569 (N_1569,In_1308,In_1123);
or U1570 (N_1570,In_1405,In_1210);
nand U1571 (N_1571,In_899,In_1478);
nor U1572 (N_1572,In_1378,In_179);
xnor U1573 (N_1573,In_1195,In_512);
nand U1574 (N_1574,In_106,In_1468);
nand U1575 (N_1575,In_1416,In_519);
nand U1576 (N_1576,In_442,In_245);
or U1577 (N_1577,In_188,In_302);
nor U1578 (N_1578,In_482,In_192);
nand U1579 (N_1579,In_419,In_856);
nand U1580 (N_1580,In_1456,In_1399);
or U1581 (N_1581,In_337,In_453);
and U1582 (N_1582,In_747,In_1247);
and U1583 (N_1583,In_232,In_1300);
or U1584 (N_1584,In_909,In_393);
or U1585 (N_1585,In_1243,In_369);
and U1586 (N_1586,In_462,In_1252);
or U1587 (N_1587,In_976,In_541);
xnor U1588 (N_1588,In_1306,In_275);
xnor U1589 (N_1589,In_1151,In_850);
and U1590 (N_1590,In_1354,In_1357);
nand U1591 (N_1591,In_414,In_234);
and U1592 (N_1592,In_1310,In_1416);
nand U1593 (N_1593,In_219,In_1326);
or U1594 (N_1594,In_1172,In_192);
nand U1595 (N_1595,In_341,In_525);
nor U1596 (N_1596,In_743,In_1032);
nor U1597 (N_1597,In_1499,In_754);
xnor U1598 (N_1598,In_735,In_62);
or U1599 (N_1599,In_47,In_1215);
xor U1600 (N_1600,In_702,In_777);
nor U1601 (N_1601,In_1100,In_837);
and U1602 (N_1602,In_1277,In_762);
nor U1603 (N_1603,In_354,In_210);
or U1604 (N_1604,In_8,In_808);
or U1605 (N_1605,In_613,In_1054);
and U1606 (N_1606,In_945,In_1025);
or U1607 (N_1607,In_110,In_671);
nand U1608 (N_1608,In_1301,In_664);
nor U1609 (N_1609,In_1386,In_271);
nor U1610 (N_1610,In_1009,In_1168);
and U1611 (N_1611,In_1145,In_406);
and U1612 (N_1612,In_1484,In_90);
nand U1613 (N_1613,In_1206,In_26);
xnor U1614 (N_1614,In_225,In_407);
nand U1615 (N_1615,In_1066,In_399);
nor U1616 (N_1616,In_105,In_324);
nor U1617 (N_1617,In_858,In_139);
and U1618 (N_1618,In_848,In_374);
xnor U1619 (N_1619,In_998,In_1335);
nand U1620 (N_1620,In_574,In_13);
nor U1621 (N_1621,In_889,In_1488);
and U1622 (N_1622,In_1261,In_1090);
or U1623 (N_1623,In_999,In_942);
or U1624 (N_1624,In_1480,In_1093);
nand U1625 (N_1625,In_1236,In_535);
and U1626 (N_1626,In_1469,In_1299);
nand U1627 (N_1627,In_1452,In_76);
or U1628 (N_1628,In_74,In_248);
nand U1629 (N_1629,In_281,In_1055);
or U1630 (N_1630,In_90,In_1393);
and U1631 (N_1631,In_213,In_1492);
or U1632 (N_1632,In_20,In_1243);
nand U1633 (N_1633,In_769,In_552);
and U1634 (N_1634,In_1300,In_1293);
or U1635 (N_1635,In_173,In_837);
and U1636 (N_1636,In_125,In_103);
and U1637 (N_1637,In_952,In_682);
nor U1638 (N_1638,In_840,In_725);
xor U1639 (N_1639,In_999,In_67);
and U1640 (N_1640,In_492,In_1434);
nor U1641 (N_1641,In_152,In_166);
and U1642 (N_1642,In_103,In_338);
or U1643 (N_1643,In_1429,In_782);
xor U1644 (N_1644,In_134,In_1395);
xnor U1645 (N_1645,In_148,In_784);
or U1646 (N_1646,In_1387,In_189);
and U1647 (N_1647,In_59,In_452);
nor U1648 (N_1648,In_491,In_1012);
nand U1649 (N_1649,In_370,In_705);
nor U1650 (N_1650,In_369,In_698);
and U1651 (N_1651,In_574,In_102);
xor U1652 (N_1652,In_363,In_1438);
and U1653 (N_1653,In_943,In_1371);
and U1654 (N_1654,In_570,In_779);
and U1655 (N_1655,In_807,In_1202);
or U1656 (N_1656,In_776,In_887);
or U1657 (N_1657,In_363,In_1047);
nand U1658 (N_1658,In_1221,In_127);
xnor U1659 (N_1659,In_31,In_1043);
nor U1660 (N_1660,In_132,In_272);
or U1661 (N_1661,In_1401,In_53);
xor U1662 (N_1662,In_527,In_403);
and U1663 (N_1663,In_514,In_550);
and U1664 (N_1664,In_896,In_1257);
or U1665 (N_1665,In_468,In_195);
or U1666 (N_1666,In_108,In_563);
nand U1667 (N_1667,In_482,In_560);
nand U1668 (N_1668,In_82,In_502);
or U1669 (N_1669,In_731,In_416);
and U1670 (N_1670,In_1479,In_750);
nand U1671 (N_1671,In_1252,In_418);
xnor U1672 (N_1672,In_852,In_796);
nand U1673 (N_1673,In_505,In_245);
nand U1674 (N_1674,In_465,In_268);
nand U1675 (N_1675,In_925,In_1030);
and U1676 (N_1676,In_549,In_1448);
nand U1677 (N_1677,In_858,In_1106);
and U1678 (N_1678,In_315,In_635);
and U1679 (N_1679,In_1004,In_1322);
and U1680 (N_1680,In_496,In_656);
nor U1681 (N_1681,In_1105,In_544);
nor U1682 (N_1682,In_1421,In_166);
xnor U1683 (N_1683,In_591,In_808);
nand U1684 (N_1684,In_736,In_743);
xor U1685 (N_1685,In_412,In_87);
nand U1686 (N_1686,In_522,In_597);
nand U1687 (N_1687,In_448,In_235);
nor U1688 (N_1688,In_556,In_814);
or U1689 (N_1689,In_1347,In_174);
nand U1690 (N_1690,In_616,In_158);
and U1691 (N_1691,In_879,In_1114);
and U1692 (N_1692,In_295,In_8);
nand U1693 (N_1693,In_484,In_397);
and U1694 (N_1694,In_748,In_1380);
nor U1695 (N_1695,In_988,In_1386);
nor U1696 (N_1696,In_912,In_1007);
or U1697 (N_1697,In_695,In_70);
nand U1698 (N_1698,In_1233,In_231);
nor U1699 (N_1699,In_584,In_1388);
or U1700 (N_1700,In_426,In_1112);
xnor U1701 (N_1701,In_56,In_92);
nor U1702 (N_1702,In_1364,In_667);
nand U1703 (N_1703,In_144,In_1199);
and U1704 (N_1704,In_246,In_641);
or U1705 (N_1705,In_387,In_1065);
and U1706 (N_1706,In_314,In_809);
nor U1707 (N_1707,In_990,In_815);
nand U1708 (N_1708,In_216,In_716);
nor U1709 (N_1709,In_34,In_20);
and U1710 (N_1710,In_189,In_1418);
nor U1711 (N_1711,In_1242,In_654);
and U1712 (N_1712,In_843,In_929);
nand U1713 (N_1713,In_1239,In_1231);
or U1714 (N_1714,In_400,In_817);
and U1715 (N_1715,In_215,In_1274);
and U1716 (N_1716,In_557,In_656);
and U1717 (N_1717,In_1323,In_1252);
xnor U1718 (N_1718,In_1235,In_1075);
or U1719 (N_1719,In_376,In_1446);
or U1720 (N_1720,In_448,In_1197);
or U1721 (N_1721,In_1153,In_189);
nand U1722 (N_1722,In_1279,In_447);
xor U1723 (N_1723,In_87,In_1247);
or U1724 (N_1724,In_736,In_299);
and U1725 (N_1725,In_674,In_1293);
xnor U1726 (N_1726,In_449,In_864);
or U1727 (N_1727,In_719,In_39);
or U1728 (N_1728,In_1185,In_321);
nor U1729 (N_1729,In_579,In_989);
nand U1730 (N_1730,In_301,In_1360);
and U1731 (N_1731,In_1357,In_695);
nand U1732 (N_1732,In_784,In_465);
nand U1733 (N_1733,In_645,In_1375);
nor U1734 (N_1734,In_416,In_272);
and U1735 (N_1735,In_837,In_997);
nand U1736 (N_1736,In_860,In_392);
nor U1737 (N_1737,In_1199,In_546);
and U1738 (N_1738,In_907,In_658);
nor U1739 (N_1739,In_881,In_279);
and U1740 (N_1740,In_92,In_785);
or U1741 (N_1741,In_807,In_233);
or U1742 (N_1742,In_489,In_1156);
nand U1743 (N_1743,In_394,In_1142);
and U1744 (N_1744,In_92,In_1109);
or U1745 (N_1745,In_1005,In_1200);
xnor U1746 (N_1746,In_265,In_1122);
nor U1747 (N_1747,In_1052,In_519);
nand U1748 (N_1748,In_574,In_1007);
nand U1749 (N_1749,In_362,In_111);
xnor U1750 (N_1750,In_182,In_779);
nand U1751 (N_1751,In_235,In_992);
nand U1752 (N_1752,In_1261,In_929);
and U1753 (N_1753,In_520,In_353);
nand U1754 (N_1754,In_798,In_298);
and U1755 (N_1755,In_1399,In_1312);
or U1756 (N_1756,In_68,In_3);
nor U1757 (N_1757,In_28,In_1353);
or U1758 (N_1758,In_1016,In_1290);
or U1759 (N_1759,In_109,In_1180);
and U1760 (N_1760,In_15,In_1107);
and U1761 (N_1761,In_247,In_824);
and U1762 (N_1762,In_277,In_1426);
nand U1763 (N_1763,In_1367,In_431);
or U1764 (N_1764,In_1054,In_181);
nor U1765 (N_1765,In_1382,In_819);
nand U1766 (N_1766,In_763,In_808);
xnor U1767 (N_1767,In_632,In_836);
nor U1768 (N_1768,In_1314,In_997);
nor U1769 (N_1769,In_18,In_1102);
or U1770 (N_1770,In_733,In_364);
nand U1771 (N_1771,In_569,In_1138);
nor U1772 (N_1772,In_407,In_570);
nor U1773 (N_1773,In_1071,In_457);
nand U1774 (N_1774,In_456,In_1304);
or U1775 (N_1775,In_85,In_353);
nor U1776 (N_1776,In_139,In_1377);
nand U1777 (N_1777,In_1146,In_393);
or U1778 (N_1778,In_403,In_1304);
and U1779 (N_1779,In_1,In_1277);
and U1780 (N_1780,In_1110,In_939);
and U1781 (N_1781,In_421,In_1207);
or U1782 (N_1782,In_798,In_1048);
nand U1783 (N_1783,In_1399,In_424);
nand U1784 (N_1784,In_297,In_1376);
nor U1785 (N_1785,In_264,In_1042);
nand U1786 (N_1786,In_680,In_422);
nor U1787 (N_1787,In_1230,In_489);
or U1788 (N_1788,In_299,In_1389);
xor U1789 (N_1789,In_1226,In_1215);
nand U1790 (N_1790,In_918,In_740);
or U1791 (N_1791,In_849,In_911);
or U1792 (N_1792,In_797,In_1265);
and U1793 (N_1793,In_731,In_1166);
and U1794 (N_1794,In_713,In_305);
nor U1795 (N_1795,In_1280,In_341);
nor U1796 (N_1796,In_120,In_103);
nand U1797 (N_1797,In_1445,In_1366);
or U1798 (N_1798,In_926,In_255);
nor U1799 (N_1799,In_1325,In_233);
and U1800 (N_1800,In_282,In_538);
nor U1801 (N_1801,In_326,In_542);
nand U1802 (N_1802,In_1433,In_852);
or U1803 (N_1803,In_1083,In_36);
and U1804 (N_1804,In_1082,In_671);
and U1805 (N_1805,In_1334,In_408);
nand U1806 (N_1806,In_107,In_264);
nor U1807 (N_1807,In_220,In_450);
nand U1808 (N_1808,In_912,In_243);
and U1809 (N_1809,In_472,In_576);
and U1810 (N_1810,In_168,In_1341);
or U1811 (N_1811,In_364,In_985);
nand U1812 (N_1812,In_266,In_635);
nand U1813 (N_1813,In_981,In_380);
and U1814 (N_1814,In_998,In_940);
or U1815 (N_1815,In_617,In_686);
nand U1816 (N_1816,In_1148,In_1230);
xor U1817 (N_1817,In_229,In_845);
or U1818 (N_1818,In_468,In_1101);
xnor U1819 (N_1819,In_1059,In_565);
nor U1820 (N_1820,In_1271,In_700);
and U1821 (N_1821,In_293,In_371);
nand U1822 (N_1822,In_1432,In_358);
nor U1823 (N_1823,In_319,In_967);
nor U1824 (N_1824,In_796,In_574);
nor U1825 (N_1825,In_736,In_493);
or U1826 (N_1826,In_24,In_407);
or U1827 (N_1827,In_1177,In_968);
nor U1828 (N_1828,In_1199,In_1086);
nand U1829 (N_1829,In_26,In_1161);
nor U1830 (N_1830,In_967,In_741);
and U1831 (N_1831,In_261,In_904);
nand U1832 (N_1832,In_1158,In_497);
or U1833 (N_1833,In_326,In_399);
and U1834 (N_1834,In_320,In_573);
nand U1835 (N_1835,In_742,In_1469);
and U1836 (N_1836,In_486,In_198);
and U1837 (N_1837,In_214,In_818);
and U1838 (N_1838,In_53,In_48);
or U1839 (N_1839,In_1470,In_1145);
and U1840 (N_1840,In_1460,In_1158);
and U1841 (N_1841,In_765,In_1117);
nand U1842 (N_1842,In_763,In_241);
or U1843 (N_1843,In_287,In_1327);
xnor U1844 (N_1844,In_1039,In_1472);
or U1845 (N_1845,In_790,In_1155);
or U1846 (N_1846,In_809,In_84);
xor U1847 (N_1847,In_1028,In_909);
nor U1848 (N_1848,In_381,In_1079);
nand U1849 (N_1849,In_415,In_596);
and U1850 (N_1850,In_539,In_80);
nand U1851 (N_1851,In_1130,In_1450);
and U1852 (N_1852,In_918,In_816);
nand U1853 (N_1853,In_110,In_126);
nand U1854 (N_1854,In_43,In_682);
nor U1855 (N_1855,In_590,In_767);
nand U1856 (N_1856,In_1116,In_1250);
and U1857 (N_1857,In_938,In_238);
or U1858 (N_1858,In_157,In_1039);
and U1859 (N_1859,In_646,In_778);
or U1860 (N_1860,In_992,In_1036);
xnor U1861 (N_1861,In_1200,In_546);
or U1862 (N_1862,In_949,In_88);
or U1863 (N_1863,In_56,In_914);
nor U1864 (N_1864,In_858,In_924);
nor U1865 (N_1865,In_462,In_355);
nor U1866 (N_1866,In_863,In_743);
xnor U1867 (N_1867,In_615,In_271);
or U1868 (N_1868,In_1447,In_664);
nand U1869 (N_1869,In_280,In_462);
or U1870 (N_1870,In_201,In_1075);
and U1871 (N_1871,In_111,In_205);
and U1872 (N_1872,In_769,In_956);
nand U1873 (N_1873,In_136,In_531);
or U1874 (N_1874,In_479,In_612);
xnor U1875 (N_1875,In_932,In_1490);
and U1876 (N_1876,In_301,In_748);
or U1877 (N_1877,In_963,In_1366);
and U1878 (N_1878,In_361,In_911);
and U1879 (N_1879,In_151,In_1159);
nor U1880 (N_1880,In_843,In_263);
nand U1881 (N_1881,In_1171,In_1486);
or U1882 (N_1882,In_1422,In_860);
nand U1883 (N_1883,In_1384,In_499);
xor U1884 (N_1884,In_859,In_934);
nor U1885 (N_1885,In_437,In_1290);
or U1886 (N_1886,In_1365,In_481);
or U1887 (N_1887,In_1099,In_1068);
nor U1888 (N_1888,In_723,In_843);
nor U1889 (N_1889,In_763,In_1493);
and U1890 (N_1890,In_752,In_1367);
and U1891 (N_1891,In_1385,In_833);
and U1892 (N_1892,In_217,In_608);
and U1893 (N_1893,In_16,In_985);
and U1894 (N_1894,In_1297,In_572);
or U1895 (N_1895,In_1399,In_752);
nor U1896 (N_1896,In_783,In_139);
xnor U1897 (N_1897,In_954,In_1230);
xnor U1898 (N_1898,In_1190,In_1431);
xor U1899 (N_1899,In_673,In_981);
xor U1900 (N_1900,In_1306,In_1138);
and U1901 (N_1901,In_536,In_1215);
or U1902 (N_1902,In_1354,In_907);
xnor U1903 (N_1903,In_173,In_641);
nor U1904 (N_1904,In_1073,In_337);
nor U1905 (N_1905,In_1399,In_644);
nand U1906 (N_1906,In_343,In_1111);
nand U1907 (N_1907,In_635,In_1381);
nand U1908 (N_1908,In_249,In_211);
xnor U1909 (N_1909,In_544,In_327);
and U1910 (N_1910,In_794,In_960);
nand U1911 (N_1911,In_250,In_114);
or U1912 (N_1912,In_348,In_291);
nand U1913 (N_1913,In_409,In_1064);
and U1914 (N_1914,In_1001,In_387);
nor U1915 (N_1915,In_250,In_1372);
nor U1916 (N_1916,In_1192,In_631);
nor U1917 (N_1917,In_778,In_1028);
nand U1918 (N_1918,In_130,In_1219);
and U1919 (N_1919,In_86,In_1239);
or U1920 (N_1920,In_4,In_767);
or U1921 (N_1921,In_1387,In_986);
or U1922 (N_1922,In_240,In_1365);
and U1923 (N_1923,In_869,In_1494);
or U1924 (N_1924,In_1056,In_922);
xor U1925 (N_1925,In_203,In_1244);
nand U1926 (N_1926,In_986,In_1351);
nor U1927 (N_1927,In_1417,In_1156);
nor U1928 (N_1928,In_1442,In_1001);
or U1929 (N_1929,In_116,In_766);
nand U1930 (N_1930,In_777,In_787);
nand U1931 (N_1931,In_52,In_497);
and U1932 (N_1932,In_5,In_47);
nor U1933 (N_1933,In_316,In_1249);
or U1934 (N_1934,In_1367,In_1448);
or U1935 (N_1935,In_582,In_240);
or U1936 (N_1936,In_1485,In_271);
nand U1937 (N_1937,In_205,In_360);
nand U1938 (N_1938,In_1274,In_1033);
and U1939 (N_1939,In_415,In_1242);
nand U1940 (N_1940,In_772,In_932);
or U1941 (N_1941,In_541,In_1189);
or U1942 (N_1942,In_694,In_774);
and U1943 (N_1943,In_630,In_380);
nor U1944 (N_1944,In_1468,In_340);
and U1945 (N_1945,In_312,In_1487);
nand U1946 (N_1946,In_115,In_800);
nand U1947 (N_1947,In_970,In_816);
and U1948 (N_1948,In_762,In_780);
or U1949 (N_1949,In_337,In_109);
or U1950 (N_1950,In_1361,In_546);
nor U1951 (N_1951,In_1400,In_1126);
and U1952 (N_1952,In_776,In_190);
nand U1953 (N_1953,In_963,In_817);
or U1954 (N_1954,In_293,In_1026);
nor U1955 (N_1955,In_1401,In_290);
or U1956 (N_1956,In_486,In_19);
nand U1957 (N_1957,In_790,In_460);
nand U1958 (N_1958,In_291,In_1012);
nand U1959 (N_1959,In_455,In_349);
nor U1960 (N_1960,In_359,In_81);
or U1961 (N_1961,In_952,In_440);
nand U1962 (N_1962,In_317,In_758);
xor U1963 (N_1963,In_210,In_1305);
or U1964 (N_1964,In_298,In_1454);
and U1965 (N_1965,In_230,In_1236);
and U1966 (N_1966,In_1148,In_1371);
nand U1967 (N_1967,In_118,In_1049);
nand U1968 (N_1968,In_1268,In_960);
nor U1969 (N_1969,In_663,In_955);
and U1970 (N_1970,In_699,In_1223);
and U1971 (N_1971,In_621,In_327);
nand U1972 (N_1972,In_1282,In_1298);
nand U1973 (N_1973,In_34,In_587);
or U1974 (N_1974,In_539,In_732);
and U1975 (N_1975,In_257,In_244);
nand U1976 (N_1976,In_977,In_1458);
nand U1977 (N_1977,In_1000,In_795);
nand U1978 (N_1978,In_1421,In_32);
nand U1979 (N_1979,In_273,In_376);
nand U1980 (N_1980,In_910,In_1137);
and U1981 (N_1981,In_1167,In_54);
nor U1982 (N_1982,In_868,In_237);
and U1983 (N_1983,In_1498,In_473);
nor U1984 (N_1984,In_761,In_426);
or U1985 (N_1985,In_439,In_837);
nor U1986 (N_1986,In_11,In_465);
nand U1987 (N_1987,In_92,In_164);
or U1988 (N_1988,In_330,In_1111);
nor U1989 (N_1989,In_1443,In_948);
nand U1990 (N_1990,In_833,In_1136);
nor U1991 (N_1991,In_1455,In_542);
and U1992 (N_1992,In_313,In_304);
and U1993 (N_1993,In_1098,In_866);
nand U1994 (N_1994,In_513,In_895);
nor U1995 (N_1995,In_1363,In_1240);
and U1996 (N_1996,In_1384,In_1466);
nand U1997 (N_1997,In_1241,In_173);
nand U1998 (N_1998,In_398,In_202);
or U1999 (N_1999,In_408,In_1147);
and U2000 (N_2000,In_1293,In_155);
nor U2001 (N_2001,In_705,In_615);
or U2002 (N_2002,In_738,In_91);
or U2003 (N_2003,In_389,In_1451);
nor U2004 (N_2004,In_1047,In_23);
and U2005 (N_2005,In_301,In_968);
nand U2006 (N_2006,In_951,In_1323);
or U2007 (N_2007,In_354,In_901);
nand U2008 (N_2008,In_597,In_391);
xnor U2009 (N_2009,In_1285,In_1410);
nand U2010 (N_2010,In_413,In_58);
nor U2011 (N_2011,In_1274,In_221);
nand U2012 (N_2012,In_1245,In_433);
nor U2013 (N_2013,In_135,In_967);
xnor U2014 (N_2014,In_1100,In_899);
and U2015 (N_2015,In_636,In_1113);
or U2016 (N_2016,In_700,In_929);
nand U2017 (N_2017,In_92,In_433);
and U2018 (N_2018,In_259,In_266);
or U2019 (N_2019,In_1415,In_415);
nor U2020 (N_2020,In_797,In_801);
or U2021 (N_2021,In_740,In_776);
nand U2022 (N_2022,In_798,In_996);
nand U2023 (N_2023,In_395,In_432);
xnor U2024 (N_2024,In_1481,In_1230);
or U2025 (N_2025,In_1329,In_1370);
or U2026 (N_2026,In_162,In_1036);
nor U2027 (N_2027,In_91,In_377);
or U2028 (N_2028,In_1191,In_1243);
nor U2029 (N_2029,In_843,In_1335);
or U2030 (N_2030,In_1468,In_755);
nand U2031 (N_2031,In_104,In_968);
and U2032 (N_2032,In_1065,In_852);
and U2033 (N_2033,In_530,In_1481);
or U2034 (N_2034,In_977,In_541);
nand U2035 (N_2035,In_1317,In_434);
xor U2036 (N_2036,In_30,In_108);
or U2037 (N_2037,In_798,In_1366);
or U2038 (N_2038,In_369,In_1182);
xor U2039 (N_2039,In_563,In_1113);
nor U2040 (N_2040,In_741,In_438);
nand U2041 (N_2041,In_1313,In_659);
or U2042 (N_2042,In_162,In_147);
xnor U2043 (N_2043,In_869,In_1398);
and U2044 (N_2044,In_1396,In_960);
nor U2045 (N_2045,In_678,In_1401);
nand U2046 (N_2046,In_654,In_176);
nor U2047 (N_2047,In_1223,In_510);
nor U2048 (N_2048,In_1013,In_1281);
and U2049 (N_2049,In_884,In_511);
nand U2050 (N_2050,In_283,In_725);
nand U2051 (N_2051,In_238,In_985);
and U2052 (N_2052,In_393,In_1454);
and U2053 (N_2053,In_842,In_1465);
nand U2054 (N_2054,In_1300,In_30);
nor U2055 (N_2055,In_720,In_696);
nor U2056 (N_2056,In_870,In_1366);
xnor U2057 (N_2057,In_238,In_82);
xnor U2058 (N_2058,In_762,In_1040);
nand U2059 (N_2059,In_402,In_1444);
nor U2060 (N_2060,In_981,In_758);
and U2061 (N_2061,In_1069,In_454);
nand U2062 (N_2062,In_1443,In_121);
nor U2063 (N_2063,In_1164,In_686);
and U2064 (N_2064,In_110,In_475);
nand U2065 (N_2065,In_1213,In_1067);
and U2066 (N_2066,In_901,In_318);
and U2067 (N_2067,In_784,In_356);
and U2068 (N_2068,In_1457,In_605);
and U2069 (N_2069,In_729,In_1196);
or U2070 (N_2070,In_486,In_1216);
xnor U2071 (N_2071,In_775,In_1104);
nor U2072 (N_2072,In_474,In_521);
nand U2073 (N_2073,In_450,In_954);
nor U2074 (N_2074,In_291,In_224);
or U2075 (N_2075,In_706,In_658);
xnor U2076 (N_2076,In_226,In_424);
or U2077 (N_2077,In_640,In_1438);
nor U2078 (N_2078,In_973,In_1182);
nand U2079 (N_2079,In_587,In_1367);
and U2080 (N_2080,In_880,In_645);
nand U2081 (N_2081,In_1029,In_1073);
xor U2082 (N_2082,In_726,In_825);
nor U2083 (N_2083,In_1484,In_995);
nor U2084 (N_2084,In_400,In_1261);
and U2085 (N_2085,In_923,In_612);
nand U2086 (N_2086,In_150,In_568);
nand U2087 (N_2087,In_210,In_1143);
or U2088 (N_2088,In_150,In_256);
nor U2089 (N_2089,In_883,In_1445);
xor U2090 (N_2090,In_980,In_766);
and U2091 (N_2091,In_1106,In_899);
nand U2092 (N_2092,In_1048,In_1303);
nand U2093 (N_2093,In_239,In_578);
nor U2094 (N_2094,In_1085,In_1378);
or U2095 (N_2095,In_1300,In_75);
and U2096 (N_2096,In_462,In_935);
xor U2097 (N_2097,In_1115,In_1406);
and U2098 (N_2098,In_1439,In_591);
xor U2099 (N_2099,In_404,In_1107);
nor U2100 (N_2100,In_87,In_1413);
nor U2101 (N_2101,In_374,In_321);
nor U2102 (N_2102,In_304,In_1342);
nor U2103 (N_2103,In_985,In_1306);
nand U2104 (N_2104,In_1345,In_1047);
nand U2105 (N_2105,In_1354,In_473);
nor U2106 (N_2106,In_85,In_164);
or U2107 (N_2107,In_1436,In_1414);
or U2108 (N_2108,In_790,In_1170);
or U2109 (N_2109,In_1386,In_526);
or U2110 (N_2110,In_530,In_818);
and U2111 (N_2111,In_1017,In_612);
and U2112 (N_2112,In_457,In_420);
or U2113 (N_2113,In_1077,In_1046);
nand U2114 (N_2114,In_366,In_90);
nand U2115 (N_2115,In_390,In_1331);
nand U2116 (N_2116,In_1000,In_1161);
and U2117 (N_2117,In_1418,In_1043);
xor U2118 (N_2118,In_1363,In_880);
nor U2119 (N_2119,In_848,In_1046);
nand U2120 (N_2120,In_1420,In_1233);
nor U2121 (N_2121,In_929,In_1359);
nor U2122 (N_2122,In_662,In_50);
nand U2123 (N_2123,In_869,In_338);
and U2124 (N_2124,In_151,In_1495);
or U2125 (N_2125,In_115,In_928);
nand U2126 (N_2126,In_487,In_1259);
and U2127 (N_2127,In_1375,In_906);
or U2128 (N_2128,In_658,In_1397);
nor U2129 (N_2129,In_86,In_1104);
or U2130 (N_2130,In_1497,In_66);
nor U2131 (N_2131,In_591,In_482);
nor U2132 (N_2132,In_1079,In_339);
nor U2133 (N_2133,In_432,In_107);
nand U2134 (N_2134,In_472,In_1148);
xnor U2135 (N_2135,In_610,In_1372);
nor U2136 (N_2136,In_1455,In_1099);
and U2137 (N_2137,In_949,In_1053);
nand U2138 (N_2138,In_901,In_1365);
nand U2139 (N_2139,In_670,In_488);
nor U2140 (N_2140,In_1271,In_223);
or U2141 (N_2141,In_246,In_1170);
xor U2142 (N_2142,In_1188,In_589);
and U2143 (N_2143,In_502,In_793);
and U2144 (N_2144,In_1107,In_522);
nor U2145 (N_2145,In_1354,In_575);
nand U2146 (N_2146,In_713,In_1302);
nor U2147 (N_2147,In_1211,In_1029);
and U2148 (N_2148,In_533,In_499);
nand U2149 (N_2149,In_727,In_1428);
nor U2150 (N_2150,In_1368,In_1061);
and U2151 (N_2151,In_15,In_1172);
and U2152 (N_2152,In_1448,In_1249);
or U2153 (N_2153,In_114,In_977);
and U2154 (N_2154,In_588,In_1034);
and U2155 (N_2155,In_1154,In_643);
nand U2156 (N_2156,In_1313,In_362);
nor U2157 (N_2157,In_222,In_90);
nor U2158 (N_2158,In_1012,In_1366);
or U2159 (N_2159,In_626,In_1059);
nand U2160 (N_2160,In_903,In_997);
xnor U2161 (N_2161,In_473,In_1326);
xor U2162 (N_2162,In_957,In_567);
or U2163 (N_2163,In_866,In_228);
or U2164 (N_2164,In_892,In_729);
and U2165 (N_2165,In_1013,In_76);
and U2166 (N_2166,In_1497,In_1346);
nand U2167 (N_2167,In_185,In_978);
and U2168 (N_2168,In_1429,In_492);
nand U2169 (N_2169,In_595,In_108);
and U2170 (N_2170,In_787,In_432);
nand U2171 (N_2171,In_722,In_900);
nor U2172 (N_2172,In_292,In_1473);
and U2173 (N_2173,In_678,In_851);
nand U2174 (N_2174,In_1467,In_38);
or U2175 (N_2175,In_48,In_671);
or U2176 (N_2176,In_9,In_1126);
and U2177 (N_2177,In_1087,In_1463);
nand U2178 (N_2178,In_1008,In_193);
nand U2179 (N_2179,In_1403,In_382);
nor U2180 (N_2180,In_1423,In_794);
nand U2181 (N_2181,In_1479,In_752);
nor U2182 (N_2182,In_766,In_784);
or U2183 (N_2183,In_842,In_320);
nand U2184 (N_2184,In_1114,In_89);
nand U2185 (N_2185,In_767,In_587);
and U2186 (N_2186,In_884,In_858);
and U2187 (N_2187,In_516,In_1);
nand U2188 (N_2188,In_541,In_500);
and U2189 (N_2189,In_859,In_1486);
and U2190 (N_2190,In_1168,In_963);
nor U2191 (N_2191,In_402,In_788);
and U2192 (N_2192,In_209,In_474);
and U2193 (N_2193,In_365,In_1411);
nor U2194 (N_2194,In_148,In_891);
nor U2195 (N_2195,In_405,In_422);
or U2196 (N_2196,In_492,In_1332);
xor U2197 (N_2197,In_600,In_583);
and U2198 (N_2198,In_437,In_1414);
nand U2199 (N_2199,In_76,In_1001);
nand U2200 (N_2200,In_407,In_56);
nor U2201 (N_2201,In_1485,In_985);
and U2202 (N_2202,In_1188,In_1125);
and U2203 (N_2203,In_688,In_1397);
and U2204 (N_2204,In_584,In_465);
or U2205 (N_2205,In_89,In_1323);
or U2206 (N_2206,In_1312,In_191);
and U2207 (N_2207,In_910,In_1436);
or U2208 (N_2208,In_1187,In_1152);
nor U2209 (N_2209,In_347,In_46);
or U2210 (N_2210,In_1010,In_758);
xnor U2211 (N_2211,In_1417,In_243);
nor U2212 (N_2212,In_540,In_579);
nor U2213 (N_2213,In_1440,In_212);
nand U2214 (N_2214,In_630,In_334);
and U2215 (N_2215,In_1014,In_242);
or U2216 (N_2216,In_844,In_88);
or U2217 (N_2217,In_73,In_376);
nand U2218 (N_2218,In_959,In_698);
or U2219 (N_2219,In_1031,In_527);
nand U2220 (N_2220,In_1367,In_781);
nand U2221 (N_2221,In_971,In_1096);
and U2222 (N_2222,In_572,In_258);
xnor U2223 (N_2223,In_197,In_802);
nor U2224 (N_2224,In_1203,In_1300);
xnor U2225 (N_2225,In_278,In_415);
or U2226 (N_2226,In_325,In_1391);
or U2227 (N_2227,In_857,In_632);
and U2228 (N_2228,In_1362,In_1238);
or U2229 (N_2229,In_1065,In_526);
nor U2230 (N_2230,In_1497,In_444);
or U2231 (N_2231,In_1094,In_950);
nor U2232 (N_2232,In_1327,In_572);
or U2233 (N_2233,In_600,In_1178);
nand U2234 (N_2234,In_212,In_698);
nor U2235 (N_2235,In_247,In_1139);
nor U2236 (N_2236,In_406,In_357);
nand U2237 (N_2237,In_882,In_1024);
or U2238 (N_2238,In_1230,In_835);
or U2239 (N_2239,In_218,In_353);
nand U2240 (N_2240,In_1072,In_964);
nor U2241 (N_2241,In_1158,In_755);
or U2242 (N_2242,In_1481,In_1413);
or U2243 (N_2243,In_809,In_16);
nand U2244 (N_2244,In_1440,In_809);
nand U2245 (N_2245,In_573,In_677);
nor U2246 (N_2246,In_666,In_45);
and U2247 (N_2247,In_233,In_830);
xnor U2248 (N_2248,In_603,In_1372);
or U2249 (N_2249,In_940,In_923);
nand U2250 (N_2250,In_781,In_694);
and U2251 (N_2251,In_555,In_1377);
and U2252 (N_2252,In_310,In_646);
or U2253 (N_2253,In_335,In_947);
nor U2254 (N_2254,In_184,In_1373);
xor U2255 (N_2255,In_1226,In_42);
nor U2256 (N_2256,In_1231,In_917);
nor U2257 (N_2257,In_1379,In_230);
nand U2258 (N_2258,In_915,In_125);
nor U2259 (N_2259,In_1230,In_539);
nor U2260 (N_2260,In_460,In_287);
nor U2261 (N_2261,In_1206,In_662);
nand U2262 (N_2262,In_139,In_365);
nor U2263 (N_2263,In_1456,In_633);
nand U2264 (N_2264,In_555,In_528);
nor U2265 (N_2265,In_577,In_235);
or U2266 (N_2266,In_1123,In_901);
or U2267 (N_2267,In_418,In_202);
nand U2268 (N_2268,In_1302,In_114);
nand U2269 (N_2269,In_1328,In_935);
nand U2270 (N_2270,In_568,In_945);
and U2271 (N_2271,In_262,In_352);
xor U2272 (N_2272,In_219,In_827);
xnor U2273 (N_2273,In_295,In_950);
xnor U2274 (N_2274,In_1355,In_149);
and U2275 (N_2275,In_1412,In_960);
and U2276 (N_2276,In_855,In_811);
or U2277 (N_2277,In_918,In_65);
and U2278 (N_2278,In_1025,In_407);
and U2279 (N_2279,In_805,In_298);
or U2280 (N_2280,In_209,In_201);
xor U2281 (N_2281,In_903,In_905);
or U2282 (N_2282,In_848,In_370);
nor U2283 (N_2283,In_413,In_1259);
nand U2284 (N_2284,In_12,In_188);
or U2285 (N_2285,In_1470,In_127);
nand U2286 (N_2286,In_263,In_1302);
nand U2287 (N_2287,In_469,In_453);
and U2288 (N_2288,In_1017,In_199);
and U2289 (N_2289,In_825,In_832);
nand U2290 (N_2290,In_1013,In_814);
nand U2291 (N_2291,In_820,In_202);
or U2292 (N_2292,In_1066,In_738);
nor U2293 (N_2293,In_806,In_1165);
nor U2294 (N_2294,In_197,In_1066);
or U2295 (N_2295,In_230,In_1433);
nand U2296 (N_2296,In_633,In_514);
or U2297 (N_2297,In_196,In_1456);
or U2298 (N_2298,In_608,In_1047);
and U2299 (N_2299,In_981,In_1162);
or U2300 (N_2300,In_1091,In_826);
nor U2301 (N_2301,In_580,In_211);
nand U2302 (N_2302,In_902,In_835);
nor U2303 (N_2303,In_1365,In_540);
xnor U2304 (N_2304,In_994,In_421);
or U2305 (N_2305,In_231,In_330);
nand U2306 (N_2306,In_588,In_1375);
xnor U2307 (N_2307,In_695,In_355);
nor U2308 (N_2308,In_1378,In_372);
nand U2309 (N_2309,In_335,In_304);
nor U2310 (N_2310,In_1152,In_762);
and U2311 (N_2311,In_654,In_1366);
or U2312 (N_2312,In_1368,In_1451);
xnor U2313 (N_2313,In_1494,In_331);
nor U2314 (N_2314,In_659,In_1320);
nand U2315 (N_2315,In_1115,In_1317);
or U2316 (N_2316,In_1448,In_1286);
and U2317 (N_2317,In_434,In_982);
and U2318 (N_2318,In_1113,In_1406);
nand U2319 (N_2319,In_245,In_60);
nor U2320 (N_2320,In_803,In_1296);
nand U2321 (N_2321,In_1043,In_670);
and U2322 (N_2322,In_724,In_258);
nor U2323 (N_2323,In_1385,In_107);
and U2324 (N_2324,In_870,In_621);
nor U2325 (N_2325,In_444,In_773);
or U2326 (N_2326,In_959,In_404);
nand U2327 (N_2327,In_1175,In_51);
xnor U2328 (N_2328,In_1117,In_1217);
nor U2329 (N_2329,In_1175,In_546);
and U2330 (N_2330,In_643,In_439);
or U2331 (N_2331,In_53,In_1466);
and U2332 (N_2332,In_1017,In_1236);
xnor U2333 (N_2333,In_1038,In_637);
nor U2334 (N_2334,In_608,In_833);
xnor U2335 (N_2335,In_55,In_165);
nand U2336 (N_2336,In_21,In_1470);
or U2337 (N_2337,In_1017,In_856);
nor U2338 (N_2338,In_449,In_731);
nor U2339 (N_2339,In_1001,In_601);
nand U2340 (N_2340,In_821,In_1149);
xor U2341 (N_2341,In_1128,In_221);
nand U2342 (N_2342,In_497,In_786);
or U2343 (N_2343,In_856,In_1201);
nand U2344 (N_2344,In_1021,In_1303);
xnor U2345 (N_2345,In_401,In_482);
nand U2346 (N_2346,In_594,In_470);
or U2347 (N_2347,In_191,In_1440);
xor U2348 (N_2348,In_1043,In_517);
nor U2349 (N_2349,In_1030,In_989);
nor U2350 (N_2350,In_831,In_524);
and U2351 (N_2351,In_1357,In_1424);
xor U2352 (N_2352,In_1206,In_1307);
nand U2353 (N_2353,In_170,In_322);
or U2354 (N_2354,In_821,In_444);
nor U2355 (N_2355,In_656,In_1008);
and U2356 (N_2356,In_759,In_0);
and U2357 (N_2357,In_1399,In_328);
or U2358 (N_2358,In_275,In_675);
nor U2359 (N_2359,In_1238,In_862);
and U2360 (N_2360,In_1001,In_147);
and U2361 (N_2361,In_89,In_969);
nor U2362 (N_2362,In_1312,In_1341);
and U2363 (N_2363,In_634,In_573);
or U2364 (N_2364,In_851,In_105);
or U2365 (N_2365,In_765,In_998);
nand U2366 (N_2366,In_1484,In_160);
and U2367 (N_2367,In_1341,In_276);
and U2368 (N_2368,In_1344,In_1282);
and U2369 (N_2369,In_1099,In_124);
xor U2370 (N_2370,In_611,In_1110);
or U2371 (N_2371,In_945,In_1026);
or U2372 (N_2372,In_1053,In_907);
and U2373 (N_2373,In_1466,In_316);
and U2374 (N_2374,In_1064,In_1055);
and U2375 (N_2375,In_1149,In_302);
nor U2376 (N_2376,In_54,In_652);
xor U2377 (N_2377,In_1326,In_755);
nor U2378 (N_2378,In_84,In_1274);
nand U2379 (N_2379,In_899,In_1369);
nand U2380 (N_2380,In_862,In_1054);
nand U2381 (N_2381,In_55,In_30);
nor U2382 (N_2382,In_1150,In_453);
nor U2383 (N_2383,In_375,In_692);
nor U2384 (N_2384,In_177,In_1236);
and U2385 (N_2385,In_39,In_246);
nor U2386 (N_2386,In_1171,In_227);
and U2387 (N_2387,In_461,In_443);
and U2388 (N_2388,In_841,In_1407);
nor U2389 (N_2389,In_888,In_434);
nand U2390 (N_2390,In_788,In_1338);
nand U2391 (N_2391,In_1372,In_1392);
or U2392 (N_2392,In_30,In_604);
nand U2393 (N_2393,In_988,In_1012);
and U2394 (N_2394,In_1376,In_1385);
nor U2395 (N_2395,In_754,In_332);
nand U2396 (N_2396,In_950,In_291);
xnor U2397 (N_2397,In_560,In_934);
or U2398 (N_2398,In_276,In_1131);
nor U2399 (N_2399,In_680,In_707);
and U2400 (N_2400,In_1159,In_700);
xnor U2401 (N_2401,In_979,In_230);
nor U2402 (N_2402,In_1400,In_914);
xor U2403 (N_2403,In_1138,In_464);
or U2404 (N_2404,In_1070,In_1307);
or U2405 (N_2405,In_571,In_1395);
nor U2406 (N_2406,In_537,In_390);
or U2407 (N_2407,In_373,In_1488);
nor U2408 (N_2408,In_751,In_223);
and U2409 (N_2409,In_986,In_1439);
nor U2410 (N_2410,In_842,In_1035);
and U2411 (N_2411,In_868,In_356);
and U2412 (N_2412,In_294,In_818);
nor U2413 (N_2413,In_443,In_1435);
or U2414 (N_2414,In_194,In_863);
xnor U2415 (N_2415,In_40,In_551);
nand U2416 (N_2416,In_471,In_1026);
nor U2417 (N_2417,In_1162,In_1178);
or U2418 (N_2418,In_1280,In_949);
xor U2419 (N_2419,In_708,In_970);
nor U2420 (N_2420,In_1136,In_1055);
or U2421 (N_2421,In_188,In_1444);
nor U2422 (N_2422,In_777,In_71);
nor U2423 (N_2423,In_699,In_194);
nand U2424 (N_2424,In_956,In_197);
and U2425 (N_2425,In_583,In_755);
xor U2426 (N_2426,In_727,In_1290);
nor U2427 (N_2427,In_1055,In_1034);
xnor U2428 (N_2428,In_14,In_1057);
or U2429 (N_2429,In_318,In_292);
or U2430 (N_2430,In_360,In_1046);
or U2431 (N_2431,In_1131,In_77);
nand U2432 (N_2432,In_672,In_1212);
and U2433 (N_2433,In_139,In_549);
nand U2434 (N_2434,In_1145,In_1248);
or U2435 (N_2435,In_725,In_38);
nand U2436 (N_2436,In_1474,In_1039);
or U2437 (N_2437,In_609,In_1071);
nor U2438 (N_2438,In_1001,In_893);
xnor U2439 (N_2439,In_1261,In_1412);
nor U2440 (N_2440,In_611,In_626);
xnor U2441 (N_2441,In_1301,In_734);
nor U2442 (N_2442,In_1108,In_228);
nor U2443 (N_2443,In_984,In_64);
nand U2444 (N_2444,In_1159,In_1408);
nor U2445 (N_2445,In_172,In_1327);
or U2446 (N_2446,In_1451,In_497);
and U2447 (N_2447,In_1094,In_1327);
or U2448 (N_2448,In_1258,In_1205);
nor U2449 (N_2449,In_913,In_141);
nand U2450 (N_2450,In_400,In_583);
and U2451 (N_2451,In_1301,In_1484);
or U2452 (N_2452,In_57,In_804);
or U2453 (N_2453,In_793,In_958);
xor U2454 (N_2454,In_837,In_193);
nor U2455 (N_2455,In_423,In_734);
nor U2456 (N_2456,In_131,In_124);
xnor U2457 (N_2457,In_781,In_1440);
xnor U2458 (N_2458,In_992,In_148);
nand U2459 (N_2459,In_1282,In_884);
or U2460 (N_2460,In_841,In_353);
or U2461 (N_2461,In_970,In_621);
nor U2462 (N_2462,In_1108,In_1287);
xor U2463 (N_2463,In_1169,In_691);
nor U2464 (N_2464,In_840,In_1041);
nor U2465 (N_2465,In_549,In_231);
nand U2466 (N_2466,In_1103,In_1472);
nand U2467 (N_2467,In_91,In_1067);
and U2468 (N_2468,In_767,In_1419);
or U2469 (N_2469,In_1278,In_893);
nand U2470 (N_2470,In_147,In_919);
or U2471 (N_2471,In_686,In_285);
and U2472 (N_2472,In_749,In_962);
nand U2473 (N_2473,In_338,In_904);
xor U2474 (N_2474,In_741,In_43);
or U2475 (N_2475,In_710,In_35);
and U2476 (N_2476,In_1458,In_666);
nor U2477 (N_2477,In_286,In_975);
or U2478 (N_2478,In_298,In_79);
and U2479 (N_2479,In_152,In_1331);
or U2480 (N_2480,In_1354,In_1257);
nand U2481 (N_2481,In_1387,In_115);
or U2482 (N_2482,In_760,In_183);
xor U2483 (N_2483,In_1102,In_777);
and U2484 (N_2484,In_791,In_308);
nand U2485 (N_2485,In_978,In_1071);
nand U2486 (N_2486,In_354,In_474);
nor U2487 (N_2487,In_365,In_1410);
nor U2488 (N_2488,In_265,In_1327);
and U2489 (N_2489,In_1256,In_851);
or U2490 (N_2490,In_1336,In_774);
xor U2491 (N_2491,In_432,In_1254);
nor U2492 (N_2492,In_976,In_110);
or U2493 (N_2493,In_1321,In_1173);
and U2494 (N_2494,In_391,In_206);
nand U2495 (N_2495,In_463,In_1294);
nor U2496 (N_2496,In_999,In_479);
and U2497 (N_2497,In_1252,In_1304);
and U2498 (N_2498,In_375,In_848);
or U2499 (N_2499,In_514,In_452);
and U2500 (N_2500,In_358,In_307);
nand U2501 (N_2501,In_780,In_838);
xor U2502 (N_2502,In_408,In_164);
nand U2503 (N_2503,In_516,In_503);
nand U2504 (N_2504,In_848,In_430);
and U2505 (N_2505,In_817,In_799);
nand U2506 (N_2506,In_553,In_883);
nand U2507 (N_2507,In_406,In_500);
and U2508 (N_2508,In_65,In_57);
nand U2509 (N_2509,In_100,In_85);
or U2510 (N_2510,In_1445,In_697);
and U2511 (N_2511,In_545,In_1277);
nor U2512 (N_2512,In_1329,In_657);
and U2513 (N_2513,In_1475,In_438);
or U2514 (N_2514,In_398,In_1080);
nor U2515 (N_2515,In_878,In_380);
nor U2516 (N_2516,In_233,In_495);
nand U2517 (N_2517,In_1286,In_979);
nor U2518 (N_2518,In_1123,In_1411);
nor U2519 (N_2519,In_996,In_209);
nor U2520 (N_2520,In_712,In_1382);
or U2521 (N_2521,In_1331,In_211);
xor U2522 (N_2522,In_71,In_888);
nand U2523 (N_2523,In_1303,In_634);
nor U2524 (N_2524,In_516,In_220);
and U2525 (N_2525,In_1273,In_1422);
or U2526 (N_2526,In_1108,In_590);
nand U2527 (N_2527,In_807,In_74);
xnor U2528 (N_2528,In_170,In_577);
and U2529 (N_2529,In_605,In_162);
or U2530 (N_2530,In_200,In_1214);
and U2531 (N_2531,In_668,In_1209);
or U2532 (N_2532,In_1052,In_301);
nand U2533 (N_2533,In_1168,In_152);
nand U2534 (N_2534,In_412,In_58);
or U2535 (N_2535,In_723,In_91);
and U2536 (N_2536,In_443,In_938);
nor U2537 (N_2537,In_1406,In_111);
nor U2538 (N_2538,In_919,In_1021);
nor U2539 (N_2539,In_10,In_996);
and U2540 (N_2540,In_1013,In_661);
nand U2541 (N_2541,In_290,In_1322);
nor U2542 (N_2542,In_569,In_196);
nor U2543 (N_2543,In_571,In_431);
nor U2544 (N_2544,In_1486,In_145);
xor U2545 (N_2545,In_285,In_669);
nor U2546 (N_2546,In_719,In_897);
or U2547 (N_2547,In_1230,In_1486);
nand U2548 (N_2548,In_9,In_1031);
or U2549 (N_2549,In_809,In_146);
nor U2550 (N_2550,In_120,In_846);
or U2551 (N_2551,In_562,In_400);
or U2552 (N_2552,In_302,In_1159);
or U2553 (N_2553,In_318,In_707);
nand U2554 (N_2554,In_796,In_885);
and U2555 (N_2555,In_295,In_814);
nor U2556 (N_2556,In_39,In_1440);
and U2557 (N_2557,In_1284,In_1425);
and U2558 (N_2558,In_677,In_973);
nor U2559 (N_2559,In_485,In_545);
or U2560 (N_2560,In_1400,In_896);
nand U2561 (N_2561,In_23,In_612);
and U2562 (N_2562,In_1263,In_1249);
nor U2563 (N_2563,In_174,In_1372);
nor U2564 (N_2564,In_864,In_41);
or U2565 (N_2565,In_658,In_248);
or U2566 (N_2566,In_518,In_488);
and U2567 (N_2567,In_1044,In_1487);
nor U2568 (N_2568,In_72,In_742);
nor U2569 (N_2569,In_320,In_1319);
or U2570 (N_2570,In_1484,In_652);
nand U2571 (N_2571,In_1166,In_259);
nor U2572 (N_2572,In_1373,In_286);
or U2573 (N_2573,In_966,In_37);
xor U2574 (N_2574,In_935,In_593);
xor U2575 (N_2575,In_713,In_1038);
and U2576 (N_2576,In_168,In_600);
nand U2577 (N_2577,In_372,In_465);
nand U2578 (N_2578,In_416,In_12);
nor U2579 (N_2579,In_343,In_1189);
nand U2580 (N_2580,In_1238,In_1187);
nand U2581 (N_2581,In_803,In_973);
or U2582 (N_2582,In_958,In_396);
or U2583 (N_2583,In_459,In_176);
nand U2584 (N_2584,In_140,In_605);
nand U2585 (N_2585,In_1317,In_4);
and U2586 (N_2586,In_522,In_668);
nor U2587 (N_2587,In_928,In_35);
and U2588 (N_2588,In_941,In_677);
or U2589 (N_2589,In_1361,In_384);
nand U2590 (N_2590,In_397,In_17);
or U2591 (N_2591,In_866,In_887);
and U2592 (N_2592,In_409,In_29);
nand U2593 (N_2593,In_1489,In_1319);
and U2594 (N_2594,In_922,In_208);
nor U2595 (N_2595,In_1441,In_1223);
or U2596 (N_2596,In_635,In_1140);
xor U2597 (N_2597,In_1490,In_1433);
nand U2598 (N_2598,In_565,In_419);
nand U2599 (N_2599,In_1279,In_238);
xnor U2600 (N_2600,In_597,In_248);
or U2601 (N_2601,In_201,In_1298);
nor U2602 (N_2602,In_929,In_1001);
xor U2603 (N_2603,In_815,In_1081);
or U2604 (N_2604,In_209,In_178);
nor U2605 (N_2605,In_879,In_168);
or U2606 (N_2606,In_825,In_1492);
and U2607 (N_2607,In_259,In_709);
nand U2608 (N_2608,In_835,In_705);
or U2609 (N_2609,In_720,In_982);
and U2610 (N_2610,In_951,In_777);
nand U2611 (N_2611,In_1439,In_1114);
nor U2612 (N_2612,In_610,In_638);
nor U2613 (N_2613,In_584,In_151);
nor U2614 (N_2614,In_975,In_212);
nand U2615 (N_2615,In_486,In_528);
nor U2616 (N_2616,In_258,In_472);
xnor U2617 (N_2617,In_843,In_94);
nand U2618 (N_2618,In_1350,In_656);
and U2619 (N_2619,In_1190,In_471);
and U2620 (N_2620,In_250,In_170);
xnor U2621 (N_2621,In_171,In_1359);
and U2622 (N_2622,In_140,In_1272);
or U2623 (N_2623,In_1370,In_1018);
nor U2624 (N_2624,In_1496,In_1428);
or U2625 (N_2625,In_640,In_391);
nand U2626 (N_2626,In_665,In_1388);
or U2627 (N_2627,In_169,In_360);
and U2628 (N_2628,In_401,In_176);
and U2629 (N_2629,In_872,In_757);
nor U2630 (N_2630,In_44,In_802);
or U2631 (N_2631,In_217,In_38);
or U2632 (N_2632,In_1102,In_799);
nand U2633 (N_2633,In_1006,In_1190);
xnor U2634 (N_2634,In_1066,In_502);
or U2635 (N_2635,In_798,In_984);
and U2636 (N_2636,In_1434,In_446);
xor U2637 (N_2637,In_1350,In_263);
nand U2638 (N_2638,In_510,In_156);
nand U2639 (N_2639,In_706,In_903);
and U2640 (N_2640,In_915,In_957);
and U2641 (N_2641,In_1341,In_615);
and U2642 (N_2642,In_396,In_719);
nand U2643 (N_2643,In_1477,In_1460);
or U2644 (N_2644,In_926,In_145);
or U2645 (N_2645,In_862,In_584);
or U2646 (N_2646,In_1435,In_1427);
nand U2647 (N_2647,In_491,In_765);
xor U2648 (N_2648,In_55,In_831);
nand U2649 (N_2649,In_255,In_1248);
or U2650 (N_2650,In_517,In_74);
or U2651 (N_2651,In_1434,In_314);
nor U2652 (N_2652,In_1154,In_366);
nand U2653 (N_2653,In_1362,In_1032);
or U2654 (N_2654,In_310,In_1191);
or U2655 (N_2655,In_821,In_577);
nand U2656 (N_2656,In_661,In_11);
nor U2657 (N_2657,In_1063,In_122);
or U2658 (N_2658,In_144,In_982);
xor U2659 (N_2659,In_1009,In_388);
or U2660 (N_2660,In_272,In_580);
or U2661 (N_2661,In_1123,In_948);
or U2662 (N_2662,In_150,In_655);
nor U2663 (N_2663,In_235,In_1084);
or U2664 (N_2664,In_38,In_1062);
nor U2665 (N_2665,In_1050,In_1341);
nor U2666 (N_2666,In_403,In_756);
nor U2667 (N_2667,In_107,In_416);
nor U2668 (N_2668,In_802,In_167);
or U2669 (N_2669,In_1376,In_385);
nand U2670 (N_2670,In_614,In_73);
nor U2671 (N_2671,In_1499,In_6);
and U2672 (N_2672,In_1219,In_327);
and U2673 (N_2673,In_256,In_596);
or U2674 (N_2674,In_222,In_439);
nand U2675 (N_2675,In_1342,In_61);
or U2676 (N_2676,In_272,In_1315);
nand U2677 (N_2677,In_834,In_1258);
or U2678 (N_2678,In_1371,In_112);
nor U2679 (N_2679,In_1135,In_544);
nand U2680 (N_2680,In_138,In_468);
nor U2681 (N_2681,In_722,In_914);
nand U2682 (N_2682,In_281,In_1153);
and U2683 (N_2683,In_505,In_404);
and U2684 (N_2684,In_556,In_713);
or U2685 (N_2685,In_1003,In_718);
nor U2686 (N_2686,In_411,In_463);
or U2687 (N_2687,In_1452,In_613);
nor U2688 (N_2688,In_294,In_859);
and U2689 (N_2689,In_165,In_885);
nand U2690 (N_2690,In_1014,In_761);
xor U2691 (N_2691,In_84,In_1435);
or U2692 (N_2692,In_959,In_807);
or U2693 (N_2693,In_777,In_172);
nand U2694 (N_2694,In_413,In_159);
or U2695 (N_2695,In_1145,In_494);
nand U2696 (N_2696,In_774,In_528);
xnor U2697 (N_2697,In_379,In_572);
nor U2698 (N_2698,In_1182,In_865);
nand U2699 (N_2699,In_1225,In_1120);
nor U2700 (N_2700,In_1241,In_262);
nor U2701 (N_2701,In_1338,In_472);
nand U2702 (N_2702,In_176,In_601);
nor U2703 (N_2703,In_84,In_158);
and U2704 (N_2704,In_931,In_1259);
nand U2705 (N_2705,In_45,In_1492);
nor U2706 (N_2706,In_749,In_684);
and U2707 (N_2707,In_1021,In_492);
nor U2708 (N_2708,In_1354,In_1300);
nand U2709 (N_2709,In_1337,In_876);
xnor U2710 (N_2710,In_170,In_1400);
and U2711 (N_2711,In_171,In_1056);
nand U2712 (N_2712,In_1073,In_712);
nand U2713 (N_2713,In_529,In_692);
and U2714 (N_2714,In_868,In_1460);
xnor U2715 (N_2715,In_763,In_905);
nor U2716 (N_2716,In_390,In_457);
nand U2717 (N_2717,In_920,In_543);
and U2718 (N_2718,In_78,In_206);
nor U2719 (N_2719,In_443,In_468);
or U2720 (N_2720,In_1450,In_775);
or U2721 (N_2721,In_789,In_224);
and U2722 (N_2722,In_176,In_57);
nand U2723 (N_2723,In_662,In_1182);
nand U2724 (N_2724,In_975,In_332);
nand U2725 (N_2725,In_926,In_434);
and U2726 (N_2726,In_597,In_312);
nor U2727 (N_2727,In_424,In_790);
nand U2728 (N_2728,In_596,In_317);
nand U2729 (N_2729,In_600,In_1002);
nor U2730 (N_2730,In_1398,In_375);
nor U2731 (N_2731,In_937,In_850);
nor U2732 (N_2732,In_279,In_1335);
and U2733 (N_2733,In_659,In_1103);
and U2734 (N_2734,In_714,In_1494);
nand U2735 (N_2735,In_1074,In_472);
or U2736 (N_2736,In_741,In_1058);
nand U2737 (N_2737,In_351,In_1301);
or U2738 (N_2738,In_436,In_973);
nor U2739 (N_2739,In_1151,In_221);
or U2740 (N_2740,In_143,In_739);
nor U2741 (N_2741,In_263,In_1472);
nor U2742 (N_2742,In_1171,In_184);
or U2743 (N_2743,In_670,In_1088);
or U2744 (N_2744,In_527,In_883);
or U2745 (N_2745,In_1115,In_2);
and U2746 (N_2746,In_929,In_215);
xnor U2747 (N_2747,In_1110,In_1346);
nor U2748 (N_2748,In_1045,In_1014);
nor U2749 (N_2749,In_1446,In_1058);
nand U2750 (N_2750,In_1499,In_400);
nor U2751 (N_2751,In_365,In_1445);
nand U2752 (N_2752,In_669,In_268);
or U2753 (N_2753,In_54,In_1408);
nor U2754 (N_2754,In_701,In_19);
nand U2755 (N_2755,In_749,In_557);
nor U2756 (N_2756,In_172,In_304);
nand U2757 (N_2757,In_1365,In_338);
nand U2758 (N_2758,In_958,In_1002);
and U2759 (N_2759,In_794,In_48);
or U2760 (N_2760,In_893,In_745);
and U2761 (N_2761,In_1425,In_781);
and U2762 (N_2762,In_1423,In_1173);
xor U2763 (N_2763,In_1380,In_8);
and U2764 (N_2764,In_187,In_1013);
xnor U2765 (N_2765,In_627,In_1223);
or U2766 (N_2766,In_174,In_972);
nand U2767 (N_2767,In_38,In_300);
nor U2768 (N_2768,In_621,In_1428);
nor U2769 (N_2769,In_395,In_984);
and U2770 (N_2770,In_952,In_659);
xor U2771 (N_2771,In_1142,In_325);
or U2772 (N_2772,In_1345,In_1467);
and U2773 (N_2773,In_763,In_1056);
or U2774 (N_2774,In_1119,In_900);
or U2775 (N_2775,In_726,In_808);
or U2776 (N_2776,In_1142,In_1446);
nor U2777 (N_2777,In_919,In_1463);
nand U2778 (N_2778,In_1476,In_804);
nand U2779 (N_2779,In_258,In_647);
or U2780 (N_2780,In_1247,In_564);
nor U2781 (N_2781,In_473,In_384);
or U2782 (N_2782,In_660,In_815);
nand U2783 (N_2783,In_251,In_1350);
and U2784 (N_2784,In_573,In_697);
or U2785 (N_2785,In_184,In_977);
or U2786 (N_2786,In_1453,In_684);
nand U2787 (N_2787,In_1087,In_139);
nor U2788 (N_2788,In_1437,In_1242);
and U2789 (N_2789,In_613,In_575);
nand U2790 (N_2790,In_409,In_907);
nor U2791 (N_2791,In_177,In_693);
nor U2792 (N_2792,In_1118,In_410);
nand U2793 (N_2793,In_315,In_1353);
xnor U2794 (N_2794,In_15,In_1437);
xor U2795 (N_2795,In_932,In_1455);
and U2796 (N_2796,In_27,In_1423);
nor U2797 (N_2797,In_2,In_786);
nor U2798 (N_2798,In_934,In_17);
and U2799 (N_2799,In_496,In_10);
and U2800 (N_2800,In_418,In_596);
nor U2801 (N_2801,In_1135,In_690);
and U2802 (N_2802,In_689,In_1158);
and U2803 (N_2803,In_396,In_1138);
nor U2804 (N_2804,In_619,In_1323);
nor U2805 (N_2805,In_961,In_357);
nor U2806 (N_2806,In_602,In_570);
and U2807 (N_2807,In_294,In_100);
nor U2808 (N_2808,In_12,In_1461);
nor U2809 (N_2809,In_811,In_815);
nand U2810 (N_2810,In_685,In_718);
or U2811 (N_2811,In_708,In_549);
nand U2812 (N_2812,In_114,In_296);
or U2813 (N_2813,In_1286,In_190);
or U2814 (N_2814,In_1283,In_171);
xor U2815 (N_2815,In_414,In_756);
and U2816 (N_2816,In_703,In_1284);
nand U2817 (N_2817,In_327,In_787);
xor U2818 (N_2818,In_822,In_1367);
and U2819 (N_2819,In_288,In_100);
or U2820 (N_2820,In_594,In_1162);
or U2821 (N_2821,In_247,In_693);
nand U2822 (N_2822,In_659,In_1259);
xor U2823 (N_2823,In_1052,In_1309);
xnor U2824 (N_2824,In_188,In_1012);
and U2825 (N_2825,In_768,In_976);
or U2826 (N_2826,In_443,In_704);
xor U2827 (N_2827,In_1388,In_605);
nor U2828 (N_2828,In_910,In_71);
and U2829 (N_2829,In_302,In_1220);
nand U2830 (N_2830,In_16,In_1407);
and U2831 (N_2831,In_122,In_452);
and U2832 (N_2832,In_112,In_703);
nand U2833 (N_2833,In_1293,In_1265);
xor U2834 (N_2834,In_102,In_1485);
nor U2835 (N_2835,In_421,In_1130);
and U2836 (N_2836,In_220,In_767);
xnor U2837 (N_2837,In_50,In_899);
nand U2838 (N_2838,In_1240,In_12);
nor U2839 (N_2839,In_173,In_1164);
nor U2840 (N_2840,In_1400,In_902);
nand U2841 (N_2841,In_851,In_605);
nand U2842 (N_2842,In_1334,In_1041);
and U2843 (N_2843,In_175,In_955);
nand U2844 (N_2844,In_1147,In_662);
or U2845 (N_2845,In_1019,In_630);
nand U2846 (N_2846,In_521,In_669);
nor U2847 (N_2847,In_69,In_689);
or U2848 (N_2848,In_1433,In_870);
and U2849 (N_2849,In_1280,In_979);
nand U2850 (N_2850,In_423,In_882);
and U2851 (N_2851,In_222,In_94);
and U2852 (N_2852,In_402,In_496);
and U2853 (N_2853,In_576,In_1189);
nor U2854 (N_2854,In_1080,In_1110);
xnor U2855 (N_2855,In_1313,In_1286);
and U2856 (N_2856,In_740,In_1341);
nor U2857 (N_2857,In_1178,In_1192);
and U2858 (N_2858,In_1289,In_271);
nand U2859 (N_2859,In_1233,In_275);
nand U2860 (N_2860,In_182,In_1374);
nand U2861 (N_2861,In_249,In_901);
nand U2862 (N_2862,In_555,In_4);
nand U2863 (N_2863,In_542,In_428);
or U2864 (N_2864,In_945,In_1474);
and U2865 (N_2865,In_691,In_1296);
and U2866 (N_2866,In_231,In_286);
and U2867 (N_2867,In_738,In_1481);
and U2868 (N_2868,In_232,In_704);
nor U2869 (N_2869,In_441,In_1312);
or U2870 (N_2870,In_225,In_632);
xor U2871 (N_2871,In_1057,In_726);
and U2872 (N_2872,In_732,In_1111);
nand U2873 (N_2873,In_524,In_925);
nand U2874 (N_2874,In_86,In_31);
xnor U2875 (N_2875,In_1368,In_905);
xor U2876 (N_2876,In_1409,In_109);
xnor U2877 (N_2877,In_767,In_1102);
and U2878 (N_2878,In_111,In_1101);
and U2879 (N_2879,In_87,In_827);
or U2880 (N_2880,In_1066,In_1057);
xnor U2881 (N_2881,In_388,In_1442);
nand U2882 (N_2882,In_20,In_823);
and U2883 (N_2883,In_608,In_1329);
and U2884 (N_2884,In_1058,In_1342);
nor U2885 (N_2885,In_1250,In_311);
nand U2886 (N_2886,In_113,In_493);
nand U2887 (N_2887,In_1453,In_1454);
nor U2888 (N_2888,In_193,In_1131);
nand U2889 (N_2889,In_945,In_867);
xnor U2890 (N_2890,In_1377,In_1351);
and U2891 (N_2891,In_792,In_873);
or U2892 (N_2892,In_404,In_1319);
and U2893 (N_2893,In_598,In_1327);
nor U2894 (N_2894,In_931,In_874);
or U2895 (N_2895,In_764,In_1445);
xnor U2896 (N_2896,In_610,In_614);
nor U2897 (N_2897,In_658,In_743);
and U2898 (N_2898,In_905,In_330);
nor U2899 (N_2899,In_243,In_1286);
nor U2900 (N_2900,In_552,In_499);
nor U2901 (N_2901,In_1145,In_153);
nor U2902 (N_2902,In_1378,In_147);
or U2903 (N_2903,In_575,In_749);
nor U2904 (N_2904,In_619,In_334);
and U2905 (N_2905,In_371,In_1427);
and U2906 (N_2906,In_173,In_120);
or U2907 (N_2907,In_513,In_824);
nor U2908 (N_2908,In_1441,In_174);
and U2909 (N_2909,In_1324,In_1495);
nand U2910 (N_2910,In_491,In_772);
nand U2911 (N_2911,In_216,In_773);
nor U2912 (N_2912,In_324,In_576);
nor U2913 (N_2913,In_1048,In_936);
and U2914 (N_2914,In_506,In_1347);
and U2915 (N_2915,In_1095,In_121);
and U2916 (N_2916,In_1181,In_239);
nand U2917 (N_2917,In_188,In_557);
nand U2918 (N_2918,In_67,In_176);
and U2919 (N_2919,In_614,In_30);
nand U2920 (N_2920,In_582,In_1029);
and U2921 (N_2921,In_1124,In_344);
nor U2922 (N_2922,In_265,In_1082);
or U2923 (N_2923,In_78,In_553);
nand U2924 (N_2924,In_1200,In_680);
nand U2925 (N_2925,In_1297,In_374);
or U2926 (N_2926,In_1189,In_949);
nand U2927 (N_2927,In_488,In_1413);
nand U2928 (N_2928,In_657,In_169);
nand U2929 (N_2929,In_738,In_769);
nand U2930 (N_2930,In_69,In_646);
or U2931 (N_2931,In_273,In_798);
and U2932 (N_2932,In_956,In_819);
and U2933 (N_2933,In_888,In_19);
and U2934 (N_2934,In_1001,In_1451);
nor U2935 (N_2935,In_409,In_214);
nor U2936 (N_2936,In_1019,In_11);
xor U2937 (N_2937,In_277,In_1123);
and U2938 (N_2938,In_185,In_1338);
or U2939 (N_2939,In_1308,In_533);
and U2940 (N_2940,In_656,In_155);
nand U2941 (N_2941,In_1471,In_692);
and U2942 (N_2942,In_500,In_1228);
or U2943 (N_2943,In_1306,In_1032);
or U2944 (N_2944,In_884,In_1430);
and U2945 (N_2945,In_682,In_591);
nor U2946 (N_2946,In_1404,In_583);
and U2947 (N_2947,In_1260,In_1494);
nand U2948 (N_2948,In_680,In_1010);
xnor U2949 (N_2949,In_900,In_587);
and U2950 (N_2950,In_1065,In_1042);
and U2951 (N_2951,In_759,In_67);
nor U2952 (N_2952,In_1345,In_443);
nand U2953 (N_2953,In_50,In_325);
nor U2954 (N_2954,In_224,In_140);
nor U2955 (N_2955,In_296,In_1005);
nor U2956 (N_2956,In_281,In_1051);
nand U2957 (N_2957,In_1063,In_73);
nor U2958 (N_2958,In_1366,In_1239);
nor U2959 (N_2959,In_918,In_125);
and U2960 (N_2960,In_1006,In_227);
nand U2961 (N_2961,In_1043,In_1423);
nand U2962 (N_2962,In_492,In_751);
xor U2963 (N_2963,In_949,In_250);
and U2964 (N_2964,In_1297,In_470);
nand U2965 (N_2965,In_746,In_881);
and U2966 (N_2966,In_78,In_205);
nand U2967 (N_2967,In_251,In_220);
or U2968 (N_2968,In_956,In_1479);
and U2969 (N_2969,In_206,In_138);
nand U2970 (N_2970,In_500,In_138);
or U2971 (N_2971,In_1182,In_76);
and U2972 (N_2972,In_1440,In_1333);
or U2973 (N_2973,In_523,In_516);
nor U2974 (N_2974,In_539,In_156);
or U2975 (N_2975,In_128,In_1483);
nand U2976 (N_2976,In_329,In_559);
nor U2977 (N_2977,In_246,In_994);
and U2978 (N_2978,In_894,In_516);
nand U2979 (N_2979,In_1285,In_144);
or U2980 (N_2980,In_1423,In_8);
and U2981 (N_2981,In_185,In_838);
and U2982 (N_2982,In_772,In_496);
nor U2983 (N_2983,In_154,In_626);
nor U2984 (N_2984,In_1298,In_484);
nand U2985 (N_2985,In_595,In_1351);
or U2986 (N_2986,In_367,In_382);
nand U2987 (N_2987,In_168,In_30);
nand U2988 (N_2988,In_1148,In_282);
or U2989 (N_2989,In_1147,In_573);
and U2990 (N_2990,In_1207,In_800);
nand U2991 (N_2991,In_393,In_807);
xnor U2992 (N_2992,In_98,In_8);
nor U2993 (N_2993,In_573,In_1312);
nand U2994 (N_2994,In_1178,In_1395);
nand U2995 (N_2995,In_902,In_679);
nor U2996 (N_2996,In_1245,In_1129);
nor U2997 (N_2997,In_511,In_207);
and U2998 (N_2998,In_233,In_1446);
and U2999 (N_2999,In_1255,In_88);
nor U3000 (N_3000,N_2759,N_364);
nor U3001 (N_3001,N_2418,N_2343);
nor U3002 (N_3002,N_996,N_1004);
and U3003 (N_3003,N_1444,N_2023);
and U3004 (N_3004,N_2241,N_2489);
or U3005 (N_3005,N_2787,N_2146);
and U3006 (N_3006,N_868,N_679);
nor U3007 (N_3007,N_2056,N_1389);
or U3008 (N_3008,N_589,N_2028);
or U3009 (N_3009,N_217,N_1912);
and U3010 (N_3010,N_289,N_1371);
nand U3011 (N_3011,N_2790,N_2424);
nand U3012 (N_3012,N_1349,N_460);
xnor U3013 (N_3013,N_801,N_1047);
or U3014 (N_3014,N_1992,N_722);
nor U3015 (N_3015,N_2553,N_2898);
or U3016 (N_3016,N_971,N_2858);
and U3017 (N_3017,N_1573,N_163);
nor U3018 (N_3018,N_1896,N_2805);
xnor U3019 (N_3019,N_317,N_287);
and U3020 (N_3020,N_958,N_814);
or U3021 (N_3021,N_13,N_892);
xor U3022 (N_3022,N_2435,N_49);
nand U3023 (N_3023,N_1510,N_1862);
and U3024 (N_3024,N_1619,N_2698);
and U3025 (N_3025,N_1676,N_1018);
and U3026 (N_3026,N_949,N_1469);
or U3027 (N_3027,N_2935,N_681);
nor U3028 (N_3028,N_2048,N_1338);
or U3029 (N_3029,N_1023,N_2860);
and U3030 (N_3030,N_1309,N_1561);
and U3031 (N_3031,N_705,N_1863);
nor U3032 (N_3032,N_296,N_639);
nand U3033 (N_3033,N_1365,N_2332);
nor U3034 (N_3034,N_7,N_1544);
or U3035 (N_3035,N_800,N_424);
xor U3036 (N_3036,N_786,N_1078);
and U3037 (N_3037,N_1195,N_1694);
nand U3038 (N_3038,N_2824,N_1315);
nor U3039 (N_3039,N_428,N_1884);
and U3040 (N_3040,N_2509,N_201);
and U3041 (N_3041,N_1011,N_1519);
or U3042 (N_3042,N_1995,N_1598);
nor U3043 (N_3043,N_1575,N_2059);
nand U3044 (N_3044,N_2287,N_1837);
nor U3045 (N_3045,N_902,N_2189);
or U3046 (N_3046,N_2673,N_816);
nor U3047 (N_3047,N_1553,N_1723);
or U3048 (N_3048,N_2411,N_2491);
or U3049 (N_3049,N_2134,N_1702);
xnor U3050 (N_3050,N_1502,N_1638);
and U3051 (N_3051,N_2062,N_2609);
or U3052 (N_3052,N_107,N_80);
nor U3053 (N_3053,N_2019,N_785);
or U3054 (N_3054,N_2667,N_1650);
and U3055 (N_3055,N_1853,N_2794);
or U3056 (N_3056,N_1043,N_1302);
and U3057 (N_3057,N_1559,N_554);
nand U3058 (N_3058,N_2502,N_2925);
or U3059 (N_3059,N_576,N_2578);
nand U3060 (N_3060,N_2686,N_1207);
nor U3061 (N_3061,N_1600,N_2469);
and U3062 (N_3062,N_2327,N_521);
nand U3063 (N_3063,N_623,N_2599);
or U3064 (N_3064,N_922,N_2363);
nor U3065 (N_3065,N_1703,N_1258);
nor U3066 (N_3066,N_2468,N_728);
nor U3067 (N_3067,N_948,N_1554);
xnor U3068 (N_3068,N_1601,N_2608);
and U3069 (N_3069,N_1669,N_947);
nor U3070 (N_3070,N_2781,N_2990);
or U3071 (N_3071,N_40,N_351);
xor U3072 (N_3072,N_952,N_1754);
nand U3073 (N_3073,N_1227,N_488);
and U3074 (N_3074,N_198,N_2516);
and U3075 (N_3075,N_1939,N_261);
nor U3076 (N_3076,N_1766,N_706);
and U3077 (N_3077,N_454,N_336);
nor U3078 (N_3078,N_2982,N_2574);
nor U3079 (N_3079,N_78,N_826);
or U3080 (N_3080,N_2693,N_1535);
nand U3081 (N_3081,N_1945,N_223);
nand U3082 (N_3082,N_2588,N_2326);
or U3083 (N_3083,N_356,N_2124);
and U3084 (N_3084,N_1759,N_2712);
and U3085 (N_3085,N_1279,N_2194);
nand U3086 (N_3086,N_2811,N_206);
nand U3087 (N_3087,N_2709,N_1073);
nor U3088 (N_3088,N_2598,N_1022);
or U3089 (N_3089,N_2835,N_2862);
nor U3090 (N_3090,N_1910,N_841);
or U3091 (N_3091,N_2967,N_2658);
or U3092 (N_3092,N_1895,N_1820);
or U3093 (N_3093,N_1928,N_8);
or U3094 (N_3094,N_2520,N_2754);
nand U3095 (N_3095,N_1570,N_1873);
and U3096 (N_3096,N_1103,N_859);
nor U3097 (N_3097,N_1495,N_1807);
and U3098 (N_3098,N_453,N_1982);
and U3099 (N_3099,N_2844,N_2104);
nand U3100 (N_3100,N_2796,N_2427);
or U3101 (N_3101,N_427,N_2071);
or U3102 (N_3102,N_349,N_2764);
nand U3103 (N_3103,N_2710,N_1101);
and U3104 (N_3104,N_1641,N_422);
nor U3105 (N_3105,N_850,N_1574);
nor U3106 (N_3106,N_2616,N_2610);
nor U3107 (N_3107,N_858,N_625);
nand U3108 (N_3108,N_669,N_2002);
nand U3109 (N_3109,N_1938,N_1900);
or U3110 (N_3110,N_608,N_2786);
nor U3111 (N_3111,N_2973,N_89);
nor U3112 (N_3112,N_2840,N_1872);
or U3113 (N_3113,N_821,N_908);
or U3114 (N_3114,N_2950,N_398);
nand U3115 (N_3115,N_653,N_2174);
xor U3116 (N_3116,N_2838,N_1359);
and U3117 (N_3117,N_419,N_2089);
nor U3118 (N_3118,N_1556,N_2482);
nor U3119 (N_3119,N_575,N_1955);
nand U3120 (N_3120,N_920,N_1647);
or U3121 (N_3121,N_1784,N_2851);
nor U3122 (N_3122,N_846,N_1094);
and U3123 (N_3123,N_1805,N_2348);
nand U3124 (N_3124,N_110,N_382);
and U3125 (N_3125,N_686,N_1527);
or U3126 (N_3126,N_1626,N_871);
nor U3127 (N_3127,N_2305,N_2666);
or U3128 (N_3128,N_166,N_1864);
xor U3129 (N_3129,N_1871,N_2321);
xor U3130 (N_3130,N_670,N_2014);
nor U3131 (N_3131,N_2908,N_284);
or U3132 (N_3132,N_2687,N_1836);
nand U3133 (N_3133,N_1317,N_2121);
nor U3134 (N_3134,N_1024,N_2442);
nor U3135 (N_3135,N_1341,N_467);
nand U3136 (N_3136,N_1140,N_2038);
and U3137 (N_3137,N_1831,N_843);
nor U3138 (N_3138,N_1525,N_512);
and U3139 (N_3139,N_2142,N_1085);
nor U3140 (N_3140,N_2974,N_2190);
nand U3141 (N_3141,N_2379,N_852);
or U3142 (N_3142,N_842,N_2619);
xor U3143 (N_3143,N_923,N_2128);
and U3144 (N_3144,N_2708,N_221);
and U3145 (N_3145,N_77,N_1367);
nor U3146 (N_3146,N_98,N_2793);
nor U3147 (N_3147,N_1891,N_644);
and U3148 (N_3148,N_1454,N_2976);
and U3149 (N_3149,N_2009,N_1460);
nor U3150 (N_3150,N_1280,N_2197);
and U3151 (N_3151,N_1456,N_1827);
xor U3152 (N_3152,N_1824,N_914);
nand U3153 (N_3153,N_1613,N_1726);
nor U3154 (N_3154,N_1737,N_924);
xnor U3155 (N_3155,N_584,N_2373);
or U3156 (N_3156,N_343,N_1223);
and U3157 (N_3157,N_141,N_854);
or U3158 (N_3158,N_657,N_2515);
and U3159 (N_3159,N_2499,N_1698);
nand U3160 (N_3160,N_762,N_2707);
nor U3161 (N_3161,N_2702,N_215);
or U3162 (N_3162,N_2409,N_1564);
nand U3163 (N_3163,N_981,N_1607);
nor U3164 (N_3164,N_399,N_1700);
and U3165 (N_3165,N_1437,N_2383);
nand U3166 (N_3166,N_2745,N_514);
nand U3167 (N_3167,N_2843,N_1966);
xnor U3168 (N_3168,N_2888,N_1648);
nor U3169 (N_3169,N_724,N_31);
xnor U3170 (N_3170,N_2521,N_1017);
nor U3171 (N_3171,N_2073,N_370);
nor U3172 (N_3172,N_911,N_1363);
nand U3173 (N_3173,N_1815,N_1247);
nand U3174 (N_3174,N_1388,N_2818);
or U3175 (N_3175,N_1132,N_2087);
nand U3176 (N_3176,N_2837,N_2152);
nor U3177 (N_3177,N_687,N_2487);
or U3178 (N_3178,N_2177,N_2369);
xor U3179 (N_3179,N_1209,N_2641);
and U3180 (N_3180,N_2041,N_1181);
or U3181 (N_3181,N_550,N_2182);
and U3182 (N_3182,N_2946,N_726);
and U3183 (N_3183,N_2983,N_671);
and U3184 (N_3184,N_769,N_2889);
nor U3185 (N_3185,N_960,N_1337);
or U3186 (N_3186,N_1596,N_2725);
or U3187 (N_3187,N_1045,N_2088);
xnor U3188 (N_3188,N_388,N_2043);
nand U3189 (N_3189,N_1305,N_1960);
nand U3190 (N_3190,N_1801,N_1649);
and U3191 (N_3191,N_596,N_1438);
or U3192 (N_3192,N_822,N_2508);
or U3193 (N_3193,N_1899,N_183);
nor U3194 (N_3194,N_998,N_1918);
nand U3195 (N_3195,N_1521,N_2085);
and U3196 (N_3196,N_2620,N_131);
or U3197 (N_3197,N_1707,N_2807);
nor U3198 (N_3198,N_233,N_115);
or U3199 (N_3199,N_1640,N_877);
and U3200 (N_3200,N_2886,N_486);
xnor U3201 (N_3201,N_585,N_367);
or U3202 (N_3202,N_2031,N_2068);
nor U3203 (N_3203,N_594,N_1933);
or U3204 (N_3204,N_2461,N_283);
nor U3205 (N_3205,N_1929,N_2443);
or U3206 (N_3206,N_1028,N_1434);
or U3207 (N_3207,N_910,N_2757);
nand U3208 (N_3208,N_1120,N_2706);
or U3209 (N_3209,N_1930,N_2446);
xor U3210 (N_3210,N_1975,N_226);
and U3211 (N_3211,N_2721,N_1328);
nor U3212 (N_3212,N_2954,N_1458);
xor U3213 (N_3213,N_230,N_2863);
nor U3214 (N_3214,N_55,N_527);
nor U3215 (N_3215,N_507,N_2711);
nor U3216 (N_3216,N_281,N_220);
nand U3217 (N_3217,N_293,N_202);
and U3218 (N_3218,N_480,N_2390);
nand U3219 (N_3219,N_130,N_340);
nor U3220 (N_3220,N_1608,N_2808);
nor U3221 (N_3221,N_2692,N_165);
xnor U3222 (N_3222,N_2755,N_1625);
nand U3223 (N_3223,N_2522,N_2015);
nor U3224 (N_3224,N_777,N_100);
nand U3225 (N_3225,N_593,N_304);
nand U3226 (N_3226,N_1961,N_2067);
nor U3227 (N_3227,N_2205,N_93);
or U3228 (N_3228,N_809,N_1397);
nand U3229 (N_3229,N_856,N_2010);
and U3230 (N_3230,N_742,N_1228);
nand U3231 (N_3231,N_936,N_1522);
nor U3232 (N_3232,N_1627,N_1962);
xor U3233 (N_3233,N_2762,N_713);
and U3234 (N_3234,N_1500,N_1362);
or U3235 (N_3235,N_2664,N_1413);
nand U3236 (N_3236,N_1289,N_2382);
xor U3237 (N_3237,N_845,N_2841);
or U3238 (N_3238,N_4,N_276);
nor U3239 (N_3239,N_406,N_2101);
nor U3240 (N_3240,N_2751,N_1287);
and U3241 (N_3241,N_232,N_2330);
nand U3242 (N_3242,N_2743,N_1179);
and U3243 (N_3243,N_1386,N_1849);
xnor U3244 (N_3244,N_2810,N_2804);
or U3245 (N_3245,N_1800,N_1686);
and U3246 (N_3246,N_2675,N_1922);
and U3247 (N_3247,N_1000,N_2984);
or U3248 (N_3248,N_207,N_921);
and U3249 (N_3249,N_203,N_271);
nand U3250 (N_3250,N_2940,N_408);
nand U3251 (N_3251,N_700,N_1746);
or U3252 (N_3252,N_1074,N_2744);
and U3253 (N_3253,N_185,N_530);
or U3254 (N_3254,N_2283,N_2568);
and U3255 (N_3255,N_666,N_2919);
or U3256 (N_3256,N_1780,N_1044);
or U3257 (N_3257,N_2219,N_1133);
and U3258 (N_3258,N_2822,N_2921);
and U3259 (N_3259,N_1672,N_757);
nor U3260 (N_3260,N_274,N_2628);
or U3261 (N_3261,N_1409,N_1377);
and U3262 (N_3262,N_1212,N_2127);
nand U3263 (N_3263,N_1885,N_1829);
nand U3264 (N_3264,N_2380,N_146);
or U3265 (N_3265,N_1920,N_1875);
or U3266 (N_3266,N_731,N_17);
nand U3267 (N_3267,N_893,N_394);
and U3268 (N_3268,N_1186,N_1282);
and U3269 (N_3269,N_1124,N_1901);
and U3270 (N_3270,N_180,N_699);
and U3271 (N_3271,N_2812,N_67);
nand U3272 (N_3272,N_2122,N_2078);
nor U3273 (N_3273,N_725,N_1446);
and U3274 (N_3274,N_1634,N_1270);
or U3275 (N_3275,N_1897,N_499);
or U3276 (N_3276,N_1790,N_2130);
nor U3277 (N_3277,N_2245,N_108);
or U3278 (N_3278,N_2154,N_1346);
nand U3279 (N_3279,N_690,N_2923);
and U3280 (N_3280,N_2934,N_919);
xor U3281 (N_3281,N_942,N_2963);
nor U3282 (N_3282,N_2259,N_1802);
xnor U3283 (N_3283,N_224,N_2906);
nand U3284 (N_3284,N_799,N_2845);
and U3285 (N_3285,N_277,N_2053);
and U3286 (N_3286,N_1696,N_708);
and U3287 (N_3287,N_117,N_443);
and U3288 (N_3288,N_2301,N_2277);
or U3289 (N_3289,N_696,N_2105);
nand U3290 (N_3290,N_255,N_2825);
nor U3291 (N_3291,N_675,N_346);
or U3292 (N_3292,N_689,N_781);
and U3293 (N_3293,N_95,N_1128);
and U3294 (N_3294,N_2880,N_1983);
and U3295 (N_3295,N_2634,N_1785);
and U3296 (N_3296,N_1567,N_2267);
and U3297 (N_3297,N_2311,N_2584);
nor U3298 (N_3298,N_1032,N_2864);
and U3299 (N_3299,N_2187,N_2514);
xnor U3300 (N_3300,N_76,N_1109);
or U3301 (N_3301,N_825,N_896);
nor U3302 (N_3302,N_802,N_564);
or U3303 (N_3303,N_864,N_127);
nor U3304 (N_3304,N_1435,N_22);
nor U3305 (N_3305,N_1134,N_1479);
or U3306 (N_3306,N_92,N_2823);
nor U3307 (N_3307,N_1597,N_2054);
and U3308 (N_3308,N_1376,N_2848);
and U3309 (N_3309,N_1169,N_1027);
nor U3310 (N_3310,N_837,N_2920);
nand U3311 (N_3311,N_565,N_860);
and U3312 (N_3312,N_2632,N_2082);
or U3313 (N_3313,N_189,N_1468);
nand U3314 (N_3314,N_2447,N_962);
nand U3315 (N_3315,N_2660,N_1667);
or U3316 (N_3316,N_105,N_212);
nand U3317 (N_3317,N_12,N_1814);
or U3318 (N_3318,N_2342,N_2614);
and U3319 (N_3319,N_693,N_531);
or U3320 (N_3320,N_231,N_522);
or U3321 (N_3321,N_747,N_1972);
and U3322 (N_3322,N_548,N_1840);
nor U3323 (N_3323,N_2907,N_2270);
and U3324 (N_3324,N_2685,N_2);
or U3325 (N_3325,N_1997,N_2756);
or U3326 (N_3326,N_2116,N_2434);
and U3327 (N_3327,N_2561,N_2218);
xor U3328 (N_3328,N_2292,N_1963);
nand U3329 (N_3329,N_963,N_2341);
or U3330 (N_3330,N_1808,N_1447);
or U3331 (N_3331,N_1691,N_2775);
nand U3332 (N_3332,N_2642,N_2758);
nand U3333 (N_3333,N_1579,N_600);
nand U3334 (N_3334,N_1332,N_238);
nor U3335 (N_3335,N_121,N_1086);
xnor U3336 (N_3336,N_967,N_2081);
nand U3337 (N_3337,N_838,N_344);
nor U3338 (N_3338,N_216,N_2039);
nor U3339 (N_3339,N_1906,N_2297);
and U3340 (N_3340,N_1750,N_2791);
nor U3341 (N_3341,N_138,N_2057);
and U3342 (N_3342,N_2419,N_1455);
and U3343 (N_3343,N_2813,N_812);
and U3344 (N_3344,N_545,N_2374);
nand U3345 (N_3345,N_2669,N_2732);
nor U3346 (N_3346,N_1476,N_1311);
and U3347 (N_3347,N_2417,N_1793);
xnor U3348 (N_3348,N_1036,N_2674);
or U3349 (N_3349,N_46,N_1879);
nand U3350 (N_3350,N_1439,N_1865);
nand U3351 (N_3351,N_1200,N_2894);
xor U3352 (N_3352,N_2396,N_1019);
and U3353 (N_3353,N_1248,N_2252);
or U3354 (N_3354,N_1082,N_1615);
and U3355 (N_3355,N_2716,N_2454);
nor U3356 (N_3356,N_2233,N_2306);
nand U3357 (N_3357,N_1313,N_844);
nor U3358 (N_3358,N_2004,N_1464);
nor U3359 (N_3359,N_1775,N_2200);
nand U3360 (N_3360,N_1919,N_2814);
or U3361 (N_3361,N_1462,N_342);
xnor U3362 (N_3362,N_1610,N_2286);
or U3363 (N_3363,N_2913,N_318);
nand U3364 (N_3364,N_2493,N_2278);
nand U3365 (N_3365,N_1505,N_204);
nand U3366 (N_3366,N_642,N_2501);
and U3367 (N_3367,N_1484,N_1273);
nand U3368 (N_3368,N_2340,N_1490);
nand U3369 (N_3369,N_2517,N_1913);
or U3370 (N_3370,N_387,N_2135);
nor U3371 (N_3371,N_1566,N_377);
nor U3372 (N_3372,N_953,N_1720);
nor U3373 (N_3373,N_905,N_310);
or U3374 (N_3374,N_439,N_682);
xnor U3375 (N_3375,N_739,N_2567);
or U3376 (N_3376,N_213,N_1180);
nand U3377 (N_3377,N_1551,N_883);
or U3378 (N_3378,N_1580,N_2627);
nor U3379 (N_3379,N_2497,N_413);
and U3380 (N_3380,N_411,N_1653);
and U3381 (N_3381,N_2579,N_470);
nor U3382 (N_3382,N_518,N_1944);
or U3383 (N_3383,N_159,N_2312);
or U3384 (N_3384,N_595,N_139);
xor U3385 (N_3385,N_2942,N_1628);
nor U3386 (N_3386,N_2868,N_791);
and U3387 (N_3387,N_214,N_2269);
xor U3388 (N_3388,N_1705,N_715);
xnor U3389 (N_3389,N_472,N_1744);
or U3390 (N_3390,N_1954,N_583);
and U3391 (N_3391,N_1984,N_265);
nor U3392 (N_3392,N_1661,N_1249);
or U3393 (N_3393,N_599,N_2885);
or U3394 (N_3394,N_1390,N_2846);
or U3395 (N_3395,N_797,N_1989);
nand U3396 (N_3396,N_79,N_2314);
or U3397 (N_3397,N_1583,N_2478);
and U3398 (N_3398,N_1218,N_1799);
xor U3399 (N_3399,N_1693,N_2542);
xnor U3400 (N_3400,N_2961,N_975);
nand U3401 (N_3401,N_2604,N_2884);
and U3402 (N_3402,N_1417,N_1893);
or U3403 (N_3403,N_2652,N_1952);
and U3404 (N_3404,N_2358,N_1701);
or U3405 (N_3405,N_2927,N_1285);
nand U3406 (N_3406,N_1967,N_327);
or U3407 (N_3407,N_48,N_2153);
and U3408 (N_3408,N_886,N_126);
nor U3409 (N_3409,N_1635,N_2145);
or U3410 (N_3410,N_2831,N_249);
nor U3411 (N_3411,N_1546,N_1630);
or U3412 (N_3412,N_2097,N_2391);
nand U3413 (N_3413,N_2318,N_976);
and U3414 (N_3414,N_1451,N_2730);
xor U3415 (N_3415,N_537,N_851);
nor U3416 (N_3416,N_2836,N_1292);
and U3417 (N_3417,N_519,N_688);
nand U3418 (N_3418,N_94,N_2556);
nand U3419 (N_3419,N_494,N_683);
or U3420 (N_3420,N_997,N_2282);
nand U3421 (N_3421,N_1237,N_2621);
xnor U3422 (N_3422,N_2914,N_177);
and U3423 (N_3423,N_248,N_1709);
and U3424 (N_3424,N_1883,N_954);
xor U3425 (N_3425,N_2849,N_2981);
or U3426 (N_3426,N_466,N_1742);
xor U3427 (N_3427,N_794,N_1908);
nand U3428 (N_3428,N_325,N_1526);
or U3429 (N_3429,N_1493,N_621);
nand U3430 (N_3430,N_116,N_347);
or U3431 (N_3431,N_1374,N_866);
or U3432 (N_3432,N_678,N_2916);
xnor U3433 (N_3433,N_2163,N_602);
xnor U3434 (N_3434,N_1448,N_1145);
and U3435 (N_3435,N_1356,N_348);
nor U3436 (N_3436,N_2668,N_211);
xnor U3437 (N_3437,N_1355,N_429);
and U3438 (N_3438,N_1274,N_2761);
or U3439 (N_3439,N_2738,N_1969);
and U3440 (N_3440,N_374,N_2962);
or U3441 (N_3441,N_2180,N_2425);
nor U3442 (N_3442,N_2315,N_1163);
nor U3443 (N_3443,N_552,N_1216);
or U3444 (N_3444,N_182,N_2581);
xnor U3445 (N_3445,N_1229,N_2049);
or U3446 (N_3446,N_2240,N_2792);
xor U3447 (N_3447,N_2902,N_880);
nor U3448 (N_3448,N_1738,N_628);
nor U3449 (N_3449,N_322,N_2202);
xnor U3450 (N_3450,N_855,N_2861);
or U3451 (N_3451,N_1231,N_1220);
xor U3452 (N_3452,N_1131,N_2086);
nand U3453 (N_3453,N_750,N_1157);
nor U3454 (N_3454,N_1183,N_1443);
and U3455 (N_3455,N_909,N_1869);
nand U3456 (N_3456,N_1318,N_2084);
nor U3457 (N_3457,N_2797,N_2557);
nor U3458 (N_3458,N_2900,N_280);
and U3459 (N_3459,N_2636,N_81);
nand U3460 (N_3460,N_1414,N_2834);
nand U3461 (N_3461,N_2830,N_848);
or U3462 (N_3462,N_28,N_2203);
or U3463 (N_3463,N_906,N_2821);
nor U3464 (N_3464,N_2904,N_1215);
nor U3465 (N_3465,N_533,N_1030);
and U3466 (N_3466,N_1143,N_912);
nand U3467 (N_3467,N_2550,N_2030);
or U3468 (N_3468,N_1902,N_601);
and U3469 (N_3469,N_2302,N_1704);
and U3470 (N_3470,N_2191,N_409);
and U3471 (N_3471,N_1106,N_1876);
nand U3472 (N_3472,N_616,N_2503);
nand U3473 (N_3473,N_1093,N_1096);
xnor U3474 (N_3474,N_1271,N_1189);
and U3475 (N_3475,N_2859,N_2631);
nand U3476 (N_3476,N_504,N_1010);
or U3477 (N_3477,N_2701,N_2365);
nand U3478 (N_3478,N_1416,N_169);
nor U3479 (N_3479,N_1867,N_2785);
xor U3480 (N_3480,N_2881,N_1167);
nand U3481 (N_3481,N_2000,N_974);
or U3482 (N_3482,N_2320,N_2696);
xnor U3483 (N_3483,N_1796,N_2734);
nand U3484 (N_3484,N_2271,N_1830);
xnor U3485 (N_3485,N_1839,N_2248);
and U3486 (N_3486,N_1540,N_1431);
nor U3487 (N_3487,N_235,N_1772);
or U3488 (N_3488,N_1735,N_1013);
nand U3489 (N_3489,N_292,N_2255);
and U3490 (N_3490,N_2159,N_452);
nand U3491 (N_3491,N_2899,N_2729);
nor U3492 (N_3492,N_2799,N_234);
and U3493 (N_3493,N_1734,N_418);
nor U3494 (N_3494,N_2648,N_604);
nand U3495 (N_3495,N_1114,N_793);
or U3496 (N_3496,N_1298,N_259);
xnor U3497 (N_3497,N_1344,N_2044);
and U3498 (N_3498,N_1364,N_1226);
nand U3499 (N_3499,N_503,N_359);
and U3500 (N_3500,N_38,N_1401);
nor U3501 (N_3501,N_775,N_1283);
nor U3502 (N_3502,N_626,N_561);
nor U3503 (N_3503,N_2387,N_2422);
xor U3504 (N_3504,N_560,N_2720);
nand U3505 (N_3505,N_766,N_939);
and U3506 (N_3506,N_30,N_2518);
nand U3507 (N_3507,N_581,N_1685);
nand U3508 (N_3508,N_2026,N_2242);
and U3509 (N_3509,N_1812,N_1199);
or U3510 (N_3510,N_1457,N_236);
xor U3511 (N_3511,N_331,N_312);
or U3512 (N_3512,N_2724,N_75);
or U3513 (N_3513,N_2865,N_1675);
and U3514 (N_3514,N_2486,N_2217);
or U3515 (N_3515,N_897,N_2257);
and U3516 (N_3516,N_1265,N_1187);
nor U3517 (N_3517,N_282,N_372);
nand U3518 (N_3518,N_1550,N_332);
nand U3519 (N_3519,N_2114,N_587);
or U3520 (N_3520,N_2749,N_733);
nand U3521 (N_3521,N_2959,N_2592);
and U3522 (N_3522,N_1111,N_2855);
or U3523 (N_3523,N_991,N_1266);
nor U3524 (N_3524,N_2186,N_250);
xnor U3525 (N_3525,N_1005,N_1655);
and U3526 (N_3526,N_1136,N_995);
or U3527 (N_3527,N_1402,N_665);
xnor U3528 (N_3528,N_1436,N_2661);
xnor U3529 (N_3529,N_1507,N_2137);
nand U3530 (N_3530,N_1925,N_1316);
nor U3531 (N_3531,N_738,N_827);
and U3532 (N_3532,N_2875,N_931);
or U3533 (N_3533,N_2776,N_2370);
or U3534 (N_3534,N_2997,N_1450);
nor U3535 (N_3535,N_2926,N_2008);
nand U3536 (N_3536,N_2994,N_339);
nand U3537 (N_3537,N_990,N_729);
or U3538 (N_3538,N_184,N_2551);
nand U3539 (N_3539,N_2571,N_102);
and U3540 (N_3540,N_1681,N_1465);
xnor U3541 (N_3541,N_2354,N_1420);
xor U3542 (N_3542,N_1924,N_607);
or U3543 (N_3543,N_2630,N_2288);
nand U3544 (N_3544,N_39,N_555);
nor U3545 (N_3545,N_1576,N_1588);
nand U3546 (N_3546,N_2024,N_2459);
or U3547 (N_3547,N_2157,N_2943);
nor U3548 (N_3548,N_1141,N_833);
nand U3549 (N_3549,N_1524,N_2386);
and U3550 (N_3550,N_535,N_651);
nor U3551 (N_3551,N_2236,N_2275);
or U3552 (N_3552,N_1297,N_2265);
nor U3553 (N_3553,N_502,N_1225);
nor U3554 (N_3554,N_2856,N_1798);
nor U3555 (N_3555,N_1463,N_556);
and U3556 (N_3556,N_1406,N_1585);
or U3557 (N_3557,N_1581,N_240);
and U3558 (N_3558,N_1471,N_1087);
nand U3559 (N_3559,N_1779,N_1841);
nand U3560 (N_3560,N_2770,N_1936);
nor U3561 (N_3561,N_869,N_654);
xnor U3562 (N_3562,N_440,N_2635);
or U3563 (N_3563,N_1129,N_889);
or U3564 (N_3564,N_1384,N_2753);
xnor U3565 (N_3565,N_884,N_1222);
nor U3566 (N_3566,N_2423,N_1089);
xnor U3567 (N_3567,N_2979,N_2966);
xnor U3568 (N_3568,N_573,N_2677);
nand U3569 (N_3569,N_1033,N_2091);
xnor U3570 (N_3570,N_2784,N_298);
or U3571 (N_3571,N_2742,N_129);
nor U3572 (N_3572,N_904,N_239);
or U3573 (N_3573,N_2465,N_813);
nand U3574 (N_3574,N_133,N_1856);
or U3575 (N_3575,N_2910,N_2480);
nor U3576 (N_3576,N_3,N_1515);
or U3577 (N_3577,N_2371,N_2151);
nand U3578 (N_3578,N_2460,N_541);
nand U3579 (N_3579,N_2466,N_200);
or U3580 (N_3580,N_160,N_1488);
nand U3581 (N_3581,N_562,N_147);
and U3582 (N_3582,N_1244,N_1278);
nand U3583 (N_3583,N_85,N_900);
and U3584 (N_3584,N_2644,N_425);
xnor U3585 (N_3585,N_2980,N_1260);
or U3586 (N_3586,N_720,N_1979);
and U3587 (N_3587,N_1104,N_326);
and U3588 (N_3588,N_103,N_1589);
nor U3589 (N_3589,N_1007,N_1325);
or U3590 (N_3590,N_2511,N_1304);
or U3591 (N_3591,N_1715,N_1810);
nand U3592 (N_3592,N_2451,N_618);
nand U3593 (N_3593,N_817,N_549);
or U3594 (N_3594,N_1898,N_568);
nand U3595 (N_3595,N_2367,N_1753);
nand U3596 (N_3596,N_376,N_396);
nor U3597 (N_3597,N_228,N_2325);
nor U3598 (N_3598,N_1404,N_787);
and U3599 (N_3599,N_2251,N_2211);
xor U3600 (N_3600,N_2229,N_1532);
and U3601 (N_3601,N_2562,N_59);
nand U3602 (N_3602,N_2603,N_2587);
and U3603 (N_3603,N_1964,N_2595);
nand U3604 (N_3604,N_2680,N_1198);
or U3605 (N_3605,N_1060,N_506);
nand U3606 (N_3606,N_2506,N_627);
or U3607 (N_3607,N_2395,N_2408);
nand U3608 (N_3608,N_903,N_2874);
nand U3609 (N_3609,N_2789,N_2239);
xor U3610 (N_3610,N_2530,N_1461);
and U3611 (N_3611,N_1217,N_64);
nand U3612 (N_3612,N_316,N_784);
and U3613 (N_3613,N_961,N_363);
and U3614 (N_3614,N_1254,N_915);
nor U3615 (N_3615,N_1684,N_1035);
nand U3616 (N_3616,N_369,N_2022);
or U3617 (N_3617,N_2298,N_727);
nand U3618 (N_3618,N_1623,N_935);
or U3619 (N_3619,N_229,N_1381);
xnor U3620 (N_3620,N_431,N_1501);
nor U3621 (N_3621,N_2911,N_1843);
xor U3622 (N_3622,N_2820,N_2679);
nand U3623 (N_3623,N_1821,N_1039);
nor U3624 (N_3624,N_150,N_2347);
and U3625 (N_3625,N_2853,N_756);
nor U3626 (N_3626,N_2324,N_2083);
nand U3627 (N_3627,N_2307,N_187);
nor U3628 (N_3628,N_523,N_1541);
nor U3629 (N_3629,N_1155,N_2398);
xor U3630 (N_3630,N_1868,N_44);
nand U3631 (N_3631,N_420,N_51);
nand U3632 (N_3632,N_2025,N_867);
nor U3633 (N_3633,N_455,N_106);
nand U3634 (N_3634,N_505,N_2334);
nor U3635 (N_3635,N_1208,N_1858);
and U3636 (N_3636,N_2879,N_482);
nand U3637 (N_3637,N_1243,N_2098);
and U3638 (N_3638,N_1182,N_2160);
or U3639 (N_3639,N_2118,N_1122);
or U3640 (N_3640,N_2998,N_1393);
nor U3641 (N_3641,N_740,N_1211);
or U3642 (N_3642,N_368,N_2213);
and U3643 (N_3643,N_194,N_1990);
and U3644 (N_3644,N_763,N_929);
nand U3645 (N_3645,N_2477,N_2847);
nand U3646 (N_3646,N_366,N_2777);
nand U3647 (N_3647,N_1822,N_43);
and U3648 (N_3648,N_2339,N_119);
nand U3649 (N_3649,N_1603,N_291);
or U3650 (N_3650,N_1817,N_2072);
or U3651 (N_3651,N_767,N_2570);
nor U3652 (N_3652,N_2136,N_188);
nor U3653 (N_3653,N_603,N_475);
nand U3654 (N_3654,N_2412,N_1860);
and U3655 (N_3655,N_389,N_1624);
nor U3656 (N_3656,N_2075,N_2032);
xnor U3657 (N_3657,N_222,N_539);
and U3658 (N_3658,N_979,N_1851);
or U3659 (N_3659,N_1774,N_2103);
and U3660 (N_3660,N_2402,N_1503);
nor U3661 (N_3661,N_624,N_631);
or U3662 (N_3662,N_677,N_1513);
or U3663 (N_3663,N_648,N_1776);
nor U3664 (N_3664,N_1529,N_1762);
xnor U3665 (N_3665,N_2254,N_442);
nor U3666 (N_3666,N_1866,N_362);
nand U3667 (N_3667,N_2768,N_2975);
nand U3668 (N_3668,N_1160,N_2523);
nand U3669 (N_3669,N_1320,N_2450);
and U3670 (N_3670,N_879,N_1826);
nand U3671 (N_3671,N_751,N_1430);
or U3672 (N_3672,N_510,N_18);
xor U3673 (N_3673,N_69,N_2129);
nand U3674 (N_3674,N_2212,N_2527);
and U3675 (N_3675,N_1714,N_2993);
xor U3676 (N_3676,N_1107,N_917);
and U3677 (N_3677,N_965,N_2498);
xor U3678 (N_3678,N_1953,N_1327);
or U3679 (N_3679,N_335,N_2826);
nand U3680 (N_3680,N_1764,N_1637);
or U3681 (N_3681,N_2633,N_2951);
nor U3682 (N_3682,N_476,N_1572);
and U3683 (N_3683,N_1803,N_91);
nor U3684 (N_3684,N_2164,N_2649);
nor U3685 (N_3685,N_2586,N_1880);
or U3686 (N_3686,N_153,N_1547);
xor U3687 (N_3687,N_2704,N_2029);
nand U3688 (N_3688,N_1769,N_1656);
or U3689 (N_3689,N_1053,N_417);
nand U3690 (N_3690,N_2170,N_643);
and U3691 (N_3691,N_2901,N_2280);
nor U3692 (N_3692,N_566,N_383);
or U3693 (N_3693,N_579,N_2876);
and U3694 (N_3694,N_2596,N_1116);
xnor U3695 (N_3695,N_140,N_135);
or U3696 (N_3696,N_577,N_307);
or U3697 (N_3697,N_1716,N_2351);
nor U3698 (N_3698,N_901,N_1760);
nand U3699 (N_3699,N_872,N_2033);
nand U3700 (N_3700,N_2662,N_1003);
xnor U3701 (N_3701,N_2705,N_798);
or U3702 (N_3702,N_2475,N_2591);
and U3703 (N_3703,N_2999,N_2051);
xnor U3704 (N_3704,N_134,N_474);
and U3705 (N_3705,N_630,N_1040);
and U3706 (N_3706,N_2185,N_477);
and U3707 (N_3707,N_392,N_1146);
or U3708 (N_3708,N_2891,N_1380);
or U3709 (N_3709,N_1097,N_1937);
xnor U3710 (N_3710,N_260,N_245);
nand U3711 (N_3711,N_1126,N_1825);
and U3712 (N_3712,N_2657,N_2594);
or U3713 (N_3713,N_1408,N_27);
nor U3714 (N_3714,N_1202,N_16);
or U3715 (N_3715,N_487,N_158);
nand U3716 (N_3716,N_973,N_1171);
nand U3717 (N_3717,N_711,N_2535);
nor U3718 (N_3718,N_196,N_964);
and U3719 (N_3719,N_1517,N_1110);
and U3720 (N_3720,N_1411,N_1663);
nand U3721 (N_3721,N_73,N_2394);
nand U3722 (N_3722,N_1959,N_2750);
nand U3723 (N_3723,N_172,N_526);
and U3724 (N_3724,N_1643,N_1245);
nand U3725 (N_3725,N_2924,N_2123);
and U3726 (N_3726,N_2890,N_114);
and U3727 (N_3727,N_1453,N_635);
nor U3728 (N_3728,N_1235,N_444);
nand U3729 (N_3729,N_916,N_1747);
or U3730 (N_3730,N_2102,N_2095);
or U3731 (N_3731,N_26,N_2948);
nor U3732 (N_3732,N_124,N_1782);
and U3733 (N_3733,N_2333,N_582);
xor U3734 (N_3734,N_2214,N_2645);
and U3735 (N_3735,N_266,N_1692);
nor U3736 (N_3736,N_1552,N_2580);
xnor U3737 (N_3737,N_640,N_2149);
nor U3738 (N_3738,N_2646,N_2106);
nand U3739 (N_3739,N_171,N_528);
nand U3740 (N_3740,N_992,N_2462);
nand U3741 (N_3741,N_2590,N_1314);
xor U3742 (N_3742,N_1269,N_1075);
nor U3743 (N_3743,N_2074,N_2801);
nor U3744 (N_3744,N_894,N_2220);
nand U3745 (N_3745,N_2079,N_534);
nand U3746 (N_3746,N_1072,N_1537);
xor U3747 (N_3747,N_2989,N_496);
nor U3748 (N_3748,N_831,N_1548);
nand U3749 (N_3749,N_571,N_2540);
nand U3750 (N_3750,N_2575,N_2047);
nor U3751 (N_3751,N_1422,N_591);
xnor U3752 (N_3752,N_704,N_2819);
and U3753 (N_3753,N_2654,N_456);
or U3754 (N_3754,N_1980,N_525);
and U3755 (N_3755,N_2345,N_353);
nand U3756 (N_3756,N_270,N_2006);
or U3757 (N_3757,N_1842,N_792);
or U3758 (N_3758,N_765,N_930);
nor U3759 (N_3759,N_761,N_60);
or U3760 (N_3760,N_1683,N_982);
nor U3761 (N_3761,N_1063,N_2472);
and U3762 (N_3762,N_1256,N_580);
or U3763 (N_3763,N_1395,N_1412);
nand U3764 (N_3764,N_2147,N_2682);
xor U3765 (N_3765,N_2944,N_1834);
xor U3766 (N_3766,N_2737,N_984);
nor U3767 (N_3767,N_1291,N_1788);
nor U3768 (N_3768,N_1894,N_1612);
or U3769 (N_3769,N_684,N_2613);
and U3770 (N_3770,N_1833,N_772);
and U3771 (N_3771,N_2181,N_2372);
nor U3772 (N_3772,N_2210,N_241);
or U3773 (N_3773,N_2545,N_500);
and U3774 (N_3774,N_1425,N_52);
nor U3775 (N_3775,N_32,N_421);
and U3776 (N_3776,N_818,N_1330);
nand U3777 (N_3777,N_2410,N_650);
and U3778 (N_3778,N_1015,N_1172);
and U3779 (N_3779,N_770,N_493);
nor U3780 (N_3780,N_303,N_1009);
or U3781 (N_3781,N_1931,N_2143);
or U3782 (N_3782,N_2569,N_2223);
or U3783 (N_3783,N_2204,N_258);
xor U3784 (N_3784,N_1445,N_2651);
xor U3785 (N_3785,N_1911,N_710);
or U3786 (N_3786,N_511,N_446);
and U3787 (N_3787,N_532,N_1850);
and U3788 (N_3788,N_161,N_162);
nand U3789 (N_3789,N_2249,N_1923);
or U3790 (N_3790,N_2261,N_714);
or U3791 (N_3791,N_609,N_2231);
nand U3792 (N_3792,N_1350,N_1699);
and U3793 (N_3793,N_2986,N_2547);
and U3794 (N_3794,N_338,N_2256);
nand U3795 (N_3795,N_2625,N_1161);
xnor U3796 (N_3796,N_1604,N_2464);
and U3797 (N_3797,N_2100,N_796);
or U3798 (N_3798,N_1861,N_2576);
nand U3799 (N_3799,N_2647,N_2295);
nor U3800 (N_3800,N_50,N_2534);
nand U3801 (N_3801,N_1264,N_2238);
nand U3802 (N_3802,N_1941,N_1741);
and U3803 (N_3803,N_498,N_668);
and U3804 (N_3804,N_2718,N_1947);
nor U3805 (N_3805,N_2828,N_1);
and U3806 (N_3806,N_795,N_1021);
xnor U3807 (N_3807,N_2296,N_2939);
or U3808 (N_3808,N_2558,N_125);
nand U3809 (N_3809,N_1934,N_2110);
and U3810 (N_3810,N_2546,N_2003);
or U3811 (N_3811,N_2001,N_709);
or U3812 (N_3812,N_253,N_1232);
nor U3813 (N_3813,N_2247,N_308);
or U3814 (N_3814,N_1342,N_1644);
nand U3815 (N_3815,N_1385,N_697);
and U3816 (N_3816,N_2650,N_1068);
and U3817 (N_3817,N_1755,N_1213);
xor U3818 (N_3818,N_2193,N_2175);
or U3819 (N_3819,N_590,N_987);
or U3820 (N_3820,N_1993,N_2310);
nand U3821 (N_3821,N_227,N_2779);
nand U3822 (N_3822,N_1516,N_2206);
and U3823 (N_3823,N_2148,N_538);
nand U3824 (N_3824,N_1432,N_1633);
or U3825 (N_3825,N_2260,N_2329);
or U3826 (N_3826,N_2065,N_1196);
nand U3827 (N_3827,N_748,N_2740);
and U3828 (N_3828,N_2560,N_2526);
or U3829 (N_3829,N_1062,N_2829);
and U3830 (N_3830,N_1852,N_2359);
or U3831 (N_3831,N_1100,N_2895);
and U3832 (N_3832,N_1398,N_529);
and U3833 (N_3833,N_2795,N_1728);
or U3834 (N_3834,N_2050,N_1299);
or U3835 (N_3835,N_1054,N_695);
nand U3836 (N_3836,N_2413,N_333);
xor U3837 (N_3837,N_2356,N_737);
or U3838 (N_3838,N_1823,N_2201);
nor U3839 (N_3839,N_2076,N_2833);
nor U3840 (N_3840,N_1158,N_2766);
and U3841 (N_3841,N_2771,N_1261);
nor U3842 (N_3842,N_2572,N_2012);
nor U3843 (N_3843,N_2872,N_2479);
and U3844 (N_3844,N_1905,N_1340);
or U3845 (N_3845,N_337,N_1323);
or U3846 (N_3846,N_84,N_2816);
nor U3847 (N_3847,N_1441,N_1470);
nor U3848 (N_3848,N_1275,N_1399);
and U3849 (N_3849,N_823,N_2289);
or U3850 (N_3850,N_2452,N_2376);
nand U3851 (N_3851,N_1577,N_2384);
xnor U3852 (N_3852,N_1331,N_2453);
or U3853 (N_3853,N_933,N_155);
and U3854 (N_3854,N_1391,N_1303);
nor U3855 (N_3855,N_1907,N_2096);
nand U3856 (N_3856,N_2896,N_2532);
nand U3857 (N_3857,N_329,N_1483);
and U3858 (N_3858,N_297,N_717);
nor U3859 (N_3859,N_2234,N_1804);
and U3860 (N_3860,N_1347,N_414);
nand U3861 (N_3861,N_1407,N_927);
and U3862 (N_3862,N_2713,N_457);
or U3863 (N_3863,N_225,N_181);
xnor U3864 (N_3864,N_1631,N_2739);
or U3865 (N_3865,N_874,N_2331);
nand U3866 (N_3866,N_2733,N_136);
or U3867 (N_3867,N_497,N_1307);
and U3868 (N_3868,N_1730,N_1251);
or U3869 (N_3869,N_1943,N_1818);
nand U3870 (N_3870,N_66,N_1162);
xnor U3871 (N_3871,N_2525,N_1125);
and U3872 (N_3872,N_2171,N_898);
or U3873 (N_3873,N_458,N_1088);
nor U3874 (N_3874,N_945,N_741);
nor U3875 (N_3875,N_2774,N_508);
nor U3876 (N_3876,N_540,N_569);
or U3877 (N_3877,N_2035,N_805);
nand U3878 (N_3878,N_559,N_242);
nand U3879 (N_3879,N_1809,N_862);
or U3880 (N_3880,N_1197,N_1562);
nand U3881 (N_3881,N_2883,N_1084);
nor U3882 (N_3882,N_1221,N_193);
and U3883 (N_3883,N_1002,N_1789);
nand U3884 (N_3884,N_2593,N_269);
nor U3885 (N_3885,N_1882,N_2629);
nor U3886 (N_3886,N_262,N_2438);
nor U3887 (N_3887,N_2937,N_2912);
nor U3888 (N_3888,N_2752,N_662);
or U3889 (N_3889,N_6,N_611);
or U3890 (N_3890,N_2034,N_1058);
or U3891 (N_3891,N_1729,N_1657);
xor U3892 (N_3892,N_1418,N_2870);
nand U3893 (N_3893,N_2406,N_2436);
nor U3894 (N_3894,N_2235,N_2199);
nor U3895 (N_3895,N_2947,N_811);
and U3896 (N_3896,N_132,N_1518);
nand U3897 (N_3897,N_2139,N_178);
nor U3898 (N_3898,N_612,N_179);
nand U3899 (N_3899,N_1680,N_1150);
or U3900 (N_3900,N_2640,N_2773);
and U3901 (N_3901,N_2415,N_659);
and U3902 (N_3902,N_2385,N_1605);
xnor U3903 (N_3903,N_68,N_2842);
nor U3904 (N_3904,N_1533,N_2728);
nor U3905 (N_3905,N_1077,N_1080);
nand U3906 (N_3906,N_1166,N_2703);
or U3907 (N_3907,N_806,N_661);
and U3908 (N_3908,N_1083,N_2458);
or U3909 (N_3909,N_1770,N_2892);
nand U3910 (N_3910,N_2854,N_1671);
nor U3911 (N_3911,N_490,N_2237);
nor U3912 (N_3912,N_1486,N_664);
nor U3913 (N_3913,N_256,N_2167);
or U3914 (N_3914,N_1660,N_2467);
and U3915 (N_3915,N_174,N_536);
xor U3916 (N_3916,N_2299,N_197);
and U3917 (N_3917,N_2782,N_2215);
or U3918 (N_3918,N_2131,N_712);
nor U3919 (N_3919,N_1971,N_173);
nand U3920 (N_3920,N_588,N_1646);
or U3921 (N_3921,N_1568,N_615);
nand U3922 (N_3922,N_2209,N_524);
nand U3923 (N_3923,N_2357,N_1144);
nand U3924 (N_3924,N_1763,N_1970);
and U3925 (N_3925,N_45,N_1542);
nand U3926 (N_3926,N_2061,N_1813);
xor U3927 (N_3927,N_1481,N_1816);
nor U3928 (N_3928,N_634,N_2470);
nor U3929 (N_3929,N_1545,N_1115);
and U3930 (N_3930,N_1306,N_2389);
nor U3931 (N_3931,N_2968,N_1855);
nor U3932 (N_3932,N_1277,N_2871);
and U3933 (N_3933,N_320,N_288);
or U3934 (N_3934,N_605,N_25);
or U3935 (N_3935,N_2284,N_1154);
nand U3936 (N_3936,N_63,N_199);
and U3937 (N_3937,N_1061,N_2021);
or U3938 (N_3938,N_2996,N_2941);
xnor U3939 (N_3939,N_2537,N_1678);
nand U3940 (N_3940,N_1006,N_2504);
or U3941 (N_3941,N_1878,N_1373);
or U3942 (N_3942,N_1139,N_875);
or U3943 (N_3943,N_1958,N_2168);
or U3944 (N_3944,N_449,N_663);
nor U3945 (N_3945,N_464,N_2138);
and U3946 (N_3946,N_1361,N_1038);
nand U3947 (N_3947,N_2027,N_365);
xnor U3948 (N_3948,N_1558,N_1560);
or U3949 (N_3949,N_2166,N_143);
nor U3950 (N_3950,N_1904,N_829);
nand U3951 (N_3951,N_1662,N_943);
nand U3952 (N_3952,N_471,N_2936);
or U3953 (N_3953,N_191,N_1838);
or U3954 (N_3954,N_1695,N_2852);
and U3955 (N_3955,N_2722,N_306);
or U3956 (N_3956,N_1426,N_1268);
nand U3957 (N_3957,N_1765,N_2972);
or U3958 (N_3958,N_1049,N_2589);
nor U3959 (N_3959,N_1288,N_2429);
nor U3960 (N_3960,N_1994,N_1294);
and U3961 (N_3961,N_328,N_2350);
nor U3962 (N_3962,N_1511,N_1081);
and U3963 (N_3963,N_944,N_2230);
xnor U3964 (N_3964,N_2225,N_2058);
and U3965 (N_3965,N_557,N_673);
and U3966 (N_3966,N_2173,N_572);
or U3967 (N_3967,N_2144,N_759);
nor U3968 (N_3968,N_1191,N_2931);
nor U3969 (N_3969,N_870,N_606);
and U3970 (N_3970,N_1366,N_782);
nand U3971 (N_3971,N_403,N_1449);
xnor U3972 (N_3972,N_629,N_1710);
or U3973 (N_3973,N_465,N_1214);
and U3974 (N_3974,N_660,N_649);
nor U3975 (N_3975,N_445,N_2309);
nor U3976 (N_3976,N_300,N_2602);
nor U3977 (N_3977,N_2094,N_2011);
or U3978 (N_3978,N_1112,N_2169);
nand U3979 (N_3979,N_11,N_1609);
nand U3980 (N_3980,N_983,N_2691);
nand U3981 (N_3981,N_2262,N_483);
nor U3982 (N_3982,N_2700,N_1666);
and U3983 (N_3983,N_2401,N_2735);
nand U3984 (N_3984,N_1926,N_1293);
nand U3985 (N_3985,N_1985,N_1310);
xor U3986 (N_3986,N_1743,N_2643);
and U3987 (N_3987,N_2928,N_1071);
and U3988 (N_3988,N_2623,N_2188);
or U3989 (N_3989,N_676,N_1056);
nand U3990 (N_3990,N_592,N_2392);
nand U3991 (N_3991,N_2607,N_437);
nor U3992 (N_3992,N_96,N_1617);
nor U3993 (N_3993,N_2800,N_674);
nand U3994 (N_3994,N_309,N_1206);
nand U3995 (N_3995,N_278,N_2399);
xor U3996 (N_3996,N_34,N_1204);
nand U3997 (N_3997,N_745,N_2407);
nand U3998 (N_3998,N_1756,N_694);
nand U3999 (N_3999,N_2017,N_2897);
nand U4000 (N_4000,N_744,N_1991);
nor U4001 (N_4001,N_1636,N_2281);
and U4002 (N_4002,N_570,N_1718);
or U4003 (N_4003,N_1203,N_2052);
nor U4004 (N_4004,N_969,N_1724);
nand U4005 (N_4005,N_2873,N_1392);
or U4006 (N_4006,N_788,N_1048);
nor U4007 (N_4007,N_553,N_622);
and U4008 (N_4008,N_1472,N_702);
xnor U4009 (N_4009,N_341,N_1835);
nand U4010 (N_4010,N_1151,N_1241);
or U4011 (N_4011,N_1514,N_1674);
nor U4012 (N_4012,N_447,N_2141);
nand U4013 (N_4013,N_2316,N_2496);
or U4014 (N_4014,N_1828,N_1467);
nand U4015 (N_4015,N_74,N_972);
and U4016 (N_4016,N_1064,N_2600);
and U4017 (N_4017,N_123,N_2695);
xnor U4018 (N_4018,N_1778,N_597);
nand U4019 (N_4019,N_810,N_1379);
xnor U4020 (N_4020,N_1632,N_950);
or U4021 (N_4021,N_2991,N_2405);
nor U4022 (N_4022,N_2196,N_1611);
and U4023 (N_4023,N_1236,N_1888);
xor U4024 (N_4024,N_2120,N_2681);
or U4025 (N_4025,N_1757,N_2541);
and U4026 (N_4026,N_2258,N_2555);
or U4027 (N_4027,N_828,N_1272);
nor U4028 (N_4028,N_1590,N_1654);
and U4029 (N_4029,N_1736,N_1117);
or U4030 (N_4030,N_656,N_2956);
nand U4031 (N_4031,N_753,N_1639);
and U4032 (N_4032,N_350,N_2869);
xor U4033 (N_4033,N_54,N_977);
and U4034 (N_4034,N_1565,N_355);
xnor U4035 (N_4035,N_2285,N_2803);
and U4036 (N_4036,N_2548,N_1255);
or U4037 (N_4037,N_1474,N_254);
or U4038 (N_4038,N_1951,N_2612);
and U4039 (N_4039,N_1357,N_1670);
and U4040 (N_4040,N_1001,N_35);
xnor U4041 (N_4041,N_1382,N_2932);
xnor U4042 (N_4042,N_279,N_2300);
nand U4043 (N_4043,N_655,N_2112);
or U4044 (N_4044,N_2930,N_152);
nor U4045 (N_4045,N_2268,N_2690);
and U4046 (N_4046,N_940,N_1050);
and U4047 (N_4047,N_122,N_2420);
and U4048 (N_4048,N_771,N_2208);
nand U4049 (N_4049,N_1594,N_2224);
or U4050 (N_4050,N_888,N_2066);
nand U4051 (N_4051,N_701,N_647);
xor U4052 (N_4052,N_314,N_718);
or U4053 (N_4053,N_393,N_1029);
nor U4054 (N_4054,N_2554,N_175);
and U4055 (N_4055,N_1192,N_41);
and U4056 (N_4056,N_2397,N_1319);
and U4057 (N_4057,N_2192,N_20);
and U4058 (N_4058,N_97,N_1042);
nor U4059 (N_4059,N_1098,N_849);
nor U4060 (N_4060,N_71,N_1333);
or U4061 (N_4061,N_1369,N_36);
xor U4062 (N_4062,N_61,N_381);
xnor U4063 (N_4063,N_1194,N_1797);
nor U4064 (N_4064,N_1156,N_1429);
nand U4065 (N_4065,N_680,N_2445);
nand U4066 (N_4066,N_37,N_1658);
xor U4067 (N_4067,N_853,N_2113);
xnor U4068 (N_4068,N_578,N_2611);
or U4069 (N_4069,N_2637,N_2080);
and U4070 (N_4070,N_613,N_2132);
or U4071 (N_4071,N_2839,N_2117);
or U4072 (N_4072,N_1965,N_19);
xor U4073 (N_4073,N_768,N_2226);
and U4074 (N_4074,N_928,N_2618);
and U4075 (N_4075,N_2933,N_2037);
or U4076 (N_4076,N_783,N_1794);
xnor U4077 (N_4077,N_1286,N_1326);
or U4078 (N_4078,N_1659,N_2798);
or U4079 (N_4079,N_925,N_1415);
nand U4080 (N_4080,N_1999,N_620);
and U4081 (N_4081,N_1442,N_2016);
or U4082 (N_4082,N_1477,N_1768);
and U4083 (N_4083,N_2780,N_2747);
or U4084 (N_4084,N_1620,N_2093);
nand U4085 (N_4085,N_789,N_1783);
or U4086 (N_4086,N_433,N_1052);
and U4087 (N_4087,N_14,N_2484);
and U4088 (N_4088,N_2322,N_2473);
or U4089 (N_4089,N_1690,N_516);
and U4090 (N_4090,N_1487,N_2909);
nor U4091 (N_4091,N_321,N_1351);
nor U4092 (N_4092,N_1246,N_1051);
or U4093 (N_4093,N_2655,N_386);
or U4094 (N_4094,N_295,N_1731);
nand U4095 (N_4095,N_2978,N_1530);
and U4096 (N_4096,N_1854,N_405);
or U4097 (N_4097,N_1065,N_2040);
or U4098 (N_4098,N_2444,N_636);
xnor U4099 (N_4099,N_2500,N_2013);
nand U4100 (N_4100,N_407,N_1777);
and U4101 (N_4101,N_957,N_21);
xor U4102 (N_4102,N_167,N_415);
and U4103 (N_4103,N_993,N_1890);
xor U4104 (N_4104,N_1732,N_1421);
nor U4105 (N_4105,N_1190,N_885);
or U4106 (N_4106,N_2162,N_730);
or U4107 (N_4107,N_2929,N_1602);
or U4108 (N_4108,N_1614,N_1372);
and U4109 (N_4109,N_5,N_1184);
and U4110 (N_4110,N_2918,N_1176);
nand U4111 (N_4111,N_2727,N_1410);
or U4112 (N_4112,N_2726,N_1582);
nor U4113 (N_4113,N_2404,N_1175);
or U4114 (N_4114,N_1014,N_1987);
and U4115 (N_4115,N_2232,N_257);
or U4116 (N_4116,N_142,N_1682);
nand U4117 (N_4117,N_2250,N_10);
nor U4118 (N_4118,N_1528,N_932);
nand U4119 (N_4119,N_1745,N_1739);
nand U4120 (N_4120,N_2474,N_2832);
nand U4121 (N_4121,N_410,N_1957);
nand U4122 (N_4122,N_721,N_764);
xor U4123 (N_4123,N_1986,N_732);
and U4124 (N_4124,N_1578,N_1400);
nand U4125 (N_4125,N_1606,N_1262);
or U4126 (N_4126,N_286,N_2362);
xor U4127 (N_4127,N_986,N_1523);
nand U4128 (N_4128,N_352,N_808);
nand U4129 (N_4129,N_164,N_479);
and U4130 (N_4130,N_2119,N_2005);
or U4131 (N_4131,N_2719,N_1159);
or U4132 (N_4132,N_1387,N_2622);
or U4133 (N_4133,N_2264,N_1090);
nand U4134 (N_4134,N_2063,N_667);
xnor U4135 (N_4135,N_2388,N_1149);
nand U4136 (N_4136,N_558,N_2360);
and U4137 (N_4137,N_2176,N_1066);
and U4138 (N_4138,N_2290,N_2877);
nand U4139 (N_4139,N_478,N_2437);
nand U4140 (N_4140,N_243,N_436);
nor U4141 (N_4141,N_2494,N_2198);
and U4142 (N_4142,N_412,N_1811);
nor U4143 (N_4143,N_156,N_895);
nand U4144 (N_4144,N_1673,N_2529);
and U4145 (N_4145,N_272,N_1177);
and U4146 (N_4146,N_430,N_1848);
nor U4147 (N_4147,N_633,N_489);
nand U4148 (N_4148,N_956,N_2416);
nor U4149 (N_4149,N_2638,N_2505);
xnor U4150 (N_4150,N_2788,N_1877);
and U4151 (N_4151,N_2274,N_2485);
and U4152 (N_4152,N_1806,N_876);
or U4153 (N_4153,N_1751,N_2140);
or U4154 (N_4154,N_736,N_2064);
or U4155 (N_4155,N_450,N_361);
nor U4156 (N_4156,N_2378,N_1348);
or U4157 (N_4157,N_2403,N_832);
nand U4158 (N_4158,N_2767,N_1749);
and U4159 (N_4159,N_2653,N_120);
xor U4160 (N_4160,N_517,N_2335);
xor U4161 (N_4161,N_2684,N_2293);
xnor U4162 (N_4162,N_2492,N_1927);
nor U4163 (N_4163,N_941,N_1419);
nand U4164 (N_4164,N_2077,N_891);
and U4165 (N_4165,N_481,N_1845);
nand U4166 (N_4166,N_1148,N_1489);
or U4167 (N_4167,N_1717,N_1956);
nor U4168 (N_4168,N_1973,N_2524);
or U4169 (N_4169,N_2222,N_1998);
or U4170 (N_4170,N_1688,N_1178);
nand U4171 (N_4171,N_426,N_2042);
nand U4172 (N_4172,N_989,N_2317);
or U4173 (N_4173,N_2765,N_1571);
and U4174 (N_4174,N_840,N_734);
or U4175 (N_4175,N_760,N_1290);
xor U4176 (N_4176,N_1105,N_285);
nand U4177 (N_4177,N_1230,N_1057);
nand U4178 (N_4178,N_2440,N_716);
and U4179 (N_4179,N_1485,N_273);
and U4180 (N_4180,N_1079,N_2346);
and U4181 (N_4181,N_1059,N_966);
and U4182 (N_4182,N_2195,N_746);
nand U4183 (N_4183,N_543,N_1452);
nand U4184 (N_4184,N_1791,N_113);
xnor U4185 (N_4185,N_1708,N_878);
nand U4186 (N_4186,N_373,N_90);
and U4187 (N_4187,N_1334,N_168);
and U4188 (N_4188,N_1123,N_2488);
or U4189 (N_4189,N_251,N_83);
or U4190 (N_4190,N_170,N_2915);
and U4191 (N_4191,N_33,N_1915);
or U4192 (N_4192,N_354,N_1563);
or U4193 (N_4193,N_2428,N_2328);
or U4194 (N_4194,N_1127,N_1201);
or U4195 (N_4195,N_1711,N_2393);
or U4196 (N_4196,N_53,N_1360);
or U4197 (N_4197,N_2495,N_2481);
nor U4198 (N_4198,N_513,N_56);
nor U4199 (N_4199,N_1070,N_1267);
and U4200 (N_4200,N_803,N_755);
and U4201 (N_4201,N_807,N_804);
nand U4202 (N_4202,N_1679,N_1719);
xnor U4203 (N_4203,N_1740,N_1358);
nor U4204 (N_4204,N_1886,N_485);
nor U4205 (N_4205,N_2866,N_2457);
and U4206 (N_4206,N_2126,N_484);
and U4207 (N_4207,N_743,N_1832);
and U4208 (N_4208,N_1263,N_2882);
nor U4209 (N_4209,N_2573,N_926);
or U4210 (N_4210,N_1618,N_263);
nor U4211 (N_4211,N_401,N_2671);
nand U4212 (N_4212,N_1713,N_1026);
nand U4213 (N_4213,N_1108,N_2179);
and U4214 (N_4214,N_2108,N_2221);
or U4215 (N_4215,N_2156,N_1480);
and U4216 (N_4216,N_2970,N_1153);
nor U4217 (N_4217,N_1428,N_980);
or U4218 (N_4218,N_148,N_23);
and U4219 (N_4219,N_790,N_1329);
or U4220 (N_4220,N_1819,N_1591);
nor U4221 (N_4221,N_2313,N_1142);
nand U4222 (N_4222,N_978,N_2676);
nor U4223 (N_4223,N_1012,N_563);
or U4224 (N_4224,N_1512,N_652);
nand U4225 (N_4225,N_2783,N_190);
nand U4226 (N_4226,N_2601,N_1354);
or U4227 (N_4227,N_946,N_1295);
and U4228 (N_4228,N_1205,N_610);
xor U4229 (N_4229,N_2531,N_2903);
or U4230 (N_4230,N_2353,N_2694);
or U4231 (N_4231,N_586,N_2400);
nand U4232 (N_4232,N_509,N_2699);
nand U4233 (N_4233,N_1903,N_1697);
and U4234 (N_4234,N_551,N_246);
or U4235 (N_4235,N_2905,N_137);
xnor U4236 (N_4236,N_1921,N_65);
and U4237 (N_4237,N_959,N_1492);
nand U4238 (N_4238,N_752,N_1792);
nand U4239 (N_4239,N_2857,N_2432);
xor U4240 (N_4240,N_2995,N_1761);
nand U4241 (N_4241,N_1284,N_1651);
or U4242 (N_4242,N_315,N_416);
xnor U4243 (N_4243,N_1942,N_0);
nor U4244 (N_4244,N_934,N_2672);
or U4245 (N_4245,N_2539,N_2155);
nand U4246 (N_4246,N_2717,N_515);
and U4247 (N_4247,N_2099,N_907);
nor U4248 (N_4248,N_1259,N_1531);
and U4249 (N_4249,N_658,N_638);
nor U4250 (N_4250,N_2510,N_994);
nor U4251 (N_4251,N_112,N_1946);
nand U4252 (N_4252,N_707,N_2178);
nor U4253 (N_4253,N_1219,N_890);
nor U4254 (N_4254,N_780,N_2344);
nor U4255 (N_4255,N_438,N_1593);
nor U4256 (N_4256,N_1536,N_1499);
or U4257 (N_4257,N_2513,N_209);
nor U4258 (N_4258,N_1652,N_1353);
xnor U4259 (N_4259,N_2455,N_244);
or U4260 (N_4260,N_2606,N_1041);
or U4261 (N_4261,N_87,N_86);
or U4262 (N_4262,N_1188,N_1130);
or U4263 (N_4263,N_546,N_319);
nor U4264 (N_4264,N_2957,N_2431);
and U4265 (N_4265,N_385,N_2549);
nand U4266 (N_4266,N_380,N_2184);
nor U4267 (N_4267,N_776,N_192);
nor U4268 (N_4268,N_1976,N_2806);
or U4269 (N_4269,N_151,N_219);
or U4270 (N_4270,N_2769,N_88);
or U4271 (N_4271,N_1137,N_2969);
nand U4272 (N_4272,N_873,N_2476);
or U4273 (N_4273,N_2490,N_491);
or U4274 (N_4274,N_1758,N_1881);
and U4275 (N_4275,N_2955,N_2055);
nand U4276 (N_4276,N_2583,N_145);
nand U4277 (N_4277,N_617,N_2543);
nand U4278 (N_4278,N_773,N_2748);
or U4279 (N_4279,N_1339,N_2741);
nand U4280 (N_4280,N_830,N_2988);
nor U4281 (N_4281,N_719,N_637);
or U4282 (N_4282,N_619,N_2253);
nor U4283 (N_4283,N_1099,N_567);
and U4284 (N_4284,N_111,N_2971);
or U4285 (N_4285,N_1396,N_1076);
nor U4286 (N_4286,N_2368,N_2421);
and U4287 (N_4287,N_2471,N_2375);
nand U4288 (N_4288,N_2364,N_371);
nand U4289 (N_4289,N_435,N_1733);
nand U4290 (N_4290,N_1170,N_462);
nand U4291 (N_4291,N_208,N_2483);
and U4292 (N_4292,N_2308,N_157);
nand U4293 (N_4293,N_1312,N_2952);
and U4294 (N_4294,N_299,N_1091);
xnor U4295 (N_4295,N_2953,N_473);
and U4296 (N_4296,N_1712,N_2597);
and U4297 (N_4297,N_2715,N_2714);
nand U4298 (N_4298,N_1748,N_1147);
nand U4299 (N_4299,N_1008,N_2850);
nor U4300 (N_4300,N_2639,N_2337);
or U4301 (N_4301,N_375,N_2266);
or U4302 (N_4302,N_2430,N_2678);
nor U4303 (N_4303,N_999,N_1586);
or U4304 (N_4304,N_492,N_2917);
or U4305 (N_4305,N_1459,N_985);
or U4306 (N_4306,N_691,N_520);
or U4307 (N_4307,N_1725,N_955);
nor U4308 (N_4308,N_379,N_1102);
xor U4309 (N_4309,N_2070,N_2303);
and U4310 (N_4310,N_2090,N_1067);
nand U4311 (N_4311,N_2893,N_1935);
nor U4312 (N_4312,N_1932,N_2381);
nor U4313 (N_4313,N_2559,N_1300);
nand U4314 (N_4314,N_672,N_1475);
or U4315 (N_4315,N_218,N_391);
and U4316 (N_4316,N_2723,N_1322);
or U4317 (N_4317,N_2987,N_1224);
and U4318 (N_4318,N_1752,N_951);
nand U4319 (N_4319,N_2566,N_988);
nor U4320 (N_4320,N_469,N_685);
and U4321 (N_4321,N_1164,N_1498);
or U4322 (N_4322,N_1786,N_2377);
nand U4323 (N_4323,N_1874,N_2585);
nand U4324 (N_4324,N_2069,N_2133);
nand U4325 (N_4325,N_1795,N_2565);
nand U4326 (N_4326,N_2617,N_82);
or U4327 (N_4327,N_2414,N_2763);
or U4328 (N_4328,N_2111,N_641);
nor U4329 (N_4329,N_1016,N_2960);
nor U4330 (N_4330,N_2150,N_1034);
nand U4331 (N_4331,N_402,N_1722);
or U4332 (N_4332,N_1664,N_2922);
and U4333 (N_4333,N_205,N_2772);
nand U4334 (N_4334,N_1509,N_1025);
and U4335 (N_4335,N_2615,N_334);
nand U4336 (N_4336,N_1974,N_1336);
xor U4337 (N_4337,N_1557,N_2294);
xnor U4338 (N_4338,N_397,N_1599);
or U4339 (N_4339,N_252,N_2243);
xnor U4340 (N_4340,N_451,N_1240);
nor U4341 (N_4341,N_632,N_2227);
nor U4342 (N_4342,N_2867,N_1174);
xnor U4343 (N_4343,N_24,N_1508);
nor U4344 (N_4344,N_2036,N_1020);
or U4345 (N_4345,N_1917,N_1721);
nor U4346 (N_4346,N_1403,N_1301);
nor U4347 (N_4347,N_820,N_448);
and U4348 (N_4348,N_698,N_1234);
nor U4349 (N_4349,N_1916,N_1239);
or U4350 (N_4350,N_1520,N_1252);
or U4351 (N_4351,N_2007,N_176);
or U4352 (N_4352,N_1621,N_2536);
nor U4353 (N_4353,N_2158,N_2577);
nor U4354 (N_4354,N_423,N_834);
or U4355 (N_4355,N_1394,N_2115);
nor U4356 (N_4356,N_1592,N_186);
or U4357 (N_4357,N_778,N_15);
nand U4358 (N_4358,N_268,N_836);
nand U4359 (N_4359,N_2887,N_1424);
xor U4360 (N_4360,N_2519,N_1988);
nor U4361 (N_4361,N_400,N_2060);
and U4362 (N_4362,N_1466,N_774);
nor U4363 (N_4363,N_2272,N_1847);
or U4364 (N_4364,N_118,N_395);
and U4365 (N_4365,N_1506,N_645);
or U4366 (N_4366,N_1569,N_1914);
nor U4367 (N_4367,N_58,N_2246);
and U4368 (N_4368,N_1482,N_2092);
nor U4369 (N_4369,N_735,N_544);
and U4370 (N_4370,N_42,N_47);
or U4371 (N_4371,N_2564,N_1978);
nor U4372 (N_4372,N_313,N_195);
and U4373 (N_4373,N_1539,N_598);
and U4374 (N_4374,N_1622,N_1584);
or U4375 (N_4375,N_2319,N_2352);
and U4376 (N_4376,N_2276,N_824);
nor U4377 (N_4377,N_1504,N_2802);
nand U4378 (N_4378,N_210,N_2449);
xor U4379 (N_4379,N_1889,N_501);
nand U4380 (N_4380,N_646,N_1135);
nand U4381 (N_4381,N_1276,N_2563);
nor U4382 (N_4382,N_1555,N_2683);
and U4383 (N_4383,N_468,N_463);
and U4384 (N_4384,N_2815,N_2355);
nand U4385 (N_4385,N_2697,N_1892);
xor U4386 (N_4386,N_2605,N_2125);
nor U4387 (N_4387,N_2626,N_2945);
nand U4388 (N_4388,N_1168,N_574);
or U4389 (N_4389,N_305,N_1352);
nand U4390 (N_4390,N_2349,N_815);
and U4391 (N_4391,N_839,N_2778);
or U4392 (N_4392,N_1940,N_1173);
or U4393 (N_4393,N_434,N_1046);
xor U4394 (N_4394,N_1037,N_2533);
nor U4395 (N_4395,N_2336,N_2439);
or U4396 (N_4396,N_264,N_1491);
xnor U4397 (N_4397,N_1665,N_1069);
nand U4398 (N_4398,N_1497,N_1767);
nor U4399 (N_4399,N_2161,N_1857);
nand U4400 (N_4400,N_323,N_1616);
or U4401 (N_4401,N_247,N_2046);
nand U4402 (N_4402,N_154,N_2817);
or U4403 (N_4403,N_1095,N_2361);
nor U4404 (N_4404,N_1981,N_2433);
nor U4405 (N_4405,N_70,N_1238);
or U4406 (N_4406,N_311,N_237);
or U4407 (N_4407,N_692,N_1335);
or U4408 (N_4408,N_1949,N_461);
and U4409 (N_4409,N_835,N_1909);
nand U4410 (N_4410,N_1193,N_2291);
xnor U4411 (N_4411,N_2183,N_1996);
and U4412 (N_4412,N_1368,N_1473);
nor U4413 (N_4413,N_1887,N_1687);
or U4414 (N_4414,N_2809,N_1645);
and U4415 (N_4415,N_1383,N_881);
nor U4416 (N_4416,N_1324,N_294);
or U4417 (N_4417,N_918,N_62);
nor U4418 (N_4418,N_495,N_29);
xnor U4419 (N_4419,N_2107,N_2304);
nor U4420 (N_4420,N_302,N_2878);
or U4421 (N_4421,N_882,N_2165);
nand U4422 (N_4422,N_2659,N_1375);
and U4423 (N_4423,N_144,N_2020);
nand U4424 (N_4424,N_1950,N_899);
or U4425 (N_4425,N_1642,N_2045);
xor U4426 (N_4426,N_2624,N_2977);
and U4427 (N_4427,N_1343,N_968);
nor U4428 (N_4428,N_1185,N_72);
and U4429 (N_4429,N_2512,N_1281);
nand U4430 (N_4430,N_390,N_128);
xor U4431 (N_4431,N_1121,N_758);
and U4432 (N_4432,N_1433,N_2538);
and U4433 (N_4433,N_149,N_2656);
nand U4434 (N_4434,N_2528,N_1668);
nor U4435 (N_4435,N_2448,N_1494);
nand U4436 (N_4436,N_2279,N_2244);
nor U4437 (N_4437,N_2018,N_441);
nor U4438 (N_4438,N_819,N_2273);
xnor U4439 (N_4439,N_938,N_2552);
or U4440 (N_4440,N_863,N_384);
and U4441 (N_4441,N_2949,N_749);
or U4442 (N_4442,N_2689,N_357);
nor U4443 (N_4443,N_1787,N_1859);
or U4444 (N_4444,N_754,N_2338);
nand U4445 (N_4445,N_1948,N_937);
nand U4446 (N_4446,N_2507,N_301);
nand U4447 (N_4447,N_1296,N_1138);
nand U4448 (N_4448,N_1629,N_1478);
or U4449 (N_4449,N_861,N_1496);
xnor U4450 (N_4450,N_1534,N_1257);
xor U4451 (N_4451,N_2958,N_1119);
or U4452 (N_4452,N_542,N_847);
xor U4453 (N_4453,N_404,N_2544);
or U4454 (N_4454,N_99,N_1781);
xnor U4455 (N_4455,N_1595,N_2263);
nor U4456 (N_4456,N_1773,N_459);
and U4457 (N_4457,N_2456,N_2736);
or U4458 (N_4458,N_779,N_1405);
nand U4459 (N_4459,N_1370,N_1543);
and U4460 (N_4460,N_2938,N_2366);
nor U4461 (N_4461,N_1549,N_1113);
nand U4462 (N_4462,N_1378,N_2731);
or U4463 (N_4463,N_9,N_1771);
xnor U4464 (N_4464,N_1440,N_614);
and U4465 (N_4465,N_267,N_1345);
or U4466 (N_4466,N_2670,N_2582);
nand U4467 (N_4467,N_2663,N_2985);
xor U4468 (N_4468,N_2228,N_1870);
or U4469 (N_4469,N_865,N_1727);
xnor U4470 (N_4470,N_1152,N_1250);
nand U4471 (N_4471,N_1427,N_358);
and U4472 (N_4472,N_432,N_1210);
or U4473 (N_4473,N_1253,N_101);
nor U4474 (N_4474,N_330,N_109);
xor U4475 (N_4475,N_723,N_1689);
nor U4476 (N_4476,N_290,N_913);
or U4477 (N_4477,N_2760,N_360);
or U4478 (N_4478,N_1233,N_2216);
nor U4479 (N_4479,N_970,N_2463);
nor U4480 (N_4480,N_1165,N_2827);
and U4481 (N_4481,N_378,N_2441);
or U4482 (N_4482,N_1242,N_1706);
or U4483 (N_4483,N_1308,N_2964);
nor U4484 (N_4484,N_1423,N_887);
and U4485 (N_4485,N_1321,N_2323);
and U4486 (N_4486,N_1844,N_703);
or U4487 (N_4487,N_1968,N_547);
nor U4488 (N_4488,N_2426,N_1677);
xor U4489 (N_4489,N_2207,N_2992);
and U4490 (N_4490,N_2109,N_1031);
or U4491 (N_4491,N_275,N_1587);
nor U4492 (N_4492,N_2965,N_2172);
nand U4493 (N_4493,N_2688,N_2665);
nand U4494 (N_4494,N_857,N_1118);
nand U4495 (N_4495,N_2746,N_324);
nor U4496 (N_4496,N_57,N_1846);
nor U4497 (N_4497,N_1538,N_345);
and U4498 (N_4498,N_1977,N_1055);
or U4499 (N_4499,N_104,N_1092);
or U4500 (N_4500,N_2304,N_1922);
nor U4501 (N_4501,N_1302,N_1804);
nor U4502 (N_4502,N_2155,N_2314);
nand U4503 (N_4503,N_1970,N_34);
nand U4504 (N_4504,N_2363,N_1235);
nor U4505 (N_4505,N_526,N_568);
or U4506 (N_4506,N_1672,N_956);
nand U4507 (N_4507,N_1182,N_611);
or U4508 (N_4508,N_1533,N_2526);
nand U4509 (N_4509,N_1961,N_1700);
xnor U4510 (N_4510,N_2908,N_771);
nor U4511 (N_4511,N_766,N_862);
or U4512 (N_4512,N_843,N_995);
or U4513 (N_4513,N_817,N_812);
and U4514 (N_4514,N_1359,N_318);
xor U4515 (N_4515,N_1182,N_1530);
nor U4516 (N_4516,N_433,N_1768);
nand U4517 (N_4517,N_211,N_2861);
nor U4518 (N_4518,N_1281,N_2804);
xor U4519 (N_4519,N_2819,N_845);
nand U4520 (N_4520,N_2776,N_2200);
nand U4521 (N_4521,N_1544,N_1350);
nand U4522 (N_4522,N_2546,N_2962);
nor U4523 (N_4523,N_69,N_2150);
and U4524 (N_4524,N_37,N_1888);
xor U4525 (N_4525,N_2528,N_61);
nand U4526 (N_4526,N_1713,N_2780);
nand U4527 (N_4527,N_2377,N_315);
nor U4528 (N_4528,N_544,N_2058);
nand U4529 (N_4529,N_1885,N_84);
and U4530 (N_4530,N_1203,N_2929);
or U4531 (N_4531,N_30,N_2663);
nor U4532 (N_4532,N_328,N_190);
nor U4533 (N_4533,N_2795,N_1096);
or U4534 (N_4534,N_1098,N_1781);
nand U4535 (N_4535,N_2588,N_1552);
xor U4536 (N_4536,N_1879,N_1142);
and U4537 (N_4537,N_2575,N_670);
nor U4538 (N_4538,N_2333,N_2551);
nand U4539 (N_4539,N_2833,N_2097);
nor U4540 (N_4540,N_1329,N_2505);
and U4541 (N_4541,N_991,N_1536);
or U4542 (N_4542,N_757,N_1818);
nand U4543 (N_4543,N_899,N_378);
nor U4544 (N_4544,N_2284,N_1635);
or U4545 (N_4545,N_1354,N_123);
xnor U4546 (N_4546,N_2514,N_2351);
nor U4547 (N_4547,N_2356,N_2045);
nand U4548 (N_4548,N_2899,N_2448);
and U4549 (N_4549,N_641,N_1772);
nand U4550 (N_4550,N_2882,N_2648);
nand U4551 (N_4551,N_2033,N_2053);
nand U4552 (N_4552,N_2513,N_1441);
nor U4553 (N_4553,N_685,N_93);
nor U4554 (N_4554,N_1902,N_287);
xor U4555 (N_4555,N_897,N_1802);
nor U4556 (N_4556,N_2427,N_1222);
nor U4557 (N_4557,N_2544,N_1522);
nor U4558 (N_4558,N_783,N_1239);
xor U4559 (N_4559,N_2933,N_1942);
nand U4560 (N_4560,N_1298,N_2368);
nand U4561 (N_4561,N_1854,N_2437);
nand U4562 (N_4562,N_512,N_1792);
and U4563 (N_4563,N_2157,N_1348);
nor U4564 (N_4564,N_2873,N_832);
or U4565 (N_4565,N_2336,N_2976);
nor U4566 (N_4566,N_648,N_2705);
nor U4567 (N_4567,N_522,N_1369);
nor U4568 (N_4568,N_2369,N_2889);
or U4569 (N_4569,N_335,N_1151);
and U4570 (N_4570,N_1906,N_487);
nand U4571 (N_4571,N_1829,N_2149);
nor U4572 (N_4572,N_1942,N_1810);
nor U4573 (N_4573,N_1236,N_1728);
nor U4574 (N_4574,N_1271,N_2807);
nand U4575 (N_4575,N_2483,N_1536);
nand U4576 (N_4576,N_2475,N_2301);
xor U4577 (N_4577,N_2197,N_2426);
nor U4578 (N_4578,N_2206,N_349);
or U4579 (N_4579,N_850,N_1965);
nor U4580 (N_4580,N_1924,N_2110);
and U4581 (N_4581,N_1840,N_2177);
and U4582 (N_4582,N_1474,N_408);
nand U4583 (N_4583,N_2034,N_2352);
nand U4584 (N_4584,N_1392,N_2145);
xor U4585 (N_4585,N_2892,N_1164);
and U4586 (N_4586,N_82,N_2787);
or U4587 (N_4587,N_920,N_1573);
nor U4588 (N_4588,N_53,N_730);
nand U4589 (N_4589,N_2920,N_572);
or U4590 (N_4590,N_1971,N_2456);
or U4591 (N_4591,N_195,N_2667);
and U4592 (N_4592,N_442,N_2386);
nor U4593 (N_4593,N_1362,N_2376);
nor U4594 (N_4594,N_2079,N_1700);
nand U4595 (N_4595,N_2495,N_1983);
or U4596 (N_4596,N_2217,N_1828);
nor U4597 (N_4597,N_1838,N_873);
xor U4598 (N_4598,N_2776,N_2846);
nand U4599 (N_4599,N_193,N_2967);
or U4600 (N_4600,N_145,N_1571);
nor U4601 (N_4601,N_1676,N_655);
and U4602 (N_4602,N_448,N_729);
and U4603 (N_4603,N_11,N_898);
nor U4604 (N_4604,N_1275,N_2095);
and U4605 (N_4605,N_527,N_2472);
xor U4606 (N_4606,N_2945,N_2874);
or U4607 (N_4607,N_331,N_1720);
and U4608 (N_4608,N_1116,N_1437);
or U4609 (N_4609,N_1470,N_311);
or U4610 (N_4610,N_2107,N_2046);
and U4611 (N_4611,N_2572,N_1210);
or U4612 (N_4612,N_2223,N_248);
or U4613 (N_4613,N_419,N_306);
nand U4614 (N_4614,N_1532,N_2024);
and U4615 (N_4615,N_896,N_994);
xnor U4616 (N_4616,N_1558,N_277);
and U4617 (N_4617,N_1549,N_618);
or U4618 (N_4618,N_478,N_355);
and U4619 (N_4619,N_1440,N_2143);
nand U4620 (N_4620,N_1126,N_2958);
nor U4621 (N_4621,N_640,N_1466);
nand U4622 (N_4622,N_496,N_2861);
or U4623 (N_4623,N_1665,N_1226);
nor U4624 (N_4624,N_1521,N_2345);
nand U4625 (N_4625,N_603,N_438);
or U4626 (N_4626,N_1449,N_1885);
and U4627 (N_4627,N_2279,N_1467);
nand U4628 (N_4628,N_1916,N_2086);
and U4629 (N_4629,N_2510,N_1450);
nand U4630 (N_4630,N_763,N_637);
or U4631 (N_4631,N_1824,N_2663);
and U4632 (N_4632,N_485,N_810);
nor U4633 (N_4633,N_2986,N_523);
or U4634 (N_4634,N_236,N_170);
or U4635 (N_4635,N_1072,N_513);
and U4636 (N_4636,N_2800,N_946);
nor U4637 (N_4637,N_1554,N_1386);
or U4638 (N_4638,N_1193,N_2444);
nor U4639 (N_4639,N_1066,N_2132);
nand U4640 (N_4640,N_170,N_293);
or U4641 (N_4641,N_1739,N_2989);
xnor U4642 (N_4642,N_2494,N_258);
nand U4643 (N_4643,N_1503,N_2179);
and U4644 (N_4644,N_2379,N_262);
nor U4645 (N_4645,N_302,N_1351);
or U4646 (N_4646,N_2156,N_1607);
nor U4647 (N_4647,N_2280,N_886);
nor U4648 (N_4648,N_2008,N_2584);
and U4649 (N_4649,N_912,N_2638);
and U4650 (N_4650,N_2654,N_2375);
or U4651 (N_4651,N_118,N_1508);
nand U4652 (N_4652,N_1954,N_1381);
nand U4653 (N_4653,N_2033,N_268);
and U4654 (N_4654,N_630,N_1592);
nand U4655 (N_4655,N_448,N_621);
nor U4656 (N_4656,N_402,N_694);
nand U4657 (N_4657,N_888,N_1667);
or U4658 (N_4658,N_738,N_2274);
nand U4659 (N_4659,N_763,N_759);
nor U4660 (N_4660,N_2487,N_884);
nor U4661 (N_4661,N_927,N_2753);
and U4662 (N_4662,N_139,N_45);
nand U4663 (N_4663,N_2623,N_1879);
and U4664 (N_4664,N_2933,N_175);
and U4665 (N_4665,N_2392,N_1806);
nor U4666 (N_4666,N_1258,N_487);
and U4667 (N_4667,N_2735,N_2903);
xnor U4668 (N_4668,N_1985,N_2725);
or U4669 (N_4669,N_950,N_2593);
and U4670 (N_4670,N_2940,N_1712);
nand U4671 (N_4671,N_586,N_1270);
nor U4672 (N_4672,N_707,N_1917);
and U4673 (N_4673,N_1216,N_2703);
or U4674 (N_4674,N_76,N_568);
nand U4675 (N_4675,N_2954,N_1081);
and U4676 (N_4676,N_326,N_2741);
nand U4677 (N_4677,N_2371,N_1185);
nand U4678 (N_4678,N_2946,N_1946);
xnor U4679 (N_4679,N_2921,N_1846);
and U4680 (N_4680,N_658,N_1171);
xor U4681 (N_4681,N_2209,N_1253);
nor U4682 (N_4682,N_1768,N_2094);
nand U4683 (N_4683,N_748,N_622);
and U4684 (N_4684,N_1709,N_2111);
nor U4685 (N_4685,N_878,N_1079);
or U4686 (N_4686,N_2589,N_1248);
nand U4687 (N_4687,N_856,N_1619);
nand U4688 (N_4688,N_1869,N_268);
nor U4689 (N_4689,N_25,N_2673);
and U4690 (N_4690,N_2726,N_2953);
nor U4691 (N_4691,N_818,N_2004);
nand U4692 (N_4692,N_639,N_2631);
or U4693 (N_4693,N_2293,N_1915);
and U4694 (N_4694,N_462,N_1825);
xor U4695 (N_4695,N_960,N_1343);
nor U4696 (N_4696,N_150,N_1663);
nand U4697 (N_4697,N_2651,N_575);
nand U4698 (N_4698,N_19,N_550);
and U4699 (N_4699,N_2421,N_1683);
nand U4700 (N_4700,N_1454,N_2916);
nand U4701 (N_4701,N_229,N_461);
and U4702 (N_4702,N_506,N_2388);
or U4703 (N_4703,N_2030,N_2045);
or U4704 (N_4704,N_1070,N_1395);
nor U4705 (N_4705,N_1575,N_1131);
or U4706 (N_4706,N_2568,N_790);
xor U4707 (N_4707,N_694,N_2653);
and U4708 (N_4708,N_1576,N_2546);
nor U4709 (N_4709,N_1933,N_1769);
and U4710 (N_4710,N_1203,N_74);
and U4711 (N_4711,N_2903,N_893);
and U4712 (N_4712,N_2801,N_2526);
nand U4713 (N_4713,N_2695,N_938);
or U4714 (N_4714,N_384,N_2630);
nor U4715 (N_4715,N_1562,N_1522);
or U4716 (N_4716,N_947,N_401);
or U4717 (N_4717,N_2257,N_2520);
xor U4718 (N_4718,N_426,N_523);
nand U4719 (N_4719,N_305,N_2068);
nand U4720 (N_4720,N_1666,N_1681);
and U4721 (N_4721,N_462,N_756);
or U4722 (N_4722,N_1852,N_1969);
nand U4723 (N_4723,N_794,N_400);
xor U4724 (N_4724,N_757,N_2382);
nand U4725 (N_4725,N_2361,N_2880);
nor U4726 (N_4726,N_2965,N_1266);
or U4727 (N_4727,N_2756,N_1891);
nor U4728 (N_4728,N_229,N_2231);
and U4729 (N_4729,N_457,N_402);
or U4730 (N_4730,N_642,N_1706);
nor U4731 (N_4731,N_2741,N_2638);
or U4732 (N_4732,N_317,N_2348);
and U4733 (N_4733,N_1701,N_2230);
or U4734 (N_4734,N_1782,N_2340);
or U4735 (N_4735,N_362,N_1417);
or U4736 (N_4736,N_1892,N_442);
and U4737 (N_4737,N_1394,N_1282);
or U4738 (N_4738,N_2198,N_158);
or U4739 (N_4739,N_2623,N_2847);
nand U4740 (N_4740,N_1054,N_1224);
nand U4741 (N_4741,N_783,N_2408);
nor U4742 (N_4742,N_732,N_1033);
or U4743 (N_4743,N_545,N_1984);
nand U4744 (N_4744,N_472,N_2989);
nand U4745 (N_4745,N_238,N_962);
and U4746 (N_4746,N_1696,N_1686);
or U4747 (N_4747,N_1542,N_2877);
nand U4748 (N_4748,N_979,N_601);
and U4749 (N_4749,N_2603,N_955);
and U4750 (N_4750,N_2571,N_853);
and U4751 (N_4751,N_1778,N_284);
xor U4752 (N_4752,N_1746,N_946);
nor U4753 (N_4753,N_2703,N_1916);
nand U4754 (N_4754,N_2409,N_1014);
nor U4755 (N_4755,N_2650,N_2047);
nand U4756 (N_4756,N_2436,N_1761);
nor U4757 (N_4757,N_24,N_573);
nor U4758 (N_4758,N_437,N_2672);
nand U4759 (N_4759,N_1213,N_1408);
xnor U4760 (N_4760,N_2394,N_58);
nor U4761 (N_4761,N_2595,N_1299);
or U4762 (N_4762,N_388,N_2357);
or U4763 (N_4763,N_2173,N_351);
nand U4764 (N_4764,N_1632,N_886);
or U4765 (N_4765,N_1712,N_1511);
nor U4766 (N_4766,N_297,N_2494);
nor U4767 (N_4767,N_699,N_2785);
xnor U4768 (N_4768,N_2927,N_1452);
xnor U4769 (N_4769,N_44,N_353);
xnor U4770 (N_4770,N_437,N_2271);
or U4771 (N_4771,N_829,N_579);
nor U4772 (N_4772,N_1489,N_1716);
and U4773 (N_4773,N_470,N_739);
or U4774 (N_4774,N_888,N_2334);
and U4775 (N_4775,N_146,N_2451);
nor U4776 (N_4776,N_2781,N_142);
or U4777 (N_4777,N_2103,N_1139);
or U4778 (N_4778,N_2954,N_2803);
xor U4779 (N_4779,N_945,N_1915);
or U4780 (N_4780,N_2177,N_841);
nand U4781 (N_4781,N_2079,N_623);
or U4782 (N_4782,N_27,N_61);
or U4783 (N_4783,N_293,N_1040);
xor U4784 (N_4784,N_705,N_2001);
xor U4785 (N_4785,N_2599,N_192);
nand U4786 (N_4786,N_390,N_2551);
nand U4787 (N_4787,N_1063,N_945);
xnor U4788 (N_4788,N_1999,N_373);
or U4789 (N_4789,N_2342,N_1347);
nand U4790 (N_4790,N_474,N_1644);
and U4791 (N_4791,N_2537,N_2271);
and U4792 (N_4792,N_1041,N_84);
nand U4793 (N_4793,N_1037,N_370);
or U4794 (N_4794,N_2590,N_2265);
nand U4795 (N_4795,N_2315,N_122);
nor U4796 (N_4796,N_2170,N_2945);
and U4797 (N_4797,N_593,N_1070);
nor U4798 (N_4798,N_546,N_1062);
and U4799 (N_4799,N_1087,N_1834);
or U4800 (N_4800,N_1504,N_124);
nor U4801 (N_4801,N_94,N_582);
xor U4802 (N_4802,N_1045,N_261);
nor U4803 (N_4803,N_2553,N_266);
and U4804 (N_4804,N_2017,N_1819);
and U4805 (N_4805,N_2058,N_1030);
nand U4806 (N_4806,N_6,N_864);
xor U4807 (N_4807,N_2956,N_1523);
or U4808 (N_4808,N_785,N_2609);
nor U4809 (N_4809,N_1797,N_1585);
and U4810 (N_4810,N_2648,N_2763);
nor U4811 (N_4811,N_1701,N_2607);
nor U4812 (N_4812,N_391,N_553);
nor U4813 (N_4813,N_2234,N_1505);
and U4814 (N_4814,N_2563,N_2657);
or U4815 (N_4815,N_2871,N_1939);
nand U4816 (N_4816,N_758,N_487);
or U4817 (N_4817,N_1115,N_2271);
or U4818 (N_4818,N_2761,N_2528);
or U4819 (N_4819,N_336,N_2857);
or U4820 (N_4820,N_1696,N_2679);
or U4821 (N_4821,N_1237,N_2944);
and U4822 (N_4822,N_281,N_2307);
nand U4823 (N_4823,N_2622,N_873);
and U4824 (N_4824,N_310,N_729);
or U4825 (N_4825,N_1721,N_2561);
xor U4826 (N_4826,N_2803,N_573);
nand U4827 (N_4827,N_89,N_1354);
nand U4828 (N_4828,N_1304,N_1360);
or U4829 (N_4829,N_1620,N_2174);
and U4830 (N_4830,N_1157,N_728);
nor U4831 (N_4831,N_1132,N_1511);
or U4832 (N_4832,N_1565,N_2277);
xor U4833 (N_4833,N_128,N_1854);
and U4834 (N_4834,N_1451,N_207);
nand U4835 (N_4835,N_778,N_1932);
nor U4836 (N_4836,N_589,N_1359);
nand U4837 (N_4837,N_795,N_583);
and U4838 (N_4838,N_812,N_2755);
and U4839 (N_4839,N_1774,N_242);
nor U4840 (N_4840,N_1710,N_1558);
or U4841 (N_4841,N_2936,N_2035);
nand U4842 (N_4842,N_2172,N_244);
or U4843 (N_4843,N_216,N_527);
and U4844 (N_4844,N_212,N_2467);
and U4845 (N_4845,N_2293,N_2205);
and U4846 (N_4846,N_1523,N_2380);
xnor U4847 (N_4847,N_2498,N_981);
and U4848 (N_4848,N_2950,N_1303);
and U4849 (N_4849,N_1786,N_245);
nand U4850 (N_4850,N_1759,N_327);
xnor U4851 (N_4851,N_1131,N_2886);
nand U4852 (N_4852,N_945,N_1983);
nand U4853 (N_4853,N_259,N_2155);
and U4854 (N_4854,N_260,N_523);
nor U4855 (N_4855,N_2211,N_1845);
or U4856 (N_4856,N_592,N_667);
or U4857 (N_4857,N_498,N_1765);
nor U4858 (N_4858,N_2944,N_705);
nor U4859 (N_4859,N_64,N_1409);
nand U4860 (N_4860,N_759,N_1057);
and U4861 (N_4861,N_2003,N_807);
nand U4862 (N_4862,N_1785,N_1898);
or U4863 (N_4863,N_5,N_1592);
nor U4864 (N_4864,N_1956,N_2258);
nor U4865 (N_4865,N_1706,N_2332);
and U4866 (N_4866,N_2013,N_2344);
nor U4867 (N_4867,N_1526,N_1730);
nor U4868 (N_4868,N_2000,N_342);
xor U4869 (N_4869,N_691,N_2379);
and U4870 (N_4870,N_1251,N_1647);
or U4871 (N_4871,N_1627,N_965);
nor U4872 (N_4872,N_1424,N_1160);
nor U4873 (N_4873,N_1690,N_2351);
or U4874 (N_4874,N_2262,N_1538);
nor U4875 (N_4875,N_669,N_2029);
xnor U4876 (N_4876,N_1251,N_32);
xor U4877 (N_4877,N_2176,N_1984);
or U4878 (N_4878,N_73,N_2967);
and U4879 (N_4879,N_2845,N_495);
nand U4880 (N_4880,N_1429,N_2940);
nand U4881 (N_4881,N_697,N_431);
and U4882 (N_4882,N_2684,N_1304);
or U4883 (N_4883,N_1205,N_1988);
nor U4884 (N_4884,N_2173,N_449);
and U4885 (N_4885,N_2046,N_105);
or U4886 (N_4886,N_2949,N_793);
or U4887 (N_4887,N_392,N_1236);
nand U4888 (N_4888,N_2254,N_2294);
xnor U4889 (N_4889,N_1687,N_834);
and U4890 (N_4890,N_1673,N_1872);
and U4891 (N_4891,N_1333,N_2149);
xnor U4892 (N_4892,N_2042,N_2681);
nand U4893 (N_4893,N_1925,N_1750);
nor U4894 (N_4894,N_2403,N_194);
or U4895 (N_4895,N_752,N_2699);
and U4896 (N_4896,N_2556,N_2364);
nor U4897 (N_4897,N_226,N_2194);
xor U4898 (N_4898,N_2877,N_1214);
and U4899 (N_4899,N_1554,N_1853);
and U4900 (N_4900,N_2829,N_490);
nand U4901 (N_4901,N_2845,N_2370);
xor U4902 (N_4902,N_1783,N_2427);
nand U4903 (N_4903,N_1061,N_1530);
and U4904 (N_4904,N_2220,N_1038);
nor U4905 (N_4905,N_1312,N_211);
nand U4906 (N_4906,N_224,N_1857);
nor U4907 (N_4907,N_2553,N_201);
and U4908 (N_4908,N_2568,N_239);
xnor U4909 (N_4909,N_1456,N_1544);
nor U4910 (N_4910,N_2584,N_2148);
or U4911 (N_4911,N_1165,N_2727);
and U4912 (N_4912,N_2671,N_1346);
and U4913 (N_4913,N_904,N_272);
nor U4914 (N_4914,N_212,N_2812);
nor U4915 (N_4915,N_525,N_2918);
or U4916 (N_4916,N_2256,N_1768);
nor U4917 (N_4917,N_1013,N_1225);
and U4918 (N_4918,N_370,N_2806);
and U4919 (N_4919,N_1315,N_2857);
nor U4920 (N_4920,N_407,N_2019);
xnor U4921 (N_4921,N_1670,N_1749);
and U4922 (N_4922,N_961,N_1773);
and U4923 (N_4923,N_884,N_465);
or U4924 (N_4924,N_1750,N_1588);
nor U4925 (N_4925,N_59,N_299);
nor U4926 (N_4926,N_1732,N_2899);
or U4927 (N_4927,N_2698,N_2154);
nor U4928 (N_4928,N_344,N_1597);
nand U4929 (N_4929,N_263,N_1643);
and U4930 (N_4930,N_2190,N_2950);
nor U4931 (N_4931,N_1423,N_2335);
xnor U4932 (N_4932,N_355,N_1329);
or U4933 (N_4933,N_2473,N_2320);
nand U4934 (N_4934,N_1386,N_2122);
nand U4935 (N_4935,N_1362,N_1463);
nand U4936 (N_4936,N_958,N_100);
or U4937 (N_4937,N_1024,N_362);
and U4938 (N_4938,N_777,N_436);
xnor U4939 (N_4939,N_2892,N_393);
or U4940 (N_4940,N_1142,N_2432);
nor U4941 (N_4941,N_2388,N_1372);
and U4942 (N_4942,N_1890,N_496);
and U4943 (N_4943,N_911,N_1992);
or U4944 (N_4944,N_1062,N_2076);
nor U4945 (N_4945,N_1763,N_1014);
and U4946 (N_4946,N_62,N_1036);
nor U4947 (N_4947,N_371,N_1520);
nand U4948 (N_4948,N_1795,N_777);
or U4949 (N_4949,N_909,N_1183);
nand U4950 (N_4950,N_2784,N_1966);
nand U4951 (N_4951,N_158,N_1926);
or U4952 (N_4952,N_603,N_2091);
and U4953 (N_4953,N_2132,N_1846);
and U4954 (N_4954,N_2988,N_2692);
nor U4955 (N_4955,N_2679,N_2031);
nor U4956 (N_4956,N_1295,N_2571);
nor U4957 (N_4957,N_2638,N_1848);
nand U4958 (N_4958,N_1655,N_2453);
and U4959 (N_4959,N_2328,N_1401);
and U4960 (N_4960,N_2317,N_2342);
nand U4961 (N_4961,N_332,N_1825);
and U4962 (N_4962,N_2149,N_924);
or U4963 (N_4963,N_1535,N_1139);
xnor U4964 (N_4964,N_2928,N_775);
or U4965 (N_4965,N_1263,N_1158);
nand U4966 (N_4966,N_1272,N_1289);
or U4967 (N_4967,N_1406,N_2243);
or U4968 (N_4968,N_2459,N_2767);
xor U4969 (N_4969,N_1576,N_1682);
nor U4970 (N_4970,N_548,N_1878);
or U4971 (N_4971,N_2694,N_2667);
nand U4972 (N_4972,N_2288,N_549);
xnor U4973 (N_4973,N_2830,N_1977);
nor U4974 (N_4974,N_2879,N_2495);
nand U4975 (N_4975,N_1585,N_1385);
xnor U4976 (N_4976,N_1513,N_1131);
nand U4977 (N_4977,N_547,N_1825);
and U4978 (N_4978,N_1856,N_62);
nand U4979 (N_4979,N_1559,N_1951);
or U4980 (N_4980,N_1191,N_1699);
nand U4981 (N_4981,N_1446,N_473);
or U4982 (N_4982,N_2042,N_890);
or U4983 (N_4983,N_419,N_295);
nand U4984 (N_4984,N_1654,N_249);
nor U4985 (N_4985,N_489,N_2067);
nand U4986 (N_4986,N_2901,N_1597);
and U4987 (N_4987,N_2488,N_2039);
or U4988 (N_4988,N_2803,N_51);
nand U4989 (N_4989,N_1496,N_956);
or U4990 (N_4990,N_669,N_1765);
and U4991 (N_4991,N_2413,N_398);
or U4992 (N_4992,N_2155,N_2098);
nor U4993 (N_4993,N_1625,N_104);
or U4994 (N_4994,N_777,N_600);
and U4995 (N_4995,N_2820,N_2263);
nand U4996 (N_4996,N_1290,N_1607);
nor U4997 (N_4997,N_2925,N_1335);
nor U4998 (N_4998,N_1966,N_1052);
nor U4999 (N_4999,N_506,N_2494);
or U5000 (N_5000,N_536,N_664);
or U5001 (N_5001,N_1828,N_2222);
nor U5002 (N_5002,N_1127,N_217);
and U5003 (N_5003,N_2973,N_759);
or U5004 (N_5004,N_86,N_2089);
xor U5005 (N_5005,N_337,N_2207);
nand U5006 (N_5006,N_1584,N_1222);
and U5007 (N_5007,N_2268,N_475);
nor U5008 (N_5008,N_1743,N_2562);
nor U5009 (N_5009,N_2346,N_2886);
nor U5010 (N_5010,N_934,N_2837);
nor U5011 (N_5011,N_582,N_2848);
nor U5012 (N_5012,N_1292,N_807);
and U5013 (N_5013,N_255,N_633);
nand U5014 (N_5014,N_1195,N_1562);
nor U5015 (N_5015,N_385,N_1838);
nor U5016 (N_5016,N_1792,N_438);
or U5017 (N_5017,N_1953,N_2003);
nand U5018 (N_5018,N_1987,N_914);
and U5019 (N_5019,N_2450,N_396);
xnor U5020 (N_5020,N_461,N_337);
nor U5021 (N_5021,N_2668,N_2391);
nor U5022 (N_5022,N_874,N_449);
nand U5023 (N_5023,N_1963,N_2936);
and U5024 (N_5024,N_448,N_2451);
nor U5025 (N_5025,N_1592,N_458);
or U5026 (N_5026,N_45,N_863);
and U5027 (N_5027,N_2470,N_998);
nor U5028 (N_5028,N_2428,N_2960);
nor U5029 (N_5029,N_2308,N_2789);
nand U5030 (N_5030,N_1141,N_1168);
nor U5031 (N_5031,N_1712,N_1205);
or U5032 (N_5032,N_1534,N_2315);
nor U5033 (N_5033,N_699,N_1452);
or U5034 (N_5034,N_1548,N_1092);
nor U5035 (N_5035,N_1924,N_989);
nor U5036 (N_5036,N_949,N_1049);
or U5037 (N_5037,N_608,N_2629);
xnor U5038 (N_5038,N_489,N_1678);
nand U5039 (N_5039,N_1083,N_2436);
nor U5040 (N_5040,N_234,N_1473);
or U5041 (N_5041,N_1585,N_2530);
nor U5042 (N_5042,N_1733,N_1457);
nand U5043 (N_5043,N_196,N_1721);
nand U5044 (N_5044,N_2606,N_2811);
xor U5045 (N_5045,N_207,N_762);
nor U5046 (N_5046,N_283,N_1881);
nand U5047 (N_5047,N_519,N_2252);
nor U5048 (N_5048,N_2231,N_255);
nor U5049 (N_5049,N_1446,N_1067);
or U5050 (N_5050,N_519,N_817);
and U5051 (N_5051,N_1545,N_1226);
nand U5052 (N_5052,N_2494,N_832);
or U5053 (N_5053,N_2489,N_2078);
or U5054 (N_5054,N_7,N_2348);
and U5055 (N_5055,N_532,N_1435);
xnor U5056 (N_5056,N_2878,N_2696);
nor U5057 (N_5057,N_1748,N_1193);
and U5058 (N_5058,N_2976,N_1854);
and U5059 (N_5059,N_1185,N_1571);
nand U5060 (N_5060,N_2226,N_120);
nor U5061 (N_5061,N_1383,N_2084);
or U5062 (N_5062,N_1443,N_2216);
and U5063 (N_5063,N_2758,N_993);
or U5064 (N_5064,N_2445,N_964);
xnor U5065 (N_5065,N_176,N_288);
xor U5066 (N_5066,N_208,N_870);
nor U5067 (N_5067,N_2360,N_1005);
and U5068 (N_5068,N_1690,N_2693);
or U5069 (N_5069,N_2029,N_1633);
or U5070 (N_5070,N_1652,N_1846);
nand U5071 (N_5071,N_1414,N_2140);
or U5072 (N_5072,N_1618,N_326);
and U5073 (N_5073,N_556,N_2341);
or U5074 (N_5074,N_1347,N_2927);
nand U5075 (N_5075,N_575,N_2982);
nand U5076 (N_5076,N_1647,N_793);
and U5077 (N_5077,N_860,N_1677);
or U5078 (N_5078,N_2511,N_982);
or U5079 (N_5079,N_490,N_1592);
or U5080 (N_5080,N_2292,N_614);
and U5081 (N_5081,N_2050,N_1054);
or U5082 (N_5082,N_2995,N_2272);
nand U5083 (N_5083,N_2175,N_1946);
nor U5084 (N_5084,N_791,N_2436);
nor U5085 (N_5085,N_1477,N_2281);
nor U5086 (N_5086,N_2857,N_1875);
nor U5087 (N_5087,N_1121,N_2329);
nand U5088 (N_5088,N_1625,N_376);
or U5089 (N_5089,N_82,N_2591);
and U5090 (N_5090,N_2518,N_1268);
nand U5091 (N_5091,N_2957,N_653);
nand U5092 (N_5092,N_1456,N_2951);
nor U5093 (N_5093,N_904,N_2633);
nor U5094 (N_5094,N_2123,N_632);
and U5095 (N_5095,N_1495,N_1068);
nand U5096 (N_5096,N_703,N_2343);
nor U5097 (N_5097,N_1851,N_2707);
and U5098 (N_5098,N_2215,N_2928);
xnor U5099 (N_5099,N_1075,N_1786);
and U5100 (N_5100,N_2044,N_54);
nand U5101 (N_5101,N_2207,N_968);
nor U5102 (N_5102,N_2105,N_2392);
nor U5103 (N_5103,N_971,N_1413);
or U5104 (N_5104,N_2293,N_1807);
xnor U5105 (N_5105,N_327,N_2970);
nand U5106 (N_5106,N_1411,N_20);
nand U5107 (N_5107,N_1896,N_1387);
or U5108 (N_5108,N_63,N_2056);
nor U5109 (N_5109,N_2359,N_837);
or U5110 (N_5110,N_1194,N_2422);
or U5111 (N_5111,N_623,N_1511);
nor U5112 (N_5112,N_2283,N_372);
and U5113 (N_5113,N_1671,N_1776);
nor U5114 (N_5114,N_371,N_619);
nand U5115 (N_5115,N_2805,N_1824);
xor U5116 (N_5116,N_1765,N_1510);
nor U5117 (N_5117,N_1229,N_874);
or U5118 (N_5118,N_998,N_2434);
and U5119 (N_5119,N_475,N_1901);
or U5120 (N_5120,N_2744,N_636);
nand U5121 (N_5121,N_2048,N_2695);
or U5122 (N_5122,N_1014,N_1168);
nand U5123 (N_5123,N_275,N_981);
nor U5124 (N_5124,N_2647,N_2107);
nand U5125 (N_5125,N_2714,N_1741);
and U5126 (N_5126,N_1180,N_2320);
and U5127 (N_5127,N_428,N_1388);
or U5128 (N_5128,N_162,N_2488);
xor U5129 (N_5129,N_188,N_1863);
xnor U5130 (N_5130,N_2177,N_135);
nor U5131 (N_5131,N_886,N_2218);
and U5132 (N_5132,N_500,N_838);
or U5133 (N_5133,N_2959,N_2788);
xnor U5134 (N_5134,N_178,N_72);
or U5135 (N_5135,N_2502,N_1432);
nor U5136 (N_5136,N_1594,N_663);
and U5137 (N_5137,N_154,N_1795);
nor U5138 (N_5138,N_270,N_1814);
nand U5139 (N_5139,N_725,N_1881);
nand U5140 (N_5140,N_2201,N_522);
nand U5141 (N_5141,N_1598,N_2595);
nand U5142 (N_5142,N_1025,N_2838);
and U5143 (N_5143,N_197,N_789);
or U5144 (N_5144,N_2358,N_1335);
nor U5145 (N_5145,N_2649,N_2580);
nor U5146 (N_5146,N_1277,N_2985);
or U5147 (N_5147,N_867,N_866);
or U5148 (N_5148,N_2174,N_1563);
nand U5149 (N_5149,N_1765,N_1625);
and U5150 (N_5150,N_680,N_2065);
nor U5151 (N_5151,N_1461,N_2043);
and U5152 (N_5152,N_2263,N_625);
and U5153 (N_5153,N_2689,N_739);
or U5154 (N_5154,N_256,N_2775);
nand U5155 (N_5155,N_2022,N_1027);
and U5156 (N_5156,N_2563,N_2997);
xor U5157 (N_5157,N_192,N_1665);
and U5158 (N_5158,N_2620,N_198);
and U5159 (N_5159,N_184,N_1537);
and U5160 (N_5160,N_2513,N_1225);
nand U5161 (N_5161,N_2506,N_2770);
nand U5162 (N_5162,N_333,N_2683);
xnor U5163 (N_5163,N_1502,N_2588);
nor U5164 (N_5164,N_418,N_350);
xor U5165 (N_5165,N_2824,N_743);
nor U5166 (N_5166,N_367,N_8);
nand U5167 (N_5167,N_984,N_328);
nor U5168 (N_5168,N_665,N_2641);
nor U5169 (N_5169,N_2678,N_2387);
or U5170 (N_5170,N_1225,N_1789);
nor U5171 (N_5171,N_117,N_668);
and U5172 (N_5172,N_2941,N_275);
nand U5173 (N_5173,N_2560,N_2821);
and U5174 (N_5174,N_1900,N_1058);
nor U5175 (N_5175,N_1385,N_1610);
and U5176 (N_5176,N_2682,N_106);
and U5177 (N_5177,N_1945,N_2161);
or U5178 (N_5178,N_2878,N_39);
or U5179 (N_5179,N_1646,N_1359);
nor U5180 (N_5180,N_1106,N_1623);
or U5181 (N_5181,N_898,N_2387);
xnor U5182 (N_5182,N_1578,N_2430);
xor U5183 (N_5183,N_811,N_1160);
nor U5184 (N_5184,N_1777,N_200);
nor U5185 (N_5185,N_1145,N_778);
or U5186 (N_5186,N_2424,N_1785);
or U5187 (N_5187,N_2360,N_525);
xnor U5188 (N_5188,N_1410,N_2451);
nand U5189 (N_5189,N_1344,N_1001);
or U5190 (N_5190,N_2096,N_2051);
nor U5191 (N_5191,N_1871,N_1587);
nand U5192 (N_5192,N_134,N_1223);
xnor U5193 (N_5193,N_1994,N_2656);
nor U5194 (N_5194,N_128,N_625);
or U5195 (N_5195,N_792,N_2335);
or U5196 (N_5196,N_2150,N_1940);
xnor U5197 (N_5197,N_1847,N_1173);
nand U5198 (N_5198,N_2044,N_907);
nor U5199 (N_5199,N_241,N_1582);
and U5200 (N_5200,N_1102,N_2025);
or U5201 (N_5201,N_2224,N_363);
nor U5202 (N_5202,N_270,N_1290);
nand U5203 (N_5203,N_2103,N_2518);
xnor U5204 (N_5204,N_2780,N_2384);
and U5205 (N_5205,N_2181,N_452);
and U5206 (N_5206,N_1915,N_2377);
nand U5207 (N_5207,N_779,N_86);
or U5208 (N_5208,N_472,N_1753);
nor U5209 (N_5209,N_744,N_413);
nor U5210 (N_5210,N_853,N_1482);
nor U5211 (N_5211,N_2404,N_121);
nand U5212 (N_5212,N_1665,N_420);
and U5213 (N_5213,N_1438,N_731);
nand U5214 (N_5214,N_2728,N_432);
nand U5215 (N_5215,N_1616,N_250);
xor U5216 (N_5216,N_2788,N_1095);
nor U5217 (N_5217,N_1843,N_1666);
and U5218 (N_5218,N_2921,N_263);
nor U5219 (N_5219,N_1144,N_831);
xnor U5220 (N_5220,N_380,N_1595);
and U5221 (N_5221,N_927,N_2242);
nand U5222 (N_5222,N_696,N_668);
nor U5223 (N_5223,N_2764,N_247);
nand U5224 (N_5224,N_204,N_2891);
nor U5225 (N_5225,N_305,N_2241);
nor U5226 (N_5226,N_1229,N_250);
nand U5227 (N_5227,N_2732,N_1943);
or U5228 (N_5228,N_1491,N_2859);
or U5229 (N_5229,N_87,N_2848);
and U5230 (N_5230,N_2672,N_700);
or U5231 (N_5231,N_1704,N_2089);
and U5232 (N_5232,N_1598,N_1727);
or U5233 (N_5233,N_1552,N_1558);
nor U5234 (N_5234,N_2668,N_614);
and U5235 (N_5235,N_966,N_2122);
and U5236 (N_5236,N_2109,N_2148);
nor U5237 (N_5237,N_2494,N_66);
or U5238 (N_5238,N_821,N_1457);
nand U5239 (N_5239,N_1033,N_759);
and U5240 (N_5240,N_1314,N_279);
and U5241 (N_5241,N_2257,N_2731);
and U5242 (N_5242,N_1744,N_207);
nor U5243 (N_5243,N_2083,N_2132);
xnor U5244 (N_5244,N_1086,N_57);
or U5245 (N_5245,N_1781,N_2876);
and U5246 (N_5246,N_380,N_2934);
and U5247 (N_5247,N_1158,N_478);
and U5248 (N_5248,N_1282,N_2883);
nand U5249 (N_5249,N_987,N_2424);
nor U5250 (N_5250,N_951,N_2931);
nor U5251 (N_5251,N_301,N_2169);
and U5252 (N_5252,N_30,N_1630);
or U5253 (N_5253,N_350,N_31);
nor U5254 (N_5254,N_207,N_588);
nor U5255 (N_5255,N_2906,N_2690);
xor U5256 (N_5256,N_1165,N_2071);
or U5257 (N_5257,N_1885,N_1473);
and U5258 (N_5258,N_2947,N_2078);
xor U5259 (N_5259,N_598,N_99);
or U5260 (N_5260,N_1842,N_478);
and U5261 (N_5261,N_580,N_1146);
and U5262 (N_5262,N_1511,N_2257);
nor U5263 (N_5263,N_620,N_1847);
nand U5264 (N_5264,N_2882,N_2697);
nand U5265 (N_5265,N_2728,N_1394);
nand U5266 (N_5266,N_2824,N_1503);
and U5267 (N_5267,N_2675,N_739);
or U5268 (N_5268,N_1499,N_2904);
and U5269 (N_5269,N_2298,N_2085);
or U5270 (N_5270,N_615,N_2117);
nand U5271 (N_5271,N_441,N_692);
nand U5272 (N_5272,N_663,N_2215);
or U5273 (N_5273,N_1802,N_1842);
or U5274 (N_5274,N_1312,N_529);
nand U5275 (N_5275,N_1068,N_62);
xor U5276 (N_5276,N_2810,N_1658);
or U5277 (N_5277,N_1153,N_1096);
and U5278 (N_5278,N_2122,N_465);
or U5279 (N_5279,N_1947,N_2179);
or U5280 (N_5280,N_1464,N_2410);
and U5281 (N_5281,N_174,N_726);
nand U5282 (N_5282,N_462,N_1523);
nand U5283 (N_5283,N_942,N_2879);
nand U5284 (N_5284,N_1932,N_2374);
nand U5285 (N_5285,N_1280,N_2203);
or U5286 (N_5286,N_2341,N_600);
nor U5287 (N_5287,N_856,N_2369);
xor U5288 (N_5288,N_1654,N_1326);
and U5289 (N_5289,N_1459,N_2778);
nor U5290 (N_5290,N_2849,N_1911);
nor U5291 (N_5291,N_1965,N_128);
nand U5292 (N_5292,N_2155,N_2034);
nand U5293 (N_5293,N_819,N_1014);
nor U5294 (N_5294,N_2529,N_2688);
and U5295 (N_5295,N_1258,N_965);
and U5296 (N_5296,N_1517,N_90);
nand U5297 (N_5297,N_863,N_641);
xor U5298 (N_5298,N_937,N_1992);
nor U5299 (N_5299,N_2448,N_1403);
nor U5300 (N_5300,N_998,N_1086);
xor U5301 (N_5301,N_2070,N_60);
nand U5302 (N_5302,N_2747,N_2103);
or U5303 (N_5303,N_1261,N_1851);
or U5304 (N_5304,N_966,N_1461);
nand U5305 (N_5305,N_1942,N_1896);
nor U5306 (N_5306,N_252,N_221);
or U5307 (N_5307,N_1310,N_272);
and U5308 (N_5308,N_54,N_1180);
nor U5309 (N_5309,N_2998,N_91);
or U5310 (N_5310,N_718,N_2109);
or U5311 (N_5311,N_181,N_1191);
or U5312 (N_5312,N_497,N_1092);
or U5313 (N_5313,N_1514,N_2232);
nand U5314 (N_5314,N_2577,N_2289);
xor U5315 (N_5315,N_51,N_2481);
and U5316 (N_5316,N_1345,N_2668);
nor U5317 (N_5317,N_1575,N_1849);
or U5318 (N_5318,N_2033,N_2045);
nor U5319 (N_5319,N_1913,N_1438);
nor U5320 (N_5320,N_1249,N_2766);
or U5321 (N_5321,N_2084,N_561);
or U5322 (N_5322,N_2409,N_810);
or U5323 (N_5323,N_167,N_2958);
xnor U5324 (N_5324,N_270,N_717);
and U5325 (N_5325,N_358,N_2524);
nor U5326 (N_5326,N_1506,N_432);
or U5327 (N_5327,N_391,N_1704);
nand U5328 (N_5328,N_2480,N_2661);
nor U5329 (N_5329,N_1985,N_568);
and U5330 (N_5330,N_2227,N_697);
and U5331 (N_5331,N_2909,N_490);
or U5332 (N_5332,N_2122,N_587);
nand U5333 (N_5333,N_1715,N_2451);
nand U5334 (N_5334,N_327,N_2880);
and U5335 (N_5335,N_345,N_74);
and U5336 (N_5336,N_2730,N_1628);
nand U5337 (N_5337,N_506,N_2157);
or U5338 (N_5338,N_1466,N_2133);
or U5339 (N_5339,N_1517,N_1454);
and U5340 (N_5340,N_2775,N_2896);
nor U5341 (N_5341,N_1478,N_1998);
nand U5342 (N_5342,N_681,N_727);
nor U5343 (N_5343,N_2042,N_999);
and U5344 (N_5344,N_1064,N_2185);
nand U5345 (N_5345,N_2734,N_1860);
nor U5346 (N_5346,N_459,N_15);
and U5347 (N_5347,N_2187,N_2758);
and U5348 (N_5348,N_1407,N_1973);
nor U5349 (N_5349,N_2203,N_1194);
and U5350 (N_5350,N_2190,N_920);
xnor U5351 (N_5351,N_632,N_2081);
and U5352 (N_5352,N_1338,N_2117);
xnor U5353 (N_5353,N_952,N_689);
nor U5354 (N_5354,N_1226,N_1643);
xnor U5355 (N_5355,N_2018,N_594);
xor U5356 (N_5356,N_781,N_2511);
and U5357 (N_5357,N_205,N_6);
and U5358 (N_5358,N_493,N_2787);
nor U5359 (N_5359,N_2658,N_976);
nand U5360 (N_5360,N_2681,N_326);
nor U5361 (N_5361,N_937,N_594);
nand U5362 (N_5362,N_2111,N_1554);
or U5363 (N_5363,N_1748,N_1081);
nand U5364 (N_5364,N_2962,N_305);
or U5365 (N_5365,N_2308,N_1792);
nor U5366 (N_5366,N_192,N_7);
nand U5367 (N_5367,N_1989,N_1113);
nor U5368 (N_5368,N_306,N_2639);
nor U5369 (N_5369,N_1555,N_82);
nand U5370 (N_5370,N_2876,N_2173);
and U5371 (N_5371,N_2394,N_1311);
and U5372 (N_5372,N_1445,N_1603);
and U5373 (N_5373,N_1256,N_1767);
or U5374 (N_5374,N_1397,N_680);
or U5375 (N_5375,N_725,N_870);
xnor U5376 (N_5376,N_2913,N_1226);
xnor U5377 (N_5377,N_104,N_2771);
nand U5378 (N_5378,N_826,N_968);
nor U5379 (N_5379,N_1942,N_338);
nand U5380 (N_5380,N_1351,N_285);
nand U5381 (N_5381,N_1322,N_1292);
nand U5382 (N_5382,N_11,N_1387);
and U5383 (N_5383,N_1257,N_2476);
nand U5384 (N_5384,N_1219,N_2887);
and U5385 (N_5385,N_215,N_1472);
nand U5386 (N_5386,N_4,N_2443);
nor U5387 (N_5387,N_2752,N_922);
and U5388 (N_5388,N_1732,N_1085);
nor U5389 (N_5389,N_2674,N_2134);
nor U5390 (N_5390,N_349,N_1300);
nand U5391 (N_5391,N_2565,N_370);
and U5392 (N_5392,N_323,N_2717);
nand U5393 (N_5393,N_1098,N_2977);
and U5394 (N_5394,N_311,N_1196);
and U5395 (N_5395,N_2337,N_2077);
nand U5396 (N_5396,N_1527,N_61);
nor U5397 (N_5397,N_965,N_1053);
or U5398 (N_5398,N_2804,N_2376);
or U5399 (N_5399,N_1125,N_1463);
nor U5400 (N_5400,N_1407,N_1444);
and U5401 (N_5401,N_29,N_2475);
or U5402 (N_5402,N_467,N_178);
and U5403 (N_5403,N_2053,N_322);
and U5404 (N_5404,N_121,N_2656);
or U5405 (N_5405,N_2326,N_1718);
or U5406 (N_5406,N_906,N_861);
and U5407 (N_5407,N_886,N_318);
or U5408 (N_5408,N_1054,N_712);
and U5409 (N_5409,N_874,N_145);
nand U5410 (N_5410,N_1347,N_1591);
or U5411 (N_5411,N_1246,N_142);
nor U5412 (N_5412,N_2146,N_2549);
nor U5413 (N_5413,N_156,N_1842);
and U5414 (N_5414,N_1104,N_2338);
or U5415 (N_5415,N_1427,N_69);
nor U5416 (N_5416,N_1687,N_2610);
and U5417 (N_5417,N_366,N_930);
nand U5418 (N_5418,N_1910,N_787);
and U5419 (N_5419,N_1521,N_377);
and U5420 (N_5420,N_2665,N_658);
nand U5421 (N_5421,N_2867,N_263);
nor U5422 (N_5422,N_1720,N_1850);
and U5423 (N_5423,N_704,N_897);
nand U5424 (N_5424,N_1352,N_490);
xor U5425 (N_5425,N_2043,N_2410);
and U5426 (N_5426,N_2907,N_2453);
and U5427 (N_5427,N_2997,N_2062);
xnor U5428 (N_5428,N_897,N_757);
or U5429 (N_5429,N_1978,N_54);
or U5430 (N_5430,N_432,N_2123);
nand U5431 (N_5431,N_1693,N_1320);
nand U5432 (N_5432,N_1473,N_2439);
nor U5433 (N_5433,N_2330,N_1097);
nand U5434 (N_5434,N_1400,N_1991);
nor U5435 (N_5435,N_896,N_126);
or U5436 (N_5436,N_2723,N_841);
nor U5437 (N_5437,N_1319,N_28);
nor U5438 (N_5438,N_2543,N_2644);
nand U5439 (N_5439,N_1656,N_2781);
and U5440 (N_5440,N_1404,N_1597);
nand U5441 (N_5441,N_904,N_394);
nor U5442 (N_5442,N_1614,N_1973);
nand U5443 (N_5443,N_270,N_2204);
nand U5444 (N_5444,N_1514,N_1321);
nand U5445 (N_5445,N_2881,N_2269);
or U5446 (N_5446,N_1805,N_198);
and U5447 (N_5447,N_1447,N_2437);
or U5448 (N_5448,N_1255,N_112);
and U5449 (N_5449,N_1361,N_847);
nor U5450 (N_5450,N_111,N_2922);
and U5451 (N_5451,N_316,N_2678);
and U5452 (N_5452,N_220,N_13);
and U5453 (N_5453,N_2786,N_656);
and U5454 (N_5454,N_2847,N_965);
or U5455 (N_5455,N_274,N_1379);
or U5456 (N_5456,N_685,N_370);
xnor U5457 (N_5457,N_577,N_2611);
or U5458 (N_5458,N_958,N_1883);
nand U5459 (N_5459,N_874,N_735);
or U5460 (N_5460,N_442,N_252);
or U5461 (N_5461,N_1446,N_350);
nand U5462 (N_5462,N_1233,N_559);
and U5463 (N_5463,N_1400,N_110);
or U5464 (N_5464,N_1897,N_1106);
or U5465 (N_5465,N_1725,N_2866);
nor U5466 (N_5466,N_2294,N_2796);
nor U5467 (N_5467,N_1300,N_924);
and U5468 (N_5468,N_1079,N_1450);
nand U5469 (N_5469,N_2588,N_1951);
nor U5470 (N_5470,N_2150,N_314);
nand U5471 (N_5471,N_744,N_2866);
and U5472 (N_5472,N_2247,N_1388);
and U5473 (N_5473,N_926,N_462);
and U5474 (N_5474,N_1953,N_2443);
nor U5475 (N_5475,N_788,N_1738);
nor U5476 (N_5476,N_2298,N_1214);
and U5477 (N_5477,N_2277,N_1405);
nand U5478 (N_5478,N_391,N_2541);
and U5479 (N_5479,N_692,N_2157);
and U5480 (N_5480,N_2418,N_1094);
and U5481 (N_5481,N_2436,N_257);
nor U5482 (N_5482,N_658,N_1010);
and U5483 (N_5483,N_1302,N_439);
nand U5484 (N_5484,N_168,N_667);
nand U5485 (N_5485,N_1969,N_2650);
or U5486 (N_5486,N_1560,N_1196);
xnor U5487 (N_5487,N_2547,N_2540);
nand U5488 (N_5488,N_2194,N_637);
and U5489 (N_5489,N_2958,N_1973);
and U5490 (N_5490,N_353,N_851);
nor U5491 (N_5491,N_511,N_2649);
and U5492 (N_5492,N_901,N_1861);
nand U5493 (N_5493,N_209,N_2500);
and U5494 (N_5494,N_2939,N_2543);
nand U5495 (N_5495,N_2738,N_1164);
or U5496 (N_5496,N_2545,N_460);
or U5497 (N_5497,N_2643,N_201);
xnor U5498 (N_5498,N_1027,N_1404);
nand U5499 (N_5499,N_1315,N_760);
nor U5500 (N_5500,N_1720,N_277);
or U5501 (N_5501,N_2788,N_0);
nor U5502 (N_5502,N_861,N_2004);
xnor U5503 (N_5503,N_1951,N_852);
and U5504 (N_5504,N_2809,N_1974);
nand U5505 (N_5505,N_51,N_667);
or U5506 (N_5506,N_1617,N_1954);
nor U5507 (N_5507,N_1954,N_233);
nor U5508 (N_5508,N_2590,N_958);
and U5509 (N_5509,N_650,N_1820);
and U5510 (N_5510,N_1027,N_2805);
or U5511 (N_5511,N_894,N_1367);
and U5512 (N_5512,N_2266,N_1136);
xor U5513 (N_5513,N_459,N_1684);
nor U5514 (N_5514,N_1708,N_831);
and U5515 (N_5515,N_13,N_338);
or U5516 (N_5516,N_359,N_1953);
or U5517 (N_5517,N_1402,N_77);
and U5518 (N_5518,N_238,N_1139);
nand U5519 (N_5519,N_1715,N_681);
and U5520 (N_5520,N_632,N_2591);
and U5521 (N_5521,N_1175,N_915);
and U5522 (N_5522,N_2208,N_1709);
xor U5523 (N_5523,N_715,N_10);
nor U5524 (N_5524,N_45,N_1478);
or U5525 (N_5525,N_632,N_1507);
nand U5526 (N_5526,N_895,N_1922);
nor U5527 (N_5527,N_1458,N_1056);
and U5528 (N_5528,N_2274,N_2229);
nand U5529 (N_5529,N_211,N_1789);
nand U5530 (N_5530,N_329,N_631);
nand U5531 (N_5531,N_2447,N_404);
and U5532 (N_5532,N_271,N_983);
xnor U5533 (N_5533,N_2893,N_2524);
nand U5534 (N_5534,N_1387,N_2656);
or U5535 (N_5535,N_2680,N_2721);
and U5536 (N_5536,N_2912,N_1141);
nor U5537 (N_5537,N_1423,N_904);
nor U5538 (N_5538,N_2319,N_2216);
and U5539 (N_5539,N_2582,N_173);
and U5540 (N_5540,N_287,N_1711);
nor U5541 (N_5541,N_1762,N_2887);
or U5542 (N_5542,N_1859,N_1744);
xor U5543 (N_5543,N_2761,N_430);
or U5544 (N_5544,N_1020,N_2919);
nand U5545 (N_5545,N_788,N_2124);
nand U5546 (N_5546,N_782,N_2251);
nand U5547 (N_5547,N_2895,N_980);
and U5548 (N_5548,N_1671,N_1969);
nor U5549 (N_5549,N_64,N_1856);
nor U5550 (N_5550,N_2885,N_1660);
nand U5551 (N_5551,N_1048,N_410);
xor U5552 (N_5552,N_597,N_2552);
nand U5553 (N_5553,N_2533,N_817);
or U5554 (N_5554,N_798,N_1086);
xnor U5555 (N_5555,N_1147,N_1574);
or U5556 (N_5556,N_2913,N_1851);
nor U5557 (N_5557,N_59,N_419);
or U5558 (N_5558,N_1332,N_1845);
and U5559 (N_5559,N_493,N_212);
nor U5560 (N_5560,N_2300,N_2446);
and U5561 (N_5561,N_2717,N_1364);
and U5562 (N_5562,N_917,N_101);
or U5563 (N_5563,N_561,N_872);
nand U5564 (N_5564,N_528,N_2648);
or U5565 (N_5565,N_410,N_1840);
xnor U5566 (N_5566,N_2587,N_378);
or U5567 (N_5567,N_1599,N_1081);
nand U5568 (N_5568,N_938,N_1449);
nand U5569 (N_5569,N_992,N_414);
xnor U5570 (N_5570,N_2180,N_379);
or U5571 (N_5571,N_901,N_2097);
nand U5572 (N_5572,N_2202,N_521);
nor U5573 (N_5573,N_1091,N_1404);
or U5574 (N_5574,N_2969,N_1286);
or U5575 (N_5575,N_153,N_461);
nand U5576 (N_5576,N_2096,N_1324);
xor U5577 (N_5577,N_2744,N_1661);
or U5578 (N_5578,N_1591,N_1145);
and U5579 (N_5579,N_1452,N_2436);
nor U5580 (N_5580,N_311,N_1758);
xor U5581 (N_5581,N_1675,N_1591);
nor U5582 (N_5582,N_1018,N_2043);
or U5583 (N_5583,N_532,N_2780);
or U5584 (N_5584,N_483,N_2452);
or U5585 (N_5585,N_1286,N_1082);
or U5586 (N_5586,N_1664,N_234);
or U5587 (N_5587,N_2370,N_35);
or U5588 (N_5588,N_540,N_2763);
nor U5589 (N_5589,N_742,N_2446);
nor U5590 (N_5590,N_995,N_194);
nor U5591 (N_5591,N_2195,N_1302);
nor U5592 (N_5592,N_2484,N_1959);
and U5593 (N_5593,N_1642,N_363);
nor U5594 (N_5594,N_2720,N_1738);
xnor U5595 (N_5595,N_2929,N_406);
nand U5596 (N_5596,N_1001,N_110);
nor U5597 (N_5597,N_1006,N_142);
xnor U5598 (N_5598,N_1902,N_2736);
nand U5599 (N_5599,N_2818,N_1706);
xor U5600 (N_5600,N_2900,N_874);
nand U5601 (N_5601,N_1411,N_1347);
nor U5602 (N_5602,N_2049,N_2206);
nor U5603 (N_5603,N_2588,N_2724);
or U5604 (N_5604,N_1759,N_724);
or U5605 (N_5605,N_58,N_1378);
or U5606 (N_5606,N_716,N_238);
nor U5607 (N_5607,N_2896,N_705);
nor U5608 (N_5608,N_358,N_2756);
xnor U5609 (N_5609,N_1353,N_2749);
xnor U5610 (N_5610,N_2242,N_875);
nand U5611 (N_5611,N_234,N_1691);
and U5612 (N_5612,N_1356,N_711);
and U5613 (N_5613,N_2970,N_907);
nand U5614 (N_5614,N_32,N_1893);
nand U5615 (N_5615,N_1067,N_2229);
and U5616 (N_5616,N_2329,N_356);
nand U5617 (N_5617,N_325,N_681);
and U5618 (N_5618,N_1358,N_1216);
nor U5619 (N_5619,N_1924,N_2881);
or U5620 (N_5620,N_763,N_984);
nand U5621 (N_5621,N_1206,N_298);
and U5622 (N_5622,N_1710,N_474);
nor U5623 (N_5623,N_2563,N_88);
and U5624 (N_5624,N_2664,N_1720);
xnor U5625 (N_5625,N_854,N_1473);
nand U5626 (N_5626,N_716,N_1692);
nor U5627 (N_5627,N_749,N_561);
nand U5628 (N_5628,N_901,N_1184);
nor U5629 (N_5629,N_1242,N_575);
or U5630 (N_5630,N_2483,N_580);
and U5631 (N_5631,N_44,N_230);
and U5632 (N_5632,N_2310,N_1590);
nor U5633 (N_5633,N_2480,N_1115);
and U5634 (N_5634,N_2401,N_539);
nor U5635 (N_5635,N_36,N_1406);
or U5636 (N_5636,N_1732,N_520);
or U5637 (N_5637,N_2098,N_2608);
xnor U5638 (N_5638,N_2815,N_421);
xnor U5639 (N_5639,N_2762,N_1382);
nand U5640 (N_5640,N_618,N_2274);
nand U5641 (N_5641,N_710,N_673);
and U5642 (N_5642,N_128,N_2091);
nor U5643 (N_5643,N_262,N_1449);
nor U5644 (N_5644,N_90,N_1903);
or U5645 (N_5645,N_2429,N_1416);
nor U5646 (N_5646,N_1331,N_1125);
nand U5647 (N_5647,N_1093,N_12);
nand U5648 (N_5648,N_2326,N_1804);
and U5649 (N_5649,N_752,N_2052);
xor U5650 (N_5650,N_2194,N_1109);
or U5651 (N_5651,N_311,N_2783);
and U5652 (N_5652,N_2092,N_842);
and U5653 (N_5653,N_1531,N_894);
nor U5654 (N_5654,N_2929,N_1723);
nor U5655 (N_5655,N_805,N_1270);
nand U5656 (N_5656,N_93,N_196);
and U5657 (N_5657,N_2235,N_2020);
or U5658 (N_5658,N_154,N_147);
and U5659 (N_5659,N_1460,N_536);
nor U5660 (N_5660,N_2817,N_2395);
xnor U5661 (N_5661,N_1247,N_749);
or U5662 (N_5662,N_2714,N_2467);
xnor U5663 (N_5663,N_2474,N_606);
or U5664 (N_5664,N_2998,N_1725);
and U5665 (N_5665,N_1719,N_848);
and U5666 (N_5666,N_1192,N_996);
nor U5667 (N_5667,N_2350,N_1187);
and U5668 (N_5668,N_2478,N_811);
nor U5669 (N_5669,N_1704,N_2893);
and U5670 (N_5670,N_2657,N_1153);
and U5671 (N_5671,N_1570,N_1887);
nand U5672 (N_5672,N_20,N_130);
nor U5673 (N_5673,N_2900,N_2472);
or U5674 (N_5674,N_1470,N_1306);
nand U5675 (N_5675,N_2426,N_2727);
or U5676 (N_5676,N_2373,N_1026);
nand U5677 (N_5677,N_91,N_1834);
nor U5678 (N_5678,N_279,N_982);
and U5679 (N_5679,N_1329,N_1842);
or U5680 (N_5680,N_2028,N_1244);
or U5681 (N_5681,N_190,N_732);
nand U5682 (N_5682,N_2031,N_246);
xor U5683 (N_5683,N_1516,N_250);
and U5684 (N_5684,N_515,N_1418);
nor U5685 (N_5685,N_866,N_1648);
or U5686 (N_5686,N_1594,N_830);
nand U5687 (N_5687,N_2969,N_1497);
nand U5688 (N_5688,N_1820,N_2842);
and U5689 (N_5689,N_1482,N_2289);
nand U5690 (N_5690,N_1643,N_96);
or U5691 (N_5691,N_2241,N_1481);
or U5692 (N_5692,N_1718,N_1120);
xnor U5693 (N_5693,N_2391,N_1769);
and U5694 (N_5694,N_1722,N_962);
xnor U5695 (N_5695,N_2383,N_430);
or U5696 (N_5696,N_1802,N_1634);
xor U5697 (N_5697,N_805,N_56);
or U5698 (N_5698,N_2321,N_184);
or U5699 (N_5699,N_1535,N_547);
or U5700 (N_5700,N_699,N_761);
and U5701 (N_5701,N_1781,N_2121);
nor U5702 (N_5702,N_865,N_2083);
nor U5703 (N_5703,N_865,N_1088);
nor U5704 (N_5704,N_1045,N_1448);
nand U5705 (N_5705,N_2528,N_259);
and U5706 (N_5706,N_2901,N_1968);
or U5707 (N_5707,N_2324,N_311);
and U5708 (N_5708,N_417,N_283);
and U5709 (N_5709,N_2199,N_1030);
and U5710 (N_5710,N_835,N_1921);
xor U5711 (N_5711,N_989,N_878);
nor U5712 (N_5712,N_331,N_2281);
xor U5713 (N_5713,N_1257,N_2309);
nand U5714 (N_5714,N_1315,N_2023);
and U5715 (N_5715,N_1940,N_1118);
or U5716 (N_5716,N_2417,N_2901);
and U5717 (N_5717,N_961,N_179);
and U5718 (N_5718,N_2663,N_69);
nand U5719 (N_5719,N_2391,N_687);
and U5720 (N_5720,N_378,N_187);
and U5721 (N_5721,N_1458,N_353);
and U5722 (N_5722,N_568,N_1784);
or U5723 (N_5723,N_1861,N_1149);
nand U5724 (N_5724,N_969,N_2885);
nor U5725 (N_5725,N_1030,N_19);
or U5726 (N_5726,N_1504,N_297);
nand U5727 (N_5727,N_1554,N_2253);
or U5728 (N_5728,N_2051,N_991);
and U5729 (N_5729,N_1746,N_1092);
nor U5730 (N_5730,N_1130,N_347);
xnor U5731 (N_5731,N_2487,N_2280);
and U5732 (N_5732,N_745,N_1617);
or U5733 (N_5733,N_706,N_2307);
nand U5734 (N_5734,N_1783,N_1899);
or U5735 (N_5735,N_487,N_1718);
or U5736 (N_5736,N_2793,N_1231);
and U5737 (N_5737,N_1134,N_1219);
and U5738 (N_5738,N_173,N_2374);
nand U5739 (N_5739,N_1562,N_1933);
and U5740 (N_5740,N_2315,N_43);
or U5741 (N_5741,N_1751,N_775);
xor U5742 (N_5742,N_778,N_629);
nand U5743 (N_5743,N_646,N_1788);
nand U5744 (N_5744,N_211,N_1174);
or U5745 (N_5745,N_1106,N_1184);
nor U5746 (N_5746,N_1586,N_1672);
nor U5747 (N_5747,N_2775,N_2942);
nand U5748 (N_5748,N_2601,N_2016);
or U5749 (N_5749,N_2403,N_1011);
or U5750 (N_5750,N_1157,N_954);
xor U5751 (N_5751,N_1484,N_2458);
or U5752 (N_5752,N_1437,N_1314);
nand U5753 (N_5753,N_951,N_2142);
nor U5754 (N_5754,N_1114,N_2468);
nand U5755 (N_5755,N_2311,N_2388);
nand U5756 (N_5756,N_2358,N_1401);
or U5757 (N_5757,N_1503,N_84);
nor U5758 (N_5758,N_1267,N_200);
xnor U5759 (N_5759,N_1981,N_1309);
and U5760 (N_5760,N_2891,N_90);
or U5761 (N_5761,N_1311,N_2423);
nand U5762 (N_5762,N_2898,N_1373);
and U5763 (N_5763,N_741,N_456);
nand U5764 (N_5764,N_508,N_1598);
nor U5765 (N_5765,N_900,N_371);
and U5766 (N_5766,N_1731,N_1375);
or U5767 (N_5767,N_24,N_2371);
nand U5768 (N_5768,N_1204,N_1889);
nand U5769 (N_5769,N_680,N_1418);
nand U5770 (N_5770,N_1991,N_2708);
and U5771 (N_5771,N_2878,N_2585);
and U5772 (N_5772,N_548,N_846);
nand U5773 (N_5773,N_2766,N_235);
or U5774 (N_5774,N_119,N_201);
nand U5775 (N_5775,N_1789,N_2270);
or U5776 (N_5776,N_2147,N_525);
and U5777 (N_5777,N_2618,N_549);
or U5778 (N_5778,N_2085,N_1074);
nor U5779 (N_5779,N_1998,N_1121);
nand U5780 (N_5780,N_1674,N_2979);
nand U5781 (N_5781,N_103,N_489);
and U5782 (N_5782,N_2038,N_1396);
or U5783 (N_5783,N_933,N_1053);
and U5784 (N_5784,N_2502,N_323);
or U5785 (N_5785,N_1829,N_335);
or U5786 (N_5786,N_223,N_1061);
and U5787 (N_5787,N_989,N_2023);
and U5788 (N_5788,N_679,N_2178);
xnor U5789 (N_5789,N_1156,N_2165);
or U5790 (N_5790,N_1611,N_1751);
nor U5791 (N_5791,N_2348,N_1437);
xor U5792 (N_5792,N_350,N_1369);
nand U5793 (N_5793,N_480,N_848);
or U5794 (N_5794,N_1421,N_2304);
nor U5795 (N_5795,N_2681,N_1791);
or U5796 (N_5796,N_368,N_1695);
nand U5797 (N_5797,N_1252,N_729);
nor U5798 (N_5798,N_2831,N_671);
or U5799 (N_5799,N_2756,N_2961);
nor U5800 (N_5800,N_1086,N_2961);
nor U5801 (N_5801,N_2809,N_1771);
or U5802 (N_5802,N_2546,N_1800);
nor U5803 (N_5803,N_165,N_420);
or U5804 (N_5804,N_998,N_885);
nand U5805 (N_5805,N_1533,N_653);
and U5806 (N_5806,N_867,N_1295);
or U5807 (N_5807,N_2405,N_1028);
or U5808 (N_5808,N_109,N_8);
nor U5809 (N_5809,N_2428,N_1686);
or U5810 (N_5810,N_1852,N_300);
nor U5811 (N_5811,N_5,N_396);
and U5812 (N_5812,N_516,N_558);
nand U5813 (N_5813,N_1605,N_2159);
xor U5814 (N_5814,N_1757,N_365);
nand U5815 (N_5815,N_2231,N_66);
and U5816 (N_5816,N_707,N_2462);
nor U5817 (N_5817,N_1903,N_667);
nand U5818 (N_5818,N_2328,N_1192);
or U5819 (N_5819,N_694,N_2604);
nor U5820 (N_5820,N_2455,N_993);
and U5821 (N_5821,N_354,N_2537);
or U5822 (N_5822,N_2019,N_918);
nor U5823 (N_5823,N_2450,N_835);
nand U5824 (N_5824,N_913,N_813);
or U5825 (N_5825,N_1375,N_2933);
or U5826 (N_5826,N_2196,N_2306);
or U5827 (N_5827,N_759,N_570);
or U5828 (N_5828,N_964,N_2734);
or U5829 (N_5829,N_1228,N_2412);
or U5830 (N_5830,N_544,N_1156);
or U5831 (N_5831,N_223,N_2782);
and U5832 (N_5832,N_2442,N_2769);
nand U5833 (N_5833,N_900,N_718);
nor U5834 (N_5834,N_2985,N_369);
xnor U5835 (N_5835,N_187,N_1599);
nor U5836 (N_5836,N_1886,N_1368);
and U5837 (N_5837,N_2842,N_2672);
nand U5838 (N_5838,N_1921,N_2940);
nand U5839 (N_5839,N_228,N_2125);
nand U5840 (N_5840,N_1157,N_1985);
and U5841 (N_5841,N_2145,N_1136);
nor U5842 (N_5842,N_2064,N_122);
nand U5843 (N_5843,N_2661,N_1130);
or U5844 (N_5844,N_48,N_890);
and U5845 (N_5845,N_272,N_1106);
and U5846 (N_5846,N_2387,N_1510);
or U5847 (N_5847,N_1380,N_2071);
and U5848 (N_5848,N_1376,N_2163);
or U5849 (N_5849,N_2778,N_1100);
nor U5850 (N_5850,N_864,N_2129);
and U5851 (N_5851,N_2167,N_1033);
nand U5852 (N_5852,N_1276,N_2438);
nor U5853 (N_5853,N_1586,N_2144);
and U5854 (N_5854,N_949,N_1022);
nand U5855 (N_5855,N_1180,N_1567);
xnor U5856 (N_5856,N_458,N_2490);
xnor U5857 (N_5857,N_827,N_636);
nand U5858 (N_5858,N_755,N_1140);
and U5859 (N_5859,N_2385,N_2985);
nand U5860 (N_5860,N_1992,N_389);
xor U5861 (N_5861,N_2769,N_1530);
xor U5862 (N_5862,N_578,N_1441);
nor U5863 (N_5863,N_340,N_347);
nand U5864 (N_5864,N_1665,N_535);
xor U5865 (N_5865,N_1890,N_620);
and U5866 (N_5866,N_1582,N_2200);
or U5867 (N_5867,N_129,N_761);
nand U5868 (N_5868,N_2041,N_1369);
or U5869 (N_5869,N_2246,N_2603);
nand U5870 (N_5870,N_1905,N_1273);
nand U5871 (N_5871,N_738,N_923);
xnor U5872 (N_5872,N_1403,N_1431);
nand U5873 (N_5873,N_2978,N_313);
nand U5874 (N_5874,N_2071,N_2251);
nor U5875 (N_5875,N_127,N_2970);
or U5876 (N_5876,N_1898,N_1158);
xnor U5877 (N_5877,N_1584,N_1977);
nor U5878 (N_5878,N_1721,N_704);
or U5879 (N_5879,N_1332,N_2900);
and U5880 (N_5880,N_814,N_2033);
and U5881 (N_5881,N_1426,N_718);
nor U5882 (N_5882,N_129,N_1979);
and U5883 (N_5883,N_673,N_149);
nand U5884 (N_5884,N_2920,N_2615);
nand U5885 (N_5885,N_187,N_2913);
nand U5886 (N_5886,N_1017,N_977);
xnor U5887 (N_5887,N_2520,N_1524);
xnor U5888 (N_5888,N_338,N_319);
nand U5889 (N_5889,N_1064,N_777);
or U5890 (N_5890,N_2101,N_2316);
nand U5891 (N_5891,N_689,N_405);
nand U5892 (N_5892,N_732,N_2508);
nand U5893 (N_5893,N_2292,N_2523);
and U5894 (N_5894,N_111,N_1909);
nor U5895 (N_5895,N_2506,N_1570);
and U5896 (N_5896,N_1163,N_2069);
nand U5897 (N_5897,N_1199,N_1205);
and U5898 (N_5898,N_317,N_232);
or U5899 (N_5899,N_883,N_1915);
xnor U5900 (N_5900,N_1125,N_2778);
nor U5901 (N_5901,N_978,N_476);
nand U5902 (N_5902,N_2111,N_1112);
xnor U5903 (N_5903,N_2377,N_1998);
xor U5904 (N_5904,N_2520,N_1674);
nor U5905 (N_5905,N_1660,N_7);
or U5906 (N_5906,N_750,N_1842);
or U5907 (N_5907,N_880,N_1542);
or U5908 (N_5908,N_458,N_49);
and U5909 (N_5909,N_2584,N_1241);
or U5910 (N_5910,N_1663,N_1522);
or U5911 (N_5911,N_521,N_1130);
and U5912 (N_5912,N_891,N_882);
nor U5913 (N_5913,N_6,N_2365);
xor U5914 (N_5914,N_1029,N_2127);
nor U5915 (N_5915,N_2994,N_2508);
or U5916 (N_5916,N_825,N_2426);
nor U5917 (N_5917,N_2386,N_2081);
xnor U5918 (N_5918,N_315,N_501);
nor U5919 (N_5919,N_2196,N_1782);
xnor U5920 (N_5920,N_259,N_1833);
nor U5921 (N_5921,N_2634,N_115);
and U5922 (N_5922,N_1207,N_2362);
nand U5923 (N_5923,N_1546,N_1646);
nand U5924 (N_5924,N_1966,N_871);
or U5925 (N_5925,N_24,N_2480);
nand U5926 (N_5926,N_342,N_1664);
nor U5927 (N_5927,N_142,N_1870);
and U5928 (N_5928,N_1796,N_69);
and U5929 (N_5929,N_194,N_2592);
and U5930 (N_5930,N_6,N_180);
nor U5931 (N_5931,N_118,N_1850);
or U5932 (N_5932,N_2563,N_54);
nand U5933 (N_5933,N_962,N_1005);
nand U5934 (N_5934,N_1674,N_2036);
or U5935 (N_5935,N_654,N_1268);
nand U5936 (N_5936,N_216,N_343);
or U5937 (N_5937,N_1860,N_1131);
and U5938 (N_5938,N_2618,N_120);
nor U5939 (N_5939,N_2280,N_1424);
or U5940 (N_5940,N_2228,N_850);
or U5941 (N_5941,N_2075,N_2040);
xnor U5942 (N_5942,N_85,N_1091);
or U5943 (N_5943,N_815,N_1979);
nor U5944 (N_5944,N_2437,N_792);
nor U5945 (N_5945,N_2150,N_506);
and U5946 (N_5946,N_968,N_1918);
nand U5947 (N_5947,N_1644,N_59);
nand U5948 (N_5948,N_2734,N_177);
nor U5949 (N_5949,N_2013,N_2504);
or U5950 (N_5950,N_641,N_789);
or U5951 (N_5951,N_2803,N_564);
nand U5952 (N_5952,N_738,N_1973);
or U5953 (N_5953,N_1997,N_2298);
or U5954 (N_5954,N_1645,N_2730);
or U5955 (N_5955,N_658,N_2330);
nor U5956 (N_5956,N_894,N_2349);
nor U5957 (N_5957,N_2206,N_1643);
or U5958 (N_5958,N_2595,N_1619);
nand U5959 (N_5959,N_1320,N_1849);
nor U5960 (N_5960,N_1371,N_160);
nor U5961 (N_5961,N_2711,N_2381);
and U5962 (N_5962,N_2364,N_748);
nor U5963 (N_5963,N_448,N_813);
and U5964 (N_5964,N_647,N_2623);
or U5965 (N_5965,N_45,N_2488);
nand U5966 (N_5966,N_514,N_2790);
nand U5967 (N_5967,N_2428,N_1815);
xor U5968 (N_5968,N_574,N_1975);
nand U5969 (N_5969,N_2556,N_1241);
nand U5970 (N_5970,N_7,N_671);
nor U5971 (N_5971,N_2172,N_310);
nor U5972 (N_5972,N_2094,N_2155);
and U5973 (N_5973,N_731,N_1957);
nor U5974 (N_5974,N_533,N_2473);
nor U5975 (N_5975,N_615,N_318);
nand U5976 (N_5976,N_997,N_2900);
nand U5977 (N_5977,N_1041,N_2983);
xor U5978 (N_5978,N_260,N_737);
nor U5979 (N_5979,N_161,N_477);
nor U5980 (N_5980,N_2328,N_660);
and U5981 (N_5981,N_2788,N_1276);
nand U5982 (N_5982,N_1946,N_2201);
and U5983 (N_5983,N_988,N_1050);
and U5984 (N_5984,N_174,N_337);
nor U5985 (N_5985,N_2824,N_2473);
nand U5986 (N_5986,N_1187,N_197);
xor U5987 (N_5987,N_425,N_749);
nand U5988 (N_5988,N_2218,N_2246);
or U5989 (N_5989,N_265,N_109);
nand U5990 (N_5990,N_2472,N_1359);
and U5991 (N_5991,N_73,N_2960);
or U5992 (N_5992,N_681,N_1644);
xor U5993 (N_5993,N_2867,N_1511);
nand U5994 (N_5994,N_2148,N_2180);
nor U5995 (N_5995,N_815,N_1962);
and U5996 (N_5996,N_2578,N_2583);
xnor U5997 (N_5997,N_1805,N_1765);
nand U5998 (N_5998,N_240,N_654);
or U5999 (N_5999,N_2251,N_1971);
and U6000 (N_6000,N_3034,N_4519);
nor U6001 (N_6001,N_5896,N_5292);
nor U6002 (N_6002,N_3093,N_3009);
xor U6003 (N_6003,N_3111,N_5123);
nor U6004 (N_6004,N_3588,N_3289);
nor U6005 (N_6005,N_5958,N_5683);
nand U6006 (N_6006,N_4776,N_3225);
nand U6007 (N_6007,N_4007,N_3191);
nand U6008 (N_6008,N_4491,N_3723);
xor U6009 (N_6009,N_3898,N_3790);
nor U6010 (N_6010,N_5024,N_4340);
and U6011 (N_6011,N_5416,N_3439);
nor U6012 (N_6012,N_5921,N_4022);
and U6013 (N_6013,N_4348,N_3695);
or U6014 (N_6014,N_3558,N_3232);
nor U6015 (N_6015,N_5441,N_3420);
xnor U6016 (N_6016,N_4009,N_5503);
xnor U6017 (N_6017,N_3564,N_4233);
and U6018 (N_6018,N_4876,N_3734);
or U6019 (N_6019,N_3958,N_3581);
and U6020 (N_6020,N_4327,N_3768);
nor U6021 (N_6021,N_3902,N_5694);
xnor U6022 (N_6022,N_5258,N_5603);
and U6023 (N_6023,N_5194,N_5628);
and U6024 (N_6024,N_4249,N_4836);
nor U6025 (N_6025,N_3976,N_3379);
xnor U6026 (N_6026,N_5315,N_5122);
nand U6027 (N_6027,N_3578,N_5547);
xor U6028 (N_6028,N_4930,N_4757);
nand U6029 (N_6029,N_4690,N_5710);
nor U6030 (N_6030,N_3281,N_5169);
or U6031 (N_6031,N_4702,N_4400);
nor U6032 (N_6032,N_4916,N_5092);
nor U6033 (N_6033,N_4948,N_3963);
and U6034 (N_6034,N_3228,N_4371);
and U6035 (N_6035,N_4864,N_3503);
nand U6036 (N_6036,N_4823,N_5418);
or U6037 (N_6037,N_5959,N_3526);
nor U6038 (N_6038,N_4449,N_4872);
or U6039 (N_6039,N_5636,N_5447);
xor U6040 (N_6040,N_3540,N_5599);
nand U6041 (N_6041,N_5652,N_3630);
or U6042 (N_6042,N_5728,N_5167);
and U6043 (N_6043,N_5867,N_3167);
and U6044 (N_6044,N_5497,N_5570);
nor U6045 (N_6045,N_3023,N_3192);
or U6046 (N_6046,N_4127,N_4708);
nor U6047 (N_6047,N_4032,N_4532);
xnor U6048 (N_6048,N_4858,N_5727);
nand U6049 (N_6049,N_4970,N_5321);
nand U6050 (N_6050,N_5675,N_4067);
nor U6051 (N_6051,N_3188,N_4723);
or U6052 (N_6052,N_5677,N_3724);
and U6053 (N_6053,N_5239,N_3886);
nor U6054 (N_6054,N_4668,N_3771);
or U6055 (N_6055,N_5500,N_4115);
xnor U6056 (N_6056,N_4407,N_3008);
and U6057 (N_6057,N_5368,N_5175);
nand U6058 (N_6058,N_3012,N_4712);
nor U6059 (N_6059,N_5528,N_4697);
or U6060 (N_6060,N_4052,N_3158);
nor U6061 (N_6061,N_3146,N_4835);
and U6062 (N_6062,N_5392,N_5772);
or U6063 (N_6063,N_4418,N_5119);
and U6064 (N_6064,N_5572,N_3374);
nand U6065 (N_6065,N_3119,N_3038);
or U6066 (N_6066,N_4066,N_5449);
nand U6067 (N_6067,N_3714,N_3626);
nand U6068 (N_6068,N_3406,N_5511);
nand U6069 (N_6069,N_5851,N_5862);
nand U6070 (N_6070,N_3601,N_5939);
nor U6071 (N_6071,N_3179,N_5670);
nor U6072 (N_6072,N_5430,N_4213);
or U6073 (N_6073,N_3229,N_4461);
nand U6074 (N_6074,N_4730,N_5909);
nand U6075 (N_6075,N_4338,N_3748);
and U6076 (N_6076,N_5546,N_4806);
nand U6077 (N_6077,N_3203,N_5007);
nor U6078 (N_6078,N_5767,N_3574);
and U6079 (N_6079,N_4499,N_5973);
nor U6080 (N_6080,N_5494,N_4011);
nor U6081 (N_6081,N_3923,N_5181);
and U6082 (N_6082,N_4214,N_4793);
nand U6083 (N_6083,N_5623,N_4259);
nor U6084 (N_6084,N_4363,N_3711);
xnor U6085 (N_6085,N_5407,N_3956);
or U6086 (N_6086,N_5176,N_4902);
or U6087 (N_6087,N_3913,N_3399);
nor U6088 (N_6088,N_3155,N_4718);
nand U6089 (N_6089,N_4749,N_5417);
xnor U6090 (N_6090,N_4647,N_3161);
and U6091 (N_6091,N_3467,N_5360);
nor U6092 (N_6092,N_5280,N_3637);
nand U6093 (N_6093,N_4493,N_5350);
nand U6094 (N_6094,N_3683,N_5041);
nand U6095 (N_6095,N_3099,N_3794);
nor U6096 (N_6096,N_5733,N_4410);
or U6097 (N_6097,N_4795,N_4291);
and U6098 (N_6098,N_3264,N_4939);
and U6099 (N_6099,N_4350,N_5211);
xor U6100 (N_6100,N_3806,N_4563);
nand U6101 (N_6101,N_3973,N_4738);
xnor U6102 (N_6102,N_5595,N_5410);
nand U6103 (N_6103,N_4859,N_4055);
and U6104 (N_6104,N_5089,N_3985);
nand U6105 (N_6105,N_3471,N_3060);
nor U6106 (N_6106,N_4497,N_4450);
nor U6107 (N_6107,N_4598,N_4705);
and U6108 (N_6108,N_4402,N_3484);
nor U6109 (N_6109,N_5855,N_3352);
nand U6110 (N_6110,N_5844,N_3194);
or U6111 (N_6111,N_5362,N_3181);
nor U6112 (N_6112,N_5965,N_3715);
nand U6113 (N_6113,N_3381,N_4991);
nor U6114 (N_6114,N_5751,N_4178);
or U6115 (N_6115,N_5653,N_4379);
and U6116 (N_6116,N_4633,N_5030);
and U6117 (N_6117,N_4269,N_4159);
nor U6118 (N_6118,N_5584,N_5544);
or U6119 (N_6119,N_3125,N_4920);
and U6120 (N_6120,N_4843,N_3665);
and U6121 (N_6121,N_4355,N_4274);
or U6122 (N_6122,N_3005,N_5289);
nand U6123 (N_6123,N_3497,N_5836);
nand U6124 (N_6124,N_3656,N_4188);
nor U6125 (N_6125,N_4604,N_3906);
nor U6126 (N_6126,N_4397,N_3443);
and U6127 (N_6127,N_3651,N_5815);
xnor U6128 (N_6128,N_5145,N_5179);
nor U6129 (N_6129,N_4404,N_4284);
nand U6130 (N_6130,N_3599,N_5228);
nand U6131 (N_6131,N_3603,N_5748);
and U6132 (N_6132,N_5359,N_5643);
nor U6133 (N_6133,N_4331,N_3693);
or U6134 (N_6134,N_3817,N_5326);
and U6135 (N_6135,N_5960,N_5765);
nand U6136 (N_6136,N_4045,N_4956);
nor U6137 (N_6137,N_4034,N_5071);
or U6138 (N_6138,N_3000,N_3045);
and U6139 (N_6139,N_4280,N_3595);
nand U6140 (N_6140,N_3178,N_5691);
nand U6141 (N_6141,N_5045,N_5843);
nand U6142 (N_6142,N_3361,N_5750);
and U6143 (N_6143,N_5199,N_4536);
and U6144 (N_6144,N_3064,N_4634);
xor U6145 (N_6145,N_3842,N_3705);
and U6146 (N_6146,N_4679,N_5891);
or U6147 (N_6147,N_3669,N_5309);
and U6148 (N_6148,N_4995,N_4834);
nor U6149 (N_6149,N_4874,N_4215);
or U6150 (N_6150,N_4114,N_3988);
and U6151 (N_6151,N_3650,N_5865);
or U6152 (N_6152,N_4720,N_5083);
and U6153 (N_6153,N_5849,N_5113);
nand U6154 (N_6154,N_4089,N_5334);
nor U6155 (N_6155,N_5817,N_3849);
nand U6156 (N_6156,N_3786,N_5496);
or U6157 (N_6157,N_5532,N_4222);
xnor U6158 (N_6158,N_5752,N_5307);
nand U6159 (N_6159,N_3943,N_5517);
and U6160 (N_6160,N_5186,N_3754);
and U6161 (N_6161,N_5795,N_4005);
and U6162 (N_6162,N_5695,N_3431);
and U6163 (N_6163,N_5768,N_4316);
nand U6164 (N_6164,N_3257,N_4674);
nor U6165 (N_6165,N_4002,N_4546);
and U6166 (N_6166,N_5882,N_3680);
nand U6167 (N_6167,N_4422,N_3123);
nor U6168 (N_6168,N_5592,N_4290);
nor U6169 (N_6169,N_5962,N_3563);
or U6170 (N_6170,N_5947,N_4556);
nand U6171 (N_6171,N_4326,N_5871);
nand U6172 (N_6172,N_4539,N_3368);
nor U6173 (N_6173,N_4100,N_4027);
xnor U6174 (N_6174,N_5336,N_4555);
or U6175 (N_6175,N_3059,N_5317);
or U6176 (N_6176,N_3197,N_3719);
or U6177 (N_6177,N_3879,N_5457);
nand U6178 (N_6178,N_4817,N_3424);
nand U6179 (N_6179,N_5645,N_5217);
nand U6180 (N_6180,N_4448,N_4377);
or U6181 (N_6181,N_4049,N_4908);
or U6182 (N_6182,N_3171,N_5074);
nor U6183 (N_6183,N_3538,N_4672);
nand U6184 (N_6184,N_3318,N_4526);
nand U6185 (N_6185,N_3239,N_5117);
and U6186 (N_6186,N_3113,N_5193);
xor U6187 (N_6187,N_5827,N_4568);
and U6188 (N_6188,N_5495,N_3885);
or U6189 (N_6189,N_4505,N_5064);
nand U6190 (N_6190,N_3363,N_3300);
nor U6191 (N_6191,N_3405,N_5605);
and U6192 (N_6192,N_3136,N_3837);
or U6193 (N_6193,N_4294,N_5773);
nand U6194 (N_6194,N_5060,N_3624);
nor U6195 (N_6195,N_3738,N_5271);
and U6196 (N_6196,N_3654,N_4945);
nand U6197 (N_6197,N_5140,N_5541);
nor U6198 (N_6198,N_4594,N_4873);
xor U6199 (N_6199,N_3580,N_4341);
nor U6200 (N_6200,N_4315,N_3168);
and U6201 (N_6201,N_3717,N_5042);
and U6202 (N_6202,N_3979,N_4932);
and U6203 (N_6203,N_3511,N_3344);
nand U6204 (N_6204,N_4965,N_4498);
nand U6205 (N_6205,N_3866,N_4727);
nand U6206 (N_6206,N_3455,N_3029);
or U6207 (N_6207,N_4030,N_3869);
nand U6208 (N_6208,N_4073,N_5026);
and U6209 (N_6209,N_4942,N_4535);
nand U6210 (N_6210,N_4642,N_5957);
nand U6211 (N_6211,N_3354,N_4860);
nor U6212 (N_6212,N_5787,N_4513);
nor U6213 (N_6213,N_3280,N_3833);
xor U6214 (N_6214,N_3250,N_3076);
xnor U6215 (N_6215,N_5143,N_3919);
nor U6216 (N_6216,N_5125,N_3917);
nand U6217 (N_6217,N_4263,N_5372);
nor U6218 (N_6218,N_5450,N_5460);
nor U6219 (N_6219,N_4518,N_5501);
and U6220 (N_6220,N_4112,N_5953);
and U6221 (N_6221,N_3860,N_4924);
nor U6222 (N_6222,N_3295,N_5571);
xor U6223 (N_6223,N_4659,N_3539);
or U6224 (N_6224,N_3508,N_5130);
nand U6225 (N_6225,N_5180,N_3635);
nand U6226 (N_6226,N_3121,N_5949);
nand U6227 (N_6227,N_5835,N_5393);
nor U6228 (N_6228,N_4116,N_4050);
or U6229 (N_6229,N_5961,N_5790);
or U6230 (N_6230,N_5162,N_4297);
nor U6231 (N_6231,N_5461,N_5219);
xnor U6232 (N_6232,N_5552,N_5367);
or U6233 (N_6233,N_3224,N_4717);
and U6234 (N_6234,N_3035,N_4212);
or U6235 (N_6235,N_3547,N_4785);
xor U6236 (N_6236,N_5684,N_5667);
xor U6237 (N_6237,N_4648,N_4166);
and U6238 (N_6238,N_3733,N_4044);
nor U6239 (N_6239,N_4682,N_3075);
and U6240 (N_6240,N_5879,N_5900);
nand U6241 (N_6241,N_4706,N_5913);
or U6242 (N_6242,N_4663,N_4842);
or U6243 (N_6243,N_4919,N_5562);
or U6244 (N_6244,N_5625,N_5897);
or U6245 (N_6245,N_3241,N_5533);
nor U6246 (N_6246,N_4574,N_4875);
nor U6247 (N_6247,N_4866,N_3706);
nand U6248 (N_6248,N_5635,N_3609);
nor U6249 (N_6249,N_4688,N_5484);
or U6250 (N_6250,N_4367,N_4788);
or U6251 (N_6251,N_3288,N_3870);
nand U6252 (N_6252,N_3910,N_5907);
and U6253 (N_6253,N_3440,N_4174);
and U6254 (N_6254,N_5823,N_3341);
and U6255 (N_6255,N_5536,N_4914);
and U6256 (N_6256,N_4586,N_5491);
or U6257 (N_6257,N_5471,N_4868);
or U6258 (N_6258,N_5888,N_5698);
nand U6259 (N_6259,N_5878,N_4311);
nand U6260 (N_6260,N_5682,N_3522);
or U6261 (N_6261,N_5222,N_4314);
and U6262 (N_6262,N_4631,N_5618);
and U6263 (N_6263,N_4888,N_4298);
and U6264 (N_6264,N_3887,N_3552);
and U6265 (N_6265,N_4509,N_3423);
nand U6266 (N_6266,N_4210,N_3623);
nand U6267 (N_6267,N_5762,N_5355);
nor U6268 (N_6268,N_3534,N_3170);
nand U6269 (N_6269,N_4388,N_5602);
nand U6270 (N_6270,N_4463,N_5606);
and U6271 (N_6271,N_5408,N_3106);
nand U6272 (N_6272,N_3980,N_5974);
or U6273 (N_6273,N_3688,N_3110);
and U6274 (N_6274,N_5068,N_5190);
nand U6275 (N_6275,N_3877,N_5246);
nor U6276 (N_6276,N_4614,N_4751);
nor U6277 (N_6277,N_5565,N_4907);
nor U6278 (N_6278,N_4299,N_3215);
or U6279 (N_6279,N_5513,N_3301);
nor U6280 (N_6280,N_3287,N_5824);
nor U6281 (N_6281,N_5740,N_3253);
or U6282 (N_6282,N_3238,N_5912);
and U6283 (N_6283,N_4091,N_3841);
nand U6284 (N_6284,N_3222,N_4025);
and U6285 (N_6285,N_5029,N_4964);
or U6286 (N_6286,N_4081,N_3961);
and U6287 (N_6287,N_5035,N_5697);
or U6288 (N_6288,N_3785,N_3741);
and U6289 (N_6289,N_5290,N_4267);
xnor U6290 (N_6290,N_4624,N_5298);
nand U6291 (N_6291,N_4275,N_4118);
or U6292 (N_6292,N_5930,N_3325);
or U6293 (N_6293,N_5111,N_5875);
xnor U6294 (N_6294,N_3260,N_3182);
or U6295 (N_6295,N_4147,N_5822);
or U6296 (N_6296,N_4272,N_3830);
or U6297 (N_6297,N_3633,N_3051);
nor U6298 (N_6298,N_4987,N_4312);
nand U6299 (N_6299,N_5825,N_4561);
nor U6300 (N_6300,N_5454,N_5210);
xor U6301 (N_6301,N_4629,N_4883);
xor U6302 (N_6302,N_5242,N_5489);
or U6303 (N_6303,N_5103,N_4478);
nor U6304 (N_6304,N_3407,N_4724);
and U6305 (N_6305,N_3872,N_4979);
and U6306 (N_6306,N_5269,N_5786);
or U6307 (N_6307,N_5166,N_3932);
nor U6308 (N_6308,N_4146,N_4958);
nor U6309 (N_6309,N_5468,N_5774);
xor U6310 (N_6310,N_5012,N_4489);
and U6311 (N_6311,N_5178,N_3080);
and U6312 (N_6312,N_4732,N_3929);
xor U6313 (N_6313,N_5088,N_4783);
nand U6314 (N_6314,N_3062,N_3904);
and U6315 (N_6315,N_5658,N_4678);
nand U6316 (N_6316,N_3636,N_4657);
xor U6317 (N_6317,N_5075,N_3784);
or U6318 (N_6318,N_3871,N_5747);
nand U6319 (N_6319,N_3915,N_3172);
and U6320 (N_6320,N_4321,N_5627);
nor U6321 (N_6321,N_5470,N_4000);
and U6322 (N_6322,N_4524,N_5828);
and U6323 (N_6323,N_5008,N_4202);
or U6324 (N_6324,N_3272,N_3415);
nand U6325 (N_6325,N_4313,N_4171);
and U6326 (N_6326,N_5522,N_3356);
and U6327 (N_6327,N_3832,N_5542);
nor U6328 (N_6328,N_4552,N_4753);
nand U6329 (N_6329,N_5525,N_5034);
and U6330 (N_6330,N_5499,N_5459);
nand U6331 (N_6331,N_3367,N_4951);
nand U6332 (N_6332,N_3951,N_4160);
and U6333 (N_6333,N_3199,N_3965);
or U6334 (N_6334,N_3114,N_4562);
or U6335 (N_6335,N_3461,N_5607);
nor U6336 (N_6336,N_5356,N_4770);
nor U6337 (N_6337,N_5956,N_4270);
nor U6338 (N_6338,N_4228,N_3509);
nand U6339 (N_6339,N_4157,N_3813);
and U6340 (N_6340,N_3357,N_5070);
nor U6341 (N_6341,N_3246,N_4940);
nand U6342 (N_6342,N_3823,N_4736);
and U6343 (N_6343,N_3897,N_4437);
and U6344 (N_6344,N_4547,N_3177);
nand U6345 (N_6345,N_4543,N_3487);
nor U6346 (N_6346,N_3970,N_5300);
nand U6347 (N_6347,N_3834,N_5412);
and U6348 (N_6348,N_5788,N_4101);
nand U6349 (N_6349,N_5714,N_5263);
xnor U6350 (N_6350,N_3071,N_5028);
or U6351 (N_6351,N_3799,N_5375);
or U6352 (N_6352,N_4317,N_3912);
nand U6353 (N_6353,N_3493,N_5633);
xnor U6354 (N_6354,N_4623,N_5903);
nor U6355 (N_6355,N_5639,N_3208);
xnor U6356 (N_6356,N_5934,N_3468);
nor U6357 (N_6357,N_4802,N_3767);
nor U6358 (N_6358,N_4058,N_3226);
nand U6359 (N_6359,N_4807,N_3425);
nor U6360 (N_6360,N_3291,N_3818);
xor U6361 (N_6361,N_4515,N_5490);
nor U6362 (N_6362,N_5794,N_4961);
or U6363 (N_6363,N_4225,N_3231);
xnor U6364 (N_6364,N_5475,N_5990);
nor U6365 (N_6365,N_4238,N_4625);
and U6366 (N_6366,N_5504,N_5574);
nand U6367 (N_6367,N_5153,N_3766);
nand U6368 (N_6368,N_3925,N_5188);
nand U6369 (N_6369,N_5719,N_4024);
nand U6370 (N_6370,N_4745,N_3305);
nand U6371 (N_6371,N_3159,N_5380);
nand U6372 (N_6372,N_5832,N_4440);
nand U6373 (N_6373,N_3364,N_3556);
nor U6374 (N_6374,N_3277,N_5308);
and U6375 (N_6375,N_4703,N_5841);
and U6376 (N_6376,N_4646,N_3560);
and U6377 (N_6377,N_3605,N_5195);
and U6378 (N_6378,N_4451,N_3084);
and U6379 (N_6379,N_5201,N_5253);
or U6380 (N_6380,N_3117,N_4975);
and U6381 (N_6381,N_3720,N_3644);
nor U6382 (N_6382,N_5527,N_5955);
nand U6383 (N_6383,N_4947,N_5480);
nand U6384 (N_6384,N_3377,N_4844);
and U6385 (N_6385,N_4181,N_3607);
or U6386 (N_6386,N_5138,N_3242);
nand U6387 (N_6387,N_4131,N_5866);
or U6388 (N_6388,N_3749,N_5873);
nor U6389 (N_6389,N_4486,N_4766);
and U6390 (N_6390,N_3236,N_3263);
or U6391 (N_6391,N_3620,N_4309);
or U6392 (N_6392,N_4018,N_3313);
xnor U6393 (N_6393,N_5739,N_3881);
nand U6394 (N_6394,N_3779,N_4988);
xnor U6395 (N_6395,N_3920,N_3143);
and U6396 (N_6396,N_4768,N_3365);
nor U6397 (N_6397,N_5109,N_5651);
or U6398 (N_6398,N_3147,N_5472);
nor U6399 (N_6399,N_4302,N_5434);
or U6400 (N_6400,N_5649,N_5976);
or U6401 (N_6401,N_3426,N_3993);
xnor U6402 (N_6402,N_4607,N_3506);
or U6403 (N_6403,N_5388,N_4514);
and U6404 (N_6404,N_3882,N_4852);
and U6405 (N_6405,N_4719,N_5040);
and U6406 (N_6406,N_5267,N_5608);
or U6407 (N_6407,N_4884,N_4145);
or U6408 (N_6408,N_5177,N_5758);
xnor U6409 (N_6409,N_4984,N_4686);
nor U6410 (N_6410,N_5400,N_3375);
xor U6411 (N_6411,N_4969,N_4458);
or U6412 (N_6412,N_5686,N_5516);
or U6413 (N_6413,N_4554,N_3995);
and U6414 (N_6414,N_3050,N_5861);
and U6415 (N_6415,N_3999,N_5371);
nand U6416 (N_6416,N_4103,N_3649);
nor U6417 (N_6417,N_5343,N_4801);
and U6418 (N_6418,N_4711,N_4928);
and U6419 (N_6419,N_3632,N_5666);
xnor U6420 (N_6420,N_5227,N_4006);
nand U6421 (N_6421,N_3243,N_4848);
nor U6422 (N_6422,N_5557,N_4699);
nand U6423 (N_6423,N_4993,N_3775);
or U6424 (N_6424,N_3800,N_4784);
and U6425 (N_6425,N_4232,N_5133);
nor U6426 (N_6426,N_4231,N_3673);
or U6427 (N_6427,N_4433,N_4401);
or U6428 (N_6428,N_5975,N_3403);
nand U6429 (N_6429,N_5032,N_3731);
xnor U6430 (N_6430,N_5174,N_3716);
nand U6431 (N_6431,N_5737,N_4370);
and U6432 (N_6432,N_5889,N_5846);
and U6433 (N_6433,N_3602,N_3645);
nor U6434 (N_6434,N_4268,N_3207);
nand U6435 (N_6435,N_5485,N_4927);
and U6436 (N_6436,N_3903,N_3952);
nor U6437 (N_6437,N_4366,N_4952);
and U6438 (N_6438,N_5207,N_3393);
or U6439 (N_6439,N_4061,N_4977);
and U6440 (N_6440,N_4618,N_5509);
nand U6441 (N_6441,N_4256,N_3728);
nor U6442 (N_6442,N_4820,N_5424);
or U6443 (N_6443,N_3745,N_3308);
nand U6444 (N_6444,N_5286,N_5325);
nand U6445 (N_6445,N_4154,N_5399);
and U6446 (N_6446,N_4808,N_5700);
and U6447 (N_6447,N_5771,N_5090);
and U6448 (N_6448,N_4307,N_3247);
and U6449 (N_6449,N_4169,N_3712);
and U6450 (N_6450,N_5847,N_4420);
and U6451 (N_6451,N_4863,N_4137);
nand U6452 (N_6452,N_3011,N_3991);
nor U6453 (N_6453,N_3303,N_4983);
or U6454 (N_6454,N_4608,N_4300);
and U6455 (N_6455,N_4305,N_3438);
or U6456 (N_6456,N_4734,N_4426);
nand U6457 (N_6457,N_5352,N_3944);
nand U6458 (N_6458,N_3722,N_3070);
nor U6459 (N_6459,N_4347,N_3974);
xnor U6460 (N_6460,N_5049,N_5077);
or U6461 (N_6461,N_4803,N_4150);
or U6462 (N_6462,N_3408,N_3582);
and U6463 (N_6463,N_3679,N_3061);
nor U6464 (N_6464,N_3049,N_3502);
nor U6465 (N_6465,N_5819,N_5821);
nand U6466 (N_6466,N_4265,N_4503);
nand U6467 (N_6467,N_5445,N_4219);
nand U6468 (N_6468,N_5936,N_5105);
nor U6469 (N_6469,N_5275,N_5048);
nand U6470 (N_6470,N_4139,N_4538);
or U6471 (N_6471,N_5146,N_5241);
xnor U6472 (N_6472,N_3165,N_3498);
or U6473 (N_6473,N_4099,N_3937);
xnor U6474 (N_6474,N_4460,N_4906);
nand U6475 (N_6475,N_5314,N_4846);
or U6476 (N_6476,N_4129,N_4949);
xor U6477 (N_6477,N_5556,N_4130);
and U6478 (N_6478,N_5419,N_4251);
and U6479 (N_6479,N_3782,N_5087);
or U6480 (N_6480,N_5659,N_4192);
nand U6481 (N_6481,N_4392,N_4710);
and U6482 (N_6482,N_4273,N_3322);
xor U6483 (N_6483,N_5988,N_4056);
and U6484 (N_6484,N_5724,N_3996);
nand U6485 (N_6485,N_5502,N_3604);
nor U6486 (N_6486,N_5100,N_3825);
or U6487 (N_6487,N_3209,N_5735);
nor U6488 (N_6488,N_5025,N_4641);
nor U6489 (N_6489,N_3320,N_4797);
and U6490 (N_6490,N_5053,N_5778);
nand U6491 (N_6491,N_3819,N_4346);
or U6492 (N_6492,N_5814,N_3612);
xor U6493 (N_6493,N_3883,N_5086);
nor U6494 (N_6494,N_5134,N_5243);
nor U6495 (N_6495,N_5634,N_5019);
nand U6496 (N_6496,N_4725,N_3349);
and U6497 (N_6497,N_5523,N_5421);
and U6498 (N_6498,N_5327,N_4336);
and U6499 (N_6499,N_4588,N_5252);
xnor U6500 (N_6500,N_3404,N_4482);
xor U6501 (N_6501,N_5059,N_3590);
and U6502 (N_6502,N_3681,N_3340);
nor U6503 (N_6503,N_5906,N_3524);
nand U6504 (N_6504,N_3332,N_4709);
nor U6505 (N_6505,N_4603,N_3444);
or U6506 (N_6506,N_5255,N_4894);
nand U6507 (N_6507,N_4597,N_5310);
and U6508 (N_6508,N_5382,N_3827);
xnor U6509 (N_6509,N_5559,N_4578);
nor U6510 (N_6510,N_4387,N_3625);
nor U6511 (N_6511,N_3546,N_5863);
or U6512 (N_6512,N_3098,N_3457);
and U6513 (N_6513,N_4733,N_4800);
or U6514 (N_6514,N_5342,N_3998);
nand U6515 (N_6515,N_3659,N_4502);
nor U6516 (N_6516,N_4840,N_4587);
and U6517 (N_6517,N_3206,N_5353);
and U6518 (N_6518,N_4164,N_4296);
nand U6519 (N_6519,N_5521,N_5184);
or U6520 (N_6520,N_4764,N_4891);
nand U6521 (N_6521,N_4643,N_4580);
xor U6522 (N_6522,N_5806,N_3691);
and U6523 (N_6523,N_5112,N_3535);
or U6524 (N_6524,N_5984,N_3290);
nor U6525 (N_6525,N_3972,N_3310);
xnor U6526 (N_6526,N_5413,N_3889);
and U6527 (N_6527,N_3610,N_5800);
and U6528 (N_6528,N_3355,N_4917);
nor U6529 (N_6529,N_3351,N_5617);
and U6530 (N_6530,N_4170,N_3366);
nor U6531 (N_6531,N_3154,N_3058);
nor U6532 (N_6532,N_5868,N_5224);
nor U6533 (N_6533,N_3648,N_5428);
or U6534 (N_6534,N_3551,N_3150);
and U6535 (N_6535,N_5295,N_4735);
xor U6536 (N_6536,N_5567,N_4209);
nor U6537 (N_6537,N_5622,N_5576);
or U6538 (N_6538,N_4905,N_5783);
or U6539 (N_6539,N_3275,N_5985);
nor U6540 (N_6540,N_5226,N_4572);
or U6541 (N_6541,N_5431,N_5374);
or U6542 (N_6542,N_3274,N_4108);
nor U6543 (N_6543,N_3103,N_4152);
xor U6544 (N_6544,N_3465,N_4658);
or U6545 (N_6545,N_3152,N_4041);
xor U6546 (N_6546,N_3573,N_3737);
nor U6547 (N_6547,N_5689,N_5152);
nand U6548 (N_6548,N_3811,N_5020);
xor U6549 (N_6549,N_3577,N_3309);
and U6550 (N_6550,N_3687,N_5121);
nand U6551 (N_6551,N_4017,N_3270);
and U6552 (N_6552,N_4323,N_4707);
xor U6553 (N_6553,N_3664,N_5196);
and U6554 (N_6554,N_5438,N_3730);
nand U6555 (N_6555,N_3735,N_5157);
and U6556 (N_6556,N_3500,N_5512);
nand U6557 (N_6557,N_5776,N_4996);
nor U6558 (N_6558,N_4086,N_4357);
nand U6559 (N_6559,N_5558,N_4845);
or U6560 (N_6560,N_4804,N_3863);
or U6561 (N_6561,N_3298,N_3187);
nand U6562 (N_6562,N_4900,N_4413);
xor U6563 (N_6563,N_5853,N_5935);
nand U6564 (N_6564,N_3598,N_5706);
and U6565 (N_6565,N_3130,N_3663);
or U6566 (N_6566,N_3388,N_5529);
nand U6567 (N_6567,N_3251,N_4827);
or U6568 (N_6568,N_5389,N_5276);
or U6569 (N_6569,N_3041,N_3888);
nand U6570 (N_6570,N_4162,N_4691);
nand U6571 (N_6571,N_4981,N_4922);
nor U6572 (N_6572,N_3959,N_3921);
or U6573 (N_6573,N_4810,N_4528);
or U6574 (N_6574,N_3616,N_3448);
or U6575 (N_6575,N_3092,N_5209);
xnor U6576 (N_6576,N_3791,N_4322);
or U6577 (N_6577,N_5126,N_5015);
xnor U6578 (N_6578,N_5277,N_5182);
nor U6579 (N_6579,N_5526,N_3981);
or U6580 (N_6580,N_3100,N_4689);
xnor U6581 (N_6581,N_4356,N_3048);
and U6582 (N_6582,N_5335,N_4522);
and U6583 (N_6583,N_5937,N_5566);
nand U6584 (N_6584,N_5160,N_3053);
and U6585 (N_6585,N_5358,N_3382);
or U6586 (N_6586,N_5661,N_5303);
and U6587 (N_6587,N_4419,N_3657);
nand U6588 (N_6588,N_5980,N_3007);
nor U6589 (N_6589,N_5807,N_5137);
or U6590 (N_6590,N_5573,N_5216);
or U6591 (N_6591,N_4609,N_5948);
nand U6592 (N_6592,N_5816,N_5995);
xor U6593 (N_6593,N_3373,N_4180);
xnor U6594 (N_6594,N_3814,N_4445);
xor U6595 (N_6595,N_3317,N_4654);
nand U6596 (N_6596,N_3046,N_4673);
nand U6597 (N_6597,N_5106,N_5208);
nor U6598 (N_6598,N_3643,N_5091);
or U6599 (N_6599,N_4809,N_3781);
nand U6600 (N_6600,N_4409,N_5676);
nor U6601 (N_6601,N_5031,N_3647);
and U6602 (N_6602,N_4780,N_5038);
and U6603 (N_6603,N_5669,N_5838);
nor U6604 (N_6604,N_4226,N_3211);
or U6605 (N_6605,N_5213,N_3078);
nor U6606 (N_6606,N_3235,N_4072);
nand U6607 (N_6607,N_4083,N_4567);
nor U6608 (N_6608,N_3437,N_4989);
nor U6609 (N_6609,N_3726,N_5601);
and U6610 (N_6610,N_3279,N_3164);
nand U6611 (N_6611,N_4798,N_4046);
or U6612 (N_6612,N_5311,N_3315);
nand U6613 (N_6613,N_4829,N_5520);
xor U6614 (N_6614,N_3019,N_5970);
xor U6615 (N_6615,N_4861,N_3851);
xor U6616 (N_6616,N_5524,N_3619);
nand U6617 (N_6617,N_5132,N_3585);
and U6618 (N_6618,N_4773,N_3934);
and U6619 (N_6619,N_4075,N_4933);
or U6620 (N_6620,N_3327,N_3252);
or U6621 (N_6621,N_5397,N_3445);
nand U6622 (N_6622,N_3334,N_4242);
or U6623 (N_6623,N_4252,N_4973);
and U6624 (N_6624,N_5240,N_3180);
nor U6625 (N_6625,N_4473,N_4098);
nand U6626 (N_6626,N_5946,N_4584);
and U6627 (N_6627,N_5549,N_3495);
and U6628 (N_6628,N_5225,N_3436);
or U6629 (N_6629,N_5223,N_4759);
nor U6630 (N_6630,N_5894,N_4790);
nor U6631 (N_6631,N_4470,N_3129);
or U6632 (N_6632,N_3613,N_4258);
or U6633 (N_6633,N_5701,N_5757);
nor U6634 (N_6634,N_5594,N_3496);
nand U6635 (N_6635,N_3732,N_5338);
nor U6636 (N_6636,N_3634,N_4019);
xnor U6637 (N_6637,N_3097,N_3328);
or U6638 (N_6638,N_4992,N_4264);
nor U6639 (N_6639,N_4063,N_5681);
nor U6640 (N_6640,N_3294,N_3751);
nor U6641 (N_6641,N_3671,N_4839);
nor U6642 (N_6642,N_5621,N_5498);
nand U6643 (N_6643,N_4120,N_3930);
and U6644 (N_6644,N_3501,N_4042);
and U6645 (N_6645,N_4791,N_3583);
or U6646 (N_6646,N_3918,N_3276);
nor U6647 (N_6647,N_5510,N_5139);
xnor U6648 (N_6648,N_3662,N_4306);
or U6649 (N_6649,N_4337,N_4047);
xor U6650 (N_6650,N_5884,N_4411);
or U6651 (N_6651,N_3614,N_5918);
xor U6652 (N_6652,N_3922,N_4261);
and U6653 (N_6653,N_5761,N_5611);
nand U6654 (N_6654,N_4378,N_5539);
nor U6655 (N_6655,N_5010,N_5781);
xnor U6656 (N_6656,N_4218,N_3116);
or U6657 (N_6657,N_3808,N_3433);
nand U6658 (N_6658,N_4376,N_4204);
and U6659 (N_6659,N_4761,N_3453);
nand U6660 (N_6660,N_5596,N_5908);
xnor U6661 (N_6661,N_5411,N_4650);
and U6662 (N_6662,N_3047,N_4500);
nand U6663 (N_6663,N_3674,N_3798);
or U6664 (N_6664,N_4469,N_3175);
nor U6665 (N_6665,N_3826,N_3086);
nor U6666 (N_6666,N_5093,N_4974);
nor U6667 (N_6667,N_5312,N_3267);
or U6668 (N_6668,N_4796,N_5678);
and U6669 (N_6669,N_4755,N_5069);
and U6670 (N_6670,N_5979,N_4446);
and U6671 (N_6671,N_4369,N_5569);
nand U6672 (N_6672,N_5730,N_3261);
nand U6673 (N_6673,N_3517,N_5690);
nor U6674 (N_6674,N_5696,N_5991);
and U6675 (N_6675,N_3617,N_5972);
xor U6676 (N_6676,N_4229,N_3063);
nor U6677 (N_6677,N_5455,N_5076);
nand U6678 (N_6678,N_3997,N_5051);
nor U6679 (N_6679,N_5050,N_4639);
nand U6680 (N_6680,N_5172,N_3470);
nand U6681 (N_6681,N_5001,N_3510);
or U6682 (N_6682,N_4506,N_3718);
nor U6683 (N_6683,N_4728,N_4878);
or U6684 (N_6684,N_4282,N_3725);
nand U6685 (N_6685,N_3037,N_5799);
nand U6686 (N_6686,N_3761,N_4847);
nand U6687 (N_6687,N_4121,N_4889);
nor U6688 (N_6688,N_4240,N_5654);
or U6689 (N_6689,N_5848,N_3043);
and U6690 (N_6690,N_3316,N_4276);
nor U6691 (N_6691,N_3537,N_3911);
and U6692 (N_6692,N_5218,N_3218);
and U6693 (N_6693,N_5766,N_3213);
and U6694 (N_6694,N_4837,N_4610);
and U6695 (N_6695,N_5924,N_4248);
nand U6696 (N_6696,N_4669,N_3824);
nor U6697 (N_6697,N_3434,N_4769);
nor U6698 (N_6698,N_3642,N_5044);
and U6699 (N_6699,N_4822,N_3935);
xor U6700 (N_6700,N_3994,N_5883);
or U6701 (N_6701,N_3987,N_3542);
xnor U6702 (N_6702,N_4071,N_3942);
nand U6703 (N_6703,N_3013,N_4361);
nor U6704 (N_6704,N_5543,N_5493);
and U6705 (N_6705,N_5721,N_3678);
and U6706 (N_6706,N_5231,N_3802);
xor U6707 (N_6707,N_3025,N_5052);
and U6708 (N_6708,N_3521,N_3618);
and U6709 (N_6709,N_3266,N_4599);
nand U6710 (N_6710,N_4167,N_4014);
nand U6711 (N_6711,N_4695,N_5919);
and U6712 (N_6712,N_4429,N_3554);
and U6713 (N_6713,N_4211,N_5487);
nand U6714 (N_6714,N_5432,N_3054);
nor U6715 (N_6715,N_5297,N_5021);
nor U6716 (N_6716,N_3265,N_3052);
nor U6717 (N_6717,N_4109,N_5163);
xor U6718 (N_6718,N_5928,N_4966);
and U6719 (N_6719,N_5705,N_5018);
nor U6720 (N_6720,N_4117,N_4511);
and U6721 (N_6721,N_5080,N_3628);
nand U6722 (N_6722,N_3402,N_4540);
and U6723 (N_6723,N_4537,N_4260);
and U6724 (N_6724,N_3347,N_5237);
and U6725 (N_6725,N_4374,N_3391);
and U6726 (N_6726,N_4153,N_3169);
and U6727 (N_6727,N_5726,N_5341);
nor U6728 (N_6728,N_4416,N_3400);
xnor U6729 (N_6729,N_3562,N_5600);
nand U6730 (N_6730,N_5626,N_3750);
or U6731 (N_6731,N_4176,N_3428);
nor U6732 (N_6732,N_5887,N_5296);
or U6733 (N_6733,N_3703,N_5361);
nand U6734 (N_6734,N_5458,N_3845);
nand U6735 (N_6735,N_3763,N_4467);
xnor U6736 (N_6736,N_4595,N_5415);
nor U6737 (N_6737,N_3982,N_3293);
or U6738 (N_6738,N_4593,N_4126);
and U6739 (N_6739,N_5304,N_4566);
and U6740 (N_6740,N_5261,N_5905);
or U6741 (N_6741,N_3492,N_3507);
xnor U6742 (N_6742,N_5648,N_4010);
nor U6743 (N_6743,N_4122,N_5283);
nand U6744 (N_6744,N_4390,N_5095);
or U6745 (N_6745,N_3072,N_5564);
xor U6746 (N_6746,N_5047,N_4885);
xnor U6747 (N_6747,N_4998,N_3262);
nand U6748 (N_6748,N_3069,N_5971);
and U6749 (N_6749,N_3836,N_3787);
nand U6750 (N_6750,N_5555,N_4324);
and U6751 (N_6751,N_5084,N_5722);
nand U6752 (N_6752,N_4415,N_4849);
or U6753 (N_6753,N_4693,N_3713);
or U6754 (N_6754,N_4683,N_4343);
nor U6755 (N_6755,N_4655,N_3145);
nand U6756 (N_6756,N_5033,N_4838);
or U6757 (N_6757,N_3968,N_5250);
and U6758 (N_6758,N_3975,N_4012);
or U6759 (N_6759,N_5185,N_5023);
or U6760 (N_6760,N_4645,N_4444);
nor U6761 (N_6761,N_5379,N_4144);
nor U6762 (N_6762,N_5775,N_5128);
xnor U6763 (N_6763,N_3016,N_5085);
nand U6764 (N_6764,N_4303,N_5850);
nor U6765 (N_6765,N_5646,N_4644);
and U6766 (N_6766,N_3807,N_5704);
or U6767 (N_6767,N_3042,N_3584);
or U6768 (N_6768,N_5479,N_3454);
and U6769 (N_6769,N_3384,N_4084);
and U6770 (N_6770,N_3677,N_5876);
nand U6771 (N_6771,N_5104,N_4605);
xnor U6772 (N_6772,N_5885,N_4760);
nor U6773 (N_6773,N_3821,N_3329);
nor U6774 (N_6774,N_5394,N_5711);
nand U6775 (N_6775,N_4142,N_4656);
nand U6776 (N_6776,N_5288,N_5901);
or U6777 (N_6777,N_4333,N_3561);
nand U6778 (N_6778,N_4774,N_5687);
or U6779 (N_6779,N_3137,N_3709);
xnor U6780 (N_6780,N_4360,N_4923);
nor U6781 (N_6781,N_5344,N_4936);
xor U6782 (N_6782,N_3875,N_3810);
nand U6783 (N_6783,N_5674,N_3520);
nor U6784 (N_6784,N_5440,N_5588);
nor U6785 (N_6785,N_5385,N_5452);
nand U6786 (N_6786,N_4926,N_5833);
or U6787 (N_6787,N_5305,N_4077);
nor U6788 (N_6788,N_5782,N_4661);
nand U6789 (N_6789,N_3237,N_5720);
nor U6790 (N_6790,N_5409,N_5808);
nor U6791 (N_6791,N_3668,N_3128);
or U6792 (N_6792,N_4971,N_5745);
nand U6793 (N_6793,N_5264,N_3233);
nand U6794 (N_6794,N_5769,N_5942);
or U6795 (N_6795,N_3323,N_4627);
and U6796 (N_6796,N_3138,N_3345);
and U6797 (N_6797,N_3418,N_5647);
nand U6798 (N_6798,N_3744,N_4078);
nor U6799 (N_6799,N_3682,N_4382);
nor U6800 (N_6800,N_5348,N_4234);
nor U6801 (N_6801,N_3087,N_5347);
nand U6802 (N_6802,N_4746,N_5124);
or U6803 (N_6803,N_5204,N_3330);
nor U6804 (N_6804,N_4244,N_4490);
nor U6805 (N_6805,N_3014,N_5892);
nor U6806 (N_6806,N_3843,N_4004);
or U6807 (N_6807,N_5183,N_5785);
and U6808 (N_6808,N_3166,N_4143);
nand U6809 (N_6809,N_4036,N_4243);
or U6810 (N_6810,N_3021,N_5620);
nor U6811 (N_6811,N_3269,N_4771);
nand U6812 (N_6812,N_3077,N_4383);
or U6813 (N_6813,N_5548,N_4534);
or U6814 (N_6814,N_5232,N_5707);
or U6815 (N_6815,N_3419,N_5723);
or U6816 (N_6816,N_5809,N_4854);
and U6817 (N_6817,N_3848,N_5383);
nand U6818 (N_6818,N_5272,N_3353);
and U6819 (N_6819,N_4048,N_3414);
xor U6820 (N_6820,N_3553,N_5151);
or U6821 (N_6821,N_4141,N_4617);
nor U6822 (N_6822,N_3450,N_5993);
and U6823 (N_6823,N_5731,N_3244);
xor U6824 (N_6824,N_5554,N_3282);
or U6825 (N_6825,N_5108,N_3479);
nor U6826 (N_6826,N_5804,N_4236);
nand U6827 (N_6827,N_3331,N_5916);
xor U6828 (N_6828,N_4742,N_5097);
nor U6829 (N_6829,N_5463,N_4677);
nand U6830 (N_6830,N_4293,N_5610);
nor U6831 (N_6831,N_3876,N_5395);
or U6832 (N_6832,N_3891,N_3565);
nor U6833 (N_6833,N_4901,N_4615);
and U6834 (N_6834,N_4069,N_4637);
or U6835 (N_6835,N_3115,N_3689);
xor U6836 (N_6836,N_5729,N_5664);
nand U6837 (N_6837,N_5759,N_4021);
nand U6838 (N_6838,N_4054,N_3868);
or U6839 (N_6839,N_3629,N_5902);
or U6840 (N_6840,N_5803,N_3597);
and U6841 (N_6841,N_4216,N_5672);
and U6842 (N_6842,N_4918,N_3387);
or U6843 (N_6843,N_5999,N_4092);
or U6844 (N_6844,N_5545,N_4664);
and U6845 (N_6845,N_3820,N_3895);
or U6846 (N_6846,N_5693,N_3108);
nand U6847 (N_6847,N_4365,N_5743);
or U6848 (N_6848,N_4479,N_5013);
nor U6849 (N_6849,N_4828,N_3776);
nand U6850 (N_6850,N_4700,N_5464);
and U6851 (N_6851,N_4758,N_3548);
nor U6852 (N_6852,N_5055,N_3002);
and U6853 (N_6853,N_3389,N_4620);
and U6854 (N_6854,N_5712,N_3512);
nand U6855 (N_6855,N_4982,N_3216);
nor U6856 (N_6856,N_4140,N_4904);
nand U6857 (N_6857,N_4474,N_5631);
or U6858 (N_6858,N_4999,N_5760);
and U6859 (N_6859,N_3234,N_5192);
nor U6860 (N_6860,N_3160,N_3945);
xor U6861 (N_6861,N_3721,N_5577);
xor U6862 (N_6862,N_3067,N_3953);
or U6863 (N_6863,N_5262,N_3447);
nor U6864 (N_6864,N_4015,N_3989);
nand U6865 (N_6865,N_3196,N_5284);
or U6866 (N_6866,N_3690,N_3326);
or U6867 (N_6867,N_5478,N_3412);
nor U6868 (N_6868,N_4704,N_5136);
or U6869 (N_6869,N_3708,N_5826);
nand U6870 (N_6870,N_3983,N_4893);
xnor U6871 (N_6871,N_5789,N_5655);
and U6872 (N_6872,N_5386,N_5805);
and U6873 (N_6873,N_3030,N_5812);
nor U6874 (N_6874,N_4023,N_4484);
nor U6875 (N_6875,N_3095,N_3195);
nor U6876 (N_6876,N_4740,N_3360);
and U6877 (N_6877,N_3854,N_4385);
nand U6878 (N_6878,N_5265,N_4093);
nand U6879 (N_6879,N_4354,N_3248);
nor U6880 (N_6880,N_4575,N_3472);
and U6881 (N_6881,N_3336,N_5285);
nand U6882 (N_6882,N_3759,N_5215);
nor U6883 (N_6883,N_5869,N_4217);
nand U6884 (N_6884,N_4799,N_3964);
xor U6885 (N_6885,N_3641,N_5818);
nand U6886 (N_6886,N_5456,N_5663);
xnor U6887 (N_6887,N_4590,N_5749);
nor U6888 (N_6888,N_5127,N_5189);
nand U6889 (N_6889,N_4960,N_5212);
or U6890 (N_6890,N_5073,N_4662);
or U6891 (N_6891,N_3864,N_5154);
nor U6892 (N_6892,N_3142,N_5245);
nor U6893 (N_6893,N_4962,N_5282);
nand U6894 (N_6894,N_3132,N_4393);
nand U6895 (N_6895,N_4135,N_5632);
nor U6896 (N_6896,N_3778,N_5650);
xor U6897 (N_6897,N_5580,N_4750);
nor U6898 (N_6898,N_4855,N_5742);
nand U6899 (N_6899,N_3176,N_3700);
and U6900 (N_6900,N_4869,N_5680);
or U6901 (N_6901,N_5792,N_5469);
or U6902 (N_6902,N_5535,N_5895);
or U6903 (N_6903,N_3091,N_5989);
nor U6904 (N_6904,N_3880,N_3907);
nand U6905 (N_6905,N_5746,N_4698);
and U6906 (N_6906,N_4332,N_3901);
nor U6907 (N_6907,N_3205,N_4391);
or U6908 (N_6908,N_3685,N_4713);
nor U6909 (N_6909,N_3463,N_4815);
or U6910 (N_6910,N_3992,N_4582);
nand U6911 (N_6911,N_4230,N_4748);
and U6912 (N_6912,N_3873,N_3701);
nand U6913 (N_6913,N_3527,N_4523);
nand U6914 (N_6914,N_3255,N_5911);
nand U6915 (N_6915,N_3370,N_4950);
and U6916 (N_6916,N_3342,N_4775);
nor U6917 (N_6917,N_4779,N_4057);
and U6918 (N_6918,N_5482,N_5120);
or U6919 (N_6919,N_3653,N_5886);
nor U6920 (N_6920,N_5078,N_3947);
nand U6921 (N_6921,N_4851,N_4271);
xnor U6922 (N_6922,N_3740,N_3449);
and U6923 (N_6923,N_5922,N_3474);
and U6924 (N_6924,N_3240,N_3829);
nand U6925 (N_6925,N_5615,N_4079);
or U6926 (N_6926,N_4227,N_4441);
nand U6927 (N_6927,N_4094,N_4890);
or U6928 (N_6928,N_3314,N_3311);
or U6929 (N_6929,N_4978,N_4507);
and U6930 (N_6930,N_4487,N_4862);
or U6931 (N_6931,N_4053,N_4898);
or U6932 (N_6932,N_4512,N_5313);
nand U6933 (N_6933,N_4986,N_5969);
and U6934 (N_6934,N_3593,N_5320);
and U6935 (N_6935,N_4897,N_3220);
and U6936 (N_6936,N_4763,N_4289);
nor U6937 (N_6937,N_3338,N_3950);
nor U6938 (N_6938,N_5581,N_5467);
nor U6939 (N_6939,N_4903,N_3022);
nand U6940 (N_6940,N_5235,N_3101);
nor U6941 (N_6941,N_3839,N_4457);
nor U6942 (N_6942,N_5187,N_4675);
nor U6943 (N_6943,N_5063,N_3621);
nand U6944 (N_6944,N_5638,N_4111);
xnor U6945 (N_6945,N_3343,N_4882);
or U6946 (N_6946,N_4636,N_4899);
nor U6947 (N_6947,N_4179,N_5830);
nand U6948 (N_6948,N_3757,N_3018);
and U6949 (N_6949,N_3652,N_4896);
or U6950 (N_6950,N_4076,N_5964);
nor U6951 (N_6951,N_4187,N_4301);
nand U6952 (N_6952,N_5238,N_5550);
nand U6953 (N_6953,N_4967,N_3319);
nor U6954 (N_6954,N_3094,N_3927);
and U6955 (N_6955,N_3924,N_3914);
xnor U6956 (N_6956,N_3024,N_3210);
and U6957 (N_6957,N_3441,N_3900);
xor U6958 (N_6958,N_3515,N_4777);
or U6959 (N_6959,N_5852,N_4910);
and U6960 (N_6960,N_4043,N_4583);
xnor U6961 (N_6961,N_3955,N_4921);
nor U6962 (N_6962,N_5270,N_4694);
nor U6963 (N_6963,N_4454,N_3036);
or U6964 (N_6964,N_4729,N_3494);
xor U6965 (N_6965,N_5404,N_3458);
nand U6966 (N_6966,N_4310,N_3337);
nor U6967 (N_6967,N_5713,N_3033);
and U6968 (N_6968,N_5144,N_5043);
or U6969 (N_6969,N_3611,N_5952);
xnor U6970 (N_6970,N_4571,N_5328);
nor U6971 (N_6971,N_5009,N_3124);
or U6972 (N_6972,N_4183,N_5363);
nand U6973 (N_6973,N_5369,N_4247);
and U6974 (N_6974,N_5831,N_5339);
and U6975 (N_6975,N_4559,N_3157);
nor U6976 (N_6976,N_3815,N_4504);
or U6977 (N_6977,N_4380,N_4816);
nand U6978 (N_6978,N_3702,N_3321);
or U6979 (N_6979,N_4352,N_4281);
or U6980 (N_6980,N_4257,N_4220);
or U6981 (N_6981,N_3202,N_3480);
nand U6982 (N_6982,N_3223,N_4424);
or U6983 (N_6983,N_5987,N_5465);
nor U6984 (N_6984,N_5619,N_5997);
nor U6985 (N_6985,N_5002,N_3928);
and U6986 (N_6986,N_3938,N_3536);
and U6987 (N_6987,N_5384,N_4494);
nand U6988 (N_6988,N_5096,N_5945);
or U6989 (N_6989,N_3028,N_4198);
nand U6990 (N_6990,N_4175,N_5230);
or U6991 (N_6991,N_4037,N_3383);
and U6992 (N_6992,N_4381,N_4105);
xnor U6993 (N_6993,N_3430,N_5642);
and U6994 (N_6994,N_4468,N_5725);
or U6995 (N_6995,N_4602,N_3746);
nand U6996 (N_6996,N_3544,N_3475);
nand U6997 (N_6997,N_4781,N_3916);
xnor U6998 (N_6998,N_5537,N_3302);
and U6999 (N_6999,N_5260,N_4483);
nor U7000 (N_7000,N_3284,N_5206);
nor U7001 (N_7001,N_4191,N_3939);
nand U7002 (N_7002,N_3055,N_3686);
nand U7003 (N_7003,N_3212,N_3855);
xor U7004 (N_7004,N_5538,N_3525);
nor U7005 (N_7005,N_5062,N_4199);
nor U7006 (N_7006,N_3017,N_4279);
and U7007 (N_7007,N_3764,N_4464);
nor U7008 (N_7008,N_4520,N_5709);
xor U7009 (N_7009,N_4119,N_3491);
nand U7010 (N_7010,N_5381,N_4968);
nand U7011 (N_7011,N_3010,N_3566);
and U7012 (N_7012,N_5248,N_3941);
or U7013 (N_7013,N_5877,N_5982);
nand U7014 (N_7014,N_4364,N_3204);
xnor U7015 (N_7015,N_4841,N_3543);
nand U7016 (N_7016,N_5996,N_4944);
nor U7017 (N_7017,N_5331,N_5986);
or U7018 (N_7018,N_3600,N_3184);
nor U7019 (N_7019,N_4814,N_3587);
nand U7020 (N_7020,N_5801,N_5234);
and U7021 (N_7021,N_4517,N_5247);
nand U7022 (N_7022,N_3082,N_3089);
or U7023 (N_7023,N_5101,N_4850);
or U7024 (N_7024,N_3772,N_4495);
xor U7025 (N_7025,N_3462,N_4476);
or U7026 (N_7026,N_4765,N_4080);
xor U7027 (N_7027,N_5203,N_4123);
and U7028 (N_7028,N_4628,N_5506);
nor U7029 (N_7029,N_4148,N_4652);
nand U7030 (N_7030,N_3376,N_5391);
or U7031 (N_7031,N_5870,N_3107);
or U7032 (N_7032,N_3131,N_3027);
nand U7033 (N_7033,N_3514,N_3044);
nand U7034 (N_7034,N_5436,N_3249);
and U7035 (N_7035,N_3395,N_3747);
nor U7036 (N_7036,N_4406,N_3667);
xor U7037 (N_7037,N_4110,N_3477);
or U7038 (N_7038,N_5505,N_3847);
or U7039 (N_7039,N_3852,N_3151);
or U7040 (N_7040,N_3892,N_3596);
xor U7041 (N_7041,N_4722,N_3675);
nor U7042 (N_7042,N_5943,N_4330);
nand U7043 (N_7043,N_5777,N_5357);
nand U7044 (N_7044,N_5254,N_5741);
and U7045 (N_7045,N_3646,N_4288);
nor U7046 (N_7046,N_4830,N_3658);
xnor U7047 (N_7047,N_4501,N_4414);
or U7048 (N_7048,N_3421,N_4831);
or U7049 (N_7049,N_3348,N_3504);
and U7050 (N_7050,N_5221,N_4224);
or U7051 (N_7051,N_3369,N_4821);
or U7052 (N_7052,N_4308,N_5319);
or U7053 (N_7053,N_4955,N_4892);
or U7054 (N_7054,N_4026,N_4762);
nor U7055 (N_7055,N_5732,N_4480);
nand U7056 (N_7056,N_4640,N_4994);
or U7057 (N_7057,N_4592,N_4190);
and U7058 (N_7058,N_3127,N_4638);
and U7059 (N_7059,N_5966,N_3844);
xnor U7060 (N_7060,N_5561,N_5433);
xor U7061 (N_7061,N_3083,N_4168);
nor U7062 (N_7062,N_3661,N_3896);
nand U7063 (N_7063,N_3483,N_3835);
and U7064 (N_7064,N_4619,N_4447);
and U7065 (N_7065,N_5738,N_4395);
and U7066 (N_7066,N_5115,N_3579);
and U7067 (N_7067,N_4328,N_3085);
or U7068 (N_7068,N_5914,N_4438);
and U7069 (N_7069,N_3221,N_4496);
nor U7070 (N_7070,N_5977,N_4912);
nor U7071 (N_7071,N_3358,N_4208);
nor U7072 (N_7072,N_4492,N_4558);
nor U7073 (N_7073,N_4957,N_5514);
nor U7074 (N_7074,N_5978,N_4879);
nand U7075 (N_7075,N_4097,N_4581);
or U7076 (N_7076,N_4443,N_5293);
xor U7077 (N_7077,N_5171,N_5585);
and U7078 (N_7078,N_3006,N_3572);
xnor U7079 (N_7079,N_4319,N_4680);
xor U7080 (N_7080,N_3694,N_5829);
nor U7081 (N_7081,N_5858,N_3190);
or U7082 (N_7082,N_4398,N_3707);
nand U7083 (N_7083,N_4016,N_4207);
nor U7084 (N_7084,N_5016,N_4887);
nor U7085 (N_7085,N_3296,N_3867);
nand U7086 (N_7086,N_5764,N_4412);
and U7087 (N_7087,N_5857,N_3978);
and U7088 (N_7088,N_5508,N_3456);
nand U7089 (N_7089,N_5579,N_4937);
nand U7090 (N_7090,N_5872,N_4068);
and U7091 (N_7091,N_4342,N_4295);
or U7092 (N_7092,N_4325,N_5820);
or U7093 (N_7093,N_4545,N_5236);
or U7094 (N_7094,N_5586,N_5333);
and U7095 (N_7095,N_3126,N_3481);
nor U7096 (N_7096,N_3073,N_3488);
nor U7097 (N_7097,N_4811,N_5612);
and U7098 (N_7098,N_4857,N_3931);
nand U7099 (N_7099,N_4943,N_4375);
xnor U7100 (N_7100,N_3378,N_3528);
and U7101 (N_7101,N_4065,N_4954);
or U7102 (N_7102,N_5420,N_3079);
or U7103 (N_7103,N_5488,N_3396);
nand U7104 (N_7104,N_5963,N_5220);
nor U7105 (N_7105,N_3567,N_4082);
nor U7106 (N_7106,N_4427,N_5486);
or U7107 (N_7107,N_4283,N_5644);
nor U7108 (N_7108,N_3541,N_3292);
or U7109 (N_7109,N_4692,N_4172);
nor U7110 (N_7110,N_5753,N_4667);
and U7111 (N_7111,N_4611,N_3736);
nor U7112 (N_7112,N_3594,N_3273);
nand U7113 (N_7113,N_5856,N_3256);
nand U7114 (N_7114,N_5387,N_4205);
nand U7115 (N_7115,N_3065,N_3259);
nand U7116 (N_7116,N_5864,N_3346);
and U7117 (N_7117,N_5898,N_3335);
nor U7118 (N_7118,N_5330,N_5893);
xor U7119 (N_7119,N_3173,N_4676);
xor U7120 (N_7120,N_3801,N_5370);
xnor U7121 (N_7121,N_5402,N_5481);
or U7122 (N_7122,N_4136,N_5056);
or U7123 (N_7123,N_5301,N_4622);
nor U7124 (N_7124,N_3105,N_5932);
or U7125 (N_7125,N_4059,N_3809);
xnor U7126 (N_7126,N_4665,N_5688);
nand U7127 (N_7127,N_5067,N_4616);
nand U7128 (N_7128,N_4564,N_3793);
and U7129 (N_7129,N_3163,N_5492);
nand U7130 (N_7130,N_3812,N_4471);
and U7131 (N_7131,N_3990,N_4600);
nor U7132 (N_7132,N_3268,N_5699);
nand U7133 (N_7133,N_3838,N_3532);
and U7134 (N_7134,N_5329,N_5462);
or U7135 (N_7135,N_5598,N_3473);
nand U7136 (N_7136,N_4551,N_4529);
or U7137 (N_7137,N_3026,N_4635);
nor U7138 (N_7138,N_3926,N_5423);
nor U7139 (N_7139,N_5170,N_5058);
nor U7140 (N_7140,N_5116,N_5110);
xnor U7141 (N_7141,N_3004,N_4871);
nor U7142 (N_7142,N_5082,N_4039);
nand U7143 (N_7143,N_5756,N_4466);
nor U7144 (N_7144,N_3850,N_3627);
nand U7145 (N_7145,N_5951,N_5780);
nand U7146 (N_7146,N_5306,N_4133);
and U7147 (N_7147,N_5589,N_4953);
xor U7148 (N_7148,N_4824,N_3729);
or U7149 (N_7149,N_3186,N_5274);
nand U7150 (N_7150,N_3796,N_3359);
or U7151 (N_7151,N_4128,N_3640);
and U7152 (N_7152,N_3516,N_4601);
nor U7153 (N_7153,N_5102,N_3422);
nand U7154 (N_7154,N_4344,N_4335);
xnor U7155 (N_7155,N_5842,N_4516);
and U7156 (N_7156,N_3141,N_3777);
nand U7157 (N_7157,N_3112,N_3769);
or U7158 (N_7158,N_5164,N_4778);
and U7159 (N_7159,N_4767,N_4596);
nor U7160 (N_7160,N_5349,N_4510);
and U7161 (N_7161,N_5014,N_5364);
or U7162 (N_7162,N_4621,N_3148);
xnor U7163 (N_7163,N_4029,N_3783);
nand U7164 (N_7164,N_4033,N_4156);
nor U7165 (N_7165,N_5197,N_3219);
nand U7166 (N_7166,N_5890,N_5904);
nor U7167 (N_7167,N_4997,N_5483);
or U7168 (N_7168,N_4359,N_5519);
or U7169 (N_7169,N_5593,N_4434);
xor U7170 (N_7170,N_3271,N_3762);
nand U7171 (N_7171,N_3410,N_5131);
and U7172 (N_7172,N_4701,N_5477);
nor U7173 (N_7173,N_3831,N_3857);
or U7174 (N_7174,N_4124,N_5668);
and U7175 (N_7175,N_3371,N_3557);
nand U7176 (N_7176,N_3459,N_4417);
or U7177 (N_7177,N_5629,N_5671);
or U7178 (N_7178,N_4028,N_3003);
or U7179 (N_7179,N_3622,N_3699);
nand U7180 (N_7180,N_4612,N_4789);
nor U7181 (N_7181,N_5435,N_4186);
and U7182 (N_7182,N_5692,N_4138);
or U7183 (N_7183,N_5094,N_5398);
or U7184 (N_7184,N_4792,N_4255);
nor U7185 (N_7185,N_5597,N_4329);
or U7186 (N_7186,N_3139,N_3122);
nor U7187 (N_7187,N_3162,N_3020);
xor U7188 (N_7188,N_4877,N_3905);
or U7189 (N_7189,N_5027,N_4334);
or U7190 (N_7190,N_4935,N_4386);
nand U7191 (N_7191,N_5518,N_3840);
and U7192 (N_7192,N_4223,N_5000);
and U7193 (N_7193,N_3698,N_5717);
nand U7194 (N_7194,N_3390,N_3967);
and U7195 (N_7195,N_3696,N_3828);
nand U7196 (N_7196,N_5437,N_3482);
xnor U7197 (N_7197,N_4368,N_4373);
nor U7198 (N_7198,N_4020,N_3940);
nor U7199 (N_7199,N_5917,N_3040);
or U7200 (N_7200,N_4339,N_4345);
or U7201 (N_7201,N_3742,N_5003);
and U7202 (N_7202,N_3283,N_4040);
nand U7203 (N_7203,N_5249,N_4853);
or U7204 (N_7204,N_5273,N_4613);
and U7205 (N_7205,N_4087,N_3755);
and U7206 (N_7206,N_3499,N_3971);
or U7207 (N_7207,N_3417,N_3756);
nand U7208 (N_7208,N_4184,N_5656);
nor U7209 (N_7209,N_3606,N_4113);
and U7210 (N_7210,N_4743,N_4051);
or U7211 (N_7211,N_4425,N_4934);
nand U7212 (N_7212,N_3523,N_4895);
nor U7213 (N_7213,N_5534,N_5560);
nor U7214 (N_7214,N_4320,N_4465);
or U7215 (N_7215,N_3570,N_5763);
xnor U7216 (N_7216,N_4744,N_3697);
nand U7217 (N_7217,N_5205,N_4195);
or U7218 (N_7218,N_3760,N_4266);
nor U7219 (N_7219,N_3104,N_5004);
and U7220 (N_7220,N_5614,N_4203);
or U7221 (N_7221,N_3874,N_3333);
nor U7222 (N_7222,N_5967,N_5531);
and U7223 (N_7223,N_3856,N_3245);
or U7224 (N_7224,N_4946,N_3464);
nor U7225 (N_7225,N_5173,N_3466);
or U7226 (N_7226,N_3156,N_4158);
nor U7227 (N_7227,N_4189,N_3858);
and U7228 (N_7228,N_4177,N_4754);
or U7229 (N_7229,N_5337,N_4074);
nor U7230 (N_7230,N_5066,N_5061);
xnor U7231 (N_7231,N_5403,N_4349);
nor U7232 (N_7232,N_5037,N_3727);
xor U7233 (N_7233,N_3986,N_5158);
nor U7234 (N_7234,N_4731,N_3655);
nand U7235 (N_7235,N_5046,N_3134);
or U7236 (N_7236,N_3217,N_3962);
nand U7237 (N_7237,N_5784,N_3960);
nand U7238 (N_7238,N_3753,N_3397);
nor U7239 (N_7239,N_3057,N_5414);
and U7240 (N_7240,N_3592,N_5839);
xnor U7241 (N_7241,N_5268,N_5278);
nand U7242 (N_7242,N_4985,N_4035);
nor U7243 (N_7243,N_5366,N_5582);
nor U7244 (N_7244,N_4772,N_4833);
and U7245 (N_7245,N_3258,N_4165);
nand U7246 (N_7246,N_4931,N_5390);
nand U7247 (N_7247,N_5324,N_5302);
or U7248 (N_7248,N_5072,N_4591);
or U7249 (N_7249,N_3230,N_3519);
and U7250 (N_7250,N_5229,N_5198);
nand U7251 (N_7251,N_3254,N_4577);
nor U7252 (N_7252,N_4405,N_4544);
xor U7253 (N_7253,N_3102,N_5200);
nand U7254 (N_7254,N_5530,N_3957);
xnor U7255 (N_7255,N_4976,N_5161);
nor U7256 (N_7256,N_5811,N_4521);
and U7257 (N_7257,N_3575,N_3056);
nor U7258 (N_7258,N_5718,N_5256);
and U7259 (N_7259,N_4782,N_3899);
nor U7260 (N_7260,N_3861,N_3788);
xnor U7261 (N_7261,N_3227,N_4632);
or U7262 (N_7262,N_3984,N_5406);
or U7263 (N_7263,N_3001,N_3144);
nor U7264 (N_7264,N_5915,N_4651);
and U7265 (N_7265,N_4626,N_3530);
and U7266 (N_7266,N_4008,N_3586);
and U7267 (N_7267,N_3090,N_5515);
nor U7268 (N_7268,N_3615,N_3969);
or U7269 (N_7269,N_4553,N_5017);
nand U7270 (N_7270,N_3432,N_4106);
nor U7271 (N_7271,N_5616,N_4362);
xor U7272 (N_7272,N_4959,N_5880);
nor U7273 (N_7273,N_4990,N_4813);
or U7274 (N_7274,N_4671,N_4786);
nor U7275 (N_7275,N_4573,N_3684);
and U7276 (N_7276,N_4173,N_4456);
or U7277 (N_7277,N_3446,N_3031);
or U7278 (N_7278,N_5859,N_4653);
nand U7279 (N_7279,N_3638,N_4155);
nor U7280 (N_7280,N_4929,N_4818);
or U7281 (N_7281,N_4716,N_5118);
or U7282 (N_7282,N_3469,N_5837);
and U7283 (N_7283,N_5779,N_4739);
nand U7284 (N_7284,N_5640,N_5135);
and U7285 (N_7285,N_3884,N_5563);
or U7286 (N_7286,N_5291,N_3392);
nor U7287 (N_7287,N_4472,N_4107);
and U7288 (N_7288,N_4570,N_3936);
and U7289 (N_7289,N_4455,N_3306);
nand U7290 (N_7290,N_4666,N_4394);
and U7291 (N_7291,N_5927,N_5448);
xor U7292 (N_7292,N_3278,N_4585);
nand U7293 (N_7293,N_5755,N_4825);
nand U7294 (N_7294,N_4403,N_5798);
and U7295 (N_7295,N_3380,N_5926);
and U7296 (N_7296,N_4001,N_4134);
or U7297 (N_7297,N_3890,N_5039);
nand U7298 (N_7298,N_3429,N_5854);
nand U7299 (N_7299,N_4318,N_5129);
nor U7300 (N_7300,N_3692,N_5925);
nor U7301 (N_7301,N_5426,N_3966);
xor U7302 (N_7302,N_3859,N_3862);
and U7303 (N_7303,N_4462,N_3513);
or U7304 (N_7304,N_3977,N_4431);
or U7305 (N_7305,N_5281,N_5641);
xnor U7306 (N_7306,N_4856,N_4104);
or U7307 (N_7307,N_3096,N_4909);
nand U7308 (N_7308,N_5005,N_5251);
and U7309 (N_7309,N_5575,N_5983);
and U7310 (N_7310,N_4246,N_4372);
and U7311 (N_7311,N_5929,N_5365);
nand U7312 (N_7312,N_4096,N_4576);
nand U7313 (N_7313,N_4794,N_4278);
or U7314 (N_7314,N_4038,N_4481);
xor U7315 (N_7315,N_5716,N_5006);
nor U7316 (N_7316,N_4239,N_4737);
nand U7317 (N_7317,N_5630,N_4384);
and U7318 (N_7318,N_3789,N_4980);
nand U7319 (N_7319,N_4250,N_3670);
nand U7320 (N_7320,N_3954,N_5266);
nor U7321 (N_7321,N_3804,N_4685);
xor U7322 (N_7322,N_5114,N_4548);
and U7323 (N_7323,N_3442,N_3545);
and U7324 (N_7324,N_3490,N_5345);
nand U7325 (N_7325,N_3893,N_5609);
nor U7326 (N_7326,N_4151,N_4221);
nor U7327 (N_7327,N_3569,N_5442);
xor U7328 (N_7328,N_3398,N_3409);
and U7329 (N_7329,N_4747,N_4194);
or U7330 (N_7330,N_4867,N_3451);
xnor U7331 (N_7331,N_5142,N_3068);
nand U7332 (N_7332,N_3386,N_4687);
nand U7333 (N_7333,N_3559,N_5796);
nor U7334 (N_7334,N_4913,N_5476);
or U7335 (N_7335,N_3362,N_5466);
and U7336 (N_7336,N_4459,N_3324);
nand U7337 (N_7337,N_4805,N_5968);
nor U7338 (N_7338,N_5439,N_4485);
nand U7339 (N_7339,N_3792,N_3853);
nor U7340 (N_7340,N_3286,N_3214);
or U7341 (N_7341,N_5377,N_4085);
and U7342 (N_7342,N_4819,N_5810);
xnor U7343 (N_7343,N_4531,N_3452);
and U7344 (N_7344,N_5323,N_5637);
or U7345 (N_7345,N_5081,N_5744);
nand U7346 (N_7346,N_5860,N_3672);
and U7347 (N_7347,N_5923,N_5451);
xor U7348 (N_7348,N_3485,N_3299);
or U7349 (N_7349,N_3088,N_4941);
and U7350 (N_7350,N_3949,N_4185);
and U7351 (N_7351,N_5992,N_4439);
xor U7352 (N_7352,N_3773,N_3752);
and U7353 (N_7353,N_3933,N_4442);
nor U7354 (N_7354,N_3032,N_3770);
or U7355 (N_7355,N_5834,N_5148);
nor U7356 (N_7356,N_4304,N_5427);
or U7357 (N_7357,N_4880,N_4452);
nand U7358 (N_7358,N_5845,N_5214);
nand U7359 (N_7359,N_3571,N_4569);
nor U7360 (N_7360,N_3739,N_3339);
nor U7361 (N_7361,N_5604,N_4549);
and U7362 (N_7362,N_4938,N_4428);
nor U7363 (N_7363,N_5590,N_4125);
nor U7364 (N_7364,N_3591,N_4560);
nor U7365 (N_7365,N_3427,N_3416);
or U7366 (N_7366,N_4832,N_5159);
xor U7367 (N_7367,N_5673,N_3639);
xnor U7368 (N_7368,N_4557,N_5299);
or U7369 (N_7369,N_3394,N_5734);
and U7370 (N_7370,N_3285,N_3304);
nor U7371 (N_7371,N_4408,N_4527);
and U7372 (N_7372,N_4421,N_4670);
nor U7373 (N_7373,N_4206,N_4262);
nor U7374 (N_7374,N_4095,N_5874);
nand U7375 (N_7375,N_4193,N_3676);
and U7376 (N_7376,N_4525,N_3201);
nand U7377 (N_7377,N_4064,N_4285);
nor U7378 (N_7378,N_5165,N_5793);
nor U7379 (N_7379,N_3795,N_4541);
xnor U7380 (N_7380,N_4287,N_4149);
or U7381 (N_7381,N_3608,N_5149);
and U7382 (N_7382,N_3200,N_4606);
xor U7383 (N_7383,N_5685,N_4756);
or U7384 (N_7384,N_5036,N_3307);
or U7385 (N_7385,N_4286,N_5011);
nand U7386 (N_7386,N_5938,N_3401);
nand U7387 (N_7387,N_3476,N_5950);
nor U7388 (N_7388,N_4396,N_4915);
nor U7389 (N_7389,N_5797,N_4589);
and U7390 (N_7390,N_5191,N_5294);
or U7391 (N_7391,N_4088,N_4200);
nor U7392 (N_7392,N_4870,N_5840);
nand U7393 (N_7393,N_5553,N_5931);
xnor U7394 (N_7394,N_5920,N_5665);
and U7395 (N_7395,N_5568,N_3505);
or U7396 (N_7396,N_4062,N_4003);
xor U7397 (N_7397,N_5583,N_3174);
or U7398 (N_7398,N_3385,N_5376);
or U7399 (N_7399,N_4488,N_4292);
nor U7400 (N_7400,N_3865,N_5079);
and U7401 (N_7401,N_5507,N_3312);
xnor U7402 (N_7402,N_5933,N_3460);
nor U7403 (N_7403,N_3193,N_5802);
or U7404 (N_7404,N_3803,N_3710);
or U7405 (N_7405,N_5679,N_4196);
xor U7406 (N_7406,N_3576,N_5754);
and U7407 (N_7407,N_4963,N_3015);
xor U7408 (N_7408,N_5332,N_3908);
xnor U7409 (N_7409,N_4253,N_5141);
xor U7410 (N_7410,N_3894,N_5708);
xor U7411 (N_7411,N_4886,N_3149);
nand U7412 (N_7412,N_4881,N_5098);
and U7413 (N_7413,N_5429,N_3066);
or U7414 (N_7414,N_3478,N_3411);
or U7415 (N_7415,N_4241,N_4399);
or U7416 (N_7416,N_3109,N_5351);
or U7417 (N_7417,N_3765,N_3350);
xnor U7418 (N_7418,N_4453,N_4649);
nand U7419 (N_7419,N_4714,N_5259);
nand U7420 (N_7420,N_5444,N_3531);
xor U7421 (N_7421,N_5657,N_3118);
or U7422 (N_7422,N_5322,N_3140);
nand U7423 (N_7423,N_5401,N_4102);
and U7424 (N_7424,N_4254,N_5346);
nand U7425 (N_7425,N_5703,N_5202);
or U7426 (N_7426,N_5244,N_3774);
or U7427 (N_7427,N_3435,N_4475);
nand U7428 (N_7428,N_4477,N_3135);
and U7429 (N_7429,N_5318,N_4070);
nor U7430 (N_7430,N_5054,N_4812);
and U7431 (N_7431,N_3185,N_5613);
nor U7432 (N_7432,N_4865,N_3878);
or U7433 (N_7433,N_5587,N_5474);
nand U7434 (N_7434,N_4565,N_3074);
and U7435 (N_7435,N_4715,N_3589);
nor U7436 (N_7436,N_3039,N_3153);
nor U7437 (N_7437,N_5340,N_3413);
nand U7438 (N_7438,N_3549,N_3183);
nor U7439 (N_7439,N_5899,N_4542);
xnor U7440 (N_7440,N_4013,N_5405);
nor U7441 (N_7441,N_5791,N_5057);
and U7442 (N_7442,N_4351,N_5940);
xnor U7443 (N_7443,N_5396,N_3297);
xor U7444 (N_7444,N_3660,N_3568);
nand U7445 (N_7445,N_4925,N_5373);
and U7446 (N_7446,N_3946,N_3704);
and U7447 (N_7447,N_3533,N_4911);
nand U7448 (N_7448,N_3805,N_4201);
nor U7449 (N_7449,N_3518,N_3133);
and U7450 (N_7450,N_4389,N_4726);
nor U7451 (N_7451,N_4245,N_4721);
nor U7452 (N_7452,N_4533,N_3120);
and U7453 (N_7453,N_5624,N_4430);
nor U7454 (N_7454,N_5881,N_4423);
and U7455 (N_7455,N_4161,N_4681);
nor U7456 (N_7456,N_5998,N_3822);
or U7457 (N_7457,N_5941,N_5233);
nand U7458 (N_7458,N_3631,N_5443);
xnor U7459 (N_7459,N_5287,N_5591);
nor U7460 (N_7460,N_4684,N_5770);
or U7461 (N_7461,N_4235,N_5422);
xnor U7462 (N_7462,N_5813,N_5107);
nor U7463 (N_7463,N_4237,N_3550);
and U7464 (N_7464,N_5425,N_5099);
and U7465 (N_7465,N_5316,N_5065);
nand U7466 (N_7466,N_3797,N_4787);
or U7467 (N_7467,N_5702,N_5279);
and U7468 (N_7468,N_4752,N_4530);
nor U7469 (N_7469,N_4031,N_5981);
xnor U7470 (N_7470,N_4132,N_5578);
and U7471 (N_7471,N_5446,N_3489);
and U7472 (N_7472,N_4353,N_3486);
nor U7473 (N_7473,N_4436,N_5551);
nand U7474 (N_7474,N_4163,N_5257);
and U7475 (N_7475,N_4277,N_3372);
nor U7476 (N_7476,N_4508,N_5022);
nor U7477 (N_7477,N_3555,N_5660);
and U7478 (N_7478,N_5910,N_5540);
or U7479 (N_7479,N_4660,N_4432);
nor U7480 (N_7480,N_3189,N_4358);
and U7481 (N_7481,N_5155,N_5453);
nor U7482 (N_7482,N_4060,N_4182);
or U7483 (N_7483,N_5662,N_4630);
or U7484 (N_7484,N_3816,N_5473);
nor U7485 (N_7485,N_5715,N_5147);
and U7486 (N_7486,N_4579,N_3198);
nand U7487 (N_7487,N_4435,N_3758);
or U7488 (N_7488,N_3666,N_4550);
nand U7489 (N_7489,N_5944,N_3529);
nor U7490 (N_7490,N_3081,N_3909);
nand U7491 (N_7491,N_4972,N_5378);
and U7492 (N_7492,N_3948,N_4741);
nand U7493 (N_7493,N_5994,N_5954);
xnor U7494 (N_7494,N_4090,N_5150);
nand U7495 (N_7495,N_3846,N_5736);
or U7496 (N_7496,N_3780,N_5354);
and U7497 (N_7497,N_3743,N_5168);
or U7498 (N_7498,N_4696,N_4197);
xnor U7499 (N_7499,N_4826,N_5156);
and U7500 (N_7500,N_5022,N_4614);
nand U7501 (N_7501,N_4123,N_3076);
and U7502 (N_7502,N_5813,N_4623);
and U7503 (N_7503,N_4091,N_3210);
nand U7504 (N_7504,N_3715,N_4766);
and U7505 (N_7505,N_5126,N_4348);
or U7506 (N_7506,N_4566,N_3573);
nand U7507 (N_7507,N_4141,N_5767);
nor U7508 (N_7508,N_5545,N_5223);
nand U7509 (N_7509,N_4838,N_3633);
or U7510 (N_7510,N_5485,N_4063);
and U7511 (N_7511,N_4360,N_3374);
nand U7512 (N_7512,N_3660,N_4494);
nor U7513 (N_7513,N_5401,N_4230);
or U7514 (N_7514,N_4979,N_4665);
and U7515 (N_7515,N_4403,N_3107);
nand U7516 (N_7516,N_3154,N_3461);
and U7517 (N_7517,N_5804,N_5486);
nor U7518 (N_7518,N_4932,N_3160);
or U7519 (N_7519,N_4082,N_5952);
nor U7520 (N_7520,N_3152,N_4236);
nor U7521 (N_7521,N_4244,N_5899);
or U7522 (N_7522,N_3048,N_5126);
nand U7523 (N_7523,N_4926,N_4734);
or U7524 (N_7524,N_3579,N_5548);
xnor U7525 (N_7525,N_3374,N_5129);
or U7526 (N_7526,N_4464,N_3241);
or U7527 (N_7527,N_4009,N_4053);
nor U7528 (N_7528,N_5265,N_4602);
nand U7529 (N_7529,N_3411,N_4084);
nand U7530 (N_7530,N_3213,N_3098);
nor U7531 (N_7531,N_3983,N_3606);
nor U7532 (N_7532,N_3647,N_3255);
nor U7533 (N_7533,N_3190,N_3987);
xor U7534 (N_7534,N_3290,N_4801);
or U7535 (N_7535,N_5024,N_4962);
or U7536 (N_7536,N_3771,N_4047);
nand U7537 (N_7537,N_5991,N_4654);
nand U7538 (N_7538,N_3461,N_3690);
or U7539 (N_7539,N_5884,N_3952);
or U7540 (N_7540,N_5083,N_5353);
or U7541 (N_7541,N_4575,N_4071);
xnor U7542 (N_7542,N_4685,N_3538);
or U7543 (N_7543,N_4075,N_5958);
nand U7544 (N_7544,N_3894,N_4492);
nand U7545 (N_7545,N_3944,N_5754);
nor U7546 (N_7546,N_3864,N_3823);
nand U7547 (N_7547,N_3544,N_4053);
or U7548 (N_7548,N_3501,N_5857);
or U7549 (N_7549,N_4560,N_3070);
and U7550 (N_7550,N_3813,N_3407);
xor U7551 (N_7551,N_5139,N_4027);
or U7552 (N_7552,N_3556,N_5911);
and U7553 (N_7553,N_5351,N_5730);
nand U7554 (N_7554,N_5566,N_5430);
nor U7555 (N_7555,N_3790,N_5975);
or U7556 (N_7556,N_5745,N_5661);
nand U7557 (N_7557,N_3152,N_5739);
nor U7558 (N_7558,N_5540,N_5431);
and U7559 (N_7559,N_5731,N_4835);
and U7560 (N_7560,N_4571,N_5426);
nand U7561 (N_7561,N_4290,N_4064);
and U7562 (N_7562,N_5490,N_5752);
nor U7563 (N_7563,N_3501,N_4134);
nor U7564 (N_7564,N_5437,N_3080);
and U7565 (N_7565,N_4036,N_3441);
or U7566 (N_7566,N_3317,N_5702);
nor U7567 (N_7567,N_5596,N_5912);
nor U7568 (N_7568,N_3822,N_3046);
nand U7569 (N_7569,N_5768,N_4567);
xnor U7570 (N_7570,N_4691,N_5774);
and U7571 (N_7571,N_3349,N_4799);
nor U7572 (N_7572,N_4686,N_3972);
or U7573 (N_7573,N_5398,N_4632);
and U7574 (N_7574,N_3224,N_4344);
and U7575 (N_7575,N_4873,N_4794);
or U7576 (N_7576,N_5448,N_3458);
and U7577 (N_7577,N_5984,N_5430);
and U7578 (N_7578,N_5380,N_5309);
and U7579 (N_7579,N_4233,N_5020);
nor U7580 (N_7580,N_3640,N_5965);
or U7581 (N_7581,N_5324,N_3379);
or U7582 (N_7582,N_4343,N_3318);
nand U7583 (N_7583,N_4864,N_3424);
nor U7584 (N_7584,N_4703,N_3464);
or U7585 (N_7585,N_5497,N_5679);
nor U7586 (N_7586,N_5250,N_5785);
nor U7587 (N_7587,N_5552,N_3406);
nand U7588 (N_7588,N_5630,N_4939);
xor U7589 (N_7589,N_5606,N_5324);
and U7590 (N_7590,N_3766,N_3341);
nand U7591 (N_7591,N_5942,N_3293);
nand U7592 (N_7592,N_3021,N_5297);
and U7593 (N_7593,N_3512,N_4854);
and U7594 (N_7594,N_4510,N_4484);
and U7595 (N_7595,N_5327,N_5824);
and U7596 (N_7596,N_5039,N_4237);
or U7597 (N_7597,N_4467,N_3011);
nor U7598 (N_7598,N_3346,N_4527);
xor U7599 (N_7599,N_4015,N_3719);
nand U7600 (N_7600,N_3591,N_3363);
nor U7601 (N_7601,N_5618,N_3470);
and U7602 (N_7602,N_3800,N_5319);
nor U7603 (N_7603,N_3006,N_5583);
nand U7604 (N_7604,N_4819,N_3415);
nor U7605 (N_7605,N_4249,N_4420);
or U7606 (N_7606,N_5655,N_3299);
or U7607 (N_7607,N_4803,N_5807);
nand U7608 (N_7608,N_4983,N_5450);
nand U7609 (N_7609,N_3427,N_4233);
xnor U7610 (N_7610,N_5314,N_5730);
nand U7611 (N_7611,N_3269,N_5260);
and U7612 (N_7612,N_5158,N_5758);
nor U7613 (N_7613,N_3169,N_5553);
nor U7614 (N_7614,N_3301,N_5225);
nand U7615 (N_7615,N_3762,N_3274);
nand U7616 (N_7616,N_4292,N_4256);
nor U7617 (N_7617,N_3288,N_5997);
nand U7618 (N_7618,N_5079,N_5277);
nor U7619 (N_7619,N_5231,N_3139);
xor U7620 (N_7620,N_5962,N_3835);
xor U7621 (N_7621,N_5244,N_5205);
nor U7622 (N_7622,N_5538,N_5407);
nor U7623 (N_7623,N_3151,N_4421);
nand U7624 (N_7624,N_4618,N_3752);
and U7625 (N_7625,N_4223,N_3281);
and U7626 (N_7626,N_3432,N_5146);
or U7627 (N_7627,N_3752,N_4157);
nor U7628 (N_7628,N_5276,N_3978);
and U7629 (N_7629,N_4310,N_3833);
or U7630 (N_7630,N_5813,N_5044);
nand U7631 (N_7631,N_4161,N_3507);
nand U7632 (N_7632,N_4306,N_5085);
nand U7633 (N_7633,N_3094,N_4013);
nor U7634 (N_7634,N_5099,N_5320);
or U7635 (N_7635,N_5752,N_5061);
nand U7636 (N_7636,N_5295,N_4909);
nor U7637 (N_7637,N_4485,N_3929);
nor U7638 (N_7638,N_4579,N_5544);
nand U7639 (N_7639,N_3786,N_5810);
nor U7640 (N_7640,N_5860,N_3050);
nand U7641 (N_7641,N_5510,N_5184);
nand U7642 (N_7642,N_3582,N_3616);
xnor U7643 (N_7643,N_3436,N_3023);
xnor U7644 (N_7644,N_3286,N_3038);
or U7645 (N_7645,N_5305,N_4811);
or U7646 (N_7646,N_3520,N_5981);
nor U7647 (N_7647,N_4221,N_4296);
and U7648 (N_7648,N_4006,N_4083);
and U7649 (N_7649,N_5622,N_4420);
nand U7650 (N_7650,N_5197,N_5790);
nor U7651 (N_7651,N_3234,N_4032);
nor U7652 (N_7652,N_3109,N_5924);
and U7653 (N_7653,N_5851,N_4210);
nor U7654 (N_7654,N_5902,N_3032);
nor U7655 (N_7655,N_5223,N_3159);
nand U7656 (N_7656,N_5077,N_4698);
or U7657 (N_7657,N_3310,N_5894);
nand U7658 (N_7658,N_3163,N_3388);
and U7659 (N_7659,N_5856,N_5374);
and U7660 (N_7660,N_4587,N_5455);
nand U7661 (N_7661,N_5271,N_5182);
or U7662 (N_7662,N_4805,N_4271);
and U7663 (N_7663,N_4860,N_5235);
and U7664 (N_7664,N_4343,N_4312);
or U7665 (N_7665,N_5340,N_4049);
nand U7666 (N_7666,N_4646,N_5859);
or U7667 (N_7667,N_4458,N_4843);
or U7668 (N_7668,N_4216,N_5592);
or U7669 (N_7669,N_5403,N_4992);
or U7670 (N_7670,N_3467,N_3697);
xnor U7671 (N_7671,N_4625,N_4372);
and U7672 (N_7672,N_3340,N_4341);
and U7673 (N_7673,N_5177,N_5376);
nand U7674 (N_7674,N_3284,N_3933);
nand U7675 (N_7675,N_4064,N_5246);
and U7676 (N_7676,N_5941,N_3177);
or U7677 (N_7677,N_5932,N_4828);
and U7678 (N_7678,N_3066,N_5733);
or U7679 (N_7679,N_3931,N_4210);
nand U7680 (N_7680,N_4570,N_5546);
nand U7681 (N_7681,N_3638,N_5434);
nand U7682 (N_7682,N_4510,N_3804);
or U7683 (N_7683,N_3507,N_5924);
or U7684 (N_7684,N_3109,N_5363);
or U7685 (N_7685,N_5602,N_5516);
and U7686 (N_7686,N_5848,N_3613);
nor U7687 (N_7687,N_4329,N_3489);
or U7688 (N_7688,N_5096,N_5754);
nor U7689 (N_7689,N_3648,N_5627);
or U7690 (N_7690,N_3829,N_5396);
and U7691 (N_7691,N_3885,N_4248);
and U7692 (N_7692,N_5304,N_5108);
nand U7693 (N_7693,N_4298,N_4642);
nor U7694 (N_7694,N_5981,N_3302);
nand U7695 (N_7695,N_4119,N_3419);
nand U7696 (N_7696,N_5344,N_4778);
nor U7697 (N_7697,N_5116,N_4221);
or U7698 (N_7698,N_3094,N_4732);
nand U7699 (N_7699,N_4225,N_5331);
or U7700 (N_7700,N_5024,N_3336);
nor U7701 (N_7701,N_3161,N_3879);
or U7702 (N_7702,N_3056,N_5760);
or U7703 (N_7703,N_5032,N_5891);
and U7704 (N_7704,N_5607,N_4667);
or U7705 (N_7705,N_4686,N_3495);
nor U7706 (N_7706,N_4077,N_4324);
nand U7707 (N_7707,N_4791,N_3899);
and U7708 (N_7708,N_4723,N_3695);
or U7709 (N_7709,N_3931,N_4377);
nor U7710 (N_7710,N_4766,N_5369);
or U7711 (N_7711,N_5309,N_3240);
or U7712 (N_7712,N_3056,N_4207);
xnor U7713 (N_7713,N_4428,N_4825);
nor U7714 (N_7714,N_4280,N_3055);
nor U7715 (N_7715,N_3866,N_5060);
or U7716 (N_7716,N_5630,N_3047);
and U7717 (N_7717,N_5568,N_4362);
nand U7718 (N_7718,N_5644,N_4841);
or U7719 (N_7719,N_5219,N_4853);
nor U7720 (N_7720,N_3643,N_3554);
or U7721 (N_7721,N_5561,N_3936);
nor U7722 (N_7722,N_4424,N_3636);
nor U7723 (N_7723,N_3115,N_3176);
nand U7724 (N_7724,N_5156,N_3728);
nor U7725 (N_7725,N_3023,N_3803);
and U7726 (N_7726,N_3551,N_4544);
nor U7727 (N_7727,N_3260,N_4356);
nand U7728 (N_7728,N_5562,N_4927);
nor U7729 (N_7729,N_4784,N_3498);
nand U7730 (N_7730,N_4501,N_3481);
and U7731 (N_7731,N_5939,N_3825);
xnor U7732 (N_7732,N_4189,N_4413);
and U7733 (N_7733,N_4296,N_5775);
nor U7734 (N_7734,N_4080,N_4719);
nor U7735 (N_7735,N_4127,N_3812);
nor U7736 (N_7736,N_4892,N_5663);
nand U7737 (N_7737,N_4895,N_5570);
nand U7738 (N_7738,N_4085,N_3942);
and U7739 (N_7739,N_3928,N_5712);
and U7740 (N_7740,N_4308,N_3442);
and U7741 (N_7741,N_3327,N_4380);
nor U7742 (N_7742,N_4767,N_5951);
xor U7743 (N_7743,N_3943,N_3297);
or U7744 (N_7744,N_3850,N_5017);
or U7745 (N_7745,N_5248,N_5908);
or U7746 (N_7746,N_4495,N_3133);
nor U7747 (N_7747,N_5096,N_5533);
nand U7748 (N_7748,N_4176,N_5256);
or U7749 (N_7749,N_3570,N_4341);
nor U7750 (N_7750,N_3624,N_3981);
or U7751 (N_7751,N_3249,N_3944);
or U7752 (N_7752,N_5346,N_4216);
nor U7753 (N_7753,N_5852,N_4988);
nand U7754 (N_7754,N_4928,N_3052);
and U7755 (N_7755,N_4678,N_4227);
or U7756 (N_7756,N_3354,N_4424);
nor U7757 (N_7757,N_5564,N_5940);
nand U7758 (N_7758,N_5022,N_3110);
xor U7759 (N_7759,N_4173,N_5492);
nor U7760 (N_7760,N_5289,N_3589);
nor U7761 (N_7761,N_4661,N_3116);
nor U7762 (N_7762,N_5979,N_5417);
and U7763 (N_7763,N_5872,N_3705);
nand U7764 (N_7764,N_5598,N_4616);
nand U7765 (N_7765,N_3093,N_3539);
nand U7766 (N_7766,N_5180,N_4243);
and U7767 (N_7767,N_4043,N_3997);
nand U7768 (N_7768,N_5186,N_3253);
or U7769 (N_7769,N_3840,N_3734);
nor U7770 (N_7770,N_4626,N_3373);
or U7771 (N_7771,N_4645,N_5397);
or U7772 (N_7772,N_3671,N_5128);
nand U7773 (N_7773,N_4175,N_4817);
xnor U7774 (N_7774,N_4768,N_3490);
or U7775 (N_7775,N_3471,N_4088);
or U7776 (N_7776,N_4569,N_4522);
xnor U7777 (N_7777,N_5999,N_5223);
nor U7778 (N_7778,N_4799,N_4323);
and U7779 (N_7779,N_3509,N_4639);
or U7780 (N_7780,N_4235,N_3466);
nand U7781 (N_7781,N_4914,N_4295);
nand U7782 (N_7782,N_4029,N_3302);
xnor U7783 (N_7783,N_4329,N_3816);
or U7784 (N_7784,N_4612,N_3835);
nor U7785 (N_7785,N_5662,N_4245);
and U7786 (N_7786,N_4268,N_4305);
and U7787 (N_7787,N_4813,N_5876);
and U7788 (N_7788,N_5405,N_3668);
xor U7789 (N_7789,N_3936,N_3726);
nor U7790 (N_7790,N_3779,N_5630);
nor U7791 (N_7791,N_5781,N_5487);
or U7792 (N_7792,N_5923,N_4478);
and U7793 (N_7793,N_4889,N_5798);
nand U7794 (N_7794,N_4560,N_3172);
nand U7795 (N_7795,N_4753,N_3759);
nor U7796 (N_7796,N_3714,N_4743);
nor U7797 (N_7797,N_3901,N_3267);
nand U7798 (N_7798,N_5968,N_3775);
nor U7799 (N_7799,N_5011,N_4283);
nand U7800 (N_7800,N_3924,N_4018);
or U7801 (N_7801,N_3571,N_3139);
xnor U7802 (N_7802,N_4950,N_3875);
nor U7803 (N_7803,N_5246,N_3709);
nand U7804 (N_7804,N_4034,N_5400);
and U7805 (N_7805,N_3890,N_3105);
xnor U7806 (N_7806,N_3651,N_3818);
nor U7807 (N_7807,N_5286,N_4594);
nor U7808 (N_7808,N_3292,N_3967);
nand U7809 (N_7809,N_5903,N_4442);
nand U7810 (N_7810,N_5430,N_3048);
nand U7811 (N_7811,N_5257,N_5642);
and U7812 (N_7812,N_3005,N_5806);
nor U7813 (N_7813,N_3191,N_5296);
nor U7814 (N_7814,N_4498,N_4105);
nor U7815 (N_7815,N_5175,N_5838);
and U7816 (N_7816,N_4951,N_5772);
and U7817 (N_7817,N_5469,N_3540);
and U7818 (N_7818,N_3163,N_3370);
and U7819 (N_7819,N_5242,N_4801);
nand U7820 (N_7820,N_5317,N_4764);
or U7821 (N_7821,N_5970,N_5431);
nor U7822 (N_7822,N_4613,N_4369);
nand U7823 (N_7823,N_4222,N_4684);
or U7824 (N_7824,N_3352,N_5229);
or U7825 (N_7825,N_5521,N_4306);
nand U7826 (N_7826,N_4184,N_5516);
or U7827 (N_7827,N_4417,N_4471);
or U7828 (N_7828,N_4896,N_3244);
nand U7829 (N_7829,N_5320,N_3899);
and U7830 (N_7830,N_5014,N_5042);
or U7831 (N_7831,N_3430,N_5223);
or U7832 (N_7832,N_5977,N_3854);
and U7833 (N_7833,N_5336,N_3730);
nand U7834 (N_7834,N_4000,N_3171);
or U7835 (N_7835,N_5924,N_5079);
xnor U7836 (N_7836,N_3672,N_4525);
and U7837 (N_7837,N_4783,N_5800);
or U7838 (N_7838,N_4798,N_4205);
or U7839 (N_7839,N_3783,N_5393);
or U7840 (N_7840,N_5094,N_3220);
and U7841 (N_7841,N_5790,N_4225);
or U7842 (N_7842,N_5044,N_4968);
nand U7843 (N_7843,N_3809,N_5649);
nor U7844 (N_7844,N_4297,N_4148);
xor U7845 (N_7845,N_4871,N_4859);
or U7846 (N_7846,N_4061,N_4698);
or U7847 (N_7847,N_4434,N_4441);
nand U7848 (N_7848,N_4821,N_5025);
or U7849 (N_7849,N_3367,N_4505);
and U7850 (N_7850,N_4925,N_4207);
nor U7851 (N_7851,N_4491,N_4955);
or U7852 (N_7852,N_4669,N_5016);
and U7853 (N_7853,N_3929,N_5877);
or U7854 (N_7854,N_5969,N_3702);
xor U7855 (N_7855,N_4506,N_5448);
and U7856 (N_7856,N_4970,N_4975);
nor U7857 (N_7857,N_5432,N_4964);
nand U7858 (N_7858,N_5800,N_3214);
nor U7859 (N_7859,N_4590,N_3681);
xnor U7860 (N_7860,N_3825,N_3407);
nor U7861 (N_7861,N_3547,N_3556);
nand U7862 (N_7862,N_4495,N_4981);
nor U7863 (N_7863,N_5324,N_4267);
or U7864 (N_7864,N_3075,N_5614);
nand U7865 (N_7865,N_5571,N_3502);
nor U7866 (N_7866,N_4017,N_4825);
xnor U7867 (N_7867,N_3747,N_5304);
nor U7868 (N_7868,N_4363,N_3198);
nor U7869 (N_7869,N_5939,N_3414);
nand U7870 (N_7870,N_4883,N_4466);
or U7871 (N_7871,N_5728,N_3430);
nor U7872 (N_7872,N_5531,N_5792);
nand U7873 (N_7873,N_3855,N_4863);
xnor U7874 (N_7874,N_5714,N_3794);
and U7875 (N_7875,N_5489,N_4783);
nand U7876 (N_7876,N_4998,N_5262);
or U7877 (N_7877,N_5127,N_4760);
nand U7878 (N_7878,N_4341,N_4680);
and U7879 (N_7879,N_4402,N_4470);
nand U7880 (N_7880,N_3285,N_3016);
or U7881 (N_7881,N_5334,N_4421);
nand U7882 (N_7882,N_4877,N_3386);
and U7883 (N_7883,N_4330,N_5742);
and U7884 (N_7884,N_3102,N_5131);
xor U7885 (N_7885,N_5564,N_3589);
and U7886 (N_7886,N_4758,N_4630);
nand U7887 (N_7887,N_3510,N_4550);
nor U7888 (N_7888,N_3538,N_5713);
or U7889 (N_7889,N_3406,N_4477);
or U7890 (N_7890,N_3480,N_5794);
nand U7891 (N_7891,N_5994,N_3630);
or U7892 (N_7892,N_4805,N_4350);
and U7893 (N_7893,N_4320,N_4590);
nor U7894 (N_7894,N_3549,N_3168);
xor U7895 (N_7895,N_5935,N_3305);
and U7896 (N_7896,N_5400,N_4056);
or U7897 (N_7897,N_3148,N_3485);
nor U7898 (N_7898,N_5311,N_3582);
nor U7899 (N_7899,N_4470,N_4245);
or U7900 (N_7900,N_3430,N_4809);
or U7901 (N_7901,N_3363,N_3287);
nor U7902 (N_7902,N_4071,N_5628);
and U7903 (N_7903,N_4021,N_5463);
and U7904 (N_7904,N_4986,N_4735);
nor U7905 (N_7905,N_3662,N_3737);
and U7906 (N_7906,N_5821,N_5022);
nand U7907 (N_7907,N_5049,N_3723);
nor U7908 (N_7908,N_4911,N_3545);
nand U7909 (N_7909,N_5353,N_5345);
nand U7910 (N_7910,N_5768,N_4496);
or U7911 (N_7911,N_5755,N_3232);
or U7912 (N_7912,N_5647,N_3866);
nor U7913 (N_7913,N_4514,N_5969);
nand U7914 (N_7914,N_4195,N_4978);
and U7915 (N_7915,N_4201,N_4349);
nor U7916 (N_7916,N_5875,N_5909);
or U7917 (N_7917,N_5271,N_4390);
nor U7918 (N_7918,N_5446,N_5889);
and U7919 (N_7919,N_4833,N_5526);
and U7920 (N_7920,N_3196,N_3047);
xor U7921 (N_7921,N_5259,N_5887);
or U7922 (N_7922,N_3277,N_5742);
nor U7923 (N_7923,N_3993,N_3429);
nor U7924 (N_7924,N_4686,N_3516);
nand U7925 (N_7925,N_3786,N_3184);
nor U7926 (N_7926,N_5811,N_4069);
or U7927 (N_7927,N_5703,N_3743);
nand U7928 (N_7928,N_5411,N_3659);
and U7929 (N_7929,N_4851,N_3549);
or U7930 (N_7930,N_4227,N_5183);
or U7931 (N_7931,N_5633,N_4399);
nor U7932 (N_7932,N_3639,N_4334);
nand U7933 (N_7933,N_5366,N_3236);
and U7934 (N_7934,N_4177,N_3013);
nand U7935 (N_7935,N_3020,N_4637);
nor U7936 (N_7936,N_4479,N_4103);
and U7937 (N_7937,N_3114,N_4924);
nand U7938 (N_7938,N_3325,N_3061);
and U7939 (N_7939,N_4015,N_5597);
and U7940 (N_7940,N_4622,N_3192);
nand U7941 (N_7941,N_5410,N_5365);
or U7942 (N_7942,N_5520,N_5739);
or U7943 (N_7943,N_4171,N_4699);
and U7944 (N_7944,N_3580,N_5460);
nand U7945 (N_7945,N_5746,N_5823);
nand U7946 (N_7946,N_3751,N_5178);
and U7947 (N_7947,N_5213,N_3466);
or U7948 (N_7948,N_5337,N_4263);
nor U7949 (N_7949,N_4450,N_3060);
nand U7950 (N_7950,N_5629,N_4315);
xnor U7951 (N_7951,N_5170,N_4783);
nand U7952 (N_7952,N_5329,N_5810);
nand U7953 (N_7953,N_3512,N_5803);
xor U7954 (N_7954,N_5790,N_3561);
nand U7955 (N_7955,N_3729,N_3717);
and U7956 (N_7956,N_4286,N_5910);
and U7957 (N_7957,N_4494,N_4397);
nand U7958 (N_7958,N_5207,N_3027);
nor U7959 (N_7959,N_4268,N_5176);
nor U7960 (N_7960,N_3846,N_5160);
nor U7961 (N_7961,N_5908,N_3253);
xor U7962 (N_7962,N_4621,N_4403);
nand U7963 (N_7963,N_3186,N_5624);
nand U7964 (N_7964,N_5664,N_5508);
or U7965 (N_7965,N_4613,N_4063);
and U7966 (N_7966,N_3413,N_4868);
nand U7967 (N_7967,N_5633,N_3606);
xnor U7968 (N_7968,N_5556,N_5444);
nand U7969 (N_7969,N_3835,N_5653);
or U7970 (N_7970,N_3898,N_4755);
xor U7971 (N_7971,N_4571,N_5583);
nor U7972 (N_7972,N_5109,N_4734);
xnor U7973 (N_7973,N_4797,N_5824);
and U7974 (N_7974,N_4296,N_3912);
and U7975 (N_7975,N_4160,N_4885);
or U7976 (N_7976,N_4843,N_4705);
nor U7977 (N_7977,N_3065,N_4117);
nor U7978 (N_7978,N_3151,N_4735);
and U7979 (N_7979,N_5267,N_4475);
and U7980 (N_7980,N_3356,N_5564);
nand U7981 (N_7981,N_3091,N_4572);
or U7982 (N_7982,N_3653,N_4347);
nand U7983 (N_7983,N_4955,N_4832);
or U7984 (N_7984,N_5561,N_5644);
and U7985 (N_7985,N_3309,N_5216);
nor U7986 (N_7986,N_3206,N_3057);
and U7987 (N_7987,N_3811,N_4396);
nor U7988 (N_7988,N_3084,N_3989);
or U7989 (N_7989,N_4414,N_4589);
or U7990 (N_7990,N_4390,N_3726);
nand U7991 (N_7991,N_4459,N_5944);
and U7992 (N_7992,N_3683,N_3579);
nor U7993 (N_7993,N_4481,N_5743);
and U7994 (N_7994,N_4104,N_4424);
nor U7995 (N_7995,N_4437,N_4366);
xnor U7996 (N_7996,N_4863,N_5462);
and U7997 (N_7997,N_4815,N_3466);
nor U7998 (N_7998,N_5712,N_4024);
nor U7999 (N_7999,N_4434,N_4301);
and U8000 (N_8000,N_3666,N_5179);
nor U8001 (N_8001,N_4939,N_3923);
nand U8002 (N_8002,N_3478,N_5123);
nand U8003 (N_8003,N_5202,N_4397);
nand U8004 (N_8004,N_3661,N_3733);
and U8005 (N_8005,N_3048,N_3190);
or U8006 (N_8006,N_4104,N_3844);
and U8007 (N_8007,N_5714,N_5027);
nor U8008 (N_8008,N_4844,N_4788);
xor U8009 (N_8009,N_4261,N_5921);
nor U8010 (N_8010,N_4007,N_5582);
nor U8011 (N_8011,N_3121,N_5760);
nor U8012 (N_8012,N_5779,N_3071);
and U8013 (N_8013,N_5231,N_5801);
xnor U8014 (N_8014,N_5223,N_5516);
nand U8015 (N_8015,N_4216,N_3650);
or U8016 (N_8016,N_3173,N_5676);
and U8017 (N_8017,N_5476,N_4552);
nand U8018 (N_8018,N_5242,N_4953);
nor U8019 (N_8019,N_4366,N_3014);
nor U8020 (N_8020,N_5728,N_5966);
and U8021 (N_8021,N_4719,N_5571);
nor U8022 (N_8022,N_5842,N_3140);
nand U8023 (N_8023,N_3400,N_4730);
nor U8024 (N_8024,N_3404,N_4378);
nand U8025 (N_8025,N_3616,N_3809);
nand U8026 (N_8026,N_5504,N_3553);
or U8027 (N_8027,N_4537,N_4566);
or U8028 (N_8028,N_3200,N_3048);
and U8029 (N_8029,N_5547,N_4195);
or U8030 (N_8030,N_3401,N_4230);
nor U8031 (N_8031,N_3545,N_5505);
nand U8032 (N_8032,N_3975,N_3900);
nor U8033 (N_8033,N_3041,N_3900);
or U8034 (N_8034,N_5268,N_4231);
or U8035 (N_8035,N_5976,N_4764);
nor U8036 (N_8036,N_4931,N_4306);
or U8037 (N_8037,N_5333,N_3768);
and U8038 (N_8038,N_3598,N_3958);
xnor U8039 (N_8039,N_4329,N_3594);
or U8040 (N_8040,N_4981,N_4063);
or U8041 (N_8041,N_3836,N_4264);
or U8042 (N_8042,N_5774,N_3373);
or U8043 (N_8043,N_5017,N_4429);
or U8044 (N_8044,N_3758,N_4734);
or U8045 (N_8045,N_5730,N_3419);
or U8046 (N_8046,N_5893,N_5631);
nand U8047 (N_8047,N_5173,N_5962);
nand U8048 (N_8048,N_3666,N_3344);
and U8049 (N_8049,N_3993,N_4936);
xnor U8050 (N_8050,N_5232,N_4540);
or U8051 (N_8051,N_4923,N_5829);
nand U8052 (N_8052,N_5733,N_5433);
and U8053 (N_8053,N_4002,N_3008);
nand U8054 (N_8054,N_4622,N_5940);
and U8055 (N_8055,N_4110,N_4889);
and U8056 (N_8056,N_4178,N_3497);
or U8057 (N_8057,N_4498,N_4196);
nand U8058 (N_8058,N_3244,N_3624);
nor U8059 (N_8059,N_3763,N_3661);
nor U8060 (N_8060,N_5177,N_4442);
nand U8061 (N_8061,N_3364,N_3122);
xnor U8062 (N_8062,N_4143,N_4629);
xor U8063 (N_8063,N_4649,N_4327);
or U8064 (N_8064,N_5622,N_5483);
and U8065 (N_8065,N_3512,N_4123);
nand U8066 (N_8066,N_5616,N_4941);
nor U8067 (N_8067,N_3956,N_5021);
nand U8068 (N_8068,N_4231,N_5613);
or U8069 (N_8069,N_5849,N_4220);
and U8070 (N_8070,N_5404,N_5782);
or U8071 (N_8071,N_4842,N_5661);
and U8072 (N_8072,N_4430,N_3143);
nand U8073 (N_8073,N_5293,N_4459);
nand U8074 (N_8074,N_4242,N_5393);
xor U8075 (N_8075,N_4848,N_3232);
nor U8076 (N_8076,N_3866,N_3738);
and U8077 (N_8077,N_5817,N_4607);
and U8078 (N_8078,N_4775,N_3499);
or U8079 (N_8079,N_5464,N_4540);
nor U8080 (N_8080,N_4224,N_5845);
or U8081 (N_8081,N_4882,N_3987);
or U8082 (N_8082,N_3957,N_4195);
and U8083 (N_8083,N_4541,N_5481);
or U8084 (N_8084,N_3314,N_3106);
nor U8085 (N_8085,N_4361,N_4279);
nor U8086 (N_8086,N_4704,N_3610);
nand U8087 (N_8087,N_3877,N_5987);
or U8088 (N_8088,N_4769,N_4554);
nand U8089 (N_8089,N_5946,N_3573);
nand U8090 (N_8090,N_3206,N_5189);
or U8091 (N_8091,N_3012,N_5512);
and U8092 (N_8092,N_5986,N_3358);
nand U8093 (N_8093,N_4099,N_3220);
nor U8094 (N_8094,N_5104,N_3133);
and U8095 (N_8095,N_5606,N_3973);
and U8096 (N_8096,N_4693,N_5876);
nor U8097 (N_8097,N_3989,N_5693);
or U8098 (N_8098,N_5754,N_5771);
nor U8099 (N_8099,N_4616,N_4078);
or U8100 (N_8100,N_3016,N_3080);
and U8101 (N_8101,N_3657,N_4677);
and U8102 (N_8102,N_3860,N_4880);
and U8103 (N_8103,N_4546,N_3226);
nor U8104 (N_8104,N_4172,N_4380);
and U8105 (N_8105,N_3648,N_3905);
or U8106 (N_8106,N_3991,N_5972);
nor U8107 (N_8107,N_4115,N_3854);
or U8108 (N_8108,N_4251,N_3229);
nand U8109 (N_8109,N_4160,N_5719);
nand U8110 (N_8110,N_3457,N_3830);
and U8111 (N_8111,N_5782,N_3838);
nor U8112 (N_8112,N_4805,N_5711);
and U8113 (N_8113,N_4142,N_4807);
nand U8114 (N_8114,N_5609,N_4769);
or U8115 (N_8115,N_5039,N_4266);
or U8116 (N_8116,N_3633,N_5940);
and U8117 (N_8117,N_4215,N_4622);
nand U8118 (N_8118,N_4147,N_3951);
xnor U8119 (N_8119,N_3844,N_3310);
nor U8120 (N_8120,N_5767,N_3646);
and U8121 (N_8121,N_5402,N_5397);
or U8122 (N_8122,N_5296,N_3454);
or U8123 (N_8123,N_5980,N_4457);
or U8124 (N_8124,N_3184,N_4630);
nor U8125 (N_8125,N_5885,N_3221);
nor U8126 (N_8126,N_5373,N_4196);
nor U8127 (N_8127,N_3763,N_5987);
or U8128 (N_8128,N_5259,N_3525);
and U8129 (N_8129,N_5676,N_3773);
nand U8130 (N_8130,N_4089,N_5711);
nor U8131 (N_8131,N_4984,N_5065);
xor U8132 (N_8132,N_3429,N_3436);
or U8133 (N_8133,N_5821,N_3023);
nor U8134 (N_8134,N_3530,N_3645);
nor U8135 (N_8135,N_4158,N_4361);
nor U8136 (N_8136,N_5926,N_3015);
and U8137 (N_8137,N_3111,N_4365);
nor U8138 (N_8138,N_3936,N_4769);
nand U8139 (N_8139,N_3027,N_5086);
xor U8140 (N_8140,N_4214,N_5466);
nand U8141 (N_8141,N_3078,N_5288);
or U8142 (N_8142,N_5677,N_3169);
or U8143 (N_8143,N_3328,N_4758);
nor U8144 (N_8144,N_5717,N_5492);
nor U8145 (N_8145,N_3769,N_5871);
or U8146 (N_8146,N_4458,N_5044);
and U8147 (N_8147,N_4518,N_5027);
nor U8148 (N_8148,N_3010,N_4646);
nand U8149 (N_8149,N_5049,N_3057);
or U8150 (N_8150,N_4701,N_3627);
nor U8151 (N_8151,N_5345,N_3462);
xnor U8152 (N_8152,N_4209,N_5254);
nand U8153 (N_8153,N_5246,N_3632);
and U8154 (N_8154,N_5692,N_5891);
and U8155 (N_8155,N_4796,N_4895);
nor U8156 (N_8156,N_3808,N_4775);
nand U8157 (N_8157,N_4752,N_4582);
nor U8158 (N_8158,N_5337,N_3496);
and U8159 (N_8159,N_4191,N_3698);
nand U8160 (N_8160,N_3490,N_5823);
nand U8161 (N_8161,N_5575,N_5107);
nand U8162 (N_8162,N_5407,N_3758);
nor U8163 (N_8163,N_5531,N_3908);
and U8164 (N_8164,N_4352,N_3241);
and U8165 (N_8165,N_4092,N_4019);
or U8166 (N_8166,N_4258,N_3180);
or U8167 (N_8167,N_3269,N_5834);
or U8168 (N_8168,N_4612,N_4987);
nand U8169 (N_8169,N_3010,N_5937);
or U8170 (N_8170,N_5929,N_5208);
or U8171 (N_8171,N_4071,N_3387);
nor U8172 (N_8172,N_4470,N_5237);
nor U8173 (N_8173,N_3067,N_3296);
or U8174 (N_8174,N_4421,N_3290);
and U8175 (N_8175,N_4003,N_3134);
nor U8176 (N_8176,N_3862,N_5643);
nand U8177 (N_8177,N_3799,N_5358);
nand U8178 (N_8178,N_4293,N_3693);
nand U8179 (N_8179,N_4157,N_3259);
nand U8180 (N_8180,N_3383,N_4599);
nand U8181 (N_8181,N_5849,N_3296);
nand U8182 (N_8182,N_3152,N_5695);
and U8183 (N_8183,N_5052,N_3631);
nor U8184 (N_8184,N_3486,N_4998);
or U8185 (N_8185,N_3993,N_5255);
and U8186 (N_8186,N_4421,N_4303);
nand U8187 (N_8187,N_4700,N_5027);
or U8188 (N_8188,N_5523,N_4909);
or U8189 (N_8189,N_3072,N_5599);
xnor U8190 (N_8190,N_4331,N_3814);
and U8191 (N_8191,N_4938,N_3300);
or U8192 (N_8192,N_5029,N_5483);
or U8193 (N_8193,N_3904,N_3213);
nand U8194 (N_8194,N_5294,N_4144);
and U8195 (N_8195,N_4361,N_4339);
or U8196 (N_8196,N_4722,N_3051);
nor U8197 (N_8197,N_3611,N_5171);
or U8198 (N_8198,N_5705,N_5880);
or U8199 (N_8199,N_4395,N_5747);
nor U8200 (N_8200,N_3135,N_5410);
and U8201 (N_8201,N_3935,N_3358);
and U8202 (N_8202,N_5090,N_3592);
xor U8203 (N_8203,N_3290,N_3520);
nor U8204 (N_8204,N_4581,N_5224);
nand U8205 (N_8205,N_4679,N_5174);
xnor U8206 (N_8206,N_3921,N_5686);
nor U8207 (N_8207,N_4082,N_4042);
nand U8208 (N_8208,N_4080,N_5968);
nand U8209 (N_8209,N_4929,N_3955);
or U8210 (N_8210,N_3522,N_4666);
nand U8211 (N_8211,N_5138,N_4070);
xnor U8212 (N_8212,N_3957,N_4934);
nor U8213 (N_8213,N_5995,N_3056);
nand U8214 (N_8214,N_4643,N_4912);
and U8215 (N_8215,N_5854,N_3841);
or U8216 (N_8216,N_3400,N_5059);
or U8217 (N_8217,N_3118,N_4675);
nor U8218 (N_8218,N_4452,N_5089);
nor U8219 (N_8219,N_4132,N_5657);
xnor U8220 (N_8220,N_5666,N_5491);
nand U8221 (N_8221,N_4256,N_4164);
or U8222 (N_8222,N_4605,N_4270);
nand U8223 (N_8223,N_4869,N_5994);
or U8224 (N_8224,N_3612,N_4942);
nand U8225 (N_8225,N_3831,N_4308);
nor U8226 (N_8226,N_3293,N_4145);
nand U8227 (N_8227,N_5239,N_4058);
xor U8228 (N_8228,N_4409,N_5985);
or U8229 (N_8229,N_3509,N_4548);
and U8230 (N_8230,N_4596,N_5301);
nor U8231 (N_8231,N_3291,N_3594);
nand U8232 (N_8232,N_3110,N_3422);
and U8233 (N_8233,N_3781,N_3046);
nand U8234 (N_8234,N_3473,N_4730);
xor U8235 (N_8235,N_4164,N_5970);
xnor U8236 (N_8236,N_4714,N_3674);
nand U8237 (N_8237,N_3269,N_5984);
xor U8238 (N_8238,N_5732,N_4309);
nand U8239 (N_8239,N_5029,N_5119);
and U8240 (N_8240,N_4451,N_3784);
nand U8241 (N_8241,N_4518,N_4291);
nand U8242 (N_8242,N_3616,N_4734);
and U8243 (N_8243,N_5917,N_4921);
nor U8244 (N_8244,N_3151,N_5230);
and U8245 (N_8245,N_4309,N_5572);
nand U8246 (N_8246,N_4928,N_3991);
and U8247 (N_8247,N_3872,N_3356);
or U8248 (N_8248,N_3928,N_5363);
xnor U8249 (N_8249,N_4422,N_5430);
and U8250 (N_8250,N_4593,N_4400);
nor U8251 (N_8251,N_3291,N_3011);
and U8252 (N_8252,N_4911,N_4848);
xnor U8253 (N_8253,N_4940,N_5306);
nand U8254 (N_8254,N_4850,N_4896);
nand U8255 (N_8255,N_4321,N_5850);
or U8256 (N_8256,N_5919,N_3666);
nand U8257 (N_8257,N_5379,N_4396);
nor U8258 (N_8258,N_4765,N_5469);
or U8259 (N_8259,N_3172,N_5346);
nand U8260 (N_8260,N_4370,N_4432);
xor U8261 (N_8261,N_3159,N_4639);
nand U8262 (N_8262,N_4216,N_3656);
xor U8263 (N_8263,N_5244,N_4218);
and U8264 (N_8264,N_3507,N_5001);
and U8265 (N_8265,N_4575,N_5546);
or U8266 (N_8266,N_3727,N_5428);
or U8267 (N_8267,N_5252,N_4076);
and U8268 (N_8268,N_5229,N_5477);
and U8269 (N_8269,N_3700,N_3461);
nand U8270 (N_8270,N_3288,N_5625);
nor U8271 (N_8271,N_3962,N_5704);
nor U8272 (N_8272,N_4474,N_5995);
nor U8273 (N_8273,N_5423,N_4127);
nand U8274 (N_8274,N_5767,N_4093);
nand U8275 (N_8275,N_5691,N_3621);
and U8276 (N_8276,N_4386,N_3324);
nor U8277 (N_8277,N_3271,N_3139);
and U8278 (N_8278,N_3344,N_5864);
or U8279 (N_8279,N_3115,N_4637);
or U8280 (N_8280,N_3652,N_3508);
or U8281 (N_8281,N_3926,N_4154);
and U8282 (N_8282,N_5572,N_3618);
or U8283 (N_8283,N_5896,N_4964);
nand U8284 (N_8284,N_5973,N_5833);
xor U8285 (N_8285,N_4731,N_5861);
nand U8286 (N_8286,N_5134,N_5922);
or U8287 (N_8287,N_5755,N_3191);
xnor U8288 (N_8288,N_3112,N_4727);
or U8289 (N_8289,N_3881,N_5422);
nor U8290 (N_8290,N_4173,N_5655);
and U8291 (N_8291,N_3307,N_3279);
and U8292 (N_8292,N_3298,N_3057);
or U8293 (N_8293,N_4097,N_3518);
nor U8294 (N_8294,N_3435,N_3861);
and U8295 (N_8295,N_4766,N_4416);
and U8296 (N_8296,N_5704,N_4143);
nand U8297 (N_8297,N_3561,N_5576);
or U8298 (N_8298,N_4256,N_5893);
and U8299 (N_8299,N_5319,N_4620);
xnor U8300 (N_8300,N_5608,N_4502);
nor U8301 (N_8301,N_5643,N_3849);
or U8302 (N_8302,N_4810,N_4659);
nor U8303 (N_8303,N_3318,N_4547);
nand U8304 (N_8304,N_3238,N_3519);
or U8305 (N_8305,N_5419,N_3644);
nor U8306 (N_8306,N_3338,N_4181);
or U8307 (N_8307,N_4306,N_5615);
and U8308 (N_8308,N_4186,N_5232);
and U8309 (N_8309,N_4065,N_5081);
and U8310 (N_8310,N_4068,N_4916);
nand U8311 (N_8311,N_5293,N_5785);
nand U8312 (N_8312,N_3703,N_3080);
xnor U8313 (N_8313,N_4798,N_3595);
or U8314 (N_8314,N_5469,N_5526);
nand U8315 (N_8315,N_3990,N_5369);
or U8316 (N_8316,N_4633,N_5724);
nor U8317 (N_8317,N_5779,N_3795);
nor U8318 (N_8318,N_3449,N_5973);
and U8319 (N_8319,N_4785,N_5272);
xor U8320 (N_8320,N_4086,N_5797);
and U8321 (N_8321,N_4060,N_4203);
nor U8322 (N_8322,N_4372,N_5101);
and U8323 (N_8323,N_4801,N_3404);
nor U8324 (N_8324,N_3474,N_5771);
nand U8325 (N_8325,N_3835,N_4813);
nor U8326 (N_8326,N_4796,N_3139);
or U8327 (N_8327,N_4467,N_3682);
xor U8328 (N_8328,N_5037,N_5347);
or U8329 (N_8329,N_4126,N_4526);
and U8330 (N_8330,N_4415,N_5053);
nand U8331 (N_8331,N_5872,N_4799);
and U8332 (N_8332,N_3967,N_5028);
xnor U8333 (N_8333,N_3219,N_5561);
or U8334 (N_8334,N_3668,N_4798);
xnor U8335 (N_8335,N_5405,N_4195);
or U8336 (N_8336,N_5273,N_3081);
xor U8337 (N_8337,N_4801,N_3042);
nand U8338 (N_8338,N_5079,N_3989);
nand U8339 (N_8339,N_4225,N_3153);
or U8340 (N_8340,N_4419,N_4678);
or U8341 (N_8341,N_3377,N_3707);
nor U8342 (N_8342,N_4143,N_3391);
nor U8343 (N_8343,N_3045,N_5086);
nand U8344 (N_8344,N_3580,N_4098);
nor U8345 (N_8345,N_4518,N_3214);
nand U8346 (N_8346,N_5592,N_5845);
and U8347 (N_8347,N_3126,N_4213);
xor U8348 (N_8348,N_5286,N_4454);
nor U8349 (N_8349,N_4142,N_4393);
nor U8350 (N_8350,N_5087,N_3843);
nor U8351 (N_8351,N_5847,N_5885);
and U8352 (N_8352,N_3302,N_5356);
nor U8353 (N_8353,N_3241,N_4311);
nor U8354 (N_8354,N_5420,N_4914);
nand U8355 (N_8355,N_3418,N_5074);
nor U8356 (N_8356,N_5474,N_3198);
nor U8357 (N_8357,N_4408,N_5170);
nand U8358 (N_8358,N_5616,N_5820);
nand U8359 (N_8359,N_5891,N_5731);
and U8360 (N_8360,N_5740,N_4008);
or U8361 (N_8361,N_5956,N_4887);
or U8362 (N_8362,N_4012,N_4023);
xnor U8363 (N_8363,N_4553,N_3539);
nor U8364 (N_8364,N_3305,N_5338);
nand U8365 (N_8365,N_5615,N_5075);
nand U8366 (N_8366,N_5230,N_4893);
nor U8367 (N_8367,N_5966,N_4379);
or U8368 (N_8368,N_4903,N_5442);
nand U8369 (N_8369,N_4448,N_5696);
and U8370 (N_8370,N_3671,N_5421);
nor U8371 (N_8371,N_3523,N_4215);
and U8372 (N_8372,N_4508,N_4282);
and U8373 (N_8373,N_3685,N_5796);
nor U8374 (N_8374,N_3417,N_5761);
and U8375 (N_8375,N_5357,N_4832);
or U8376 (N_8376,N_3723,N_3523);
and U8377 (N_8377,N_3460,N_4956);
nor U8378 (N_8378,N_4431,N_4235);
nor U8379 (N_8379,N_4862,N_5571);
nand U8380 (N_8380,N_3174,N_3413);
or U8381 (N_8381,N_4625,N_5393);
nor U8382 (N_8382,N_4585,N_3304);
nand U8383 (N_8383,N_5376,N_5929);
or U8384 (N_8384,N_3989,N_5493);
and U8385 (N_8385,N_5343,N_5654);
nor U8386 (N_8386,N_4102,N_4344);
nand U8387 (N_8387,N_3710,N_5527);
or U8388 (N_8388,N_4348,N_4695);
xnor U8389 (N_8389,N_5473,N_5801);
xnor U8390 (N_8390,N_4310,N_3357);
nand U8391 (N_8391,N_4039,N_5828);
or U8392 (N_8392,N_3762,N_4782);
xnor U8393 (N_8393,N_4666,N_5006);
and U8394 (N_8394,N_3347,N_3981);
nand U8395 (N_8395,N_3385,N_3333);
or U8396 (N_8396,N_5773,N_4857);
nor U8397 (N_8397,N_5032,N_5827);
nand U8398 (N_8398,N_3624,N_5719);
nor U8399 (N_8399,N_5234,N_5645);
and U8400 (N_8400,N_4755,N_3931);
or U8401 (N_8401,N_5852,N_3801);
nor U8402 (N_8402,N_3328,N_4522);
xnor U8403 (N_8403,N_3619,N_3598);
or U8404 (N_8404,N_3139,N_3624);
nand U8405 (N_8405,N_3703,N_3917);
or U8406 (N_8406,N_3867,N_3719);
nand U8407 (N_8407,N_3820,N_4329);
and U8408 (N_8408,N_3325,N_4222);
or U8409 (N_8409,N_5171,N_3689);
nand U8410 (N_8410,N_5147,N_4294);
or U8411 (N_8411,N_3810,N_4334);
nor U8412 (N_8412,N_5712,N_5059);
nor U8413 (N_8413,N_5249,N_5846);
nor U8414 (N_8414,N_3476,N_5716);
nor U8415 (N_8415,N_4365,N_4578);
or U8416 (N_8416,N_4278,N_5170);
or U8417 (N_8417,N_5987,N_3864);
or U8418 (N_8418,N_3303,N_5733);
nand U8419 (N_8419,N_5340,N_3907);
nor U8420 (N_8420,N_4681,N_4052);
or U8421 (N_8421,N_4231,N_4942);
and U8422 (N_8422,N_3050,N_5907);
or U8423 (N_8423,N_3751,N_5365);
or U8424 (N_8424,N_3266,N_3855);
and U8425 (N_8425,N_3609,N_3169);
or U8426 (N_8426,N_5575,N_4389);
nand U8427 (N_8427,N_5990,N_4381);
xor U8428 (N_8428,N_4266,N_5996);
or U8429 (N_8429,N_5708,N_3243);
and U8430 (N_8430,N_5592,N_5374);
nor U8431 (N_8431,N_5587,N_5385);
nor U8432 (N_8432,N_3834,N_3180);
or U8433 (N_8433,N_3851,N_5094);
nor U8434 (N_8434,N_4378,N_4596);
nor U8435 (N_8435,N_5985,N_4798);
nand U8436 (N_8436,N_4614,N_4562);
nand U8437 (N_8437,N_4152,N_5134);
nor U8438 (N_8438,N_4527,N_5706);
or U8439 (N_8439,N_3785,N_4281);
nand U8440 (N_8440,N_5503,N_5337);
and U8441 (N_8441,N_5963,N_5659);
nand U8442 (N_8442,N_4521,N_4885);
nand U8443 (N_8443,N_3309,N_3194);
xnor U8444 (N_8444,N_4019,N_4886);
nand U8445 (N_8445,N_3738,N_5719);
xnor U8446 (N_8446,N_3908,N_5259);
and U8447 (N_8447,N_4815,N_4761);
or U8448 (N_8448,N_3640,N_5153);
xnor U8449 (N_8449,N_5708,N_3318);
and U8450 (N_8450,N_4882,N_5776);
nor U8451 (N_8451,N_4896,N_4328);
nand U8452 (N_8452,N_3505,N_3424);
nor U8453 (N_8453,N_3029,N_5604);
and U8454 (N_8454,N_5371,N_5634);
and U8455 (N_8455,N_5585,N_5587);
and U8456 (N_8456,N_4328,N_4418);
nor U8457 (N_8457,N_5179,N_5608);
and U8458 (N_8458,N_3498,N_3192);
nor U8459 (N_8459,N_3622,N_4758);
and U8460 (N_8460,N_5013,N_5416);
nor U8461 (N_8461,N_4793,N_3303);
and U8462 (N_8462,N_5897,N_4634);
or U8463 (N_8463,N_4660,N_5739);
or U8464 (N_8464,N_3692,N_3347);
or U8465 (N_8465,N_3118,N_5556);
nor U8466 (N_8466,N_3906,N_5156);
and U8467 (N_8467,N_5089,N_5317);
xor U8468 (N_8468,N_4938,N_4849);
nand U8469 (N_8469,N_4012,N_4946);
nand U8470 (N_8470,N_5326,N_5155);
nor U8471 (N_8471,N_4412,N_3499);
or U8472 (N_8472,N_5945,N_5719);
xor U8473 (N_8473,N_3564,N_3406);
and U8474 (N_8474,N_4389,N_4681);
or U8475 (N_8475,N_4707,N_3839);
and U8476 (N_8476,N_3748,N_5596);
and U8477 (N_8477,N_3405,N_3662);
nand U8478 (N_8478,N_5329,N_5356);
or U8479 (N_8479,N_4655,N_5317);
or U8480 (N_8480,N_4631,N_4611);
nand U8481 (N_8481,N_5646,N_5944);
nand U8482 (N_8482,N_5741,N_4641);
or U8483 (N_8483,N_3425,N_5192);
or U8484 (N_8484,N_3127,N_4965);
or U8485 (N_8485,N_3083,N_5026);
nor U8486 (N_8486,N_3663,N_5956);
and U8487 (N_8487,N_4590,N_3607);
nor U8488 (N_8488,N_5660,N_5922);
nand U8489 (N_8489,N_4802,N_4783);
nor U8490 (N_8490,N_4432,N_3640);
nor U8491 (N_8491,N_3270,N_5905);
and U8492 (N_8492,N_5370,N_4977);
nand U8493 (N_8493,N_5723,N_3319);
xor U8494 (N_8494,N_5275,N_4181);
nand U8495 (N_8495,N_5683,N_3559);
nor U8496 (N_8496,N_5720,N_5344);
nor U8497 (N_8497,N_3705,N_3909);
nor U8498 (N_8498,N_4329,N_4108);
and U8499 (N_8499,N_3284,N_4218);
nor U8500 (N_8500,N_3058,N_5455);
or U8501 (N_8501,N_4534,N_4166);
and U8502 (N_8502,N_5782,N_4490);
nand U8503 (N_8503,N_4362,N_5495);
or U8504 (N_8504,N_4013,N_3739);
nor U8505 (N_8505,N_4412,N_3065);
nand U8506 (N_8506,N_3183,N_5855);
and U8507 (N_8507,N_4208,N_5273);
and U8508 (N_8508,N_5607,N_4547);
nor U8509 (N_8509,N_5108,N_4304);
or U8510 (N_8510,N_5421,N_4155);
xor U8511 (N_8511,N_5820,N_4696);
nand U8512 (N_8512,N_5877,N_4873);
xnor U8513 (N_8513,N_3105,N_4728);
nand U8514 (N_8514,N_4685,N_4644);
and U8515 (N_8515,N_3266,N_3207);
xnor U8516 (N_8516,N_4234,N_3061);
xor U8517 (N_8517,N_5513,N_3116);
nor U8518 (N_8518,N_3422,N_5256);
and U8519 (N_8519,N_4925,N_3418);
or U8520 (N_8520,N_5155,N_4126);
xor U8521 (N_8521,N_3968,N_4986);
and U8522 (N_8522,N_3408,N_5454);
and U8523 (N_8523,N_5480,N_5108);
or U8524 (N_8524,N_3969,N_5188);
or U8525 (N_8525,N_4699,N_5880);
nand U8526 (N_8526,N_5601,N_5182);
or U8527 (N_8527,N_4344,N_5778);
nand U8528 (N_8528,N_5034,N_4415);
or U8529 (N_8529,N_4699,N_4727);
nand U8530 (N_8530,N_3332,N_3161);
nor U8531 (N_8531,N_3090,N_5108);
nor U8532 (N_8532,N_5529,N_3415);
or U8533 (N_8533,N_4843,N_4304);
or U8534 (N_8534,N_5089,N_3636);
or U8535 (N_8535,N_3685,N_3027);
nand U8536 (N_8536,N_4695,N_4832);
and U8537 (N_8537,N_4612,N_4822);
or U8538 (N_8538,N_3226,N_4702);
nand U8539 (N_8539,N_4229,N_5937);
or U8540 (N_8540,N_3973,N_3722);
nor U8541 (N_8541,N_4882,N_4372);
or U8542 (N_8542,N_4968,N_5355);
nor U8543 (N_8543,N_3282,N_5852);
nor U8544 (N_8544,N_4717,N_4301);
nand U8545 (N_8545,N_5558,N_4170);
nor U8546 (N_8546,N_3050,N_3513);
and U8547 (N_8547,N_4010,N_5896);
nand U8548 (N_8548,N_5901,N_3301);
and U8549 (N_8549,N_3132,N_4183);
and U8550 (N_8550,N_3019,N_5001);
nor U8551 (N_8551,N_4981,N_3035);
or U8552 (N_8552,N_3255,N_5002);
nand U8553 (N_8553,N_5456,N_5159);
and U8554 (N_8554,N_5288,N_4941);
and U8555 (N_8555,N_4327,N_3689);
nand U8556 (N_8556,N_4090,N_5495);
and U8557 (N_8557,N_5316,N_5120);
and U8558 (N_8558,N_5313,N_5317);
or U8559 (N_8559,N_3506,N_3372);
xor U8560 (N_8560,N_5142,N_5545);
nor U8561 (N_8561,N_3449,N_5796);
nand U8562 (N_8562,N_5840,N_5456);
or U8563 (N_8563,N_4749,N_5541);
nor U8564 (N_8564,N_5892,N_4503);
and U8565 (N_8565,N_5189,N_5441);
and U8566 (N_8566,N_4996,N_4668);
nor U8567 (N_8567,N_3746,N_5748);
nor U8568 (N_8568,N_4082,N_4197);
and U8569 (N_8569,N_5636,N_4040);
nand U8570 (N_8570,N_4633,N_4741);
or U8571 (N_8571,N_3451,N_3530);
nand U8572 (N_8572,N_3015,N_5403);
or U8573 (N_8573,N_4986,N_5893);
or U8574 (N_8574,N_5791,N_4689);
and U8575 (N_8575,N_3328,N_5053);
or U8576 (N_8576,N_5086,N_5108);
nor U8577 (N_8577,N_3217,N_3852);
and U8578 (N_8578,N_3099,N_5264);
or U8579 (N_8579,N_3227,N_3264);
nand U8580 (N_8580,N_4940,N_3431);
and U8581 (N_8581,N_3194,N_3837);
nand U8582 (N_8582,N_5991,N_3157);
nand U8583 (N_8583,N_4349,N_4592);
xor U8584 (N_8584,N_3159,N_3033);
and U8585 (N_8585,N_4788,N_3301);
or U8586 (N_8586,N_3724,N_4155);
nor U8587 (N_8587,N_5087,N_3937);
nor U8588 (N_8588,N_3756,N_3136);
or U8589 (N_8589,N_4881,N_5226);
nor U8590 (N_8590,N_5331,N_3023);
xor U8591 (N_8591,N_5687,N_4602);
xor U8592 (N_8592,N_5978,N_4163);
or U8593 (N_8593,N_5186,N_3908);
nand U8594 (N_8594,N_4860,N_4152);
or U8595 (N_8595,N_3183,N_5815);
nand U8596 (N_8596,N_5244,N_4231);
nor U8597 (N_8597,N_5218,N_3225);
nor U8598 (N_8598,N_4871,N_4923);
and U8599 (N_8599,N_3929,N_3190);
and U8600 (N_8600,N_5488,N_3928);
nand U8601 (N_8601,N_5541,N_5400);
xnor U8602 (N_8602,N_5330,N_5734);
xor U8603 (N_8603,N_5578,N_5689);
and U8604 (N_8604,N_3173,N_4928);
and U8605 (N_8605,N_4447,N_4899);
nor U8606 (N_8606,N_3436,N_4716);
nor U8607 (N_8607,N_3860,N_3599);
xor U8608 (N_8608,N_4375,N_4397);
nor U8609 (N_8609,N_5865,N_4575);
nand U8610 (N_8610,N_3554,N_3218);
nor U8611 (N_8611,N_5233,N_3479);
and U8612 (N_8612,N_5408,N_4100);
nand U8613 (N_8613,N_5488,N_3162);
nand U8614 (N_8614,N_5732,N_5578);
or U8615 (N_8615,N_4996,N_4968);
nand U8616 (N_8616,N_4022,N_5187);
or U8617 (N_8617,N_5855,N_4838);
and U8618 (N_8618,N_3158,N_5831);
nand U8619 (N_8619,N_3402,N_5748);
nor U8620 (N_8620,N_5148,N_4987);
nor U8621 (N_8621,N_4079,N_4087);
and U8622 (N_8622,N_3284,N_5312);
nand U8623 (N_8623,N_4804,N_5214);
and U8624 (N_8624,N_4547,N_3614);
xnor U8625 (N_8625,N_5909,N_4197);
nor U8626 (N_8626,N_5443,N_5646);
xor U8627 (N_8627,N_4380,N_3653);
or U8628 (N_8628,N_3504,N_5157);
nor U8629 (N_8629,N_3356,N_3790);
xnor U8630 (N_8630,N_5820,N_5109);
nor U8631 (N_8631,N_4201,N_4557);
nand U8632 (N_8632,N_3926,N_5907);
or U8633 (N_8633,N_5181,N_3155);
or U8634 (N_8634,N_4711,N_5433);
nor U8635 (N_8635,N_3741,N_3015);
nor U8636 (N_8636,N_3664,N_5539);
nor U8637 (N_8637,N_4858,N_5669);
nor U8638 (N_8638,N_5736,N_4581);
nand U8639 (N_8639,N_4189,N_4969);
nand U8640 (N_8640,N_3525,N_4985);
or U8641 (N_8641,N_3012,N_5168);
and U8642 (N_8642,N_5087,N_4224);
nor U8643 (N_8643,N_4874,N_4060);
and U8644 (N_8644,N_4362,N_5515);
nand U8645 (N_8645,N_3869,N_3854);
nor U8646 (N_8646,N_4146,N_5630);
or U8647 (N_8647,N_4704,N_3826);
or U8648 (N_8648,N_5148,N_5618);
or U8649 (N_8649,N_4420,N_5786);
or U8650 (N_8650,N_5816,N_5387);
nand U8651 (N_8651,N_5858,N_3426);
xor U8652 (N_8652,N_3060,N_5358);
and U8653 (N_8653,N_4098,N_3308);
or U8654 (N_8654,N_4767,N_3487);
nor U8655 (N_8655,N_4439,N_4009);
nand U8656 (N_8656,N_3416,N_5524);
or U8657 (N_8657,N_3092,N_5465);
and U8658 (N_8658,N_3369,N_3587);
and U8659 (N_8659,N_4668,N_4820);
xor U8660 (N_8660,N_4422,N_4538);
or U8661 (N_8661,N_4057,N_3821);
and U8662 (N_8662,N_4357,N_3040);
or U8663 (N_8663,N_3904,N_3823);
or U8664 (N_8664,N_5674,N_4042);
or U8665 (N_8665,N_3496,N_5748);
nand U8666 (N_8666,N_3343,N_4503);
or U8667 (N_8667,N_4601,N_4571);
xnor U8668 (N_8668,N_3808,N_4427);
and U8669 (N_8669,N_4324,N_4805);
or U8670 (N_8670,N_5046,N_4740);
and U8671 (N_8671,N_4824,N_5714);
and U8672 (N_8672,N_4314,N_5810);
xnor U8673 (N_8673,N_4156,N_5779);
or U8674 (N_8674,N_5424,N_3323);
or U8675 (N_8675,N_4622,N_4861);
xor U8676 (N_8676,N_5217,N_3627);
and U8677 (N_8677,N_3770,N_4311);
or U8678 (N_8678,N_5868,N_3498);
xor U8679 (N_8679,N_4604,N_5559);
and U8680 (N_8680,N_3919,N_3270);
nand U8681 (N_8681,N_4964,N_4378);
and U8682 (N_8682,N_5240,N_4409);
nor U8683 (N_8683,N_5000,N_4909);
xor U8684 (N_8684,N_4159,N_5815);
or U8685 (N_8685,N_4760,N_4809);
nand U8686 (N_8686,N_5057,N_4647);
and U8687 (N_8687,N_4742,N_3406);
or U8688 (N_8688,N_4636,N_3123);
xnor U8689 (N_8689,N_4937,N_3006);
nand U8690 (N_8690,N_5382,N_5067);
nor U8691 (N_8691,N_5397,N_3505);
or U8692 (N_8692,N_5212,N_3391);
or U8693 (N_8693,N_5258,N_3647);
or U8694 (N_8694,N_3032,N_5699);
and U8695 (N_8695,N_3267,N_5577);
nand U8696 (N_8696,N_3261,N_4897);
xnor U8697 (N_8697,N_5021,N_5205);
or U8698 (N_8698,N_3700,N_5279);
or U8699 (N_8699,N_3038,N_5479);
or U8700 (N_8700,N_3543,N_3180);
and U8701 (N_8701,N_3566,N_4485);
nand U8702 (N_8702,N_4263,N_3744);
or U8703 (N_8703,N_5141,N_3112);
nor U8704 (N_8704,N_5329,N_3678);
or U8705 (N_8705,N_4079,N_3093);
nand U8706 (N_8706,N_3750,N_4919);
nor U8707 (N_8707,N_3817,N_3345);
and U8708 (N_8708,N_4781,N_4079);
and U8709 (N_8709,N_5778,N_4375);
xnor U8710 (N_8710,N_5492,N_5791);
and U8711 (N_8711,N_4236,N_3477);
nand U8712 (N_8712,N_4171,N_5579);
or U8713 (N_8713,N_5273,N_5137);
nor U8714 (N_8714,N_3118,N_4286);
and U8715 (N_8715,N_5752,N_4711);
or U8716 (N_8716,N_3141,N_3341);
nor U8717 (N_8717,N_5760,N_5721);
nor U8718 (N_8718,N_5639,N_3519);
nand U8719 (N_8719,N_4569,N_3882);
and U8720 (N_8720,N_4373,N_5976);
or U8721 (N_8721,N_5143,N_3557);
nand U8722 (N_8722,N_5607,N_4518);
or U8723 (N_8723,N_5417,N_5938);
nand U8724 (N_8724,N_4247,N_4545);
nand U8725 (N_8725,N_5470,N_4578);
and U8726 (N_8726,N_5548,N_3060);
nor U8727 (N_8727,N_4717,N_4376);
or U8728 (N_8728,N_4766,N_3348);
and U8729 (N_8729,N_3907,N_4916);
nand U8730 (N_8730,N_3954,N_4372);
and U8731 (N_8731,N_3479,N_4759);
nor U8732 (N_8732,N_4770,N_4254);
nor U8733 (N_8733,N_4231,N_5487);
or U8734 (N_8734,N_5142,N_3892);
and U8735 (N_8735,N_3349,N_3843);
nor U8736 (N_8736,N_3285,N_5800);
nor U8737 (N_8737,N_3177,N_3835);
or U8738 (N_8738,N_5693,N_3382);
nand U8739 (N_8739,N_4058,N_5142);
nor U8740 (N_8740,N_4096,N_5957);
nand U8741 (N_8741,N_3543,N_4022);
nand U8742 (N_8742,N_4317,N_4612);
nor U8743 (N_8743,N_4353,N_5151);
and U8744 (N_8744,N_5144,N_4589);
or U8745 (N_8745,N_5020,N_4893);
nand U8746 (N_8746,N_3983,N_5237);
nand U8747 (N_8747,N_3928,N_4673);
nand U8748 (N_8748,N_4824,N_5070);
nor U8749 (N_8749,N_4714,N_3731);
nor U8750 (N_8750,N_4099,N_4916);
nand U8751 (N_8751,N_5136,N_3838);
or U8752 (N_8752,N_4612,N_5724);
or U8753 (N_8753,N_4423,N_5084);
nor U8754 (N_8754,N_3552,N_4599);
nor U8755 (N_8755,N_3085,N_3409);
or U8756 (N_8756,N_3298,N_4025);
nand U8757 (N_8757,N_3688,N_5203);
or U8758 (N_8758,N_3128,N_3475);
nor U8759 (N_8759,N_5618,N_3076);
or U8760 (N_8760,N_3564,N_3414);
nor U8761 (N_8761,N_3440,N_4368);
or U8762 (N_8762,N_4760,N_3892);
nand U8763 (N_8763,N_5424,N_4374);
and U8764 (N_8764,N_4244,N_4265);
or U8765 (N_8765,N_5741,N_3742);
xor U8766 (N_8766,N_4019,N_3473);
or U8767 (N_8767,N_3300,N_5513);
or U8768 (N_8768,N_5218,N_3747);
or U8769 (N_8769,N_5353,N_4329);
and U8770 (N_8770,N_3278,N_4464);
nand U8771 (N_8771,N_4782,N_3061);
xor U8772 (N_8772,N_4255,N_3580);
or U8773 (N_8773,N_5728,N_4044);
or U8774 (N_8774,N_3876,N_5203);
nand U8775 (N_8775,N_5885,N_5483);
nand U8776 (N_8776,N_4662,N_5028);
nand U8777 (N_8777,N_3468,N_4555);
nand U8778 (N_8778,N_5330,N_3528);
or U8779 (N_8779,N_4226,N_4179);
nand U8780 (N_8780,N_5419,N_4406);
and U8781 (N_8781,N_4394,N_3418);
nor U8782 (N_8782,N_3410,N_4970);
or U8783 (N_8783,N_5437,N_5919);
or U8784 (N_8784,N_3966,N_5379);
xnor U8785 (N_8785,N_3086,N_4354);
or U8786 (N_8786,N_4352,N_5168);
nand U8787 (N_8787,N_4872,N_3563);
nand U8788 (N_8788,N_5217,N_3386);
nand U8789 (N_8789,N_5332,N_4643);
and U8790 (N_8790,N_3212,N_5200);
or U8791 (N_8791,N_5687,N_3142);
xnor U8792 (N_8792,N_5383,N_4727);
nand U8793 (N_8793,N_5718,N_5039);
or U8794 (N_8794,N_3254,N_4250);
and U8795 (N_8795,N_3526,N_5814);
nor U8796 (N_8796,N_3348,N_4017);
and U8797 (N_8797,N_4782,N_3871);
nor U8798 (N_8798,N_4874,N_4441);
and U8799 (N_8799,N_4870,N_4490);
or U8800 (N_8800,N_5197,N_5036);
nor U8801 (N_8801,N_4565,N_4462);
or U8802 (N_8802,N_4026,N_3258);
or U8803 (N_8803,N_3680,N_4961);
and U8804 (N_8804,N_3874,N_5118);
and U8805 (N_8805,N_5235,N_5000);
or U8806 (N_8806,N_5035,N_4850);
xor U8807 (N_8807,N_4192,N_4942);
and U8808 (N_8808,N_5770,N_4492);
xor U8809 (N_8809,N_4752,N_3390);
nor U8810 (N_8810,N_4608,N_3994);
xor U8811 (N_8811,N_3879,N_3738);
xor U8812 (N_8812,N_3435,N_4645);
nor U8813 (N_8813,N_4010,N_5691);
and U8814 (N_8814,N_3725,N_4267);
and U8815 (N_8815,N_5607,N_4128);
nand U8816 (N_8816,N_4542,N_3072);
and U8817 (N_8817,N_4021,N_4526);
and U8818 (N_8818,N_3819,N_5112);
or U8819 (N_8819,N_4595,N_4519);
nor U8820 (N_8820,N_5213,N_4168);
nand U8821 (N_8821,N_4240,N_3426);
nand U8822 (N_8822,N_5743,N_5502);
or U8823 (N_8823,N_3794,N_3295);
or U8824 (N_8824,N_4191,N_3039);
nor U8825 (N_8825,N_3389,N_5446);
and U8826 (N_8826,N_3659,N_3997);
or U8827 (N_8827,N_5929,N_3842);
nand U8828 (N_8828,N_4792,N_4160);
nor U8829 (N_8829,N_4343,N_3791);
nor U8830 (N_8830,N_5266,N_4841);
and U8831 (N_8831,N_5859,N_4282);
nor U8832 (N_8832,N_5622,N_4598);
nor U8833 (N_8833,N_3678,N_3808);
xor U8834 (N_8834,N_3763,N_5669);
and U8835 (N_8835,N_5212,N_5605);
nand U8836 (N_8836,N_5399,N_5815);
and U8837 (N_8837,N_4430,N_5593);
or U8838 (N_8838,N_3373,N_4592);
xnor U8839 (N_8839,N_5899,N_5529);
nor U8840 (N_8840,N_3459,N_4831);
or U8841 (N_8841,N_3161,N_4578);
and U8842 (N_8842,N_4430,N_3447);
and U8843 (N_8843,N_5780,N_5215);
and U8844 (N_8844,N_4951,N_3705);
nor U8845 (N_8845,N_3941,N_4476);
and U8846 (N_8846,N_5141,N_3797);
nor U8847 (N_8847,N_5335,N_4349);
nor U8848 (N_8848,N_5234,N_5751);
nor U8849 (N_8849,N_3193,N_3181);
nand U8850 (N_8850,N_4698,N_3318);
or U8851 (N_8851,N_5609,N_3094);
nand U8852 (N_8852,N_4398,N_3862);
or U8853 (N_8853,N_4293,N_5425);
or U8854 (N_8854,N_5536,N_4771);
and U8855 (N_8855,N_5794,N_5960);
or U8856 (N_8856,N_4808,N_5918);
and U8857 (N_8857,N_4625,N_4816);
or U8858 (N_8858,N_5506,N_5115);
nand U8859 (N_8859,N_3249,N_5532);
nor U8860 (N_8860,N_4720,N_3012);
and U8861 (N_8861,N_3305,N_4340);
and U8862 (N_8862,N_3739,N_5920);
nor U8863 (N_8863,N_5935,N_5580);
nand U8864 (N_8864,N_5220,N_3473);
xnor U8865 (N_8865,N_4233,N_5138);
nor U8866 (N_8866,N_3470,N_3102);
and U8867 (N_8867,N_4519,N_3703);
or U8868 (N_8868,N_3886,N_3515);
and U8869 (N_8869,N_3144,N_5150);
or U8870 (N_8870,N_4490,N_3664);
nand U8871 (N_8871,N_3740,N_5832);
or U8872 (N_8872,N_4203,N_3942);
or U8873 (N_8873,N_3870,N_3835);
nor U8874 (N_8874,N_5217,N_3316);
nor U8875 (N_8875,N_4637,N_5297);
and U8876 (N_8876,N_5537,N_5722);
or U8877 (N_8877,N_4092,N_5990);
or U8878 (N_8878,N_3851,N_4716);
and U8879 (N_8879,N_3755,N_4599);
xor U8880 (N_8880,N_5689,N_5336);
or U8881 (N_8881,N_3020,N_4481);
xor U8882 (N_8882,N_3383,N_3446);
nand U8883 (N_8883,N_3055,N_3342);
or U8884 (N_8884,N_4831,N_4691);
and U8885 (N_8885,N_3501,N_4724);
nand U8886 (N_8886,N_4320,N_4319);
nand U8887 (N_8887,N_5288,N_4555);
or U8888 (N_8888,N_5329,N_3661);
or U8889 (N_8889,N_3887,N_3271);
and U8890 (N_8890,N_4654,N_3100);
and U8891 (N_8891,N_5757,N_3471);
xor U8892 (N_8892,N_4486,N_5666);
nor U8893 (N_8893,N_5901,N_4558);
xnor U8894 (N_8894,N_4360,N_3638);
or U8895 (N_8895,N_4260,N_3994);
nand U8896 (N_8896,N_5637,N_4620);
or U8897 (N_8897,N_3086,N_4368);
or U8898 (N_8898,N_5487,N_5853);
and U8899 (N_8899,N_5374,N_4414);
or U8900 (N_8900,N_5759,N_4926);
nor U8901 (N_8901,N_3356,N_5288);
nor U8902 (N_8902,N_4073,N_5374);
or U8903 (N_8903,N_4857,N_3908);
nor U8904 (N_8904,N_4283,N_4157);
nor U8905 (N_8905,N_5115,N_5270);
nor U8906 (N_8906,N_4013,N_5460);
nor U8907 (N_8907,N_4958,N_4117);
nand U8908 (N_8908,N_5405,N_5795);
or U8909 (N_8909,N_5906,N_5605);
nand U8910 (N_8910,N_4508,N_3184);
nor U8911 (N_8911,N_3883,N_3058);
and U8912 (N_8912,N_5452,N_3382);
nand U8913 (N_8913,N_3991,N_3627);
and U8914 (N_8914,N_3135,N_4947);
nand U8915 (N_8915,N_5574,N_3195);
and U8916 (N_8916,N_3457,N_3640);
nand U8917 (N_8917,N_5908,N_3975);
nor U8918 (N_8918,N_4760,N_4774);
or U8919 (N_8919,N_3927,N_5268);
nor U8920 (N_8920,N_3943,N_3559);
nor U8921 (N_8921,N_5313,N_5948);
xor U8922 (N_8922,N_4608,N_3756);
nor U8923 (N_8923,N_4022,N_4780);
nor U8924 (N_8924,N_3783,N_4648);
nor U8925 (N_8925,N_4531,N_3399);
nor U8926 (N_8926,N_4674,N_3923);
or U8927 (N_8927,N_3855,N_4404);
nor U8928 (N_8928,N_3010,N_5703);
and U8929 (N_8929,N_5826,N_3261);
and U8930 (N_8930,N_3073,N_5104);
or U8931 (N_8931,N_4874,N_5049);
or U8932 (N_8932,N_4510,N_3030);
xnor U8933 (N_8933,N_4550,N_4074);
nand U8934 (N_8934,N_5425,N_5856);
xnor U8935 (N_8935,N_4704,N_4856);
xor U8936 (N_8936,N_4118,N_3866);
and U8937 (N_8937,N_5933,N_5078);
and U8938 (N_8938,N_3062,N_3004);
nand U8939 (N_8939,N_5287,N_5816);
nand U8940 (N_8940,N_5153,N_4968);
xnor U8941 (N_8941,N_3203,N_4681);
nor U8942 (N_8942,N_3045,N_4324);
nor U8943 (N_8943,N_5687,N_5149);
nor U8944 (N_8944,N_4398,N_3050);
and U8945 (N_8945,N_5695,N_4041);
or U8946 (N_8946,N_5063,N_4746);
and U8947 (N_8947,N_5065,N_4450);
xor U8948 (N_8948,N_3324,N_3233);
nor U8949 (N_8949,N_5301,N_4977);
or U8950 (N_8950,N_4684,N_5112);
nand U8951 (N_8951,N_4707,N_3945);
or U8952 (N_8952,N_5051,N_4678);
nand U8953 (N_8953,N_5102,N_5261);
nor U8954 (N_8954,N_3232,N_4618);
nand U8955 (N_8955,N_3307,N_3541);
nor U8956 (N_8956,N_5157,N_5287);
nand U8957 (N_8957,N_3095,N_3328);
or U8958 (N_8958,N_3127,N_3133);
nor U8959 (N_8959,N_3621,N_5104);
nor U8960 (N_8960,N_4090,N_4695);
nor U8961 (N_8961,N_5247,N_5842);
or U8962 (N_8962,N_4772,N_5152);
nor U8963 (N_8963,N_5515,N_5132);
or U8964 (N_8964,N_4995,N_5016);
nand U8965 (N_8965,N_5384,N_3674);
and U8966 (N_8966,N_4663,N_5086);
and U8967 (N_8967,N_5278,N_3736);
xor U8968 (N_8968,N_3959,N_4776);
and U8969 (N_8969,N_3416,N_4766);
and U8970 (N_8970,N_3149,N_5468);
xor U8971 (N_8971,N_4707,N_3907);
nand U8972 (N_8972,N_5894,N_5975);
nand U8973 (N_8973,N_4416,N_4650);
or U8974 (N_8974,N_3705,N_4716);
and U8975 (N_8975,N_5099,N_4806);
and U8976 (N_8976,N_4299,N_3016);
or U8977 (N_8977,N_3963,N_5652);
or U8978 (N_8978,N_4923,N_3282);
and U8979 (N_8979,N_3693,N_3228);
or U8980 (N_8980,N_4400,N_3316);
nor U8981 (N_8981,N_4747,N_4405);
nand U8982 (N_8982,N_3051,N_4396);
and U8983 (N_8983,N_5439,N_3620);
nand U8984 (N_8984,N_3572,N_5786);
xnor U8985 (N_8985,N_5251,N_5440);
and U8986 (N_8986,N_3748,N_4128);
or U8987 (N_8987,N_4039,N_3914);
nand U8988 (N_8988,N_4914,N_5921);
or U8989 (N_8989,N_5052,N_5019);
nor U8990 (N_8990,N_5587,N_3783);
nor U8991 (N_8991,N_5593,N_5868);
nand U8992 (N_8992,N_3239,N_3500);
nand U8993 (N_8993,N_4225,N_5740);
nor U8994 (N_8994,N_3405,N_5436);
xnor U8995 (N_8995,N_3527,N_5207);
or U8996 (N_8996,N_5039,N_3673);
xnor U8997 (N_8997,N_3635,N_5640);
xor U8998 (N_8998,N_4494,N_5069);
nand U8999 (N_8999,N_4688,N_4154);
and U9000 (N_9000,N_8504,N_8202);
and U9001 (N_9001,N_7945,N_7658);
and U9002 (N_9002,N_6701,N_7519);
and U9003 (N_9003,N_6567,N_8076);
nand U9004 (N_9004,N_8345,N_8502);
and U9005 (N_9005,N_7647,N_8271);
or U9006 (N_9006,N_7791,N_8252);
nor U9007 (N_9007,N_7286,N_8874);
xnor U9008 (N_9008,N_8259,N_6821);
nand U9009 (N_9009,N_8421,N_8021);
nor U9010 (N_9010,N_7645,N_8849);
xor U9011 (N_9011,N_8553,N_7199);
nor U9012 (N_9012,N_7513,N_6325);
nand U9013 (N_9013,N_6921,N_7481);
nand U9014 (N_9014,N_6077,N_8125);
xnor U9015 (N_9015,N_7242,N_7599);
xnor U9016 (N_9016,N_6303,N_8028);
nor U9017 (N_9017,N_8172,N_6984);
nand U9018 (N_9018,N_7902,N_7412);
and U9019 (N_9019,N_6496,N_8101);
nand U9020 (N_9020,N_7657,N_6495);
nor U9021 (N_9021,N_8393,N_6735);
and U9022 (N_9022,N_8280,N_7471);
nor U9023 (N_9023,N_8499,N_8639);
or U9024 (N_9024,N_7179,N_8495);
nor U9025 (N_9025,N_7121,N_8425);
nand U9026 (N_9026,N_8936,N_7558);
or U9027 (N_9027,N_6319,N_8550);
and U9028 (N_9028,N_8452,N_8012);
nand U9029 (N_9029,N_7730,N_7810);
and U9030 (N_9030,N_6071,N_6279);
or U9031 (N_9031,N_6963,N_8194);
or U9032 (N_9032,N_8337,N_7542);
or U9033 (N_9033,N_8303,N_6060);
nor U9034 (N_9034,N_6847,N_6753);
or U9035 (N_9035,N_7058,N_7014);
or U9036 (N_9036,N_7153,N_7280);
nand U9037 (N_9037,N_6056,N_7928);
or U9038 (N_9038,N_8606,N_7890);
and U9039 (N_9039,N_6273,N_7588);
nor U9040 (N_9040,N_7722,N_6391);
xor U9041 (N_9041,N_6783,N_8689);
or U9042 (N_9042,N_7719,N_6520);
xnor U9043 (N_9043,N_6591,N_8927);
nand U9044 (N_9044,N_8179,N_8363);
nor U9045 (N_9045,N_6212,N_6599);
or U9046 (N_9046,N_6021,N_8230);
nand U9047 (N_9047,N_8679,N_6517);
or U9048 (N_9048,N_7463,N_6888);
or U9049 (N_9049,N_6694,N_7566);
nand U9050 (N_9050,N_6018,N_6923);
and U9051 (N_9051,N_7414,N_8124);
xor U9052 (N_9052,N_8264,N_7649);
nand U9053 (N_9053,N_8435,N_7748);
and U9054 (N_9054,N_7825,N_7541);
nand U9055 (N_9055,N_6390,N_7528);
nor U9056 (N_9056,N_8890,N_6868);
or U9057 (N_9057,N_6014,N_6122);
nor U9058 (N_9058,N_7422,N_7630);
nor U9059 (N_9059,N_8070,N_8098);
and U9060 (N_9060,N_6399,N_7025);
and U9061 (N_9061,N_6320,N_6815);
xnor U9062 (N_9062,N_6543,N_8790);
or U9063 (N_9063,N_6975,N_7036);
nor U9064 (N_9064,N_6779,N_8901);
or U9065 (N_9065,N_6778,N_6628);
and U9066 (N_9066,N_8919,N_6463);
xnor U9067 (N_9067,N_8604,N_7064);
or U9068 (N_9068,N_8103,N_7336);
or U9069 (N_9069,N_8857,N_6448);
or U9070 (N_9070,N_6756,N_6149);
or U9071 (N_9071,N_7554,N_8605);
and U9072 (N_9072,N_8294,N_8488);
or U9073 (N_9073,N_7237,N_6811);
or U9074 (N_9074,N_7339,N_6434);
or U9075 (N_9075,N_6968,N_7456);
nor U9076 (N_9076,N_8327,N_6416);
nor U9077 (N_9077,N_8834,N_8400);
and U9078 (N_9078,N_8551,N_8150);
nor U9079 (N_9079,N_8462,N_7869);
or U9080 (N_9080,N_7778,N_7202);
and U9081 (N_9081,N_8286,N_7685);
and U9082 (N_9082,N_8586,N_6950);
nand U9083 (N_9083,N_6177,N_8626);
and U9084 (N_9084,N_7849,N_6057);
nand U9085 (N_9085,N_8977,N_8965);
nor U9086 (N_9086,N_6262,N_7495);
nand U9087 (N_9087,N_6015,N_6394);
or U9088 (N_9088,N_8422,N_6827);
and U9089 (N_9089,N_6108,N_8651);
or U9090 (N_9090,N_6803,N_8732);
and U9091 (N_9091,N_6630,N_6314);
nor U9092 (N_9092,N_6876,N_7430);
or U9093 (N_9093,N_6079,N_8270);
or U9094 (N_9094,N_7668,N_7054);
nand U9095 (N_9095,N_6248,N_6220);
or U9096 (N_9096,N_6493,N_6267);
and U9097 (N_9097,N_8723,N_6016);
nand U9098 (N_9098,N_6310,N_7538);
or U9099 (N_9099,N_6557,N_7671);
nor U9100 (N_9100,N_7888,N_7651);
and U9101 (N_9101,N_8968,N_8596);
nand U9102 (N_9102,N_7874,N_8691);
and U9103 (N_9103,N_8443,N_8432);
or U9104 (N_9104,N_8290,N_6252);
nor U9105 (N_9105,N_6810,N_7881);
and U9106 (N_9106,N_6441,N_6569);
nor U9107 (N_9107,N_8917,N_6937);
or U9108 (N_9108,N_8897,N_6193);
nor U9109 (N_9109,N_8001,N_6622);
or U9110 (N_9110,N_7909,N_7401);
nor U9111 (N_9111,N_7355,N_7589);
nor U9112 (N_9112,N_7823,N_6405);
xor U9113 (N_9113,N_8372,N_7906);
and U9114 (N_9114,N_6996,N_7619);
or U9115 (N_9115,N_8380,N_8269);
or U9116 (N_9116,N_6052,N_6710);
xnor U9117 (N_9117,N_6788,N_6846);
nor U9118 (N_9118,N_7806,N_8835);
and U9119 (N_9119,N_6328,N_7992);
or U9120 (N_9120,N_8705,N_6718);
or U9121 (N_9121,N_7785,N_8141);
and U9122 (N_9122,N_6908,N_8126);
or U9123 (N_9123,N_7260,N_7988);
nor U9124 (N_9124,N_8559,N_6476);
or U9125 (N_9125,N_6955,N_7073);
and U9126 (N_9126,N_6420,N_6528);
nand U9127 (N_9127,N_6263,N_8880);
or U9128 (N_9128,N_6832,N_7451);
nor U9129 (N_9129,N_7195,N_8404);
nand U9130 (N_9130,N_8644,N_7290);
nand U9131 (N_9131,N_7109,N_6335);
and U9132 (N_9132,N_8715,N_7374);
and U9133 (N_9133,N_6137,N_8884);
and U9134 (N_9134,N_6489,N_6726);
xnor U9135 (N_9135,N_6171,N_8784);
xor U9136 (N_9136,N_7027,N_6411);
nor U9137 (N_9137,N_7600,N_8780);
or U9138 (N_9138,N_8584,N_6118);
xor U9139 (N_9139,N_8506,N_6227);
nor U9140 (N_9140,N_7830,N_8189);
nand U9141 (N_9141,N_6451,N_8467);
nand U9142 (N_9142,N_6860,N_6259);
nand U9143 (N_9143,N_7099,N_8240);
nor U9144 (N_9144,N_6749,N_8456);
nor U9145 (N_9145,N_7230,N_6112);
or U9146 (N_9146,N_6045,N_8091);
nand U9147 (N_9147,N_6764,N_6854);
nand U9148 (N_9148,N_7532,N_8077);
and U9149 (N_9149,N_6813,N_8044);
nor U9150 (N_9150,N_8489,N_7434);
nor U9151 (N_9151,N_6902,N_8468);
and U9152 (N_9152,N_6246,N_7580);
nand U9153 (N_9153,N_8397,N_7677);
or U9154 (N_9154,N_8867,N_6419);
nand U9155 (N_9155,N_6047,N_7104);
nand U9156 (N_9156,N_8072,N_8951);
nand U9157 (N_9157,N_7498,N_7922);
nor U9158 (N_9158,N_8318,N_7643);
and U9159 (N_9159,N_6090,N_6017);
or U9160 (N_9160,N_7585,N_7060);
nor U9161 (N_9161,N_8576,N_6377);
nor U9162 (N_9162,N_7586,N_8983);
or U9163 (N_9163,N_6992,N_7026);
nand U9164 (N_9164,N_6928,N_8587);
nand U9165 (N_9165,N_7170,N_6871);
nand U9166 (N_9166,N_6671,N_8075);
and U9167 (N_9167,N_7937,N_7051);
and U9168 (N_9168,N_8683,N_6147);
and U9169 (N_9169,N_7112,N_6487);
and U9170 (N_9170,N_6432,N_6229);
or U9171 (N_9171,N_6375,N_7961);
or U9172 (N_9172,N_6799,N_8094);
or U9173 (N_9173,N_8210,N_6761);
and U9174 (N_9174,N_6022,N_6930);
and U9175 (N_9175,N_7892,N_8907);
and U9176 (N_9176,N_8619,N_6596);
nand U9177 (N_9177,N_6197,N_7614);
nand U9178 (N_9178,N_7946,N_8307);
xor U9179 (N_9179,N_6505,N_8391);
nor U9180 (N_9180,N_6070,N_7682);
xor U9181 (N_9181,N_7052,N_8356);
and U9182 (N_9182,N_6877,N_7860);
nor U9183 (N_9183,N_6673,N_6115);
nor U9184 (N_9184,N_6576,N_8281);
or U9185 (N_9185,N_7088,N_8967);
xnor U9186 (N_9186,N_7033,N_6893);
nand U9187 (N_9187,N_6750,N_7145);
xor U9188 (N_9188,N_8184,N_8537);
nand U9189 (N_9189,N_6953,N_8810);
or U9190 (N_9190,N_8726,N_8825);
and U9191 (N_9191,N_6833,N_6550);
or U9192 (N_9192,N_8065,N_8038);
and U9193 (N_9193,N_8417,N_7844);
nand U9194 (N_9194,N_7704,N_6474);
and U9195 (N_9195,N_6105,N_6379);
or U9196 (N_9196,N_6793,N_8196);
and U9197 (N_9197,N_8465,N_6980);
xnor U9198 (N_9198,N_6317,N_6271);
and U9199 (N_9199,N_8292,N_7159);
nand U9200 (N_9200,N_8326,N_7505);
nor U9201 (N_9201,N_6402,N_8197);
nand U9202 (N_9202,N_7009,N_6538);
or U9203 (N_9203,N_6480,N_7897);
nand U9204 (N_9204,N_6678,N_7255);
nor U9205 (N_9205,N_6770,N_6195);
and U9206 (N_9206,N_6425,N_7267);
or U9207 (N_9207,N_7817,N_6798);
nand U9208 (N_9208,N_6777,N_8058);
nand U9209 (N_9209,N_6703,N_7470);
nand U9210 (N_9210,N_7572,N_6527);
and U9211 (N_9211,N_7822,N_6027);
and U9212 (N_9212,N_7512,N_7592);
nor U9213 (N_9213,N_8446,N_6362);
nand U9214 (N_9214,N_8224,N_7072);
nor U9215 (N_9215,N_6397,N_8416);
nand U9216 (N_9216,N_6326,N_6019);
nand U9217 (N_9217,N_6180,N_8128);
and U9218 (N_9218,N_7217,N_7755);
or U9219 (N_9219,N_7919,N_8974);
or U9220 (N_9220,N_8140,N_7689);
nand U9221 (N_9221,N_6958,N_7150);
or U9222 (N_9222,N_7871,N_6597);
or U9223 (N_9223,N_7077,N_7085);
or U9224 (N_9224,N_7916,N_7969);
nand U9225 (N_9225,N_6670,N_6545);
and U9226 (N_9226,N_8132,N_8831);
nor U9227 (N_9227,N_7421,N_7587);
or U9228 (N_9228,N_8568,N_6780);
nor U9229 (N_9229,N_8785,N_8144);
nand U9230 (N_9230,N_7898,N_8673);
and U9231 (N_9231,N_6625,N_8401);
or U9232 (N_9232,N_8203,N_8932);
and U9233 (N_9233,N_8820,N_6007);
xor U9234 (N_9234,N_8105,N_7761);
and U9235 (N_9235,N_8807,N_7924);
or U9236 (N_9236,N_6169,N_6393);
nor U9237 (N_9237,N_6605,N_6521);
and U9238 (N_9238,N_6892,N_6037);
and U9239 (N_9239,N_7577,N_7269);
nand U9240 (N_9240,N_6824,N_6305);
nor U9241 (N_9241,N_6348,N_7758);
or U9242 (N_9242,N_6618,N_6050);
nor U9243 (N_9243,N_8390,N_6296);
and U9244 (N_9244,N_6743,N_8593);
nand U9245 (N_9245,N_8242,N_8866);
and U9246 (N_9246,N_7034,N_8888);
xor U9247 (N_9247,N_8876,N_8585);
and U9248 (N_9248,N_6737,N_7624);
nand U9249 (N_9249,N_8655,N_8061);
nor U9250 (N_9250,N_7131,N_8321);
nor U9251 (N_9251,N_6188,N_8449);
nor U9252 (N_9252,N_7674,N_6525);
nor U9253 (N_9253,N_8153,N_7895);
and U9254 (N_9254,N_7189,N_7661);
or U9255 (N_9255,N_8082,N_8274);
or U9256 (N_9256,N_6174,N_7807);
xor U9257 (N_9257,N_6617,N_8178);
xnor U9258 (N_9258,N_7363,N_6251);
nor U9259 (N_9259,N_8209,N_6454);
nand U9260 (N_9260,N_7763,N_8223);
nand U9261 (N_9261,N_6429,N_7876);
and U9262 (N_9262,N_7067,N_6554);
nand U9263 (N_9263,N_8768,N_6604);
or U9264 (N_9264,N_7057,N_6791);
nand U9265 (N_9265,N_8433,N_8622);
or U9266 (N_9266,N_8842,N_8751);
xnor U9267 (N_9267,N_8323,N_7894);
nor U9268 (N_9268,N_7493,N_6140);
and U9269 (N_9269,N_8067,N_7246);
and U9270 (N_9270,N_8746,N_7344);
and U9271 (N_9271,N_6106,N_6082);
or U9272 (N_9272,N_7773,N_8385);
or U9273 (N_9273,N_8000,N_7819);
or U9274 (N_9274,N_8332,N_8913);
or U9275 (N_9275,N_6184,N_8675);
nand U9276 (N_9276,N_7662,N_8251);
nor U9277 (N_9277,N_8371,N_7116);
nor U9278 (N_9278,N_6991,N_8250);
and U9279 (N_9279,N_6468,N_6960);
nand U9280 (N_9280,N_7450,N_8118);
xor U9281 (N_9281,N_8032,N_7990);
xnor U9282 (N_9282,N_6616,N_7068);
nor U9283 (N_9283,N_7136,N_8163);
nor U9284 (N_9284,N_8826,N_8187);
and U9285 (N_9285,N_8361,N_8764);
and U9286 (N_9286,N_8343,N_8561);
nor U9287 (N_9287,N_7602,N_7779);
or U9288 (N_9288,N_7347,N_7211);
and U9289 (N_9289,N_8515,N_8309);
nor U9290 (N_9290,N_8472,N_8466);
xnor U9291 (N_9291,N_8518,N_6512);
or U9292 (N_9292,N_6818,N_6318);
or U9293 (N_9293,N_8293,N_7163);
or U9294 (N_9294,N_7385,N_7288);
nand U9295 (N_9295,N_6152,N_6688);
nor U9296 (N_9296,N_7155,N_8633);
or U9297 (N_9297,N_6068,N_8713);
nand U9298 (N_9298,N_6843,N_6638);
and U9299 (N_9299,N_6182,N_7837);
and U9300 (N_9300,N_7023,N_8582);
or U9301 (N_9301,N_6336,N_6542);
or U9302 (N_9302,N_6654,N_6054);
or U9303 (N_9303,N_6594,N_7375);
nand U9304 (N_9304,N_7555,N_6461);
and U9305 (N_9305,N_7277,N_8516);
nor U9306 (N_9306,N_7501,N_6502);
xor U9307 (N_9307,N_7413,N_6927);
nand U9308 (N_9308,N_7606,N_6974);
nand U9309 (N_9309,N_7356,N_8228);
nand U9310 (N_9310,N_7846,N_6931);
nor U9311 (N_9311,N_8903,N_6136);
or U9312 (N_9312,N_8775,N_8761);
and U9313 (N_9313,N_6484,N_6825);
nand U9314 (N_9314,N_7843,N_8154);
and U9315 (N_9315,N_7490,N_8454);
nand U9316 (N_9316,N_6219,N_8064);
nand U9317 (N_9317,N_7194,N_6933);
and U9318 (N_9318,N_6396,N_6615);
or U9319 (N_9319,N_8860,N_6154);
nor U9320 (N_9320,N_6245,N_6883);
nand U9321 (N_9321,N_7573,N_6181);
nor U9322 (N_9322,N_7642,N_6210);
nor U9323 (N_9323,N_6922,N_6870);
or U9324 (N_9324,N_6342,N_8868);
nor U9325 (N_9325,N_7182,N_6460);
or U9326 (N_9326,N_7582,N_7103);
or U9327 (N_9327,N_8226,N_6413);
or U9328 (N_9328,N_6566,N_6491);
xnor U9329 (N_9329,N_8025,N_8700);
nand U9330 (N_9330,N_8944,N_7521);
nor U9331 (N_9331,N_8737,N_8672);
nand U9332 (N_9332,N_6947,N_6849);
xnor U9333 (N_9333,N_7929,N_6697);
or U9334 (N_9334,N_7842,N_6059);
nand U9335 (N_9335,N_7313,N_7133);
or U9336 (N_9336,N_7623,N_7087);
nand U9337 (N_9337,N_6672,N_8352);
or U9338 (N_9338,N_8182,N_8912);
and U9339 (N_9339,N_6561,N_7224);
nand U9340 (N_9340,N_7388,N_6510);
and U9341 (N_9341,N_6661,N_7066);
or U9342 (N_9342,N_6266,N_8762);
xnor U9343 (N_9343,N_7708,N_7633);
nor U9344 (N_9344,N_8015,N_8262);
nand U9345 (N_9345,N_6041,N_7128);
and U9346 (N_9346,N_8086,N_8265);
nor U9347 (N_9347,N_8946,N_8883);
nand U9348 (N_9348,N_8313,N_6530);
nand U9349 (N_9349,N_8523,N_7256);
nand U9350 (N_9350,N_8734,N_8996);
or U9351 (N_9351,N_7265,N_7648);
xnor U9352 (N_9352,N_8354,N_7002);
nand U9353 (N_9353,N_8317,N_6952);
nor U9354 (N_9354,N_6498,N_8003);
and U9355 (N_9355,N_8779,N_8632);
and U9356 (N_9356,N_7770,N_7850);
nand U9357 (N_9357,N_7010,N_6686);
or U9358 (N_9358,N_6848,N_8666);
or U9359 (N_9359,N_8546,N_6675);
xor U9360 (N_9360,N_7784,N_8685);
xnor U9361 (N_9361,N_6986,N_6053);
nor U9362 (N_9362,N_7438,N_8589);
nor U9363 (N_9363,N_7972,N_7392);
and U9364 (N_9364,N_6095,N_8459);
nor U9365 (N_9365,N_7613,N_6702);
nor U9366 (N_9366,N_8056,N_6819);
nand U9367 (N_9367,N_6745,N_6157);
nand U9368 (N_9368,N_7764,N_8512);
xnor U9369 (N_9369,N_8073,N_8167);
nor U9370 (N_9370,N_7973,N_7035);
nor U9371 (N_9371,N_6570,N_6709);
xor U9372 (N_9372,N_8852,N_7877);
and U9373 (N_9373,N_7759,N_7122);
or U9374 (N_9374,N_7040,N_8158);
nor U9375 (N_9375,N_6005,N_6636);
and U9376 (N_9376,N_8957,N_6398);
nand U9377 (N_9377,N_8279,N_7458);
nor U9378 (N_9378,N_6715,N_6354);
or U9379 (N_9379,N_8009,N_7631);
xor U9380 (N_9380,N_6533,N_6064);
and U9381 (N_9381,N_8902,N_7251);
xnor U9382 (N_9382,N_8846,N_7183);
nand U9383 (N_9383,N_6565,N_8724);
or U9384 (N_9384,N_6339,N_7132);
xnor U9385 (N_9385,N_6150,N_8205);
xor U9386 (N_9386,N_8319,N_7681);
and U9387 (N_9387,N_6728,N_8096);
and U9388 (N_9388,N_8249,N_6903);
or U9389 (N_9389,N_6073,N_7640);
xnor U9390 (N_9390,N_7612,N_7208);
and U9391 (N_9391,N_8148,N_6312);
or U9392 (N_9392,N_6404,N_8749);
nand U9393 (N_9393,N_6055,N_7031);
and U9394 (N_9394,N_6131,N_6741);
xnor U9395 (N_9395,N_7177,N_7792);
and U9396 (N_9396,N_6250,N_7905);
nor U9397 (N_9397,N_8641,N_7095);
nand U9398 (N_9398,N_8398,N_8816);
nor U9399 (N_9399,N_7149,N_6641);
nand U9400 (N_9400,N_8873,N_6198);
nor U9401 (N_9401,N_6967,N_6657);
xor U9402 (N_9402,N_8198,N_6524);
nor U9403 (N_9403,N_8207,N_6293);
nand U9404 (N_9404,N_6300,N_7571);
nor U9405 (N_9405,N_8438,N_8680);
nor U9406 (N_9406,N_7598,N_6916);
or U9407 (N_9407,N_7976,N_8068);
and U9408 (N_9408,N_8862,N_8110);
and U9409 (N_9409,N_6444,N_6241);
nand U9410 (N_9410,N_6024,N_6719);
nor U9411 (N_9411,N_8538,N_8419);
nand U9412 (N_9412,N_6869,N_8199);
nand U9413 (N_9413,N_6361,N_6101);
nor U9414 (N_9414,N_8953,N_8299);
and U9415 (N_9415,N_6817,N_6886);
or U9416 (N_9416,N_7728,N_6584);
and U9417 (N_9417,N_6985,N_7565);
and U9418 (N_9418,N_7169,N_6117);
or U9419 (N_9419,N_6286,N_7480);
nand U9420 (N_9420,N_6176,N_7100);
and U9421 (N_9421,N_7848,N_8282);
xnor U9422 (N_9422,N_6532,N_8099);
nor U9423 (N_9423,N_8778,N_7167);
and U9424 (N_9424,N_6431,N_8253);
and U9425 (N_9425,N_8349,N_8809);
or U9426 (N_9426,N_6768,N_8239);
and U9427 (N_9427,N_7814,N_8827);
nor U9428 (N_9428,N_8336,N_8706);
and U9429 (N_9429,N_8678,N_7574);
nor U9430 (N_9430,N_8838,N_8402);
and U9431 (N_9431,N_6679,N_8273);
nand U9432 (N_9432,N_8413,N_7694);
or U9433 (N_9433,N_8601,N_6836);
nor U9434 (N_9434,N_8513,N_8915);
or U9435 (N_9435,N_6765,N_6588);
or U9436 (N_9436,N_8029,N_8630);
nand U9437 (N_9437,N_6573,N_6544);
and U9438 (N_9438,N_7882,N_6882);
xnor U9439 (N_9439,N_7464,N_8939);
nand U9440 (N_9440,N_6951,N_6546);
and U9441 (N_9441,N_6013,N_7098);
or U9442 (N_9442,N_6729,N_7611);
and U9443 (N_9443,N_8389,N_7717);
and U9444 (N_9444,N_6043,N_8989);
and U9445 (N_9445,N_6653,N_8916);
nand U9446 (N_9446,N_8865,N_6168);
nand U9447 (N_9447,N_8844,N_8578);
xor U9448 (N_9448,N_7084,N_7408);
and U9449 (N_9449,N_7774,N_8514);
xor U9450 (N_9450,N_8079,N_7366);
nand U9451 (N_9451,N_7552,N_6478);
and U9452 (N_9452,N_7944,N_7338);
nand U9453 (N_9453,N_8366,N_8934);
and U9454 (N_9454,N_8621,N_8027);
or U9455 (N_9455,N_8374,N_6580);
nand U9456 (N_9456,N_6255,N_6352);
nor U9457 (N_9457,N_8213,N_6215);
nand U9458 (N_9458,N_7457,N_8174);
and U9459 (N_9459,N_6374,N_6156);
nand U9460 (N_9460,N_6809,N_8129);
or U9461 (N_9461,N_6134,N_8486);
nand U9462 (N_9462,N_7665,N_8219);
nor U9463 (N_9463,N_6072,N_7446);
nand U9464 (N_9464,N_6917,N_7912);
nand U9465 (N_9465,N_6976,N_7735);
nor U9466 (N_9466,N_6295,N_7931);
nand U9467 (N_9467,N_7680,N_8333);
and U9468 (N_9468,N_6757,N_6069);
or U9469 (N_9469,N_7402,N_7380);
and U9470 (N_9470,N_6660,N_7731);
and U9471 (N_9471,N_6065,N_6587);
or U9472 (N_9472,N_6471,N_7635);
and U9473 (N_9473,N_8288,N_6627);
nor U9474 (N_9474,N_8221,N_7678);
and U9475 (N_9475,N_8891,N_6620);
and U9476 (N_9476,N_6682,N_6107);
and U9477 (N_9477,N_7274,N_6001);
xnor U9478 (N_9478,N_6839,N_6531);
nand U9479 (N_9479,N_7516,N_7839);
nor U9480 (N_9480,N_6595,N_7325);
nand U9481 (N_9481,N_8696,N_8926);
nand U9482 (N_9482,N_7497,N_8699);
or U9483 (N_9483,N_6746,N_8526);
nand U9484 (N_9484,N_7080,N_8440);
nand U9485 (N_9485,N_7377,N_8853);
and U9486 (N_9486,N_7423,N_8010);
and U9487 (N_9487,N_7301,N_6924);
xnor U9488 (N_9488,N_7768,N_7790);
or U9489 (N_9489,N_7016,N_7711);
nor U9490 (N_9490,N_6285,N_7569);
or U9491 (N_9491,N_7082,N_6277);
nand U9492 (N_9492,N_8961,N_7448);
or U9493 (N_9493,N_7901,N_8115);
nor U9494 (N_9494,N_6631,N_8690);
or U9495 (N_9495,N_8415,N_7296);
and U9496 (N_9496,N_8405,N_6635);
or U9497 (N_9497,N_7621,N_6455);
and U9498 (N_9498,N_6206,N_8954);
or U9499 (N_9499,N_6600,N_8276);
nand U9500 (N_9500,N_6945,N_7370);
or U9501 (N_9501,N_7854,N_6380);
nand U9502 (N_9502,N_7117,N_6943);
nand U9503 (N_9503,N_6674,N_6051);
nor U9504 (N_9504,N_8471,N_7171);
nand U9505 (N_9505,N_8436,N_6861);
nand U9506 (N_9506,N_6837,N_6619);
or U9507 (N_9507,N_7397,N_7013);
or U9508 (N_9508,N_8930,N_6733);
nand U9509 (N_9509,N_7734,N_8671);
nor U9510 (N_9510,N_6164,N_8870);
or U9511 (N_9511,N_8171,N_6540);
and U9512 (N_9512,N_7838,N_6831);
nor U9513 (N_9513,N_6372,N_8758);
and U9514 (N_9514,N_8896,N_6829);
nand U9515 (N_9515,N_7632,N_7015);
nor U9516 (N_9516,N_6677,N_8485);
nand U9517 (N_9517,N_7174,N_7856);
nor U9518 (N_9518,N_7308,N_8406);
nand U9519 (N_9519,N_8815,N_7204);
nor U9520 (N_9520,N_8060,N_8730);
nand U9521 (N_9521,N_7297,N_6033);
or U9522 (N_9522,N_8200,N_7028);
or U9523 (N_9523,N_7878,N_6564);
nor U9524 (N_9524,N_7479,N_7568);
or U9525 (N_9525,N_6754,N_8407);
and U9526 (N_9526,N_7326,N_7382);
nor U9527 (N_9527,N_6151,N_6170);
xor U9528 (N_9528,N_8709,N_8367);
nand U9529 (N_9529,N_7815,N_7652);
xor U9530 (N_9530,N_7921,N_7219);
or U9531 (N_9531,N_6091,N_7889);
nor U9532 (N_9532,N_6324,N_6822);
and U9533 (N_9533,N_7861,N_7168);
nor U9534 (N_9534,N_7176,N_7281);
xnor U9535 (N_9535,N_8940,N_7210);
and U9536 (N_9536,N_8947,N_6359);
or U9537 (N_9537,N_6349,N_7736);
nand U9538 (N_9538,N_6522,N_8135);
and U9539 (N_9539,N_7707,N_7886);
and U9540 (N_9540,N_8763,N_8695);
nand U9541 (N_9541,N_6655,N_7579);
nor U9542 (N_9542,N_6997,N_7941);
nand U9543 (N_9543,N_8972,N_7322);
and U9544 (N_9544,N_8987,N_7918);
nand U9545 (N_9545,N_6563,N_8937);
nor U9546 (N_9546,N_7469,N_7386);
nor U9547 (N_9547,N_6488,N_6987);
nand U9548 (N_9548,N_6284,N_6651);
or U9549 (N_9549,N_8920,N_6485);
xor U9550 (N_9550,N_7192,N_8752);
nor U9551 (N_9551,N_6370,N_8905);
and U9552 (N_9552,N_8581,N_8591);
nand U9553 (N_9553,N_7746,N_8134);
xnor U9554 (N_9554,N_6887,N_6915);
nand U9555 (N_9555,N_7804,N_6479);
nand U9556 (N_9556,N_8295,N_8772);
nor U9557 (N_9557,N_8636,N_6972);
nand U9558 (N_9558,N_7517,N_6256);
nor U9559 (N_9559,N_6683,N_8160);
nor U9560 (N_9560,N_8002,N_7314);
nand U9561 (N_9561,N_7445,N_8575);
nand U9562 (N_9562,N_7346,N_7190);
or U9563 (N_9563,N_6023,N_8225);
nor U9564 (N_9564,N_8991,N_7597);
or U9565 (N_9565,N_8611,N_7995);
xnor U9566 (N_9566,N_8748,N_8681);
or U9567 (N_9567,N_8237,N_7323);
and U9568 (N_9568,N_7917,N_7670);
nand U9569 (N_9569,N_8770,N_6239);
and U9570 (N_9570,N_8640,N_6637);
xor U9571 (N_9571,N_6738,N_7315);
or U9572 (N_9572,N_6012,N_6592);
nand U9573 (N_9573,N_8886,N_8052);
xnor U9574 (N_9574,N_7750,N_8244);
nor U9575 (N_9575,N_7244,N_6503);
nor U9576 (N_9576,N_6078,N_8133);
and U9577 (N_9577,N_7557,N_7319);
nand U9578 (N_9578,N_6841,N_6360);
or U9579 (N_9579,N_6353,N_8268);
or U9580 (N_9580,N_8508,N_7903);
nor U9581 (N_9581,N_6513,N_6418);
or U9582 (N_9582,N_7559,N_6690);
xor U9583 (N_9583,N_6130,N_8647);
nand U9584 (N_9584,N_8353,N_8744);
or U9585 (N_9585,N_6119,N_8981);
nor U9586 (N_9586,N_6744,N_7723);
and U9587 (N_9587,N_7324,N_8439);
xor U9588 (N_9588,N_6648,N_8477);
and U9589 (N_9589,N_6036,N_8137);
or U9590 (N_9590,N_6684,N_8973);
nand U9591 (N_9591,N_6534,N_7684);
nor U9592 (N_9592,N_7884,N_6890);
xnor U9593 (N_9593,N_7486,N_8102);
or U9594 (N_9594,N_7766,N_7616);
or U9595 (N_9595,N_7115,N_8193);
nand U9596 (N_9596,N_6747,N_8756);
or U9597 (N_9597,N_8817,N_8423);
xnor U9598 (N_9598,N_6500,N_8121);
nor U9599 (N_9599,N_6447,N_6196);
or U9600 (N_9600,N_6965,N_6581);
and U9601 (N_9601,N_8453,N_7958);
nand U9602 (N_9602,N_6662,N_7799);
xor U9603 (N_9603,N_7553,N_6389);
xor U9604 (N_9604,N_6804,N_8801);
xor U9605 (N_9605,N_7818,N_7855);
or U9606 (N_9606,N_7415,N_6203);
nor U9607 (N_9607,N_8832,N_6946);
nand U9608 (N_9608,N_6127,N_7212);
xor U9609 (N_9609,N_7709,N_7872);
nand U9610 (N_9610,N_6010,N_6233);
xor U9611 (N_9611,N_8434,N_8161);
or U9612 (N_9612,N_6378,N_6066);
xnor U9613 (N_9613,N_7775,N_6640);
and U9614 (N_9614,N_8994,N_8175);
nor U9615 (N_9615,N_8008,N_6649);
nand U9616 (N_9616,N_7518,N_7537);
nand U9617 (N_9617,N_6548,N_7820);
xnor U9618 (N_9618,N_8168,N_7429);
nand U9619 (N_9619,N_8821,N_7690);
xnor U9620 (N_9620,N_6769,N_8177);
and U9621 (N_9621,N_7046,N_7828);
nand U9622 (N_9622,N_7904,N_7341);
nor U9623 (N_9623,N_7596,N_8564);
nand U9624 (N_9624,N_8600,N_6509);
or U9625 (N_9625,N_8236,N_6593);
nand U9626 (N_9626,N_6748,N_6042);
xor U9627 (N_9627,N_8738,N_7357);
nor U9628 (N_9628,N_7294,N_8754);
and U9629 (N_9629,N_6794,N_8487);
nor U9630 (N_9630,N_6853,N_8041);
nor U9631 (N_9631,N_6321,N_6458);
or U9632 (N_9632,N_7259,N_6141);
nand U9633 (N_9633,N_7811,N_8788);
and U9634 (N_9634,N_7911,N_7113);
and U9635 (N_9635,N_8505,N_7700);
and U9636 (N_9636,N_6891,N_7691);
or U9637 (N_9637,N_8045,N_7556);
and U9638 (N_9638,N_6650,N_7548);
or U9639 (N_9639,N_6322,N_8653);
or U9640 (N_9640,N_6820,N_7419);
nor U9641 (N_9641,N_8509,N_6632);
or U9642 (N_9642,N_7368,N_8005);
nor U9643 (N_9643,N_8481,N_7835);
and U9644 (N_9644,N_7226,N_7459);
nand U9645 (N_9645,N_7130,N_7012);
nor U9646 (N_9646,N_8583,N_7173);
or U9647 (N_9647,N_7732,N_8712);
and U9648 (N_9648,N_6506,N_7782);
and U9649 (N_9649,N_8069,N_6940);
nand U9650 (N_9650,N_8714,N_6183);
and U9651 (N_9651,N_8802,N_6920);
xor U9652 (N_9652,N_6878,N_7261);
and U9653 (N_9653,N_6237,N_7982);
and U9654 (N_9654,N_6061,N_6687);
xnor U9655 (N_9655,N_8324,N_8652);
or U9656 (N_9656,N_6449,N_7638);
nand U9657 (N_9657,N_7011,N_7654);
or U9658 (N_9658,N_6428,N_8348);
or U9659 (N_9659,N_8424,N_6583);
xor U9660 (N_9660,N_7800,N_7348);
xnor U9661 (N_9661,N_7999,N_6280);
and U9662 (N_9662,N_8037,N_8624);
nor U9663 (N_9663,N_7942,N_6961);
nor U9664 (N_9664,N_7047,N_7161);
nand U9665 (N_9665,N_8580,N_8941);
or U9666 (N_9666,N_8612,N_6708);
xor U9667 (N_9667,N_7545,N_8095);
nor U9668 (N_9668,N_8183,N_8074);
or U9669 (N_9669,N_7997,N_8463);
and U9670 (N_9670,N_6166,N_7634);
nand U9671 (N_9671,N_7740,N_7186);
and U9672 (N_9672,N_6739,N_8717);
or U9673 (N_9673,N_7048,N_8854);
nor U9674 (N_9674,N_8617,N_6230);
and U9675 (N_9675,N_6035,N_8990);
and U9676 (N_9676,N_6421,N_7966);
or U9677 (N_9677,N_7305,N_8054);
nor U9678 (N_9678,N_7824,N_8034);
and U9679 (N_9679,N_8662,N_6347);
nand U9680 (N_9680,N_8043,N_6483);
nand U9681 (N_9681,N_6302,N_6939);
and U9682 (N_9682,N_8190,N_6165);
and U9683 (N_9683,N_8750,N_7989);
and U9684 (N_9684,N_6213,N_7417);
and U9685 (N_9685,N_7225,N_7510);
and U9686 (N_9686,N_8808,N_7468);
nor U9687 (N_9687,N_7178,N_7712);
nor U9688 (N_9688,N_6242,N_8450);
nand U9689 (N_9689,N_8195,N_8603);
nor U9690 (N_9690,N_8569,N_8962);
or U9691 (N_9691,N_7243,N_7795);
nand U9692 (N_9692,N_7393,N_6406);
nor U9693 (N_9693,N_7968,N_8759);
nor U9694 (N_9694,N_7108,N_7070);
nand U9695 (N_9695,N_6291,N_7461);
or U9696 (N_9696,N_7306,N_6062);
or U9697 (N_9697,N_8080,N_8757);
nor U9698 (N_9698,N_6423,N_7583);
nand U9699 (N_9699,N_6132,N_7857);
and U9700 (N_9700,N_8684,N_7832);
and U9701 (N_9701,N_7959,N_6707);
and U9702 (N_9702,N_8322,N_8992);
nand U9703 (N_9703,N_8006,N_8496);
and U9704 (N_9704,N_6459,N_6232);
and U9705 (N_9705,N_7776,N_7499);
nand U9706 (N_9706,N_8985,N_7008);
nand U9707 (N_9707,N_8176,N_8263);
nor U9708 (N_9708,N_7193,N_6899);
or U9709 (N_9709,N_8162,N_8192);
nor U9710 (N_9710,N_8929,N_6081);
nor U9711 (N_9711,N_7913,N_8057);
nand U9712 (N_9712,N_6556,N_6201);
nand U9713 (N_9713,N_6858,N_8016);
or U9714 (N_9714,N_8386,N_8260);
nand U9715 (N_9715,N_7093,N_6977);
nor U9716 (N_9716,N_6004,N_6789);
or U9717 (N_9717,N_8186,N_8688);
and U9718 (N_9718,N_8476,N_7851);
or U9719 (N_9719,N_6333,N_8243);
nand U9720 (N_9720,N_8721,N_7692);
nor U9721 (N_9721,N_6124,N_7949);
xnor U9722 (N_9722,N_6514,N_8229);
or U9723 (N_9723,N_8528,N_6482);
nand U9724 (N_9724,N_6547,N_7134);
and U9725 (N_9725,N_8794,N_8649);
nor U9726 (N_9726,N_6752,N_6161);
xor U9727 (N_9727,N_8351,N_8682);
or U9728 (N_9728,N_7829,N_8786);
and U9729 (N_9729,N_8039,N_7687);
nor U9730 (N_9730,N_6272,N_8165);
nor U9731 (N_9731,N_7157,N_7936);
nor U9732 (N_9732,N_7641,N_8590);
and U9733 (N_9733,N_7866,N_6247);
or U9734 (N_9734,N_7221,N_7191);
nand U9735 (N_9735,N_8216,N_8618);
nand U9736 (N_9736,N_7042,N_6038);
and U9737 (N_9737,N_7258,N_8933);
nand U9738 (N_9738,N_8011,N_7547);
nand U9739 (N_9739,N_6995,N_6403);
xor U9740 (N_9740,N_8898,N_8441);
nand U9741 (N_9741,N_6466,N_6721);
or U9742 (N_9742,N_8791,N_7520);
and U9743 (N_9743,N_8517,N_8800);
and U9744 (N_9744,N_7432,N_7669);
and U9745 (N_9745,N_8558,N_6585);
or U9746 (N_9746,N_6656,N_6881);
or U9747 (N_9747,N_7805,N_7729);
or U9748 (N_9748,N_7345,N_8623);
nand U9749 (N_9749,N_8375,N_8152);
or U9750 (N_9750,N_6962,N_6551);
and U9751 (N_9751,N_7358,N_7387);
or U9752 (N_9752,N_6541,N_8733);
nand U9753 (N_9753,N_6113,N_8339);
or U9754 (N_9754,N_8157,N_7865);
nand U9755 (N_9755,N_8799,N_7710);
nand U9756 (N_9756,N_6712,N_7551);
and U9757 (N_9757,N_7934,N_8863);
xor U9758 (N_9758,N_7276,N_7151);
and U9759 (N_9759,N_8277,N_7119);
nand U9760 (N_9760,N_8097,N_8208);
or U9761 (N_9761,N_7715,N_7252);
or U9762 (N_9762,N_7650,N_8627);
nor U9763 (N_9763,N_6103,N_6763);
nor U9764 (N_9764,N_8869,N_6417);
nor U9765 (N_9765,N_6442,N_8945);
xor U9766 (N_9766,N_6722,N_8480);
or U9767 (N_9767,N_6555,N_8048);
nor U9768 (N_9768,N_8218,N_7460);
nor U9769 (N_9769,N_7576,N_6109);
or U9770 (N_9770,N_8725,N_7744);
and U9771 (N_9771,N_6190,N_7549);
nor U9772 (N_9772,N_8491,N_8119);
nor U9773 (N_9773,N_7816,N_6214);
and U9774 (N_9774,N_7821,N_6194);
and U9775 (N_9775,N_7786,N_6135);
nand U9776 (N_9776,N_6146,N_7777);
nand U9777 (N_9777,N_6412,N_7299);
nand U9778 (N_9778,N_6261,N_7796);
nand U9779 (N_9779,N_8078,N_7318);
nor U9780 (N_9780,N_8494,N_6942);
nand U9781 (N_9781,N_7714,N_6453);
nand U9782 (N_9782,N_8437,N_8461);
nor U9783 (N_9783,N_7974,N_6189);
xor U9784 (N_9784,N_7188,N_8531);
nor U9785 (N_9785,N_8878,N_6910);
nor U9786 (N_9786,N_8858,N_7769);
nand U9787 (N_9787,N_7270,N_7462);
xor U9788 (N_9788,N_7235,N_7747);
nor U9789 (N_9789,N_7209,N_8819);
or U9790 (N_9790,N_6249,N_8573);
nor U9791 (N_9791,N_6304,N_8871);
nor U9792 (N_9792,N_8776,N_8830);
nand U9793 (N_9793,N_7410,N_7262);
xor U9794 (N_9794,N_8539,N_6774);
and U9795 (N_9795,N_8740,N_7765);
or U9796 (N_9796,N_8824,N_7091);
and U9797 (N_9797,N_6634,N_6574);
nor U9798 (N_9798,N_8050,N_6639);
nand U9799 (N_9799,N_7655,N_6204);
or U9800 (N_9800,N_8117,N_8597);
xnor U9801 (N_9801,N_6936,N_7328);
and U9802 (N_9802,N_8492,N_7952);
nor U9803 (N_9803,N_8116,N_6185);
nor U9804 (N_9804,N_6260,N_7017);
nor U9805 (N_9805,N_8241,N_8329);
nand U9806 (N_9806,N_6758,N_6094);
and U9807 (N_9807,N_8533,N_6138);
nor U9808 (N_9808,N_7158,N_8022);
nand U9809 (N_9809,N_8112,N_6435);
and U9810 (N_9810,N_8837,N_8151);
xor U9811 (N_9811,N_6606,N_6087);
or U9812 (N_9812,N_8409,N_8217);
or U9813 (N_9813,N_6734,N_6730);
xnor U9814 (N_9814,N_7594,N_8377);
nand U9815 (N_9815,N_8718,N_7311);
or U9816 (N_9816,N_7672,N_8365);
nand U9817 (N_9817,N_8143,N_7331);
nor U9818 (N_9818,N_7138,N_6120);
or U9819 (N_9819,N_8572,N_6497);
nand U9820 (N_9820,N_6499,N_6796);
and U9821 (N_9821,N_7213,N_8342);
and U9822 (N_9822,N_8031,N_8544);
xnor U9823 (N_9823,N_7404,N_6373);
or U9824 (N_9824,N_6560,N_7231);
and U9825 (N_9825,N_6046,N_7751);
nand U9826 (N_9826,N_6844,N_6376);
nor U9827 (N_9827,N_6327,N_7601);
and U9828 (N_9828,N_6918,N_8731);
or U9829 (N_9829,N_7074,N_7207);
or U9830 (N_9830,N_6225,N_8851);
xor U9831 (N_9831,N_7453,N_7227);
or U9832 (N_9832,N_8490,N_7907);
nor U9833 (N_9833,N_7673,N_7337);
nand U9834 (N_9834,N_7361,N_7019);
nand U9835 (N_9835,N_7407,N_8287);
or U9836 (N_9836,N_6501,N_6647);
nand U9837 (N_9837,N_6211,N_8845);
and U9838 (N_9838,N_7376,N_6623);
xnor U9839 (N_9839,N_6075,N_7218);
or U9840 (N_9840,N_8571,N_6098);
and U9841 (N_9841,N_8997,N_8474);
nand U9842 (N_9842,N_6209,N_6786);
nor U9843 (N_9843,N_8448,N_6422);
or U9844 (N_9844,N_7492,N_7840);
xnor U9845 (N_9845,N_8093,N_7487);
and U9846 (N_9846,N_6669,N_6299);
and U9847 (N_9847,N_6981,N_7291);
nor U9848 (N_9848,N_7004,N_7249);
and U9849 (N_9849,N_6784,N_7625);
and U9850 (N_9850,N_6695,N_7496);
nor U9851 (N_9851,N_8334,N_8999);
and U9852 (N_9852,N_8661,N_8298);
nand U9853 (N_9853,N_7762,N_6971);
nand U9854 (N_9854,N_6614,N_6572);
or U9855 (N_9855,N_7426,N_8180);
and U9856 (N_9856,N_8975,N_7530);
nor U9857 (N_9857,N_7196,N_6693);
nand U9858 (N_9858,N_7214,N_6367);
xnor U9859 (N_9859,N_7420,N_7365);
or U9860 (N_9860,N_8071,N_8444);
nor U9861 (N_9861,N_6257,N_8475);
nand U9862 (N_9862,N_6332,N_7351);
or U9863 (N_9863,N_8795,N_6275);
xnor U9864 (N_9864,N_6601,N_8500);
and U9865 (N_9865,N_8191,N_8812);
or U9866 (N_9866,N_8359,N_7232);
or U9867 (N_9867,N_8727,N_6607);
or U9868 (N_9868,N_6290,N_6486);
nor U9869 (N_9869,N_6516,N_7847);
nand U9870 (N_9870,N_8501,N_7564);
and U9871 (N_9871,N_7515,N_6477);
or U9872 (N_9872,N_6009,N_6395);
nor U9873 (N_9873,N_7140,N_6452);
nor U9874 (N_9874,N_7124,N_8956);
nor U9875 (N_9875,N_7923,N_7491);
nor U9876 (N_9876,N_8331,N_6329);
nor U9877 (N_9877,N_8092,N_8521);
nor U9878 (N_9878,N_6470,N_7639);
xnor U9879 (N_9879,N_8382,N_8395);
nand U9880 (N_9880,N_7720,N_7627);
or U9881 (N_9881,N_6092,N_6885);
nor U9882 (N_9882,N_6828,N_6159);
xnor U9883 (N_9883,N_7476,N_7914);
nand U9884 (N_9884,N_8470,N_8928);
nor U9885 (N_9885,N_7303,N_6571);
or U9886 (N_9886,N_6254,N_8145);
or U9887 (N_9887,N_6663,N_8634);
nor U9888 (N_9888,N_7398,N_6911);
nor U9889 (N_9889,N_7135,N_6313);
and U9890 (N_9890,N_8650,N_8484);
nor U9891 (N_9891,N_7247,N_7287);
and U9892 (N_9892,N_6802,N_7925);
or U9893 (N_9893,N_6949,N_8767);
or U9894 (N_9894,N_7215,N_7022);
or U9895 (N_9895,N_7676,N_7220);
nor U9896 (N_9896,N_7079,N_7043);
or U9897 (N_9897,N_7697,N_7440);
and U9898 (N_9898,N_8789,N_8257);
nor U9899 (N_9899,N_6199,N_6288);
nand U9900 (N_9900,N_7275,N_8960);
or U9901 (N_9901,N_6287,N_8411);
nor U9902 (N_9902,N_6970,N_6906);
and U9903 (N_9903,N_7646,N_6202);
nand U9904 (N_9904,N_8328,N_8798);
nand U9905 (N_9905,N_8894,N_6044);
and U9906 (N_9906,N_6643,N_8525);
or U9907 (N_9907,N_8004,N_7321);
nand U9908 (N_9908,N_7984,N_8686);
nand U9909 (N_9909,N_7059,N_8935);
and U9910 (N_9910,N_7834,N_8955);
or U9911 (N_9911,N_6830,N_7529);
and U9912 (N_9912,N_8950,N_8783);
nor U9913 (N_9913,N_8657,N_7742);
nor U9914 (N_9914,N_8055,N_6856);
or U9915 (N_9915,N_8510,N_8777);
and U9916 (N_9916,N_8173,N_6755);
xnor U9917 (N_9917,N_7561,N_7142);
or U9918 (N_9918,N_7005,N_6099);
or U9919 (N_9919,N_8900,N_7536);
nor U9920 (N_9920,N_8155,N_8577);
or U9921 (N_9921,N_6652,N_6704);
xor U9922 (N_9922,N_6067,N_6392);
and U9923 (N_9923,N_8879,N_8548);
or U9924 (N_9924,N_7793,N_8833);
xor U9925 (N_9925,N_7605,N_6366);
nand U9926 (N_9926,N_8412,N_8017);
or U9927 (N_9927,N_7724,N_8146);
xor U9928 (N_9928,N_6384,N_7038);
nor U9929 (N_9929,N_8669,N_8392);
xnor U9930 (N_9930,N_7926,N_7075);
or U9931 (N_9931,N_8676,N_6433);
nor U9932 (N_9932,N_7637,N_7893);
and U9933 (N_9933,N_7935,N_6696);
or U9934 (N_9934,N_7411,N_8147);
nand U9935 (N_9935,N_6030,N_7300);
nor U9936 (N_9936,N_6668,N_7757);
and U9937 (N_9937,N_8308,N_7273);
xor U9938 (N_9938,N_7981,N_8910);
nor U9939 (N_9939,N_6446,N_6034);
nand U9940 (N_9940,N_7439,N_8729);
and U9941 (N_9941,N_8410,N_8373);
nand U9942 (N_9942,N_6731,N_7384);
and U9943 (N_9943,N_7978,N_8836);
and U9944 (N_9944,N_8013,N_8289);
nand U9945 (N_9945,N_6895,N_6025);
and U9946 (N_9946,N_8036,N_8984);
nand U9947 (N_9947,N_6553,N_7248);
nor U9948 (N_9948,N_7910,N_7030);
xnor U9949 (N_9949,N_6350,N_8261);
nand U9950 (N_9950,N_8949,N_8018);
nand U9951 (N_9951,N_7474,N_8566);
nor U9952 (N_9952,N_6385,N_7360);
and U9953 (N_9953,N_6223,N_7745);
or U9954 (N_9954,N_6806,N_7436);
nand U9955 (N_9955,N_8166,N_7041);
nor U9956 (N_9956,N_8291,N_7663);
nor U9957 (N_9957,N_7603,N_7437);
nand U9958 (N_9958,N_6982,N_7760);
nor U9959 (N_9959,N_6129,N_6969);
nor U9960 (N_9960,N_7029,N_7332);
or U9961 (N_9961,N_7879,N_8087);
xor U9962 (N_9962,N_8364,N_7044);
nor U9963 (N_9963,N_7932,N_7915);
nand U9964 (N_9964,N_6253,N_8245);
nor U9965 (N_9965,N_7550,N_8340);
nor U9966 (N_9966,N_8275,N_7695);
nand U9967 (N_9967,N_7263,N_8083);
or U9968 (N_9968,N_6880,N_6148);
nand U9969 (N_9969,N_6011,N_6494);
or U9970 (N_9970,N_7097,N_8549);
nand U9971 (N_9971,N_8310,N_7139);
or U9972 (N_9972,N_6387,N_8963);
nor U9973 (N_9973,N_6472,N_7431);
nand U9974 (N_9974,N_6031,N_7378);
nand U9975 (N_9975,N_8084,N_8659);
or U9976 (N_9976,N_7409,N_6408);
or U9977 (N_9977,N_6355,N_8532);
nand U9978 (N_9978,N_8704,N_7101);
and U9979 (N_9979,N_8895,N_8227);
or U9980 (N_9980,N_7285,N_6427);
nor U9981 (N_9981,N_6155,N_7198);
or U9982 (N_9982,N_7143,N_7160);
and U9983 (N_9983,N_7660,N_6481);
or U9984 (N_9984,N_8524,N_8881);
or U9985 (N_9985,N_7092,N_6613);
or U9986 (N_9986,N_7049,N_6340);
and U9987 (N_9987,N_7688,N_6598);
nor U9988 (N_9988,N_6282,N_8616);
nor U9989 (N_9989,N_8608,N_7359);
and U9990 (N_9990,N_6088,N_8106);
and U9991 (N_9991,N_7123,N_7125);
or U9992 (N_9992,N_8429,N_8529);
nand U9993 (N_9993,N_6954,N_6897);
nand U9994 (N_9994,N_8760,N_6879);
or U9995 (N_9995,N_6518,N_6989);
xor U9996 (N_9996,N_8381,N_8703);
nor U9997 (N_9997,N_8427,N_7021);
or U9998 (N_9998,N_6192,N_8847);
or U9999 (N_9999,N_6032,N_6988);
nor U10000 (N_10000,N_8958,N_7399);
xor U10001 (N_10001,N_8545,N_6771);
nor U10002 (N_10002,N_7086,N_8445);
nand U10003 (N_10003,N_8020,N_7316);
nor U10004 (N_10004,N_7102,N_6093);
or U10005 (N_10005,N_7078,N_6872);
and U10006 (N_10006,N_6691,N_6139);
or U10007 (N_10007,N_7527,N_8822);
nand U10008 (N_10008,N_7504,N_6834);
or U10009 (N_10009,N_8948,N_6226);
nand U10010 (N_10010,N_8687,N_6175);
or U10011 (N_10011,N_6244,N_7772);
xor U10012 (N_10012,N_6121,N_7575);
or U10013 (N_10013,N_6178,N_7870);
nand U10014 (N_10014,N_7703,N_8302);
and U10015 (N_10015,N_7743,N_6665);
or U10016 (N_10016,N_6706,N_8362);
or U10017 (N_10017,N_6998,N_8766);
nand U10018 (N_10018,N_7506,N_7753);
xnor U10019 (N_10019,N_7787,N_6040);
and U10020 (N_10020,N_6633,N_6646);
or U10021 (N_10021,N_7896,N_8993);
and U10022 (N_10022,N_6450,N_6698);
and U10023 (N_10023,N_8442,N_8850);
nand U10024 (N_10024,N_6102,N_7543);
nor U10025 (N_10025,N_6383,N_6205);
or U10026 (N_10026,N_6283,N_8399);
xor U10027 (N_10027,N_8387,N_8478);
nand U10028 (N_10028,N_7333,N_7696);
and U10029 (N_10029,N_7175,N_7234);
or U10030 (N_10030,N_7292,N_6440);
xnor U10031 (N_10031,N_8774,N_7197);
and U10032 (N_10032,N_6705,N_8909);
nor U10033 (N_10033,N_7257,N_6048);
nand U10034 (N_10034,N_7478,N_6801);
xnor U10035 (N_10035,N_6862,N_6875);
and U10036 (N_10036,N_8278,N_7686);
nor U10037 (N_10037,N_8710,N_8320);
and U10038 (N_10038,N_8797,N_8388);
nand U10039 (N_10039,N_8266,N_6983);
nand U10040 (N_10040,N_7024,N_7570);
nor U10041 (N_10041,N_8966,N_8511);
and U10042 (N_10042,N_8376,N_7228);
xor U10043 (N_10043,N_6457,N_7617);
nor U10044 (N_10044,N_8698,N_7391);
nor U10045 (N_10045,N_8358,N_8893);
and U10046 (N_10046,N_6944,N_6867);
or U10047 (N_10047,N_6941,N_8745);
nor U10048 (N_10048,N_8610,N_8875);
and U10049 (N_10049,N_6492,N_7885);
xor U10050 (N_10050,N_7418,N_8120);
and U10051 (N_10051,N_7141,N_7381);
and U10052 (N_10052,N_7063,N_8579);
nand U10053 (N_10053,N_6003,N_7433);
and U10054 (N_10054,N_7442,N_7636);
and U10055 (N_10055,N_6179,N_8557);
and U10056 (N_10056,N_8908,N_7526);
and U10057 (N_10057,N_6465,N_7546);
and U10058 (N_10058,N_8394,N_6128);
or U10059 (N_10059,N_7452,N_7607);
or U10060 (N_10060,N_8024,N_8663);
and U10061 (N_10061,N_7309,N_7137);
and U10062 (N_10062,N_8643,N_8355);
nand U10063 (N_10063,N_6823,N_6713);
nand U10064 (N_10064,N_7295,N_6111);
nand U10065 (N_10065,N_6711,N_7739);
and U10066 (N_10066,N_6368,N_8081);
nor U10067 (N_10067,N_7284,N_8460);
or U10068 (N_10068,N_8285,N_6577);
nand U10069 (N_10069,N_8231,N_6104);
nor U10070 (N_10070,N_6934,N_8931);
nor U10071 (N_10071,N_7693,N_7164);
and U10072 (N_10072,N_6873,N_6464);
and U10073 (N_10073,N_6508,N_6445);
and U10074 (N_10074,N_8925,N_7939);
and U10075 (N_10075,N_6097,N_8464);
nand U10076 (N_10076,N_7081,N_8995);
nand U10077 (N_10077,N_7129,N_7500);
nor U10078 (N_10078,N_8628,N_8964);
xnor U10079 (N_10079,N_6959,N_7831);
nand U10080 (N_10080,N_7721,N_7482);
or U10081 (N_10081,N_6388,N_8677);
or U10082 (N_10082,N_7593,N_8062);
nand U10083 (N_10083,N_7511,N_7977);
or U10084 (N_10084,N_7335,N_6243);
nor U10085 (N_10085,N_7180,N_8887);
and U10086 (N_10086,N_6805,N_6716);
nor U10087 (N_10087,N_7618,N_7425);
or U10088 (N_10088,N_7447,N_6415);
or U10089 (N_10089,N_7615,N_6797);
or U10090 (N_10090,N_8457,N_6274);
and U10091 (N_10091,N_7389,N_6790);
or U10092 (N_10092,N_8877,N_8357);
nor U10093 (N_10093,N_7007,N_7726);
or U10094 (N_10094,N_7238,N_8418);
nand U10095 (N_10095,N_8497,N_6659);
and U10096 (N_10096,N_8814,N_8554);
and U10097 (N_10097,N_7118,N_7733);
or U10098 (N_10098,N_8547,N_7349);
and U10099 (N_10099,N_7354,N_8567);
and U10100 (N_10100,N_6990,N_8841);
nand U10101 (N_10101,N_7020,N_6490);
and U10102 (N_10102,N_6268,N_8565);
nand U10103 (N_10103,N_7522,N_7435);
nand U10104 (N_10104,N_7236,N_7996);
nor U10105 (N_10105,N_6889,N_8360);
or U10106 (N_10106,N_6238,N_7887);
nand U10107 (N_10107,N_6558,N_8090);
nor U10108 (N_10108,N_6371,N_6076);
nor U10109 (N_10109,N_8615,N_8848);
and U10110 (N_10110,N_7126,N_7970);
nand U10111 (N_10111,N_7390,N_6133);
xor U10112 (N_10112,N_7781,N_7154);
nand U10113 (N_10113,N_6343,N_6020);
xnor U10114 (N_10114,N_6049,N_8707);
xnor U10115 (N_10115,N_7334,N_6306);
or U10116 (N_10116,N_8127,N_8859);
nor U10117 (N_10117,N_6341,N_7679);
and U10118 (N_10118,N_8828,N_6381);
nand U10119 (N_10119,N_7987,N_8222);
nor U10120 (N_10120,N_7329,N_6767);
nand U10121 (N_10121,N_8536,N_7604);
nand U10122 (N_10122,N_8379,N_8638);
or U10123 (N_10123,N_7788,N_7524);
or U10124 (N_10124,N_8645,N_6430);
nor U10125 (N_10125,N_6162,N_7069);
xor U10126 (N_10126,N_8431,N_8769);
xnor U10127 (N_10127,N_8430,N_6143);
nand U10128 (N_10128,N_7938,N_6629);
nor U10129 (N_10129,N_8426,N_7864);
and U10130 (N_10130,N_6294,N_6224);
nor U10131 (N_10131,N_7254,N_7184);
or U10132 (N_10132,N_7089,N_6835);
nor U10133 (N_10133,N_8914,N_8316);
nand U10134 (N_10134,N_8765,N_7229);
and U10135 (N_10135,N_7373,N_6163);
and U10136 (N_10136,N_8451,N_6603);
and U10137 (N_10137,N_7953,N_8104);
nor U10138 (N_10138,N_6173,N_8131);
nand U10139 (N_10139,N_7975,N_6400);
or U10140 (N_10140,N_6278,N_6401);
or U10141 (N_10141,N_7394,N_7056);
nand U10142 (N_10142,N_6443,N_6409);
and U10143 (N_10143,N_6973,N_6852);
nor U10144 (N_10144,N_6913,N_8959);
or U10145 (N_10145,N_6863,N_6338);
and U10146 (N_10146,N_8033,N_8922);
nor U10147 (N_10147,N_8042,N_7675);
nand U10148 (N_10148,N_8384,N_6228);
nor U10149 (N_10149,N_7165,N_8743);
and U10150 (N_10150,N_6200,N_6307);
nor U10151 (N_10151,N_6167,N_6365);
and U10152 (N_10152,N_8212,N_7201);
and U10153 (N_10153,N_6218,N_7808);
and U10154 (N_10154,N_8206,N_7239);
nand U10155 (N_10155,N_7664,N_6281);
and U10156 (N_10156,N_8482,N_8297);
or U10157 (N_10157,N_6664,N_7455);
xor U10158 (N_10158,N_7798,N_6356);
nand U10159 (N_10159,N_7200,N_6787);
nor U10160 (N_10160,N_7827,N_8139);
nand U10161 (N_10161,N_7927,N_7006);
or U10162 (N_10162,N_8665,N_7350);
nand U10163 (N_10163,N_7037,N_6426);
or U10164 (N_10164,N_7312,N_7427);
nor U10165 (N_10165,N_8455,N_7473);
nor U10166 (N_10166,N_7899,N_7626);
nor U10167 (N_10167,N_8114,N_8635);
or U10168 (N_10168,N_8648,N_7863);
nand U10169 (N_10169,N_8108,N_6642);
or U10170 (N_10170,N_6114,N_8306);
or U10171 (N_10171,N_6058,N_6006);
xnor U10172 (N_10172,N_8560,N_7920);
or U10173 (N_10173,N_6187,N_7699);
and U10174 (N_10174,N_8805,N_8555);
and U10175 (N_10175,N_7282,N_7591);
nand U10176 (N_10176,N_7868,N_8602);
or U10177 (N_10177,N_6894,N_6345);
nor U10178 (N_10178,N_6901,N_8314);
or U10179 (N_10179,N_8796,N_7858);
nand U10180 (N_10180,N_6909,N_7342);
nand U10181 (N_10181,N_8414,N_7994);
nor U10182 (N_10182,N_7147,N_7279);
or U10183 (N_10183,N_8330,N_7756);
nor U10184 (N_10184,N_7383,N_6725);
nor U10185 (N_10185,N_6424,N_8138);
or U10186 (N_10186,N_7609,N_8370);
and U10187 (N_10187,N_7862,N_6626);
nand U10188 (N_10188,N_8856,N_8254);
or U10189 (N_10189,N_6158,N_7400);
and U10190 (N_10190,N_6938,N_7172);
and U10191 (N_10191,N_7562,N_7000);
nand U10192 (N_10192,N_6658,N_8818);
nor U10193 (N_10193,N_6144,N_7443);
and U10194 (N_10194,N_7653,N_8344);
or U10195 (N_10195,N_7659,N_8019);
nor U10196 (N_10196,N_7353,N_6568);
nor U10197 (N_10197,N_7628,N_7727);
nand U10198 (N_10198,N_6732,N_6994);
nor U10199 (N_10199,N_8978,N_6907);
nor U10200 (N_10200,N_7967,N_7055);
xor U10201 (N_10201,N_6002,N_7629);
or U10202 (N_10202,N_6978,N_7698);
nor U10203 (N_10203,N_8736,N_8540);
xnor U10204 (N_10204,N_8542,N_6851);
nand U10205 (N_10205,N_7960,N_7003);
nand U10206 (N_10206,N_8085,N_6153);
and U10207 (N_10207,N_7289,N_7780);
nand U10208 (N_10208,N_6612,N_6240);
or U10209 (N_10209,N_7485,N_8256);
nand U10210 (N_10210,N_8159,N_7071);
or U10211 (N_10211,N_6579,N_6515);
nor U10212 (N_10212,N_6826,N_7563);
or U10213 (N_10213,N_8595,N_8918);
nor U10214 (N_10214,N_6000,N_7250);
or U10215 (N_10215,N_7340,N_6912);
or U10216 (N_10216,N_7867,N_8035);
nand U10217 (N_10217,N_6610,N_6590);
or U10218 (N_10218,N_8267,N_7991);
and U10219 (N_10219,N_7107,N_6699);
or U10220 (N_10220,N_7610,N_8556);
nand U10221 (N_10221,N_6207,N_6504);
nand U10222 (N_10222,N_6582,N_6473);
or U10223 (N_10223,N_7622,N_8047);
nor U10224 (N_10224,N_7466,N_6331);
nand U10225 (N_10225,N_7754,N_6624);
nand U10226 (N_10226,N_7127,N_8971);
or U10227 (N_10227,N_8829,N_8629);
nand U10228 (N_10228,N_6186,N_7406);
nand U10229 (N_10229,N_6437,N_6759);
nand U10230 (N_10230,N_7203,N_8889);
nand U10231 (N_10231,N_6602,N_6334);
or U10232 (N_10232,N_6160,N_7114);
or U10233 (N_10233,N_7222,N_7971);
or U10234 (N_10234,N_7317,N_6838);
and U10235 (N_10235,N_8493,N_6549);
nand U10236 (N_10236,N_7253,N_7475);
and U10237 (N_10237,N_8026,N_7090);
nand U10238 (N_10238,N_8483,N_6315);
or U10239 (N_10239,N_7416,N_7880);
xor U10240 (N_10240,N_8613,N_6896);
and U10241 (N_10241,N_6083,N_6644);
and U10242 (N_10242,N_6776,N_7233);
nand U10243 (N_10243,N_6855,N_6932);
and U10244 (N_10244,N_6410,N_6258);
nor U10245 (N_10245,N_8541,N_8839);
and U10246 (N_10246,N_6865,N_6874);
or U10247 (N_10247,N_7836,N_7320);
nand U10248 (N_10248,N_8188,N_7801);
nand U10249 (N_10249,N_6364,N_6172);
nand U10250 (N_10250,N_6884,N_7930);
and U10251 (N_10251,N_8522,N_6234);
or U10252 (N_10252,N_8614,N_7144);
or U10253 (N_10253,N_8970,N_8988);
nor U10254 (N_10254,N_8719,N_7032);
or U10255 (N_10255,N_6269,N_6008);
or U10256 (N_10256,N_6816,N_7560);
or U10257 (N_10257,N_8315,N_8204);
or U10258 (N_10258,N_7245,N_7106);
or U10259 (N_10259,N_8169,N_6382);
nand U10260 (N_10260,N_7094,N_8892);
nor U10261 (N_10261,N_6919,N_6270);
nor U10262 (N_10262,N_6308,N_8692);
nor U10263 (N_10263,N_7797,N_6864);
nand U10264 (N_10264,N_6222,N_7396);
nor U10265 (N_10265,N_8051,N_7581);
xnor U10266 (N_10266,N_8864,N_6842);
nor U10267 (N_10267,N_7018,N_8943);
nor U10268 (N_10268,N_8469,N_6309);
nand U10269 (N_10269,N_8787,N_7985);
and U10270 (N_10270,N_8111,N_7957);
and U10271 (N_10271,N_8089,N_7185);
or U10272 (N_10272,N_7428,N_7152);
nand U10273 (N_10273,N_8164,N_6221);
and U10274 (N_10274,N_7705,N_8066);
or U10275 (N_10275,N_7364,N_6191);
or U10276 (N_10276,N_6084,N_7216);
nand U10277 (N_10277,N_8594,N_7472);
or U10278 (N_10278,N_7803,N_7813);
or U10279 (N_10279,N_8220,N_8234);
or U10280 (N_10280,N_8088,N_7535);
or U10281 (N_10281,N_7272,N_7534);
nor U10282 (N_10282,N_8170,N_7933);
nor U10283 (N_10283,N_8609,N_7713);
or U10284 (N_10284,N_7488,N_8040);
nor U10285 (N_10285,N_8693,N_7205);
nand U10286 (N_10286,N_6529,N_6814);
and U10287 (N_10287,N_8347,N_6438);
or U10288 (N_10288,N_8498,N_7950);
nor U10289 (N_10289,N_6609,N_6536);
and U10290 (N_10290,N_8899,N_8014);
or U10291 (N_10291,N_8702,N_7156);
nand U10292 (N_10292,N_8637,N_6301);
nand U10293 (N_10293,N_6526,N_6904);
nand U10294 (N_10294,N_7716,N_8300);
and U10295 (N_10295,N_7955,N_7741);
or U10296 (N_10296,N_7223,N_6929);
and U10297 (N_10297,N_7162,N_7531);
and U10298 (N_10298,N_6645,N_8708);
nor U10299 (N_10299,N_7484,N_8806);
nand U10300 (N_10300,N_8100,N_8296);
nand U10301 (N_10301,N_7900,N_8969);
and U10302 (N_10302,N_6344,N_7809);
nor U10303 (N_10303,N_6676,N_7369);
or U10304 (N_10304,N_8923,N_7367);
xnor U10305 (N_10305,N_6116,N_7110);
or U10306 (N_10306,N_6736,N_8535);
and U10307 (N_10307,N_8741,N_6812);
and U10308 (N_10308,N_6123,N_6926);
nor U10309 (N_10309,N_7302,N_8520);
nand U10310 (N_10310,N_8403,N_8771);
and U10311 (N_10311,N_8861,N_7187);
or U10312 (N_10312,N_7001,N_8755);
or U10313 (N_10313,N_8258,N_7525);
xor U10314 (N_10314,N_8952,N_6231);
and U10315 (N_10315,N_6781,N_7738);
nor U10316 (N_10316,N_8711,N_6539);
and U10317 (N_10317,N_8701,N_6956);
nand U10318 (N_10318,N_7268,N_7841);
or U10319 (N_10319,N_6772,N_7964);
or U10320 (N_10320,N_6762,N_7065);
nor U10321 (N_10321,N_6386,N_7053);
and U10322 (N_10322,N_7833,N_7352);
nand U10323 (N_10323,N_7330,N_8976);
nor U10324 (N_10324,N_6727,N_7372);
or U10325 (N_10325,N_8238,N_6742);
nor U10326 (N_10326,N_6145,N_7507);
and U10327 (N_10327,N_6800,N_6456);
and U10328 (N_10328,N_7062,N_8428);
xnor U10329 (N_10329,N_6519,N_8255);
and U10330 (N_10330,N_7523,N_7783);
or U10331 (N_10331,N_6898,N_8301);
xnor U10332 (N_10332,N_6957,N_7620);
nor U10333 (N_10333,N_8246,N_8046);
nor U10334 (N_10334,N_7166,N_7883);
or U10335 (N_10335,N_7307,N_6795);
nor U10336 (N_10336,N_7962,N_8855);
xnor U10337 (N_10337,N_8543,N_7590);
and U10338 (N_10338,N_7963,N_6407);
nand U10339 (N_10339,N_8813,N_8181);
nand U10340 (N_10340,N_7718,N_8793);
nand U10341 (N_10341,N_6724,N_7293);
and U10342 (N_10342,N_8396,N_7656);
nor U10343 (N_10343,N_6096,N_7477);
nor U10344 (N_10344,N_6357,N_8938);
nor U10345 (N_10345,N_6039,N_6216);
and U10346 (N_10346,N_7940,N_6782);
and U10347 (N_10347,N_7061,N_7111);
nor U10348 (N_10348,N_7533,N_7752);
nand U10349 (N_10349,N_8304,N_8063);
nand U10350 (N_10350,N_8911,N_6507);
xnor U10351 (N_10351,N_6845,N_6346);
and U10352 (N_10352,N_6792,N_6714);
and U10353 (N_10353,N_7424,N_7873);
nor U10354 (N_10354,N_8059,N_7852);
nand U10355 (N_10355,N_8023,N_8007);
nor U10356 (N_10356,N_7584,N_8534);
nand U10357 (N_10357,N_8942,N_8654);
nor U10358 (N_10358,N_8592,N_8747);
and U10359 (N_10359,N_7298,N_6766);
or U10360 (N_10360,N_8773,N_8674);
and U10361 (N_10361,N_7449,N_8185);
nor U10362 (N_10362,N_6264,N_8625);
nor U10363 (N_10363,N_7343,N_7206);
and U10364 (N_10364,N_6537,N_7812);
nor U10365 (N_10365,N_6323,N_8519);
or U10366 (N_10366,N_7240,N_8305);
nor U10367 (N_10367,N_8670,N_8697);
and U10368 (N_10368,N_7327,N_8843);
and U10369 (N_10369,N_6289,N_7509);
nand U10370 (N_10370,N_8420,N_7483);
and U10371 (N_10371,N_8473,N_7444);
nor U10372 (N_10372,N_7514,N_8503);
nor U10373 (N_10373,N_7405,N_7737);
or U10374 (N_10374,N_6700,N_6126);
nand U10375 (N_10375,N_6773,N_6578);
nor U10376 (N_10376,N_7794,N_8660);
nand U10377 (N_10377,N_7749,N_7702);
nor U10378 (N_10378,N_7826,N_7271);
nand U10379 (N_10379,N_7948,N_7083);
and U10380 (N_10380,N_7441,N_6086);
nor U10381 (N_10381,N_6074,N_7503);
nand U10382 (N_10382,N_6462,N_7667);
and U10383 (N_10383,N_8722,N_8479);
or U10384 (N_10384,N_8782,N_6298);
nand U10385 (N_10385,N_6063,N_7310);
and U10386 (N_10386,N_8350,N_6775);
nand U10387 (N_10387,N_7045,N_6723);
nand U10388 (N_10388,N_8904,N_6236);
and U10389 (N_10389,N_7540,N_6080);
nand U10390 (N_10390,N_6808,N_8840);
xnor U10391 (N_10391,N_7467,N_7489);
nor U10392 (N_10392,N_7465,N_6142);
and U10393 (N_10393,N_6689,N_8804);
nand U10394 (N_10394,N_6467,N_7039);
nor U10395 (N_10395,N_8980,N_6966);
nand U10396 (N_10396,N_8924,N_8201);
and U10397 (N_10397,N_8507,N_6511);
xor U10398 (N_10398,N_6311,N_6608);
nor U10399 (N_10399,N_8735,N_8109);
nor U10400 (N_10400,N_7403,N_8720);
and U10401 (N_10401,N_7146,N_6575);
and U10402 (N_10402,N_6692,N_7980);
and U10403 (N_10403,N_6085,N_6217);
and U10404 (N_10404,N_6026,N_8753);
nor U10405 (N_10405,N_6859,N_6363);
nor U10406 (N_10406,N_8232,N_8214);
nor U10407 (N_10407,N_7998,N_8325);
and U10408 (N_10408,N_8311,N_6586);
nor U10409 (N_10409,N_8122,N_7454);
and U10410 (N_10410,N_6589,N_6611);
nand U10411 (N_10411,N_7666,N_6439);
nor U10412 (N_10412,N_8781,N_8338);
or U10413 (N_10413,N_8742,N_6857);
nor U10414 (N_10414,N_6235,N_7379);
xnor U10415 (N_10415,N_8998,N_7395);
nand U10416 (N_10416,N_8107,N_8642);
nand U10417 (N_10417,N_7608,N_6469);
xnor U10418 (N_10418,N_7802,N_6208);
nand U10419 (N_10419,N_7264,N_7241);
nor U10420 (N_10420,N_7789,N_7148);
nand U10421 (N_10421,N_6751,N_8149);
and U10422 (N_10422,N_7050,N_8235);
or U10423 (N_10423,N_7567,N_6666);
and U10424 (N_10424,N_8211,N_6028);
and U10425 (N_10425,N_7578,N_8574);
xor U10426 (N_10426,N_7096,N_7859);
and U10427 (N_10427,N_6029,N_8136);
nor U10428 (N_10428,N_6276,N_8113);
and U10429 (N_10429,N_8335,N_7986);
nand U10430 (N_10430,N_6760,N_6993);
or U10431 (N_10431,N_7508,N_7539);
nor U10432 (N_10432,N_6351,N_8882);
or U10433 (N_10433,N_8215,N_8982);
nand U10434 (N_10434,N_8123,N_7266);
nand U10435 (N_10435,N_8130,N_6523);
xnor U10436 (N_10436,N_6925,N_7725);
or U10437 (N_10437,N_8142,N_6717);
nand U10438 (N_10438,N_6562,N_8607);
or U10439 (N_10439,N_8872,N_7908);
and U10440 (N_10440,N_7181,N_6089);
and U10441 (N_10441,N_6475,N_7875);
and U10442 (N_10442,N_7771,N_7105);
and U10443 (N_10443,N_8458,N_6866);
or U10444 (N_10444,N_6979,N_7120);
nand U10445 (N_10445,N_6680,N_8530);
and U10446 (N_10446,N_8383,N_8284);
nor U10447 (N_10447,N_6292,N_8885);
xor U10448 (N_10448,N_8620,N_6337);
nor U10449 (N_10449,N_6100,N_7983);
nand U10450 (N_10450,N_6935,N_7076);
and U10451 (N_10451,N_8716,N_7683);
and U10452 (N_10452,N_8408,N_8156);
and U10453 (N_10453,N_6840,N_6552);
or U10454 (N_10454,N_7951,N_8272);
and U10455 (N_10455,N_8341,N_7362);
and U10456 (N_10456,N_6414,N_7701);
xor U10457 (N_10457,N_8906,N_7278);
nand U10458 (N_10458,N_8368,N_8656);
and U10459 (N_10459,N_8588,N_7954);
nor U10460 (N_10460,N_6850,N_8646);
or U10461 (N_10461,N_8921,N_8247);
or U10462 (N_10462,N_7943,N_6785);
nor U10463 (N_10463,N_6125,N_6999);
nand U10464 (N_10464,N_8030,N_8631);
or U10465 (N_10465,N_7891,N_8283);
xnor U10466 (N_10466,N_6914,N_8811);
nand U10467 (N_10467,N_6535,N_6436);
nor U10468 (N_10468,N_7644,N_8739);
and U10469 (N_10469,N_7706,N_8312);
and U10470 (N_10470,N_6265,N_6559);
or U10471 (N_10471,N_8447,N_7965);
nor U10472 (N_10472,N_6900,N_7283);
and U10473 (N_10473,N_6964,N_8664);
or U10474 (N_10474,N_6948,N_6369);
and U10475 (N_10475,N_8527,N_8563);
and U10476 (N_10476,N_8378,N_8667);
or U10477 (N_10477,N_8049,N_8552);
nor U10478 (N_10478,N_7544,N_8053);
nor U10479 (N_10479,N_7371,N_8658);
and U10480 (N_10480,N_8668,N_7767);
xor U10481 (N_10481,N_8694,N_7993);
or U10482 (N_10482,N_6667,N_8248);
nand U10483 (N_10483,N_6720,N_6621);
or U10484 (N_10484,N_7947,N_8986);
or U10485 (N_10485,N_7956,N_8233);
or U10486 (N_10486,N_6297,N_6110);
nand U10487 (N_10487,N_7845,N_7502);
nor U10488 (N_10488,N_8979,N_8570);
xor U10489 (N_10489,N_6358,N_7494);
or U10490 (N_10490,N_6330,N_6681);
nor U10491 (N_10491,N_8792,N_6316);
and U10492 (N_10492,N_8599,N_7595);
nor U10493 (N_10493,N_7304,N_8803);
or U10494 (N_10494,N_6685,N_8369);
nor U10495 (N_10495,N_8598,N_8346);
or U10496 (N_10496,N_7979,N_6740);
nor U10497 (N_10497,N_8728,N_6905);
nand U10498 (N_10498,N_8562,N_7853);
xnor U10499 (N_10499,N_8823,N_6807);
nor U10500 (N_10500,N_7199,N_6255);
nor U10501 (N_10501,N_6395,N_6553);
or U10502 (N_10502,N_8245,N_6053);
or U10503 (N_10503,N_8456,N_7022);
nand U10504 (N_10504,N_6934,N_8582);
nor U10505 (N_10505,N_7709,N_7804);
nor U10506 (N_10506,N_7998,N_7392);
and U10507 (N_10507,N_7145,N_8800);
nor U10508 (N_10508,N_7837,N_6532);
or U10509 (N_10509,N_8736,N_6411);
nand U10510 (N_10510,N_7005,N_8568);
nor U10511 (N_10511,N_6009,N_6544);
nor U10512 (N_10512,N_7941,N_7591);
nor U10513 (N_10513,N_7624,N_8049);
nor U10514 (N_10514,N_7120,N_6930);
and U10515 (N_10515,N_7301,N_8810);
xnor U10516 (N_10516,N_6320,N_6114);
nand U10517 (N_10517,N_7801,N_6273);
nor U10518 (N_10518,N_6701,N_8781);
and U10519 (N_10519,N_8298,N_7462);
nor U10520 (N_10520,N_7768,N_7040);
and U10521 (N_10521,N_7857,N_8344);
nand U10522 (N_10522,N_8120,N_6901);
nor U10523 (N_10523,N_6495,N_7768);
and U10524 (N_10524,N_8806,N_8611);
nor U10525 (N_10525,N_8627,N_6938);
nand U10526 (N_10526,N_8410,N_7086);
or U10527 (N_10527,N_7411,N_8901);
nor U10528 (N_10528,N_8458,N_6820);
nor U10529 (N_10529,N_7786,N_7863);
nor U10530 (N_10530,N_8697,N_7523);
or U10531 (N_10531,N_7180,N_6160);
or U10532 (N_10532,N_7799,N_8117);
or U10533 (N_10533,N_8144,N_6764);
and U10534 (N_10534,N_8617,N_7430);
nand U10535 (N_10535,N_8091,N_6692);
and U10536 (N_10536,N_7964,N_8277);
and U10537 (N_10537,N_6028,N_8344);
nand U10538 (N_10538,N_8584,N_8788);
nand U10539 (N_10539,N_7735,N_6681);
and U10540 (N_10540,N_6454,N_7413);
nand U10541 (N_10541,N_8421,N_6994);
nand U10542 (N_10542,N_8896,N_6880);
and U10543 (N_10543,N_7801,N_8733);
or U10544 (N_10544,N_7487,N_8529);
or U10545 (N_10545,N_8020,N_6162);
and U10546 (N_10546,N_7009,N_6050);
nor U10547 (N_10547,N_8858,N_6751);
or U10548 (N_10548,N_6633,N_6970);
or U10549 (N_10549,N_6335,N_6812);
nand U10550 (N_10550,N_8132,N_6608);
and U10551 (N_10551,N_8157,N_7130);
or U10552 (N_10552,N_8912,N_7226);
and U10553 (N_10553,N_6850,N_6294);
nor U10554 (N_10554,N_6807,N_6448);
or U10555 (N_10555,N_7557,N_8861);
xnor U10556 (N_10556,N_8379,N_7202);
and U10557 (N_10557,N_8637,N_7019);
nor U10558 (N_10558,N_7740,N_7060);
nor U10559 (N_10559,N_8195,N_8213);
and U10560 (N_10560,N_8957,N_6707);
or U10561 (N_10561,N_8538,N_8504);
or U10562 (N_10562,N_7205,N_8756);
and U10563 (N_10563,N_8340,N_8641);
and U10564 (N_10564,N_6366,N_7526);
xnor U10565 (N_10565,N_8773,N_7872);
and U10566 (N_10566,N_8120,N_7419);
nand U10567 (N_10567,N_6108,N_7732);
nand U10568 (N_10568,N_6552,N_7230);
xor U10569 (N_10569,N_8901,N_7911);
or U10570 (N_10570,N_6893,N_6390);
nor U10571 (N_10571,N_8849,N_8132);
xor U10572 (N_10572,N_8115,N_7179);
nor U10573 (N_10573,N_6039,N_7772);
nand U10574 (N_10574,N_6125,N_8802);
or U10575 (N_10575,N_7269,N_6702);
or U10576 (N_10576,N_6463,N_7078);
nand U10577 (N_10577,N_6701,N_6633);
nand U10578 (N_10578,N_6487,N_6685);
xor U10579 (N_10579,N_6088,N_6789);
and U10580 (N_10580,N_6290,N_6274);
nand U10581 (N_10581,N_8771,N_6186);
or U10582 (N_10582,N_6042,N_6314);
nor U10583 (N_10583,N_8777,N_8810);
nand U10584 (N_10584,N_6300,N_7269);
or U10585 (N_10585,N_8448,N_8128);
nand U10586 (N_10586,N_6622,N_6314);
and U10587 (N_10587,N_6640,N_6448);
or U10588 (N_10588,N_7099,N_7031);
and U10589 (N_10589,N_6838,N_6400);
nand U10590 (N_10590,N_8249,N_8038);
nand U10591 (N_10591,N_7661,N_8831);
nand U10592 (N_10592,N_6340,N_6063);
and U10593 (N_10593,N_8526,N_6706);
or U10594 (N_10594,N_6608,N_7641);
xnor U10595 (N_10595,N_6769,N_6830);
nor U10596 (N_10596,N_6901,N_8576);
or U10597 (N_10597,N_8276,N_7289);
xor U10598 (N_10598,N_8467,N_8022);
nor U10599 (N_10599,N_7945,N_7840);
or U10600 (N_10600,N_7228,N_8490);
nor U10601 (N_10601,N_7935,N_7665);
and U10602 (N_10602,N_7509,N_7508);
nand U10603 (N_10603,N_6042,N_8762);
nand U10604 (N_10604,N_8716,N_8001);
nor U10605 (N_10605,N_6883,N_6967);
nand U10606 (N_10606,N_7984,N_6122);
nor U10607 (N_10607,N_8632,N_6999);
or U10608 (N_10608,N_7563,N_8688);
nand U10609 (N_10609,N_6985,N_7807);
nand U10610 (N_10610,N_8904,N_8449);
nor U10611 (N_10611,N_8692,N_7208);
nand U10612 (N_10612,N_6474,N_7356);
and U10613 (N_10613,N_6217,N_7443);
nor U10614 (N_10614,N_8781,N_6771);
or U10615 (N_10615,N_7469,N_7500);
xor U10616 (N_10616,N_8572,N_6074);
nor U10617 (N_10617,N_8694,N_7606);
xnor U10618 (N_10618,N_7213,N_6516);
or U10619 (N_10619,N_6358,N_8349);
xor U10620 (N_10620,N_8964,N_8315);
and U10621 (N_10621,N_8731,N_6040);
xnor U10622 (N_10622,N_6268,N_6667);
nor U10623 (N_10623,N_6310,N_6614);
xor U10624 (N_10624,N_7343,N_8524);
nor U10625 (N_10625,N_6604,N_7088);
nand U10626 (N_10626,N_6458,N_6157);
nor U10627 (N_10627,N_7338,N_8584);
xnor U10628 (N_10628,N_7062,N_8849);
xor U10629 (N_10629,N_8786,N_6187);
and U10630 (N_10630,N_6801,N_6385);
nand U10631 (N_10631,N_7605,N_8322);
xnor U10632 (N_10632,N_7919,N_8465);
nand U10633 (N_10633,N_6496,N_7889);
xor U10634 (N_10634,N_7219,N_6452);
nand U10635 (N_10635,N_6496,N_8009);
or U10636 (N_10636,N_6753,N_8647);
and U10637 (N_10637,N_7940,N_6305);
or U10638 (N_10638,N_7370,N_6620);
nor U10639 (N_10639,N_7757,N_6970);
or U10640 (N_10640,N_7988,N_8338);
xnor U10641 (N_10641,N_8716,N_7153);
nor U10642 (N_10642,N_8029,N_6215);
xor U10643 (N_10643,N_7516,N_8455);
nor U10644 (N_10644,N_6492,N_6364);
and U10645 (N_10645,N_8075,N_7463);
nor U10646 (N_10646,N_7639,N_7615);
or U10647 (N_10647,N_8882,N_6371);
nand U10648 (N_10648,N_7604,N_8720);
or U10649 (N_10649,N_7571,N_7780);
and U10650 (N_10650,N_6118,N_7201);
or U10651 (N_10651,N_7263,N_7065);
nor U10652 (N_10652,N_6329,N_8941);
nor U10653 (N_10653,N_6380,N_7083);
nand U10654 (N_10654,N_8710,N_6048);
xnor U10655 (N_10655,N_8914,N_6517);
or U10656 (N_10656,N_7412,N_6814);
nand U10657 (N_10657,N_7341,N_8646);
nor U10658 (N_10658,N_8894,N_8813);
nor U10659 (N_10659,N_8144,N_6427);
and U10660 (N_10660,N_6644,N_7855);
and U10661 (N_10661,N_8034,N_7966);
nor U10662 (N_10662,N_8998,N_6123);
and U10663 (N_10663,N_6468,N_6605);
nor U10664 (N_10664,N_8024,N_8964);
xnor U10665 (N_10665,N_8851,N_8670);
and U10666 (N_10666,N_8182,N_8997);
and U10667 (N_10667,N_8320,N_7591);
xnor U10668 (N_10668,N_8477,N_6833);
nand U10669 (N_10669,N_6760,N_8096);
nand U10670 (N_10670,N_7374,N_6682);
nand U10671 (N_10671,N_7893,N_8862);
nand U10672 (N_10672,N_7947,N_7888);
or U10673 (N_10673,N_7281,N_6559);
xnor U10674 (N_10674,N_8292,N_8589);
and U10675 (N_10675,N_8046,N_8308);
nand U10676 (N_10676,N_6623,N_7282);
and U10677 (N_10677,N_8369,N_7363);
or U10678 (N_10678,N_7793,N_7155);
or U10679 (N_10679,N_7511,N_6127);
or U10680 (N_10680,N_8217,N_8544);
xnor U10681 (N_10681,N_7300,N_6139);
nor U10682 (N_10682,N_6076,N_7497);
nand U10683 (N_10683,N_7203,N_7156);
or U10684 (N_10684,N_8002,N_8590);
and U10685 (N_10685,N_6843,N_6417);
and U10686 (N_10686,N_6603,N_6707);
xor U10687 (N_10687,N_8761,N_8971);
nor U10688 (N_10688,N_6279,N_6615);
and U10689 (N_10689,N_8650,N_8181);
nor U10690 (N_10690,N_7317,N_6004);
nand U10691 (N_10691,N_6665,N_8191);
nand U10692 (N_10692,N_8632,N_7958);
xnor U10693 (N_10693,N_8037,N_7892);
or U10694 (N_10694,N_6830,N_8496);
or U10695 (N_10695,N_7472,N_8931);
nor U10696 (N_10696,N_8606,N_7995);
nor U10697 (N_10697,N_7874,N_7569);
nand U10698 (N_10698,N_8363,N_7685);
and U10699 (N_10699,N_6288,N_8800);
or U10700 (N_10700,N_6903,N_7211);
nand U10701 (N_10701,N_6937,N_6597);
or U10702 (N_10702,N_7705,N_6998);
or U10703 (N_10703,N_6021,N_6597);
nor U10704 (N_10704,N_8104,N_6782);
and U10705 (N_10705,N_7936,N_8053);
or U10706 (N_10706,N_6874,N_8757);
or U10707 (N_10707,N_7786,N_8994);
and U10708 (N_10708,N_6040,N_6420);
or U10709 (N_10709,N_6252,N_8021);
or U10710 (N_10710,N_7348,N_8363);
and U10711 (N_10711,N_6015,N_8965);
or U10712 (N_10712,N_8350,N_6628);
and U10713 (N_10713,N_8062,N_8102);
xnor U10714 (N_10714,N_8830,N_8533);
xor U10715 (N_10715,N_6246,N_6947);
nor U10716 (N_10716,N_8548,N_6206);
nor U10717 (N_10717,N_7656,N_8324);
and U10718 (N_10718,N_8741,N_7948);
or U10719 (N_10719,N_6248,N_7333);
nand U10720 (N_10720,N_8889,N_7414);
nor U10721 (N_10721,N_8513,N_8334);
nor U10722 (N_10722,N_8045,N_6228);
nor U10723 (N_10723,N_7736,N_6612);
nand U10724 (N_10724,N_7030,N_7021);
nor U10725 (N_10725,N_7417,N_8042);
or U10726 (N_10726,N_8626,N_8835);
xor U10727 (N_10727,N_8991,N_6613);
nand U10728 (N_10728,N_7313,N_8230);
or U10729 (N_10729,N_8359,N_6225);
xnor U10730 (N_10730,N_6574,N_6373);
and U10731 (N_10731,N_7095,N_6445);
nand U10732 (N_10732,N_6240,N_8802);
nor U10733 (N_10733,N_8823,N_7434);
and U10734 (N_10734,N_6868,N_7244);
or U10735 (N_10735,N_8892,N_7826);
or U10736 (N_10736,N_7021,N_7357);
or U10737 (N_10737,N_8653,N_6439);
nand U10738 (N_10738,N_7881,N_7103);
and U10739 (N_10739,N_8839,N_6040);
or U10740 (N_10740,N_6636,N_8167);
nor U10741 (N_10741,N_7147,N_6159);
and U10742 (N_10742,N_8294,N_7679);
xor U10743 (N_10743,N_7202,N_7447);
and U10744 (N_10744,N_6414,N_8495);
nor U10745 (N_10745,N_8128,N_7732);
nor U10746 (N_10746,N_8323,N_7565);
and U10747 (N_10747,N_7465,N_6436);
nand U10748 (N_10748,N_7772,N_6608);
and U10749 (N_10749,N_8395,N_8523);
nand U10750 (N_10750,N_7376,N_7975);
nor U10751 (N_10751,N_8851,N_7674);
nand U10752 (N_10752,N_6378,N_6640);
nor U10753 (N_10753,N_8407,N_7480);
or U10754 (N_10754,N_7350,N_6530);
xor U10755 (N_10755,N_8357,N_6719);
nand U10756 (N_10756,N_6414,N_7691);
xnor U10757 (N_10757,N_8360,N_6774);
and U10758 (N_10758,N_8412,N_8922);
nand U10759 (N_10759,N_8970,N_6201);
or U10760 (N_10760,N_8682,N_7778);
nand U10761 (N_10761,N_8899,N_8565);
or U10762 (N_10762,N_8743,N_6687);
and U10763 (N_10763,N_6387,N_6097);
or U10764 (N_10764,N_7758,N_6863);
nor U10765 (N_10765,N_8399,N_6571);
nand U10766 (N_10766,N_7256,N_8139);
nor U10767 (N_10767,N_7940,N_6688);
nor U10768 (N_10768,N_7619,N_8275);
nand U10769 (N_10769,N_7363,N_7473);
nand U10770 (N_10770,N_8422,N_6989);
or U10771 (N_10771,N_8857,N_8674);
and U10772 (N_10772,N_7161,N_6384);
nand U10773 (N_10773,N_6990,N_8419);
or U10774 (N_10774,N_8412,N_6350);
and U10775 (N_10775,N_6111,N_8621);
nand U10776 (N_10776,N_7905,N_6881);
and U10777 (N_10777,N_7660,N_6143);
nor U10778 (N_10778,N_6527,N_6822);
or U10779 (N_10779,N_8197,N_8431);
nand U10780 (N_10780,N_7630,N_6287);
and U10781 (N_10781,N_7432,N_6275);
nand U10782 (N_10782,N_6222,N_6197);
nor U10783 (N_10783,N_7514,N_8064);
nand U10784 (N_10784,N_6962,N_7523);
or U10785 (N_10785,N_7952,N_6280);
nand U10786 (N_10786,N_7908,N_7554);
nand U10787 (N_10787,N_7662,N_7388);
nand U10788 (N_10788,N_8620,N_8244);
or U10789 (N_10789,N_8424,N_6834);
nand U10790 (N_10790,N_8485,N_6487);
nor U10791 (N_10791,N_6461,N_7309);
or U10792 (N_10792,N_6261,N_6587);
or U10793 (N_10793,N_8675,N_8738);
or U10794 (N_10794,N_8657,N_6606);
nand U10795 (N_10795,N_8214,N_6341);
nor U10796 (N_10796,N_6503,N_6048);
nor U10797 (N_10797,N_7322,N_8231);
xnor U10798 (N_10798,N_6212,N_7136);
and U10799 (N_10799,N_6363,N_7328);
nor U10800 (N_10800,N_6644,N_8591);
or U10801 (N_10801,N_7249,N_7410);
nor U10802 (N_10802,N_7350,N_7314);
xor U10803 (N_10803,N_6211,N_7820);
and U10804 (N_10804,N_7618,N_6931);
nand U10805 (N_10805,N_7336,N_7609);
nand U10806 (N_10806,N_7872,N_8256);
or U10807 (N_10807,N_7881,N_7486);
xnor U10808 (N_10808,N_8712,N_6757);
or U10809 (N_10809,N_6424,N_7296);
nor U10810 (N_10810,N_7739,N_7007);
and U10811 (N_10811,N_6316,N_8203);
nand U10812 (N_10812,N_8840,N_8430);
or U10813 (N_10813,N_6109,N_6196);
xnor U10814 (N_10814,N_8817,N_8812);
xnor U10815 (N_10815,N_6695,N_8224);
nand U10816 (N_10816,N_8068,N_7647);
nand U10817 (N_10817,N_7631,N_8558);
and U10818 (N_10818,N_7594,N_7940);
nand U10819 (N_10819,N_6516,N_6717);
and U10820 (N_10820,N_7312,N_6781);
xnor U10821 (N_10821,N_7874,N_6540);
nor U10822 (N_10822,N_7755,N_7873);
nand U10823 (N_10823,N_8730,N_7068);
and U10824 (N_10824,N_8751,N_7072);
nor U10825 (N_10825,N_7854,N_7221);
nor U10826 (N_10826,N_7964,N_7212);
or U10827 (N_10827,N_8884,N_8652);
nand U10828 (N_10828,N_6190,N_6381);
nand U10829 (N_10829,N_6602,N_6148);
nor U10830 (N_10830,N_8603,N_7260);
or U10831 (N_10831,N_6158,N_6352);
or U10832 (N_10832,N_7840,N_6811);
xnor U10833 (N_10833,N_7633,N_7459);
xnor U10834 (N_10834,N_8677,N_7414);
or U10835 (N_10835,N_8439,N_8326);
or U10836 (N_10836,N_7431,N_7044);
nor U10837 (N_10837,N_8672,N_6181);
and U10838 (N_10838,N_8877,N_8710);
xor U10839 (N_10839,N_6697,N_6780);
or U10840 (N_10840,N_7818,N_8454);
nor U10841 (N_10841,N_6358,N_7054);
and U10842 (N_10842,N_7898,N_6619);
and U10843 (N_10843,N_6874,N_6875);
or U10844 (N_10844,N_8649,N_6854);
or U10845 (N_10845,N_6682,N_6916);
or U10846 (N_10846,N_6161,N_6660);
nor U10847 (N_10847,N_8720,N_7896);
nor U10848 (N_10848,N_8977,N_6189);
nor U10849 (N_10849,N_6447,N_8486);
nand U10850 (N_10850,N_8186,N_8277);
xor U10851 (N_10851,N_6772,N_8337);
nand U10852 (N_10852,N_6876,N_7576);
nor U10853 (N_10853,N_8764,N_7907);
nand U10854 (N_10854,N_7679,N_6071);
xnor U10855 (N_10855,N_6476,N_7528);
and U10856 (N_10856,N_6473,N_8978);
or U10857 (N_10857,N_7331,N_8042);
and U10858 (N_10858,N_6797,N_7408);
and U10859 (N_10859,N_8069,N_7806);
nand U10860 (N_10860,N_7723,N_8094);
and U10861 (N_10861,N_8279,N_6665);
and U10862 (N_10862,N_8461,N_8240);
nor U10863 (N_10863,N_6617,N_8481);
nand U10864 (N_10864,N_6329,N_7945);
nor U10865 (N_10865,N_8867,N_6829);
nand U10866 (N_10866,N_6575,N_8394);
nor U10867 (N_10867,N_7253,N_8489);
nand U10868 (N_10868,N_8903,N_7092);
and U10869 (N_10869,N_8420,N_6331);
xnor U10870 (N_10870,N_6093,N_8358);
nor U10871 (N_10871,N_6218,N_6661);
and U10872 (N_10872,N_7598,N_6208);
nand U10873 (N_10873,N_7440,N_7955);
nand U10874 (N_10874,N_8049,N_8326);
or U10875 (N_10875,N_8081,N_7695);
nor U10876 (N_10876,N_6009,N_8448);
or U10877 (N_10877,N_8723,N_6537);
xor U10878 (N_10878,N_7904,N_6707);
or U10879 (N_10879,N_7002,N_6644);
nand U10880 (N_10880,N_7783,N_6520);
or U10881 (N_10881,N_8435,N_6045);
xor U10882 (N_10882,N_8699,N_7189);
xnor U10883 (N_10883,N_7876,N_6367);
and U10884 (N_10884,N_6599,N_6746);
and U10885 (N_10885,N_8386,N_8637);
or U10886 (N_10886,N_7918,N_6742);
and U10887 (N_10887,N_6774,N_6822);
and U10888 (N_10888,N_8253,N_8897);
nor U10889 (N_10889,N_7651,N_7480);
and U10890 (N_10890,N_6380,N_6285);
or U10891 (N_10891,N_6196,N_7018);
xor U10892 (N_10892,N_8928,N_6772);
nand U10893 (N_10893,N_6797,N_6150);
and U10894 (N_10894,N_8792,N_6486);
and U10895 (N_10895,N_7811,N_7088);
nand U10896 (N_10896,N_6404,N_7757);
and U10897 (N_10897,N_8752,N_6271);
and U10898 (N_10898,N_7459,N_7359);
nor U10899 (N_10899,N_8899,N_8908);
xor U10900 (N_10900,N_6394,N_7497);
and U10901 (N_10901,N_7559,N_7175);
nand U10902 (N_10902,N_7986,N_6656);
nand U10903 (N_10903,N_8595,N_7261);
and U10904 (N_10904,N_6144,N_7710);
and U10905 (N_10905,N_6684,N_6440);
nand U10906 (N_10906,N_7201,N_8550);
or U10907 (N_10907,N_7373,N_6049);
nand U10908 (N_10908,N_8507,N_7101);
nor U10909 (N_10909,N_8340,N_6775);
and U10910 (N_10910,N_6348,N_8578);
or U10911 (N_10911,N_8755,N_6955);
or U10912 (N_10912,N_8657,N_8829);
nor U10913 (N_10913,N_8446,N_7647);
nand U10914 (N_10914,N_7224,N_7839);
or U10915 (N_10915,N_8848,N_6544);
or U10916 (N_10916,N_7835,N_8736);
and U10917 (N_10917,N_6650,N_6324);
or U10918 (N_10918,N_7085,N_7093);
and U10919 (N_10919,N_6519,N_6274);
and U10920 (N_10920,N_6498,N_7838);
or U10921 (N_10921,N_8894,N_8149);
nor U10922 (N_10922,N_7196,N_6521);
or U10923 (N_10923,N_6515,N_6168);
nand U10924 (N_10924,N_6067,N_8727);
and U10925 (N_10925,N_8923,N_6183);
nor U10926 (N_10926,N_8898,N_8209);
and U10927 (N_10927,N_8613,N_8178);
nor U10928 (N_10928,N_8657,N_8265);
or U10929 (N_10929,N_8386,N_8915);
or U10930 (N_10930,N_8439,N_6917);
or U10931 (N_10931,N_8499,N_8399);
nor U10932 (N_10932,N_6183,N_8539);
and U10933 (N_10933,N_6203,N_6252);
and U10934 (N_10934,N_6783,N_8195);
and U10935 (N_10935,N_7264,N_7212);
and U10936 (N_10936,N_8372,N_7989);
xnor U10937 (N_10937,N_8231,N_7793);
and U10938 (N_10938,N_7689,N_7160);
nand U10939 (N_10939,N_8856,N_7067);
nand U10940 (N_10940,N_6671,N_6150);
and U10941 (N_10941,N_7213,N_6420);
or U10942 (N_10942,N_6612,N_7281);
and U10943 (N_10943,N_7202,N_7368);
and U10944 (N_10944,N_7945,N_8798);
nand U10945 (N_10945,N_8325,N_6665);
nand U10946 (N_10946,N_6067,N_8726);
or U10947 (N_10947,N_8102,N_8080);
nand U10948 (N_10948,N_8345,N_7062);
nand U10949 (N_10949,N_7720,N_8948);
xnor U10950 (N_10950,N_6300,N_8672);
nor U10951 (N_10951,N_7671,N_7112);
xor U10952 (N_10952,N_7261,N_6193);
and U10953 (N_10953,N_8409,N_7692);
nor U10954 (N_10954,N_7535,N_8694);
nand U10955 (N_10955,N_7892,N_7491);
or U10956 (N_10956,N_8258,N_8924);
and U10957 (N_10957,N_8481,N_8786);
or U10958 (N_10958,N_8876,N_6388);
or U10959 (N_10959,N_7707,N_7817);
nand U10960 (N_10960,N_7794,N_8138);
xor U10961 (N_10961,N_6557,N_8311);
and U10962 (N_10962,N_6321,N_6093);
nor U10963 (N_10963,N_7749,N_6485);
nor U10964 (N_10964,N_8761,N_8475);
or U10965 (N_10965,N_7573,N_6691);
and U10966 (N_10966,N_8241,N_7634);
and U10967 (N_10967,N_7662,N_6361);
nor U10968 (N_10968,N_8060,N_6697);
nor U10969 (N_10969,N_8311,N_7124);
nor U10970 (N_10970,N_8138,N_7367);
nand U10971 (N_10971,N_8375,N_8591);
or U10972 (N_10972,N_7811,N_7232);
nand U10973 (N_10973,N_8038,N_7570);
and U10974 (N_10974,N_8498,N_8345);
and U10975 (N_10975,N_7775,N_6617);
xnor U10976 (N_10976,N_7977,N_8069);
and U10977 (N_10977,N_6391,N_7437);
or U10978 (N_10978,N_8169,N_8710);
nor U10979 (N_10979,N_8488,N_6842);
xnor U10980 (N_10980,N_8432,N_6225);
nand U10981 (N_10981,N_6144,N_8021);
and U10982 (N_10982,N_8073,N_8463);
or U10983 (N_10983,N_8170,N_7612);
nor U10984 (N_10984,N_7878,N_8338);
or U10985 (N_10985,N_7279,N_6828);
and U10986 (N_10986,N_8096,N_6038);
and U10987 (N_10987,N_8507,N_7196);
xnor U10988 (N_10988,N_7000,N_8733);
or U10989 (N_10989,N_6318,N_6692);
and U10990 (N_10990,N_7663,N_7205);
or U10991 (N_10991,N_8502,N_8672);
nand U10992 (N_10992,N_8490,N_6613);
nor U10993 (N_10993,N_7457,N_6827);
and U10994 (N_10994,N_8650,N_7382);
and U10995 (N_10995,N_6808,N_6829);
and U10996 (N_10996,N_7101,N_7645);
nand U10997 (N_10997,N_6226,N_8502);
and U10998 (N_10998,N_7548,N_6110);
nand U10999 (N_10999,N_7205,N_6299);
and U11000 (N_11000,N_8910,N_7816);
or U11001 (N_11001,N_8551,N_7086);
or U11002 (N_11002,N_8608,N_7803);
and U11003 (N_11003,N_6536,N_6211);
nand U11004 (N_11004,N_7928,N_7112);
and U11005 (N_11005,N_7400,N_8723);
nor U11006 (N_11006,N_8483,N_8803);
nand U11007 (N_11007,N_7178,N_6001);
or U11008 (N_11008,N_8336,N_8047);
and U11009 (N_11009,N_6229,N_7731);
nand U11010 (N_11010,N_8007,N_6362);
nand U11011 (N_11011,N_6090,N_8499);
nor U11012 (N_11012,N_6780,N_8800);
nand U11013 (N_11013,N_7028,N_6464);
or U11014 (N_11014,N_8969,N_8851);
xor U11015 (N_11015,N_7200,N_8510);
nor U11016 (N_11016,N_7146,N_6124);
or U11017 (N_11017,N_6127,N_6361);
or U11018 (N_11018,N_7416,N_7791);
nor U11019 (N_11019,N_7397,N_6800);
nand U11020 (N_11020,N_6607,N_8115);
nor U11021 (N_11021,N_8154,N_6112);
and U11022 (N_11022,N_6415,N_6577);
and U11023 (N_11023,N_8459,N_8705);
nor U11024 (N_11024,N_6249,N_7362);
or U11025 (N_11025,N_7821,N_8509);
or U11026 (N_11026,N_8849,N_6916);
or U11027 (N_11027,N_7710,N_7143);
and U11028 (N_11028,N_8926,N_6232);
or U11029 (N_11029,N_6801,N_8254);
nand U11030 (N_11030,N_7434,N_6629);
nor U11031 (N_11031,N_8692,N_7407);
or U11032 (N_11032,N_8874,N_7016);
nand U11033 (N_11033,N_8722,N_7101);
and U11034 (N_11034,N_8168,N_8297);
nor U11035 (N_11035,N_6415,N_6786);
xnor U11036 (N_11036,N_8237,N_8973);
nor U11037 (N_11037,N_8276,N_6569);
nor U11038 (N_11038,N_6551,N_8768);
and U11039 (N_11039,N_6804,N_8893);
or U11040 (N_11040,N_8672,N_6709);
nor U11041 (N_11041,N_8903,N_6354);
nand U11042 (N_11042,N_6031,N_6993);
nor U11043 (N_11043,N_8091,N_8114);
or U11044 (N_11044,N_8597,N_6827);
or U11045 (N_11045,N_7311,N_6593);
nor U11046 (N_11046,N_7740,N_6337);
xor U11047 (N_11047,N_7736,N_6560);
nand U11048 (N_11048,N_8439,N_8683);
nor U11049 (N_11049,N_7167,N_8364);
or U11050 (N_11050,N_8775,N_7503);
nand U11051 (N_11051,N_8742,N_7474);
nor U11052 (N_11052,N_6424,N_7614);
nor U11053 (N_11053,N_6955,N_7932);
nor U11054 (N_11054,N_7146,N_6780);
or U11055 (N_11055,N_7557,N_7754);
and U11056 (N_11056,N_7481,N_7685);
nand U11057 (N_11057,N_8973,N_6727);
nand U11058 (N_11058,N_6763,N_7480);
or U11059 (N_11059,N_8442,N_7234);
or U11060 (N_11060,N_7458,N_7104);
nand U11061 (N_11061,N_7054,N_8187);
nand U11062 (N_11062,N_7418,N_8842);
and U11063 (N_11063,N_7217,N_6678);
and U11064 (N_11064,N_7556,N_6571);
and U11065 (N_11065,N_8227,N_7722);
nor U11066 (N_11066,N_7343,N_7140);
and U11067 (N_11067,N_6234,N_7990);
nand U11068 (N_11068,N_6351,N_6834);
and U11069 (N_11069,N_7166,N_7190);
nand U11070 (N_11070,N_6179,N_7129);
or U11071 (N_11071,N_7463,N_7179);
nor U11072 (N_11072,N_8097,N_8553);
and U11073 (N_11073,N_8131,N_6581);
nand U11074 (N_11074,N_8566,N_7940);
nand U11075 (N_11075,N_6381,N_7787);
or U11076 (N_11076,N_7382,N_7075);
xnor U11077 (N_11077,N_7103,N_6744);
and U11078 (N_11078,N_8084,N_6265);
or U11079 (N_11079,N_6795,N_8927);
or U11080 (N_11080,N_7321,N_6206);
xor U11081 (N_11081,N_6177,N_7562);
and U11082 (N_11082,N_7318,N_8358);
nand U11083 (N_11083,N_8714,N_8630);
nor U11084 (N_11084,N_6348,N_8471);
nand U11085 (N_11085,N_8867,N_8852);
and U11086 (N_11086,N_7109,N_7083);
nor U11087 (N_11087,N_7613,N_7786);
nor U11088 (N_11088,N_7070,N_6757);
and U11089 (N_11089,N_7574,N_6960);
or U11090 (N_11090,N_6203,N_8849);
nand U11091 (N_11091,N_7267,N_6802);
nand U11092 (N_11092,N_6898,N_6546);
and U11093 (N_11093,N_6090,N_7275);
nor U11094 (N_11094,N_6005,N_6223);
nand U11095 (N_11095,N_7088,N_6684);
xnor U11096 (N_11096,N_8473,N_6864);
or U11097 (N_11097,N_7207,N_8207);
nand U11098 (N_11098,N_8104,N_8981);
and U11099 (N_11099,N_8741,N_6807);
or U11100 (N_11100,N_7667,N_6796);
nor U11101 (N_11101,N_6940,N_8749);
nor U11102 (N_11102,N_7324,N_8890);
nor U11103 (N_11103,N_6448,N_8696);
and U11104 (N_11104,N_8340,N_8412);
nor U11105 (N_11105,N_6294,N_6997);
or U11106 (N_11106,N_6713,N_6109);
nor U11107 (N_11107,N_8994,N_7050);
or U11108 (N_11108,N_6592,N_7350);
nand U11109 (N_11109,N_7704,N_7552);
nor U11110 (N_11110,N_8124,N_6819);
nor U11111 (N_11111,N_7640,N_6101);
or U11112 (N_11112,N_7088,N_8078);
nand U11113 (N_11113,N_6301,N_7847);
nor U11114 (N_11114,N_6565,N_7534);
and U11115 (N_11115,N_6469,N_8599);
or U11116 (N_11116,N_6951,N_6441);
nand U11117 (N_11117,N_8496,N_6923);
or U11118 (N_11118,N_6401,N_7859);
nor U11119 (N_11119,N_7217,N_8395);
nor U11120 (N_11120,N_7952,N_8139);
nor U11121 (N_11121,N_6724,N_7205);
or U11122 (N_11122,N_7167,N_7706);
or U11123 (N_11123,N_7043,N_7223);
nor U11124 (N_11124,N_8592,N_7445);
or U11125 (N_11125,N_6404,N_7569);
or U11126 (N_11126,N_7489,N_8288);
nor U11127 (N_11127,N_6868,N_6918);
nor U11128 (N_11128,N_8854,N_8842);
or U11129 (N_11129,N_8029,N_7871);
xnor U11130 (N_11130,N_8295,N_8486);
nor U11131 (N_11131,N_7068,N_6578);
nor U11132 (N_11132,N_7250,N_8128);
nand U11133 (N_11133,N_8399,N_7008);
or U11134 (N_11134,N_6810,N_8710);
or U11135 (N_11135,N_7082,N_6463);
xor U11136 (N_11136,N_8740,N_7914);
and U11137 (N_11137,N_8254,N_8755);
nand U11138 (N_11138,N_8058,N_8528);
xor U11139 (N_11139,N_7119,N_6087);
nand U11140 (N_11140,N_6966,N_6485);
nor U11141 (N_11141,N_7232,N_8090);
nor U11142 (N_11142,N_6939,N_6181);
xnor U11143 (N_11143,N_7675,N_6661);
or U11144 (N_11144,N_6901,N_7192);
nor U11145 (N_11145,N_7083,N_7003);
nand U11146 (N_11146,N_7774,N_6442);
and U11147 (N_11147,N_8371,N_7269);
and U11148 (N_11148,N_7472,N_7812);
nor U11149 (N_11149,N_6549,N_7283);
or U11150 (N_11150,N_6193,N_8927);
or U11151 (N_11151,N_8184,N_8362);
nor U11152 (N_11152,N_6827,N_7956);
nand U11153 (N_11153,N_6208,N_7543);
xor U11154 (N_11154,N_7666,N_8928);
and U11155 (N_11155,N_6098,N_8234);
xor U11156 (N_11156,N_6850,N_8344);
and U11157 (N_11157,N_7135,N_7297);
nand U11158 (N_11158,N_7121,N_6993);
nor U11159 (N_11159,N_7426,N_8872);
and U11160 (N_11160,N_7363,N_7056);
nand U11161 (N_11161,N_8385,N_8206);
nand U11162 (N_11162,N_6949,N_8753);
or U11163 (N_11163,N_6714,N_8052);
or U11164 (N_11164,N_7096,N_8136);
nand U11165 (N_11165,N_7340,N_7907);
nand U11166 (N_11166,N_7447,N_6797);
nand U11167 (N_11167,N_6531,N_7675);
or U11168 (N_11168,N_8548,N_7038);
nand U11169 (N_11169,N_8287,N_7963);
nor U11170 (N_11170,N_8614,N_8628);
and U11171 (N_11171,N_7353,N_8636);
nor U11172 (N_11172,N_8785,N_6906);
or U11173 (N_11173,N_6203,N_6516);
nor U11174 (N_11174,N_8369,N_7058);
and U11175 (N_11175,N_6251,N_6214);
nand U11176 (N_11176,N_6924,N_7906);
or U11177 (N_11177,N_6628,N_8551);
xnor U11178 (N_11178,N_8176,N_8423);
and U11179 (N_11179,N_6731,N_6387);
nand U11180 (N_11180,N_7408,N_7760);
and U11181 (N_11181,N_7564,N_7980);
and U11182 (N_11182,N_6107,N_6590);
nor U11183 (N_11183,N_8689,N_6692);
or U11184 (N_11184,N_7084,N_8023);
or U11185 (N_11185,N_8107,N_8174);
nand U11186 (N_11186,N_8701,N_7353);
or U11187 (N_11187,N_7629,N_6519);
nand U11188 (N_11188,N_6145,N_8045);
xor U11189 (N_11189,N_7780,N_6673);
or U11190 (N_11190,N_8780,N_8767);
nor U11191 (N_11191,N_6677,N_7549);
and U11192 (N_11192,N_6202,N_7870);
nor U11193 (N_11193,N_7164,N_6430);
nor U11194 (N_11194,N_6424,N_7173);
and U11195 (N_11195,N_7335,N_7187);
or U11196 (N_11196,N_6996,N_7876);
or U11197 (N_11197,N_6604,N_8045);
nor U11198 (N_11198,N_8594,N_8826);
nor U11199 (N_11199,N_7780,N_6639);
nor U11200 (N_11200,N_7286,N_6390);
and U11201 (N_11201,N_7631,N_6156);
nor U11202 (N_11202,N_8201,N_6232);
and U11203 (N_11203,N_7894,N_8144);
and U11204 (N_11204,N_7358,N_7383);
or U11205 (N_11205,N_7806,N_6851);
nor U11206 (N_11206,N_7800,N_8967);
nand U11207 (N_11207,N_7000,N_8477);
nand U11208 (N_11208,N_6999,N_6744);
nor U11209 (N_11209,N_6605,N_7118);
nor U11210 (N_11210,N_6726,N_8051);
nor U11211 (N_11211,N_6449,N_7938);
and U11212 (N_11212,N_6986,N_6831);
and U11213 (N_11213,N_8316,N_7710);
and U11214 (N_11214,N_6610,N_7370);
or U11215 (N_11215,N_8816,N_6362);
nor U11216 (N_11216,N_8850,N_6517);
and U11217 (N_11217,N_6395,N_6668);
or U11218 (N_11218,N_6430,N_8464);
or U11219 (N_11219,N_8665,N_6146);
or U11220 (N_11220,N_6826,N_8924);
or U11221 (N_11221,N_8052,N_8035);
nand U11222 (N_11222,N_8985,N_6933);
or U11223 (N_11223,N_8950,N_6516);
and U11224 (N_11224,N_8819,N_7450);
or U11225 (N_11225,N_7556,N_6413);
and U11226 (N_11226,N_8412,N_8021);
nor U11227 (N_11227,N_8239,N_8643);
or U11228 (N_11228,N_8458,N_7955);
nor U11229 (N_11229,N_7580,N_6886);
nand U11230 (N_11230,N_6226,N_6920);
and U11231 (N_11231,N_8019,N_7500);
nor U11232 (N_11232,N_7346,N_7363);
nand U11233 (N_11233,N_7158,N_7236);
nor U11234 (N_11234,N_6821,N_7438);
nand U11235 (N_11235,N_6023,N_6991);
nor U11236 (N_11236,N_8196,N_6142);
nand U11237 (N_11237,N_8828,N_6323);
nand U11238 (N_11238,N_7730,N_8300);
nand U11239 (N_11239,N_8847,N_7033);
nand U11240 (N_11240,N_8305,N_6896);
nand U11241 (N_11241,N_7276,N_7308);
nor U11242 (N_11242,N_8067,N_7115);
xnor U11243 (N_11243,N_6281,N_7485);
nand U11244 (N_11244,N_7184,N_7784);
or U11245 (N_11245,N_6337,N_7938);
xnor U11246 (N_11246,N_8649,N_6435);
or U11247 (N_11247,N_8975,N_8294);
nand U11248 (N_11248,N_6945,N_8090);
xor U11249 (N_11249,N_6853,N_8629);
and U11250 (N_11250,N_8639,N_7236);
and U11251 (N_11251,N_6759,N_7874);
nand U11252 (N_11252,N_8369,N_8620);
or U11253 (N_11253,N_8464,N_7991);
xnor U11254 (N_11254,N_7999,N_7096);
nand U11255 (N_11255,N_6291,N_6840);
nand U11256 (N_11256,N_6473,N_7231);
and U11257 (N_11257,N_7093,N_6124);
nand U11258 (N_11258,N_8126,N_7942);
and U11259 (N_11259,N_6277,N_8593);
xor U11260 (N_11260,N_7816,N_8102);
and U11261 (N_11261,N_8207,N_6350);
and U11262 (N_11262,N_8789,N_7904);
nor U11263 (N_11263,N_7747,N_6987);
and U11264 (N_11264,N_8415,N_7435);
and U11265 (N_11265,N_8782,N_7220);
nand U11266 (N_11266,N_7655,N_7511);
nor U11267 (N_11267,N_6257,N_8397);
nor U11268 (N_11268,N_8092,N_8957);
xor U11269 (N_11269,N_6778,N_8460);
or U11270 (N_11270,N_6284,N_7984);
or U11271 (N_11271,N_8955,N_6839);
nand U11272 (N_11272,N_7840,N_8634);
or U11273 (N_11273,N_8204,N_7760);
and U11274 (N_11274,N_7607,N_8565);
or U11275 (N_11275,N_8035,N_8723);
and U11276 (N_11276,N_8504,N_8047);
nor U11277 (N_11277,N_8523,N_8459);
and U11278 (N_11278,N_8855,N_6811);
xnor U11279 (N_11279,N_8092,N_8527);
nand U11280 (N_11280,N_7754,N_7663);
and U11281 (N_11281,N_7551,N_6206);
or U11282 (N_11282,N_8094,N_8886);
nor U11283 (N_11283,N_8961,N_7341);
or U11284 (N_11284,N_6486,N_8684);
nor U11285 (N_11285,N_7214,N_6025);
or U11286 (N_11286,N_8902,N_6544);
nor U11287 (N_11287,N_7290,N_8590);
or U11288 (N_11288,N_6128,N_7818);
nor U11289 (N_11289,N_7313,N_8630);
nand U11290 (N_11290,N_8653,N_7534);
and U11291 (N_11291,N_8679,N_7252);
nand U11292 (N_11292,N_7106,N_8712);
nand U11293 (N_11293,N_8887,N_8231);
xnor U11294 (N_11294,N_8941,N_6526);
and U11295 (N_11295,N_6696,N_8830);
and U11296 (N_11296,N_7151,N_8318);
xnor U11297 (N_11297,N_8278,N_6178);
nor U11298 (N_11298,N_6054,N_6225);
or U11299 (N_11299,N_6588,N_6087);
or U11300 (N_11300,N_7244,N_7921);
or U11301 (N_11301,N_7687,N_7393);
nand U11302 (N_11302,N_6131,N_6221);
nand U11303 (N_11303,N_6514,N_6879);
and U11304 (N_11304,N_8877,N_6142);
and U11305 (N_11305,N_7775,N_7027);
nor U11306 (N_11306,N_6227,N_8882);
nor U11307 (N_11307,N_6090,N_6503);
and U11308 (N_11308,N_8661,N_8501);
nor U11309 (N_11309,N_6577,N_8374);
nand U11310 (N_11310,N_8630,N_6593);
nand U11311 (N_11311,N_7700,N_7092);
and U11312 (N_11312,N_8282,N_8749);
nor U11313 (N_11313,N_8806,N_6256);
nand U11314 (N_11314,N_6508,N_7466);
nor U11315 (N_11315,N_6253,N_8778);
and U11316 (N_11316,N_6098,N_8311);
nand U11317 (N_11317,N_8165,N_7615);
nor U11318 (N_11318,N_8170,N_6146);
nor U11319 (N_11319,N_6449,N_8450);
nor U11320 (N_11320,N_7619,N_8696);
nor U11321 (N_11321,N_6798,N_8639);
and U11322 (N_11322,N_7518,N_7998);
xor U11323 (N_11323,N_7518,N_8287);
xor U11324 (N_11324,N_7914,N_7999);
nand U11325 (N_11325,N_7245,N_8687);
nand U11326 (N_11326,N_8376,N_8960);
nor U11327 (N_11327,N_7939,N_7318);
nor U11328 (N_11328,N_6087,N_6144);
and U11329 (N_11329,N_8986,N_7604);
and U11330 (N_11330,N_8187,N_6186);
or U11331 (N_11331,N_7668,N_6458);
nand U11332 (N_11332,N_7833,N_6742);
nor U11333 (N_11333,N_7834,N_8481);
nand U11334 (N_11334,N_8562,N_7204);
or U11335 (N_11335,N_7537,N_8235);
or U11336 (N_11336,N_6930,N_8841);
nor U11337 (N_11337,N_8953,N_7164);
nor U11338 (N_11338,N_8214,N_6483);
or U11339 (N_11339,N_6923,N_8708);
xnor U11340 (N_11340,N_7648,N_8793);
xor U11341 (N_11341,N_8775,N_8935);
and U11342 (N_11342,N_6850,N_8380);
and U11343 (N_11343,N_7203,N_6899);
and U11344 (N_11344,N_6963,N_6823);
xnor U11345 (N_11345,N_7480,N_8252);
or U11346 (N_11346,N_7968,N_6757);
or U11347 (N_11347,N_7149,N_7546);
or U11348 (N_11348,N_6329,N_6432);
and U11349 (N_11349,N_6000,N_8331);
and U11350 (N_11350,N_8357,N_7381);
and U11351 (N_11351,N_7930,N_7347);
xor U11352 (N_11352,N_7606,N_7425);
and U11353 (N_11353,N_8683,N_6414);
and U11354 (N_11354,N_6939,N_7144);
or U11355 (N_11355,N_8263,N_6009);
xor U11356 (N_11356,N_8864,N_8609);
and U11357 (N_11357,N_8778,N_6977);
nor U11358 (N_11358,N_6959,N_7610);
or U11359 (N_11359,N_8148,N_6459);
nor U11360 (N_11360,N_8042,N_8404);
and U11361 (N_11361,N_7063,N_8476);
or U11362 (N_11362,N_8194,N_8189);
xor U11363 (N_11363,N_8875,N_7681);
nor U11364 (N_11364,N_6797,N_7265);
xor U11365 (N_11365,N_7920,N_7072);
nand U11366 (N_11366,N_7668,N_8557);
nor U11367 (N_11367,N_6138,N_6353);
nand U11368 (N_11368,N_6484,N_8137);
or U11369 (N_11369,N_7095,N_6197);
or U11370 (N_11370,N_6643,N_6195);
or U11371 (N_11371,N_8304,N_6663);
or U11372 (N_11372,N_7421,N_8835);
and U11373 (N_11373,N_6019,N_7841);
nand U11374 (N_11374,N_7766,N_7795);
or U11375 (N_11375,N_8401,N_8154);
and U11376 (N_11376,N_8787,N_7225);
nand U11377 (N_11377,N_7444,N_7547);
nand U11378 (N_11378,N_7513,N_6689);
nor U11379 (N_11379,N_6816,N_8773);
nand U11380 (N_11380,N_8485,N_6663);
and U11381 (N_11381,N_7703,N_7875);
xnor U11382 (N_11382,N_6983,N_8174);
and U11383 (N_11383,N_8391,N_7830);
nand U11384 (N_11384,N_8989,N_7564);
or U11385 (N_11385,N_6927,N_6716);
nand U11386 (N_11386,N_7727,N_7157);
nand U11387 (N_11387,N_6789,N_8585);
xor U11388 (N_11388,N_6006,N_8691);
and U11389 (N_11389,N_7033,N_6055);
and U11390 (N_11390,N_7115,N_8788);
or U11391 (N_11391,N_8653,N_6560);
or U11392 (N_11392,N_6835,N_8067);
nor U11393 (N_11393,N_6306,N_7943);
xnor U11394 (N_11394,N_7758,N_7270);
nand U11395 (N_11395,N_8109,N_8839);
or U11396 (N_11396,N_7822,N_8952);
or U11397 (N_11397,N_7432,N_8489);
nand U11398 (N_11398,N_6185,N_7407);
and U11399 (N_11399,N_6669,N_7525);
xor U11400 (N_11400,N_7784,N_6251);
nor U11401 (N_11401,N_6821,N_7350);
nand U11402 (N_11402,N_6433,N_8369);
and U11403 (N_11403,N_8752,N_7619);
nor U11404 (N_11404,N_7599,N_6209);
and U11405 (N_11405,N_6325,N_6764);
nand U11406 (N_11406,N_8162,N_8871);
and U11407 (N_11407,N_6655,N_6400);
or U11408 (N_11408,N_8063,N_6911);
nand U11409 (N_11409,N_7512,N_8360);
nand U11410 (N_11410,N_7330,N_6129);
nor U11411 (N_11411,N_8894,N_6653);
or U11412 (N_11412,N_8633,N_7735);
nand U11413 (N_11413,N_8801,N_8566);
nand U11414 (N_11414,N_8735,N_8691);
xnor U11415 (N_11415,N_7151,N_6250);
nand U11416 (N_11416,N_8282,N_7322);
and U11417 (N_11417,N_6880,N_6896);
nor U11418 (N_11418,N_7308,N_7361);
and U11419 (N_11419,N_7265,N_8745);
nand U11420 (N_11420,N_8702,N_8367);
nand U11421 (N_11421,N_6711,N_7319);
nand U11422 (N_11422,N_6777,N_8044);
xnor U11423 (N_11423,N_8114,N_7172);
nor U11424 (N_11424,N_8975,N_8285);
nor U11425 (N_11425,N_8672,N_7262);
xor U11426 (N_11426,N_7363,N_6114);
and U11427 (N_11427,N_6806,N_8063);
and U11428 (N_11428,N_8764,N_7759);
and U11429 (N_11429,N_6640,N_6361);
nor U11430 (N_11430,N_8390,N_6683);
and U11431 (N_11431,N_8542,N_6969);
and U11432 (N_11432,N_6440,N_8344);
nor U11433 (N_11433,N_8064,N_7630);
xor U11434 (N_11434,N_6655,N_7152);
nor U11435 (N_11435,N_8203,N_6709);
nor U11436 (N_11436,N_8943,N_7279);
and U11437 (N_11437,N_6576,N_6193);
xnor U11438 (N_11438,N_7682,N_6619);
nor U11439 (N_11439,N_6136,N_8575);
and U11440 (N_11440,N_8295,N_8438);
nand U11441 (N_11441,N_6927,N_7627);
nor U11442 (N_11442,N_6002,N_7187);
nor U11443 (N_11443,N_7292,N_7209);
and U11444 (N_11444,N_8008,N_6318);
nand U11445 (N_11445,N_7752,N_8123);
and U11446 (N_11446,N_7136,N_8272);
xor U11447 (N_11447,N_8231,N_7731);
and U11448 (N_11448,N_8330,N_8852);
nor U11449 (N_11449,N_6290,N_7740);
nor U11450 (N_11450,N_7895,N_8953);
and U11451 (N_11451,N_6394,N_8573);
or U11452 (N_11452,N_6500,N_6035);
or U11453 (N_11453,N_7500,N_7181);
nand U11454 (N_11454,N_8459,N_6086);
or U11455 (N_11455,N_6903,N_6789);
nand U11456 (N_11456,N_8786,N_8943);
and U11457 (N_11457,N_7351,N_8929);
nand U11458 (N_11458,N_6008,N_6937);
and U11459 (N_11459,N_7136,N_7300);
and U11460 (N_11460,N_8221,N_7258);
nand U11461 (N_11461,N_7220,N_6097);
nand U11462 (N_11462,N_6865,N_6867);
nand U11463 (N_11463,N_7060,N_6748);
or U11464 (N_11464,N_7607,N_7255);
nand U11465 (N_11465,N_6700,N_8795);
xnor U11466 (N_11466,N_8556,N_8099);
nor U11467 (N_11467,N_6349,N_8273);
or U11468 (N_11468,N_7117,N_8572);
or U11469 (N_11469,N_7825,N_6133);
or U11470 (N_11470,N_6038,N_8754);
nor U11471 (N_11471,N_7969,N_6562);
nand U11472 (N_11472,N_7993,N_6798);
or U11473 (N_11473,N_8774,N_7693);
and U11474 (N_11474,N_8531,N_7297);
nor U11475 (N_11475,N_7832,N_6527);
and U11476 (N_11476,N_6619,N_8874);
or U11477 (N_11477,N_7938,N_7350);
nand U11478 (N_11478,N_7332,N_7679);
nand U11479 (N_11479,N_6862,N_6448);
nand U11480 (N_11480,N_8012,N_6998);
nor U11481 (N_11481,N_6898,N_8836);
nand U11482 (N_11482,N_8061,N_6018);
and U11483 (N_11483,N_6921,N_8779);
nand U11484 (N_11484,N_8862,N_6512);
nor U11485 (N_11485,N_7944,N_8147);
and U11486 (N_11486,N_8101,N_6122);
and U11487 (N_11487,N_8262,N_8817);
and U11488 (N_11488,N_6242,N_6465);
nor U11489 (N_11489,N_6383,N_6174);
nand U11490 (N_11490,N_6658,N_7044);
nand U11491 (N_11491,N_8794,N_6619);
nand U11492 (N_11492,N_8772,N_6813);
xor U11493 (N_11493,N_7372,N_8315);
and U11494 (N_11494,N_7063,N_8137);
and U11495 (N_11495,N_6646,N_8648);
and U11496 (N_11496,N_7603,N_8297);
nand U11497 (N_11497,N_7233,N_8546);
nand U11498 (N_11498,N_7576,N_7273);
and U11499 (N_11499,N_6224,N_8147);
xor U11500 (N_11500,N_6357,N_7901);
and U11501 (N_11501,N_8733,N_7332);
nor U11502 (N_11502,N_7901,N_6037);
or U11503 (N_11503,N_7452,N_8591);
nand U11504 (N_11504,N_6413,N_7474);
nand U11505 (N_11505,N_7071,N_8108);
and U11506 (N_11506,N_8961,N_7954);
or U11507 (N_11507,N_8381,N_8737);
and U11508 (N_11508,N_6903,N_8374);
nand U11509 (N_11509,N_7600,N_8897);
nand U11510 (N_11510,N_8288,N_7961);
nor U11511 (N_11511,N_8435,N_8347);
nor U11512 (N_11512,N_8431,N_6856);
or U11513 (N_11513,N_6214,N_6558);
or U11514 (N_11514,N_7587,N_6025);
nor U11515 (N_11515,N_7693,N_8008);
or U11516 (N_11516,N_8399,N_7937);
nand U11517 (N_11517,N_7913,N_8557);
or U11518 (N_11518,N_6390,N_7793);
nand U11519 (N_11519,N_7287,N_6119);
or U11520 (N_11520,N_6428,N_8772);
or U11521 (N_11521,N_6487,N_6463);
xnor U11522 (N_11522,N_7512,N_6069);
xor U11523 (N_11523,N_6625,N_6743);
and U11524 (N_11524,N_8206,N_6643);
and U11525 (N_11525,N_8692,N_6767);
and U11526 (N_11526,N_7937,N_7325);
xor U11527 (N_11527,N_6710,N_8983);
xor U11528 (N_11528,N_8895,N_7530);
and U11529 (N_11529,N_8786,N_8677);
nand U11530 (N_11530,N_8868,N_8517);
or U11531 (N_11531,N_8935,N_6803);
nor U11532 (N_11532,N_7462,N_8173);
nor U11533 (N_11533,N_8086,N_8286);
and U11534 (N_11534,N_7253,N_6203);
nor U11535 (N_11535,N_7576,N_6515);
nand U11536 (N_11536,N_7901,N_7465);
nand U11537 (N_11537,N_7507,N_8343);
or U11538 (N_11538,N_8983,N_6239);
or U11539 (N_11539,N_7905,N_6754);
xnor U11540 (N_11540,N_8785,N_7383);
and U11541 (N_11541,N_7561,N_8466);
nand U11542 (N_11542,N_7164,N_8318);
or U11543 (N_11543,N_7633,N_7775);
or U11544 (N_11544,N_7769,N_8097);
nor U11545 (N_11545,N_6900,N_6276);
nor U11546 (N_11546,N_6493,N_7171);
and U11547 (N_11547,N_6514,N_6281);
nor U11548 (N_11548,N_6620,N_6748);
nor U11549 (N_11549,N_7998,N_8160);
and U11550 (N_11550,N_7855,N_8162);
nor U11551 (N_11551,N_6752,N_8149);
and U11552 (N_11552,N_7906,N_6546);
or U11553 (N_11553,N_7234,N_7264);
or U11554 (N_11554,N_8692,N_7694);
and U11555 (N_11555,N_6901,N_8008);
nor U11556 (N_11556,N_7909,N_8199);
or U11557 (N_11557,N_6245,N_8300);
and U11558 (N_11558,N_6443,N_8067);
nor U11559 (N_11559,N_6599,N_8880);
or U11560 (N_11560,N_6639,N_6582);
nand U11561 (N_11561,N_6937,N_8425);
and U11562 (N_11562,N_8495,N_6336);
and U11563 (N_11563,N_6415,N_8510);
nand U11564 (N_11564,N_8642,N_8646);
nand U11565 (N_11565,N_7515,N_8119);
nor U11566 (N_11566,N_7198,N_8939);
and U11567 (N_11567,N_8607,N_8180);
nand U11568 (N_11568,N_6345,N_6237);
nand U11569 (N_11569,N_6929,N_8295);
or U11570 (N_11570,N_8564,N_8825);
xnor U11571 (N_11571,N_7384,N_8557);
nand U11572 (N_11572,N_7187,N_8363);
nand U11573 (N_11573,N_7693,N_8594);
and U11574 (N_11574,N_8279,N_6161);
or U11575 (N_11575,N_6200,N_7999);
or U11576 (N_11576,N_6987,N_6230);
nand U11577 (N_11577,N_8047,N_7699);
or U11578 (N_11578,N_6709,N_6553);
nand U11579 (N_11579,N_6889,N_8310);
nor U11580 (N_11580,N_7524,N_7722);
nand U11581 (N_11581,N_7939,N_8898);
xor U11582 (N_11582,N_8677,N_8391);
and U11583 (N_11583,N_8047,N_6249);
nand U11584 (N_11584,N_8198,N_8875);
or U11585 (N_11585,N_8739,N_7951);
nand U11586 (N_11586,N_6000,N_8553);
nand U11587 (N_11587,N_8916,N_6343);
and U11588 (N_11588,N_8904,N_6290);
or U11589 (N_11589,N_7765,N_8118);
and U11590 (N_11590,N_7641,N_7376);
or U11591 (N_11591,N_8317,N_8321);
and U11592 (N_11592,N_7983,N_8562);
nor U11593 (N_11593,N_8381,N_6991);
and U11594 (N_11594,N_6700,N_7767);
xnor U11595 (N_11595,N_7573,N_7719);
nor U11596 (N_11596,N_8950,N_7297);
and U11597 (N_11597,N_7878,N_6385);
or U11598 (N_11598,N_8792,N_8180);
nand U11599 (N_11599,N_7482,N_6364);
or U11600 (N_11600,N_8769,N_8458);
nand U11601 (N_11601,N_7196,N_8161);
or U11602 (N_11602,N_8679,N_7521);
or U11603 (N_11603,N_6160,N_8094);
nor U11604 (N_11604,N_6511,N_6725);
nand U11605 (N_11605,N_8530,N_7976);
or U11606 (N_11606,N_6704,N_7293);
xnor U11607 (N_11607,N_7694,N_8332);
nor U11608 (N_11608,N_8347,N_8419);
xor U11609 (N_11609,N_7452,N_8479);
and U11610 (N_11610,N_8183,N_6200);
nor U11611 (N_11611,N_6036,N_8109);
xnor U11612 (N_11612,N_6334,N_8803);
and U11613 (N_11613,N_8413,N_8957);
nor U11614 (N_11614,N_6486,N_8398);
and U11615 (N_11615,N_6990,N_7208);
nor U11616 (N_11616,N_7481,N_8155);
or U11617 (N_11617,N_8558,N_7876);
or U11618 (N_11618,N_7501,N_6542);
nor U11619 (N_11619,N_7451,N_8418);
xor U11620 (N_11620,N_8735,N_6891);
nor U11621 (N_11621,N_6407,N_7411);
nand U11622 (N_11622,N_6167,N_6749);
or U11623 (N_11623,N_6036,N_6709);
and U11624 (N_11624,N_8611,N_7157);
xor U11625 (N_11625,N_8981,N_6385);
and U11626 (N_11626,N_6639,N_7006);
nor U11627 (N_11627,N_6109,N_8031);
nor U11628 (N_11628,N_6864,N_8562);
xor U11629 (N_11629,N_7623,N_8223);
and U11630 (N_11630,N_6029,N_8826);
or U11631 (N_11631,N_7102,N_7226);
nand U11632 (N_11632,N_7303,N_7873);
nor U11633 (N_11633,N_8963,N_8055);
and U11634 (N_11634,N_7461,N_8168);
xor U11635 (N_11635,N_6271,N_6218);
nand U11636 (N_11636,N_7495,N_8015);
and U11637 (N_11637,N_6020,N_8171);
nand U11638 (N_11638,N_7590,N_7510);
nand U11639 (N_11639,N_7500,N_8621);
xnor U11640 (N_11640,N_8857,N_7472);
or U11641 (N_11641,N_7630,N_7413);
or U11642 (N_11642,N_7074,N_8202);
or U11643 (N_11643,N_6582,N_6166);
nor U11644 (N_11644,N_7213,N_7131);
or U11645 (N_11645,N_8779,N_8296);
and U11646 (N_11646,N_7710,N_7777);
nor U11647 (N_11647,N_7692,N_7446);
nor U11648 (N_11648,N_8416,N_7664);
and U11649 (N_11649,N_6148,N_6456);
and U11650 (N_11650,N_8958,N_6528);
nand U11651 (N_11651,N_6652,N_8208);
nor U11652 (N_11652,N_7624,N_8019);
nand U11653 (N_11653,N_6204,N_8206);
xnor U11654 (N_11654,N_6533,N_7282);
and U11655 (N_11655,N_7451,N_8722);
and U11656 (N_11656,N_6885,N_7373);
or U11657 (N_11657,N_6631,N_7918);
nand U11658 (N_11658,N_7183,N_7901);
or U11659 (N_11659,N_8402,N_8364);
nand U11660 (N_11660,N_6954,N_7107);
or U11661 (N_11661,N_7414,N_6578);
nor U11662 (N_11662,N_7239,N_7248);
nand U11663 (N_11663,N_7330,N_8506);
nand U11664 (N_11664,N_7969,N_6251);
nor U11665 (N_11665,N_6183,N_8246);
nor U11666 (N_11666,N_7368,N_6091);
xnor U11667 (N_11667,N_8859,N_7464);
or U11668 (N_11668,N_8463,N_7709);
nand U11669 (N_11669,N_7172,N_7889);
or U11670 (N_11670,N_7225,N_7499);
nor U11671 (N_11671,N_8391,N_6686);
nor U11672 (N_11672,N_8636,N_7000);
nand U11673 (N_11673,N_6769,N_6096);
or U11674 (N_11674,N_7602,N_8212);
and U11675 (N_11675,N_7201,N_6179);
xor U11676 (N_11676,N_7642,N_7026);
and U11677 (N_11677,N_6783,N_8788);
nand U11678 (N_11678,N_7373,N_6340);
or U11679 (N_11679,N_6073,N_6814);
nand U11680 (N_11680,N_8716,N_7078);
xnor U11681 (N_11681,N_6163,N_7609);
or U11682 (N_11682,N_7125,N_6848);
or U11683 (N_11683,N_8332,N_7524);
and U11684 (N_11684,N_7776,N_7765);
nand U11685 (N_11685,N_6725,N_6153);
and U11686 (N_11686,N_8725,N_7644);
or U11687 (N_11687,N_6535,N_6728);
and U11688 (N_11688,N_6074,N_6965);
nor U11689 (N_11689,N_7186,N_6136);
nand U11690 (N_11690,N_8608,N_8770);
xor U11691 (N_11691,N_7696,N_6734);
and U11692 (N_11692,N_7023,N_7773);
nand U11693 (N_11693,N_7625,N_7091);
nand U11694 (N_11694,N_7783,N_6595);
or U11695 (N_11695,N_8407,N_6136);
xor U11696 (N_11696,N_6420,N_7194);
or U11697 (N_11697,N_6609,N_7637);
nand U11698 (N_11698,N_7603,N_6471);
and U11699 (N_11699,N_8173,N_6156);
or U11700 (N_11700,N_6506,N_7972);
or U11701 (N_11701,N_6208,N_7612);
nor U11702 (N_11702,N_6696,N_8555);
xnor U11703 (N_11703,N_6489,N_6809);
and U11704 (N_11704,N_6986,N_8701);
or U11705 (N_11705,N_6354,N_8819);
and U11706 (N_11706,N_8884,N_6871);
and U11707 (N_11707,N_8018,N_7632);
nor U11708 (N_11708,N_7215,N_6355);
or U11709 (N_11709,N_6329,N_6682);
nand U11710 (N_11710,N_6379,N_6972);
nand U11711 (N_11711,N_7715,N_7595);
nor U11712 (N_11712,N_6368,N_6936);
nor U11713 (N_11713,N_6137,N_8994);
or U11714 (N_11714,N_7737,N_6775);
and U11715 (N_11715,N_7186,N_8299);
or U11716 (N_11716,N_7988,N_6240);
nand U11717 (N_11717,N_7367,N_8811);
nand U11718 (N_11718,N_6230,N_7811);
nand U11719 (N_11719,N_6984,N_8790);
xor U11720 (N_11720,N_6135,N_6986);
nor U11721 (N_11721,N_6860,N_6605);
nor U11722 (N_11722,N_7761,N_8673);
or U11723 (N_11723,N_7200,N_6727);
and U11724 (N_11724,N_6078,N_6707);
nand U11725 (N_11725,N_7745,N_7060);
and U11726 (N_11726,N_6220,N_6335);
nor U11727 (N_11727,N_8209,N_6267);
nor U11728 (N_11728,N_8662,N_8034);
nand U11729 (N_11729,N_7108,N_8837);
nand U11730 (N_11730,N_8087,N_8582);
nand U11731 (N_11731,N_7428,N_7584);
nor U11732 (N_11732,N_7160,N_6004);
or U11733 (N_11733,N_8634,N_7053);
or U11734 (N_11734,N_6886,N_6303);
or U11735 (N_11735,N_6768,N_6032);
xnor U11736 (N_11736,N_8517,N_8913);
nand U11737 (N_11737,N_7296,N_6618);
and U11738 (N_11738,N_6863,N_7831);
or U11739 (N_11739,N_8061,N_7913);
nor U11740 (N_11740,N_6164,N_7926);
nor U11741 (N_11741,N_7908,N_6765);
nor U11742 (N_11742,N_6923,N_8446);
or U11743 (N_11743,N_7437,N_8168);
nor U11744 (N_11744,N_8373,N_7930);
nor U11745 (N_11745,N_8295,N_8355);
or U11746 (N_11746,N_7495,N_6716);
xnor U11747 (N_11747,N_8821,N_6783);
nor U11748 (N_11748,N_8741,N_6513);
and U11749 (N_11749,N_6403,N_7927);
nand U11750 (N_11750,N_7597,N_7350);
nor U11751 (N_11751,N_7939,N_6238);
nand U11752 (N_11752,N_7706,N_7303);
or U11753 (N_11753,N_7196,N_6613);
and U11754 (N_11754,N_6288,N_7576);
nand U11755 (N_11755,N_7787,N_8759);
nor U11756 (N_11756,N_8318,N_6823);
and U11757 (N_11757,N_8952,N_8332);
and U11758 (N_11758,N_8029,N_8768);
or U11759 (N_11759,N_6251,N_6817);
nor U11760 (N_11760,N_6754,N_8355);
nor U11761 (N_11761,N_8009,N_8983);
nor U11762 (N_11762,N_8423,N_8629);
or U11763 (N_11763,N_6214,N_8532);
nor U11764 (N_11764,N_6448,N_6698);
and U11765 (N_11765,N_7041,N_8415);
and U11766 (N_11766,N_8630,N_8553);
and U11767 (N_11767,N_6394,N_7078);
nor U11768 (N_11768,N_8530,N_8353);
and U11769 (N_11769,N_8292,N_6505);
or U11770 (N_11770,N_6245,N_8724);
nand U11771 (N_11771,N_8047,N_8404);
nand U11772 (N_11772,N_6227,N_8457);
nand U11773 (N_11773,N_6237,N_7108);
and U11774 (N_11774,N_8331,N_8324);
or U11775 (N_11775,N_6935,N_7740);
nand U11776 (N_11776,N_6919,N_8545);
nor U11777 (N_11777,N_7140,N_6902);
nand U11778 (N_11778,N_8112,N_6635);
or U11779 (N_11779,N_6590,N_8602);
or U11780 (N_11780,N_7362,N_7719);
and U11781 (N_11781,N_7664,N_6294);
and U11782 (N_11782,N_6578,N_6084);
nor U11783 (N_11783,N_7840,N_8213);
nor U11784 (N_11784,N_6592,N_7826);
nand U11785 (N_11785,N_8268,N_6225);
or U11786 (N_11786,N_7701,N_8034);
nor U11787 (N_11787,N_7945,N_7926);
and U11788 (N_11788,N_6545,N_6127);
and U11789 (N_11789,N_8241,N_8063);
and U11790 (N_11790,N_7376,N_6969);
nand U11791 (N_11791,N_8117,N_6359);
or U11792 (N_11792,N_8580,N_7704);
xnor U11793 (N_11793,N_7825,N_6177);
or U11794 (N_11794,N_6473,N_7060);
or U11795 (N_11795,N_8440,N_8527);
nor U11796 (N_11796,N_6651,N_7232);
nor U11797 (N_11797,N_8516,N_8897);
and U11798 (N_11798,N_7290,N_7149);
xnor U11799 (N_11799,N_6077,N_8861);
or U11800 (N_11800,N_7698,N_6141);
xnor U11801 (N_11801,N_7072,N_7656);
nor U11802 (N_11802,N_6616,N_8022);
nor U11803 (N_11803,N_8490,N_8444);
or U11804 (N_11804,N_8234,N_6861);
nor U11805 (N_11805,N_8340,N_7293);
and U11806 (N_11806,N_6320,N_6991);
nand U11807 (N_11807,N_6237,N_7850);
nor U11808 (N_11808,N_8364,N_7365);
and U11809 (N_11809,N_7981,N_7425);
or U11810 (N_11810,N_8497,N_7551);
nand U11811 (N_11811,N_6973,N_6448);
and U11812 (N_11812,N_6169,N_8309);
nor U11813 (N_11813,N_8626,N_8644);
and U11814 (N_11814,N_7554,N_8025);
nand U11815 (N_11815,N_6549,N_8757);
nand U11816 (N_11816,N_8035,N_8649);
and U11817 (N_11817,N_6444,N_6547);
nand U11818 (N_11818,N_6306,N_6602);
or U11819 (N_11819,N_6456,N_7256);
nor U11820 (N_11820,N_6060,N_6862);
nor U11821 (N_11821,N_8129,N_7254);
or U11822 (N_11822,N_6738,N_8345);
nand U11823 (N_11823,N_6812,N_8172);
nand U11824 (N_11824,N_6582,N_7802);
nor U11825 (N_11825,N_6040,N_7410);
and U11826 (N_11826,N_6647,N_7557);
nand U11827 (N_11827,N_6603,N_8066);
or U11828 (N_11828,N_7546,N_7272);
nor U11829 (N_11829,N_6881,N_8088);
or U11830 (N_11830,N_6605,N_7646);
nor U11831 (N_11831,N_7590,N_6135);
nor U11832 (N_11832,N_7865,N_6338);
xnor U11833 (N_11833,N_8314,N_7509);
nor U11834 (N_11834,N_6829,N_7604);
or U11835 (N_11835,N_7023,N_6710);
or U11836 (N_11836,N_8908,N_7262);
nor U11837 (N_11837,N_6359,N_7525);
nor U11838 (N_11838,N_7353,N_7971);
and U11839 (N_11839,N_8764,N_8298);
or U11840 (N_11840,N_6422,N_7369);
nor U11841 (N_11841,N_6693,N_8344);
or U11842 (N_11842,N_6426,N_6923);
xor U11843 (N_11843,N_8070,N_7480);
nor U11844 (N_11844,N_6440,N_8724);
xor U11845 (N_11845,N_6147,N_8766);
nand U11846 (N_11846,N_8239,N_6289);
or U11847 (N_11847,N_7079,N_6745);
nand U11848 (N_11848,N_7499,N_7751);
or U11849 (N_11849,N_8306,N_7672);
nand U11850 (N_11850,N_8461,N_6846);
and U11851 (N_11851,N_6646,N_7174);
or U11852 (N_11852,N_8619,N_7939);
or U11853 (N_11853,N_8148,N_8725);
nand U11854 (N_11854,N_8276,N_6670);
and U11855 (N_11855,N_8837,N_6653);
and U11856 (N_11856,N_6287,N_7241);
nand U11857 (N_11857,N_6342,N_6096);
nand U11858 (N_11858,N_6899,N_8432);
nand U11859 (N_11859,N_6260,N_6254);
nor U11860 (N_11860,N_6045,N_6136);
nor U11861 (N_11861,N_7851,N_8267);
and U11862 (N_11862,N_6777,N_8331);
nand U11863 (N_11863,N_8024,N_8705);
nor U11864 (N_11864,N_8193,N_7961);
nor U11865 (N_11865,N_8677,N_8945);
xnor U11866 (N_11866,N_7435,N_6126);
nor U11867 (N_11867,N_6290,N_6207);
nor U11868 (N_11868,N_6063,N_6460);
nor U11869 (N_11869,N_6107,N_8222);
or U11870 (N_11870,N_6134,N_6375);
nor U11871 (N_11871,N_7440,N_8781);
nor U11872 (N_11872,N_8846,N_7933);
nor U11873 (N_11873,N_8678,N_7533);
nor U11874 (N_11874,N_6910,N_7632);
and U11875 (N_11875,N_7855,N_7368);
or U11876 (N_11876,N_7034,N_7381);
nor U11877 (N_11877,N_6295,N_6678);
nor U11878 (N_11878,N_8918,N_6181);
or U11879 (N_11879,N_7368,N_6443);
nand U11880 (N_11880,N_8807,N_6443);
and U11881 (N_11881,N_7550,N_7949);
nand U11882 (N_11882,N_6616,N_7944);
nor U11883 (N_11883,N_6915,N_6811);
or U11884 (N_11884,N_8694,N_6782);
or U11885 (N_11885,N_6311,N_6368);
or U11886 (N_11886,N_7951,N_8241);
or U11887 (N_11887,N_6795,N_6592);
and U11888 (N_11888,N_8480,N_8150);
nor U11889 (N_11889,N_7720,N_6090);
and U11890 (N_11890,N_6807,N_6321);
nor U11891 (N_11891,N_6332,N_8390);
nand U11892 (N_11892,N_7298,N_6830);
xnor U11893 (N_11893,N_6255,N_6288);
nor U11894 (N_11894,N_6807,N_7382);
and U11895 (N_11895,N_7282,N_6302);
nor U11896 (N_11896,N_6385,N_7374);
and U11897 (N_11897,N_6939,N_8383);
or U11898 (N_11898,N_7866,N_6722);
or U11899 (N_11899,N_8534,N_6677);
and U11900 (N_11900,N_8254,N_6744);
nor U11901 (N_11901,N_8067,N_7624);
nand U11902 (N_11902,N_6305,N_6473);
nand U11903 (N_11903,N_6363,N_6453);
and U11904 (N_11904,N_8785,N_8371);
nor U11905 (N_11905,N_8599,N_8277);
nand U11906 (N_11906,N_8281,N_6360);
and U11907 (N_11907,N_7725,N_6897);
or U11908 (N_11908,N_7952,N_8628);
nor U11909 (N_11909,N_7324,N_6630);
and U11910 (N_11910,N_7098,N_7210);
nand U11911 (N_11911,N_7459,N_8474);
nor U11912 (N_11912,N_7314,N_8208);
or U11913 (N_11913,N_7289,N_8932);
and U11914 (N_11914,N_7267,N_6574);
and U11915 (N_11915,N_6363,N_6029);
and U11916 (N_11916,N_8525,N_7271);
or U11917 (N_11917,N_6782,N_8905);
xnor U11918 (N_11918,N_7068,N_7411);
or U11919 (N_11919,N_7189,N_6380);
nor U11920 (N_11920,N_6575,N_7257);
and U11921 (N_11921,N_6852,N_7335);
nand U11922 (N_11922,N_8877,N_7450);
and U11923 (N_11923,N_6987,N_8341);
nand U11924 (N_11924,N_8759,N_6553);
or U11925 (N_11925,N_7260,N_8290);
and U11926 (N_11926,N_6526,N_7735);
nor U11927 (N_11927,N_7790,N_6024);
and U11928 (N_11928,N_7780,N_7058);
nand U11929 (N_11929,N_6957,N_7108);
xor U11930 (N_11930,N_6912,N_6477);
or U11931 (N_11931,N_6016,N_6382);
nand U11932 (N_11932,N_8314,N_6358);
nand U11933 (N_11933,N_6675,N_8696);
and U11934 (N_11934,N_6940,N_7893);
and U11935 (N_11935,N_8716,N_8743);
or U11936 (N_11936,N_7448,N_7792);
and U11937 (N_11937,N_7709,N_7664);
nand U11938 (N_11938,N_6366,N_7478);
nand U11939 (N_11939,N_6502,N_6576);
and U11940 (N_11940,N_8104,N_6202);
nor U11941 (N_11941,N_8095,N_6664);
or U11942 (N_11942,N_8375,N_8713);
or U11943 (N_11943,N_8600,N_6706);
or U11944 (N_11944,N_8817,N_6215);
nand U11945 (N_11945,N_8097,N_8276);
or U11946 (N_11946,N_6821,N_8447);
xnor U11947 (N_11947,N_8866,N_6859);
xnor U11948 (N_11948,N_7152,N_8853);
and U11949 (N_11949,N_6785,N_8938);
or U11950 (N_11950,N_6265,N_6936);
or U11951 (N_11951,N_8588,N_6494);
nor U11952 (N_11952,N_6133,N_8206);
or U11953 (N_11953,N_7458,N_8483);
and U11954 (N_11954,N_8366,N_8485);
nor U11955 (N_11955,N_8176,N_6555);
xor U11956 (N_11956,N_7825,N_8330);
and U11957 (N_11957,N_7335,N_6037);
and U11958 (N_11958,N_8348,N_8294);
or U11959 (N_11959,N_7317,N_6106);
or U11960 (N_11960,N_6438,N_7416);
or U11961 (N_11961,N_6515,N_8258);
and U11962 (N_11962,N_6116,N_8137);
nor U11963 (N_11963,N_7229,N_7263);
and U11964 (N_11964,N_6605,N_7178);
nand U11965 (N_11965,N_6571,N_8245);
nand U11966 (N_11966,N_8699,N_8519);
nor U11967 (N_11967,N_6190,N_6174);
nand U11968 (N_11968,N_8297,N_6437);
or U11969 (N_11969,N_8291,N_7957);
and U11970 (N_11970,N_8870,N_7089);
nand U11971 (N_11971,N_6764,N_6794);
and U11972 (N_11972,N_7567,N_7109);
nor U11973 (N_11973,N_8175,N_8667);
nand U11974 (N_11974,N_6121,N_7351);
nor U11975 (N_11975,N_7686,N_8230);
or U11976 (N_11976,N_8763,N_7993);
and U11977 (N_11977,N_7139,N_8334);
nor U11978 (N_11978,N_7148,N_7609);
nor U11979 (N_11979,N_8628,N_6483);
and U11980 (N_11980,N_7409,N_6624);
and U11981 (N_11981,N_7414,N_7635);
nand U11982 (N_11982,N_8751,N_7810);
nor U11983 (N_11983,N_7211,N_8106);
xnor U11984 (N_11984,N_7842,N_8462);
and U11985 (N_11985,N_7077,N_6124);
xnor U11986 (N_11986,N_6341,N_7714);
and U11987 (N_11987,N_7245,N_6269);
and U11988 (N_11988,N_6071,N_7186);
xnor U11989 (N_11989,N_7930,N_8673);
and U11990 (N_11990,N_6665,N_7417);
nor U11991 (N_11991,N_8313,N_6938);
xor U11992 (N_11992,N_6101,N_8096);
nor U11993 (N_11993,N_8042,N_8414);
nand U11994 (N_11994,N_8245,N_8586);
xnor U11995 (N_11995,N_7172,N_6304);
or U11996 (N_11996,N_8370,N_8598);
nand U11997 (N_11997,N_7069,N_6637);
nor U11998 (N_11998,N_8255,N_7945);
nor U11999 (N_11999,N_8891,N_6783);
and U12000 (N_12000,N_9689,N_11119);
and U12001 (N_12001,N_9198,N_9555);
nor U12002 (N_12002,N_9662,N_9974);
or U12003 (N_12003,N_9395,N_9569);
nor U12004 (N_12004,N_9730,N_9201);
nand U12005 (N_12005,N_9603,N_10334);
or U12006 (N_12006,N_9690,N_10291);
nor U12007 (N_12007,N_11920,N_10381);
nand U12008 (N_12008,N_10131,N_9746);
nand U12009 (N_12009,N_9670,N_11616);
and U12010 (N_12010,N_11514,N_9303);
and U12011 (N_12011,N_9350,N_11880);
or U12012 (N_12012,N_9669,N_10156);
nand U12013 (N_12013,N_10403,N_10915);
nor U12014 (N_12014,N_10786,N_11744);
nand U12015 (N_12015,N_9728,N_9848);
nor U12016 (N_12016,N_11445,N_11135);
xnor U12017 (N_12017,N_11216,N_11888);
or U12018 (N_12018,N_9786,N_9164);
nor U12019 (N_12019,N_10204,N_9561);
or U12020 (N_12020,N_11309,N_9267);
nor U12021 (N_12021,N_9089,N_11193);
nand U12022 (N_12022,N_10867,N_11863);
and U12023 (N_12023,N_11368,N_10388);
xnor U12024 (N_12024,N_10792,N_10329);
nand U12025 (N_12025,N_9487,N_11221);
and U12026 (N_12026,N_9485,N_10695);
and U12027 (N_12027,N_10583,N_11894);
nor U12028 (N_12028,N_10872,N_11025);
nand U12029 (N_12029,N_9191,N_9241);
and U12030 (N_12030,N_10449,N_10524);
and U12031 (N_12031,N_10154,N_11434);
nand U12032 (N_12032,N_10511,N_11364);
or U12033 (N_12033,N_10039,N_10272);
or U12034 (N_12034,N_10262,N_9006);
or U12035 (N_12035,N_10495,N_11977);
or U12036 (N_12036,N_10557,N_11294);
nand U12037 (N_12037,N_9770,N_10653);
xor U12038 (N_12038,N_11254,N_11873);
nor U12039 (N_12039,N_9927,N_9389);
nor U12040 (N_12040,N_10116,N_10554);
nor U12041 (N_12041,N_10103,N_11029);
nand U12042 (N_12042,N_11056,N_9245);
nand U12043 (N_12043,N_9254,N_10568);
or U12044 (N_12044,N_9323,N_9454);
and U12045 (N_12045,N_11592,N_10913);
nand U12046 (N_12046,N_10151,N_11341);
and U12047 (N_12047,N_9217,N_11027);
and U12048 (N_12048,N_11844,N_9824);
and U12049 (N_12049,N_9257,N_10491);
nand U12050 (N_12050,N_9192,N_9953);
nand U12051 (N_12051,N_11186,N_9731);
and U12052 (N_12052,N_10532,N_9322);
nor U12053 (N_12053,N_11635,N_11628);
and U12054 (N_12054,N_9070,N_10119);
nand U12055 (N_12055,N_10161,N_11022);
xnor U12056 (N_12056,N_11702,N_9744);
nor U12057 (N_12057,N_10207,N_9961);
nor U12058 (N_12058,N_11982,N_11596);
xor U12059 (N_12059,N_9204,N_10410);
xnor U12060 (N_12060,N_9686,N_10470);
and U12061 (N_12061,N_10299,N_10167);
nand U12062 (N_12062,N_11480,N_9931);
and U12063 (N_12063,N_10603,N_10916);
and U12064 (N_12064,N_10307,N_10331);
nand U12065 (N_12065,N_9993,N_9171);
or U12066 (N_12066,N_10973,N_11741);
nand U12067 (N_12067,N_9236,N_10644);
nand U12068 (N_12068,N_9610,N_9720);
or U12069 (N_12069,N_9685,N_11330);
and U12070 (N_12070,N_11849,N_10084);
nand U12071 (N_12071,N_11952,N_9157);
and U12072 (N_12072,N_10674,N_10088);
and U12073 (N_12073,N_10178,N_11639);
and U12074 (N_12074,N_11542,N_9562);
and U12075 (N_12075,N_10337,N_9664);
and U12076 (N_12076,N_11381,N_11013);
and U12077 (N_12077,N_10621,N_11566);
nor U12078 (N_12078,N_10487,N_11719);
nand U12079 (N_12079,N_11537,N_9736);
and U12080 (N_12080,N_10046,N_9626);
nor U12081 (N_12081,N_11290,N_10360);
and U12082 (N_12082,N_9873,N_10545);
nor U12083 (N_12083,N_10268,N_11005);
or U12084 (N_12084,N_10666,N_10997);
and U12085 (N_12085,N_10376,N_9379);
or U12086 (N_12086,N_9392,N_10591);
nand U12087 (N_12087,N_10816,N_9806);
nor U12088 (N_12088,N_11520,N_11436);
nor U12089 (N_12089,N_9028,N_10781);
nor U12090 (N_12090,N_10411,N_10966);
nand U12091 (N_12091,N_11040,N_10009);
nand U12092 (N_12092,N_10395,N_10089);
nor U12093 (N_12093,N_9694,N_11021);
or U12094 (N_12094,N_10054,N_9699);
or U12095 (N_12095,N_11404,N_9503);
and U12096 (N_12096,N_11804,N_10122);
or U12097 (N_12097,N_11623,N_11041);
nand U12098 (N_12098,N_11107,N_10308);
nand U12099 (N_12099,N_11337,N_10121);
nor U12100 (N_12100,N_10622,N_9166);
nor U12101 (N_12101,N_11698,N_11223);
xor U12102 (N_12102,N_10830,N_10118);
and U12103 (N_12103,N_9834,N_11806);
nand U12104 (N_12104,N_10418,N_10798);
and U12105 (N_12105,N_9879,N_10908);
nor U12106 (N_12106,N_9889,N_9698);
nor U12107 (N_12107,N_10412,N_9176);
or U12108 (N_12108,N_11609,N_10738);
nor U12109 (N_12109,N_9839,N_10964);
or U12110 (N_12110,N_9109,N_10726);
nor U12111 (N_12111,N_10895,N_10928);
nand U12112 (N_12112,N_10701,N_11078);
and U12113 (N_12113,N_10098,N_11438);
nor U12114 (N_12114,N_10139,N_9156);
and U12115 (N_12115,N_11295,N_9572);
or U12116 (N_12116,N_9384,N_9570);
xnor U12117 (N_12117,N_10101,N_10157);
nor U12118 (N_12118,N_11509,N_9508);
and U12119 (N_12119,N_11482,N_11988);
nor U12120 (N_12120,N_9058,N_10905);
and U12121 (N_12121,N_11594,N_10092);
nand U12122 (N_12122,N_11811,N_9712);
and U12123 (N_12123,N_11731,N_9039);
or U12124 (N_12124,N_9856,N_11046);
and U12125 (N_12125,N_9059,N_11069);
and U12126 (N_12126,N_10043,N_9026);
or U12127 (N_12127,N_9009,N_11419);
xnor U12128 (N_12128,N_9130,N_11978);
and U12129 (N_12129,N_9695,N_10227);
or U12130 (N_12130,N_10011,N_10649);
nand U12131 (N_12131,N_9709,N_10069);
nand U12132 (N_12132,N_9423,N_11966);
xnor U12133 (N_12133,N_10284,N_10764);
nor U12134 (N_12134,N_11817,N_10359);
nor U12135 (N_12135,N_11389,N_11864);
or U12136 (N_12136,N_11053,N_9901);
or U12137 (N_12137,N_10193,N_11211);
or U12138 (N_12138,N_10454,N_9148);
and U12139 (N_12139,N_10680,N_11585);
nand U12140 (N_12140,N_11410,N_11933);
nand U12141 (N_12141,N_10433,N_9511);
or U12142 (N_12142,N_11887,N_11174);
or U12143 (N_12143,N_9928,N_10091);
xnor U12144 (N_12144,N_11175,N_11802);
or U12145 (N_12145,N_9776,N_9755);
nand U12146 (N_12146,N_9173,N_9808);
nand U12147 (N_12147,N_9894,N_10825);
or U12148 (N_12148,N_10108,N_9683);
or U12149 (N_12149,N_11260,N_11365);
nand U12150 (N_12150,N_9718,N_9262);
nor U12151 (N_12151,N_10006,N_11975);
and U12152 (N_12152,N_10063,N_11197);
and U12153 (N_12153,N_9319,N_9134);
or U12154 (N_12154,N_9108,N_9781);
nand U12155 (N_12155,N_11536,N_10828);
xor U12156 (N_12156,N_11421,N_11766);
nor U12157 (N_12157,N_10215,N_11997);
or U12158 (N_12158,N_9253,N_10181);
nand U12159 (N_12159,N_11296,N_9172);
nor U12160 (N_12160,N_10717,N_11976);
nor U12161 (N_12161,N_9393,N_9499);
or U12162 (N_12162,N_10507,N_11753);
xnor U12163 (N_12163,N_10567,N_9643);
or U12164 (N_12164,N_10796,N_10897);
nand U12165 (N_12165,N_11358,N_11469);
or U12166 (N_12166,N_11557,N_10014);
and U12167 (N_12167,N_11406,N_9126);
or U12168 (N_12168,N_9283,N_11108);
and U12169 (N_12169,N_9490,N_11904);
nor U12170 (N_12170,N_11762,N_10348);
or U12171 (N_12171,N_10580,N_9729);
nand U12172 (N_12172,N_9999,N_9275);
or U12173 (N_12173,N_9002,N_9910);
and U12174 (N_12174,N_11048,N_11556);
nand U12175 (N_12175,N_10851,N_11467);
xor U12176 (N_12176,N_9819,N_10080);
nor U12177 (N_12177,N_10049,N_9365);
nor U12178 (N_12178,N_11477,N_10559);
and U12179 (N_12179,N_9850,N_10231);
xor U12180 (N_12180,N_10102,N_9483);
nor U12181 (N_12181,N_11986,N_9977);
xnor U12182 (N_12182,N_10310,N_10956);
nor U12183 (N_12183,N_10140,N_9525);
nand U12184 (N_12184,N_10561,N_11170);
and U12185 (N_12185,N_11209,N_11552);
nor U12186 (N_12186,N_10222,N_11889);
nor U12187 (N_12187,N_10074,N_10574);
nand U12188 (N_12188,N_9722,N_11739);
or U12189 (N_12189,N_10317,N_11336);
or U12190 (N_12190,N_10247,N_11190);
nand U12191 (N_12191,N_11661,N_9015);
nand U12192 (N_12192,N_10045,N_11716);
xor U12193 (N_12193,N_11265,N_10078);
and U12194 (N_12194,N_9587,N_9925);
nor U12195 (N_12195,N_10129,N_11916);
and U12196 (N_12196,N_9450,N_11924);
nor U12197 (N_12197,N_9445,N_10171);
nor U12198 (N_12198,N_10489,N_9593);
nor U12199 (N_12199,N_11014,N_10893);
nand U12200 (N_12200,N_9214,N_11906);
nand U12201 (N_12201,N_11574,N_11865);
nand U12202 (N_12202,N_9747,N_9964);
and U12203 (N_12203,N_11447,N_11637);
and U12204 (N_12204,N_10233,N_11163);
nor U12205 (N_12205,N_9601,N_9589);
and U12206 (N_12206,N_9252,N_10292);
nand U12207 (N_12207,N_9458,N_11625);
nor U12208 (N_12208,N_9578,N_10048);
and U12209 (N_12209,N_9622,N_10585);
nand U12210 (N_12210,N_10326,N_11159);
nor U12211 (N_12211,N_9213,N_11981);
nor U12212 (N_12212,N_10994,N_9631);
or U12213 (N_12213,N_10052,N_9372);
or U12214 (N_12214,N_11302,N_11738);
nand U12215 (N_12215,N_9543,N_11036);
and U12216 (N_12216,N_9607,N_11973);
xnor U12217 (N_12217,N_10422,N_9829);
nor U12218 (N_12218,N_11416,N_10221);
nor U12219 (N_12219,N_11532,N_10976);
nand U12220 (N_12220,N_9051,N_9361);
and U12221 (N_12221,N_9835,N_11782);
and U12222 (N_12222,N_11886,N_9138);
nor U12223 (N_12223,N_11922,N_9987);
nand U12224 (N_12224,N_10390,N_10345);
or U12225 (N_12225,N_11602,N_10393);
nor U12226 (N_12226,N_10279,N_9674);
or U12227 (N_12227,N_10939,N_9069);
or U12228 (N_12228,N_9795,N_9875);
nor U12229 (N_12229,N_11508,N_11359);
or U12230 (N_12230,N_10197,N_9628);
nand U12231 (N_12231,N_11678,N_11343);
xor U12232 (N_12232,N_10703,N_10175);
nand U12233 (N_12233,N_11736,N_10737);
or U12234 (N_12234,N_11052,N_11909);
nand U12235 (N_12235,N_11481,N_10216);
nor U12236 (N_12236,N_10620,N_9491);
or U12237 (N_12237,N_11881,N_11286);
or U12238 (N_12238,N_10025,N_10068);
and U12239 (N_12239,N_10773,N_11009);
xor U12240 (N_12240,N_11861,N_10637);
or U12241 (N_12241,N_9013,N_10278);
nand U12242 (N_12242,N_9595,N_11092);
nor U12243 (N_12243,N_9853,N_10484);
nand U12244 (N_12244,N_10750,N_9778);
nor U12245 (N_12245,N_11905,N_9012);
or U12246 (N_12246,N_11100,N_9400);
xnor U12247 (N_12247,N_9549,N_9453);
nor U12248 (N_12248,N_9190,N_10318);
and U12249 (N_12249,N_11824,N_11113);
nand U12250 (N_12250,N_11323,N_9513);
and U12251 (N_12251,N_11554,N_11334);
and U12252 (N_12252,N_9957,N_10691);
and U12253 (N_12253,N_11696,N_11506);
and U12254 (N_12254,N_9340,N_10041);
nor U12255 (N_12255,N_9127,N_10423);
and U12256 (N_12256,N_9004,N_10671);
or U12257 (N_12257,N_9331,N_11312);
nor U12258 (N_12258,N_10364,N_10768);
and U12259 (N_12259,N_10351,N_11161);
nor U12260 (N_12260,N_11649,N_9019);
or U12261 (N_12261,N_10571,N_10944);
xnor U12262 (N_12262,N_11152,N_9760);
or U12263 (N_12263,N_10625,N_9202);
or U12264 (N_12264,N_10237,N_9588);
nand U12265 (N_12265,N_9300,N_11394);
and U12266 (N_12266,N_11533,N_11812);
nor U12267 (N_12267,N_11491,N_9355);
nand U12268 (N_12268,N_10904,N_9655);
or U12269 (N_12269,N_11856,N_11183);
nor U12270 (N_12270,N_10142,N_11495);
or U12271 (N_12271,N_11023,N_10022);
and U12272 (N_12272,N_10001,N_10341);
and U12273 (N_12273,N_9529,N_9212);
or U12274 (N_12274,N_9510,N_11751);
and U12275 (N_12275,N_9658,N_9633);
and U12276 (N_12276,N_10060,N_9207);
and U12277 (N_12277,N_10678,N_9412);
nor U12278 (N_12278,N_9542,N_11130);
nand U12279 (N_12279,N_9544,N_9494);
xor U12280 (N_12280,N_11417,N_11051);
nor U12281 (N_12281,N_11383,N_10479);
and U12282 (N_12282,N_9992,N_10981);
xor U12283 (N_12283,N_10255,N_10465);
and U12284 (N_12284,N_11167,N_9823);
nand U12285 (N_12285,N_11611,N_11391);
nor U12286 (N_12286,N_10455,N_11985);
or U12287 (N_12287,N_9291,N_9660);
and U12288 (N_12288,N_9014,N_10898);
nand U12289 (N_12289,N_11274,N_9566);
or U12290 (N_12290,N_10642,N_11665);
and U12291 (N_12291,N_10824,N_9251);
nor U12292 (N_12292,N_11143,N_9584);
or U12293 (N_12293,N_11805,N_10028);
nor U12294 (N_12294,N_9264,N_11188);
or U12295 (N_12295,N_10126,N_10055);
or U12296 (N_12296,N_9041,N_11354);
and U12297 (N_12297,N_9533,N_11489);
or U12298 (N_12298,N_9536,N_11243);
nand U12299 (N_12299,N_10845,N_10784);
nand U12300 (N_12300,N_10040,N_10841);
xor U12301 (N_12301,N_9416,N_10361);
and U12302 (N_12302,N_9055,N_9863);
and U12303 (N_12303,N_9946,N_10076);
nor U12304 (N_12304,N_9713,N_10529);
or U12305 (N_12305,N_10244,N_9318);
or U12306 (N_12306,N_10117,N_11387);
xnor U12307 (N_12307,N_11499,N_11786);
or U12308 (N_12308,N_9272,N_11775);
and U12309 (N_12309,N_10270,N_9527);
and U12310 (N_12310,N_11821,N_9723);
and U12311 (N_12311,N_9305,N_10837);
xor U12312 (N_12312,N_11373,N_10606);
and U12313 (N_12313,N_11422,N_10544);
nand U12314 (N_12314,N_10892,N_10431);
or U12315 (N_12315,N_9313,N_9158);
nor U12316 (N_12316,N_11995,N_9937);
nand U12317 (N_12317,N_10473,N_9955);
nor U12318 (N_12318,N_9500,N_11194);
and U12319 (N_12319,N_9609,N_9507);
and U12320 (N_12320,N_11385,N_9103);
and U12321 (N_12321,N_9452,N_11897);
and U12322 (N_12322,N_11727,N_11384);
nand U12323 (N_12323,N_10772,N_9758);
nand U12324 (N_12324,N_9401,N_11043);
nor U12325 (N_12325,N_9209,N_10120);
nand U12326 (N_12326,N_11693,N_9611);
xnor U12327 (N_12327,N_11841,N_10609);
nor U12328 (N_12328,N_10300,N_11714);
and U12329 (N_12329,N_9606,N_11362);
nand U12330 (N_12330,N_10462,N_10400);
or U12331 (N_12331,N_9552,N_10296);
and U12332 (N_12332,N_10718,N_9762);
or U12333 (N_12333,N_9440,N_9288);
nor U12334 (N_12334,N_11768,N_9676);
or U12335 (N_12335,N_11031,N_9310);
nand U12336 (N_12336,N_9700,N_10560);
xnor U12337 (N_12337,N_10767,N_9942);
nor U12338 (N_12338,N_9205,N_11610);
and U12339 (N_12339,N_9738,N_11112);
or U12340 (N_12340,N_10812,N_9558);
or U12341 (N_12341,N_10763,N_11346);
nor U12342 (N_12342,N_10790,N_9515);
nor U12343 (N_12343,N_11285,N_9680);
or U12344 (N_12344,N_9667,N_9968);
or U12345 (N_12345,N_9276,N_9696);
or U12346 (N_12346,N_11672,N_11444);
nor U12347 (N_12347,N_11063,N_10371);
nand U12348 (N_12348,N_10230,N_11129);
or U12349 (N_12349,N_9029,N_10182);
nor U12350 (N_12350,N_10205,N_10506);
or U12351 (N_12351,N_11634,N_11452);
or U12352 (N_12352,N_9421,N_9329);
nor U12353 (N_12353,N_9080,N_9324);
xnor U12354 (N_12354,N_10192,N_9582);
xor U12355 (N_12355,N_10152,N_11272);
and U12356 (N_12356,N_10459,N_11002);
or U12357 (N_12357,N_11972,N_9597);
or U12358 (N_12358,N_11626,N_11244);
xor U12359 (N_12359,N_9887,N_10373);
or U12360 (N_12360,N_9362,N_11248);
and U12361 (N_12361,N_11748,N_11195);
nor U12362 (N_12362,N_10782,N_11870);
nor U12363 (N_12363,N_11456,N_10107);
nand U12364 (N_12364,N_10385,N_10632);
or U12365 (N_12365,N_11466,N_11879);
or U12366 (N_12366,N_10936,N_9299);
or U12367 (N_12367,N_11987,N_9710);
or U12368 (N_12368,N_11049,N_10271);
and U12369 (N_12369,N_9949,N_10200);
and U12370 (N_12370,N_9088,N_11613);
nor U12371 (N_12371,N_11034,N_10190);
nand U12372 (N_12372,N_10518,N_9818);
xor U12373 (N_12373,N_10293,N_9016);
or U12374 (N_12374,N_11529,N_9085);
nand U12375 (N_12375,N_10443,N_11640);
nor U12376 (N_12376,N_9492,N_11517);
xor U12377 (N_12377,N_11430,N_9040);
nand U12378 (N_12378,N_11237,N_10732);
nor U12379 (N_12379,N_9225,N_10934);
or U12380 (N_12380,N_9404,N_10514);
xor U12381 (N_12381,N_10413,N_10747);
or U12382 (N_12382,N_11468,N_11131);
nand U12383 (N_12383,N_9419,N_10807);
nand U12384 (N_12384,N_10212,N_10971);
nor U12385 (N_12385,N_10987,N_9789);
or U12386 (N_12386,N_9197,N_10010);
nor U12387 (N_12387,N_10809,N_9281);
or U12388 (N_12388,N_10957,N_9801);
and U12389 (N_12389,N_9477,N_9470);
and U12390 (N_12390,N_11019,N_11086);
nand U12391 (N_12391,N_10409,N_11356);
or U12392 (N_12392,N_10087,N_11307);
nor U12393 (N_12393,N_10819,N_9541);
or U12394 (N_12394,N_11726,N_10958);
nand U12395 (N_12395,N_10970,N_10508);
nor U12396 (N_12396,N_9017,N_11701);
and U12397 (N_12397,N_11728,N_9495);
and U12398 (N_12398,N_10760,N_9433);
nor U12399 (N_12399,N_10705,N_10498);
or U12400 (N_12400,N_11098,N_9258);
nand U12401 (N_12401,N_9153,N_11379);
or U12402 (N_12402,N_11217,N_9708);
or U12403 (N_12403,N_9881,N_10275);
nor U12404 (N_12404,N_10594,N_11443);
nor U12405 (N_12405,N_10616,N_10922);
or U12406 (N_12406,N_10062,N_11154);
or U12407 (N_12407,N_9360,N_9346);
nor U12408 (N_12408,N_9897,N_10196);
and U12409 (N_12409,N_10176,N_9864);
and U12410 (N_12410,N_11746,N_10150);
nand U12411 (N_12411,N_11666,N_11671);
and U12412 (N_12412,N_9199,N_10093);
nor U12413 (N_12413,N_9571,N_10864);
and U12414 (N_12414,N_10287,N_10871);
or U12415 (N_12415,N_9037,N_9074);
nor U12416 (N_12416,N_10327,N_11965);
or U12417 (N_12417,N_9087,N_9091);
nor U12418 (N_12418,N_10739,N_11488);
and U12419 (N_12419,N_10505,N_11968);
and U12420 (N_12420,N_9739,N_10111);
nor U12421 (N_12421,N_9915,N_10562);
nand U12422 (N_12422,N_10914,N_10324);
and U12423 (N_12423,N_11471,N_9046);
and U12424 (N_12424,N_11771,N_9586);
and U12425 (N_12425,N_11835,N_9327);
nand U12426 (N_12426,N_11442,N_9926);
or U12427 (N_12427,N_10408,N_11939);
and U12428 (N_12428,N_11273,N_9996);
nor U12429 (N_12429,N_9282,N_11589);
nor U12430 (N_12430,N_9556,N_10597);
xor U12431 (N_12431,N_11721,N_11655);
nand U12432 (N_12432,N_10463,N_9725);
or U12433 (N_12433,N_11711,N_11549);
or U12434 (N_12434,N_11527,N_9785);
nand U12435 (N_12435,N_10382,N_9733);
nand U12436 (N_12436,N_11038,N_10984);
and U12437 (N_12437,N_9304,N_10810);
xor U12438 (N_12438,N_11277,N_10829);
and U12439 (N_12439,N_9005,N_10047);
xnor U12440 (N_12440,N_10659,N_10995);
nor U12441 (N_12441,N_10607,N_9090);
or U12442 (N_12442,N_11572,N_11578);
nor U12443 (N_12443,N_10015,N_11951);
nor U12444 (N_12444,N_10243,N_10700);
nor U12445 (N_12445,N_11629,N_9938);
nand U12446 (N_12446,N_10124,N_9737);
nand U12447 (N_12447,N_9001,N_10269);
and U12448 (N_12448,N_9576,N_11949);
and U12449 (N_12449,N_9751,N_9451);
or U12450 (N_12450,N_11937,N_9383);
and U12451 (N_12451,N_9519,N_11010);
nor U12452 (N_12452,N_9054,N_10234);
or U12453 (N_12453,N_11658,N_11868);
nor U12454 (N_12454,N_10058,N_9973);
xnor U12455 (N_12455,N_10744,N_11301);
nand U12456 (N_12456,N_11929,N_10723);
nand U12457 (N_12457,N_11297,N_10902);
xnor U12458 (N_12458,N_9101,N_9935);
nand U12459 (N_12459,N_10213,N_11134);
nand U12460 (N_12460,N_10826,N_10467);
nand U12461 (N_12461,N_11462,N_9547);
and U12462 (N_12462,N_10840,N_11180);
xnor U12463 (N_12463,N_10657,N_9625);
nor U12464 (N_12464,N_10950,N_11440);
and U12465 (N_12465,N_10662,N_11411);
and U12466 (N_12466,N_9128,N_9447);
or U12467 (N_12467,N_10512,N_10194);
or U12468 (N_12468,N_9446,N_10123);
nor U12469 (N_12469,N_11798,N_10394);
and U12470 (N_12470,N_9902,N_10881);
xnor U12471 (N_12471,N_9098,N_11843);
nand U12472 (N_12472,N_11355,N_11528);
xor U12473 (N_12473,N_9271,N_10766);
or U12474 (N_12474,N_9203,N_10004);
nor U12475 (N_12475,N_9971,N_9025);
xor U12476 (N_12476,N_11245,N_9697);
or U12477 (N_12477,N_9124,N_10785);
and U12478 (N_12478,N_9984,N_9514);
nor U12479 (N_12479,N_10249,N_9430);
nand U12480 (N_12480,N_9408,N_11024);
and U12481 (N_12481,N_11213,N_9684);
nor U12482 (N_12482,N_10309,N_11374);
nand U12483 (N_12483,N_9208,N_9765);
or U12484 (N_12484,N_10406,N_9820);
nor U12485 (N_12485,N_11316,N_11974);
and U12486 (N_12486,N_10754,N_9261);
nand U12487 (N_12487,N_11901,N_9704);
and U12488 (N_12488,N_11115,N_10177);
nand U12489 (N_12489,N_11559,N_9121);
and U12490 (N_12490,N_11765,N_9285);
and U12491 (N_12491,N_11016,N_11749);
nand U12492 (N_12492,N_10064,N_11291);
nand U12493 (N_12493,N_9979,N_10668);
or U12494 (N_12494,N_10099,N_9232);
or U12495 (N_12495,N_9443,N_9076);
xor U12496 (N_12496,N_10502,N_11000);
nand U12497 (N_12497,N_9356,N_10709);
nand U12498 (N_12498,N_11020,N_11867);
and U12499 (N_12499,N_9010,N_10547);
xnor U12500 (N_12500,N_11651,N_11058);
and U12501 (N_12501,N_9096,N_11799);
and U12502 (N_12502,N_10734,N_11282);
nor U12503 (N_12503,N_11278,N_10918);
nor U12504 (N_12504,N_10745,N_9229);
xnor U12505 (N_12505,N_10073,N_11750);
nand U12506 (N_12506,N_10127,N_10855);
or U12507 (N_12507,N_9888,N_11007);
nand U12508 (N_12508,N_9613,N_10702);
or U12509 (N_12509,N_9526,N_11090);
nor U12510 (N_12510,N_10096,N_11455);
xor U12511 (N_12511,N_11641,N_11118);
or U12512 (N_12512,N_11032,N_10930);
xnor U12513 (N_12513,N_10982,N_9255);
nand U12514 (N_12514,N_10619,N_9193);
nor U12515 (N_12515,N_11697,N_9954);
nand U12516 (N_12516,N_9211,N_11247);
nor U12517 (N_12517,N_11268,N_11133);
nor U12518 (N_12518,N_9706,N_10294);
and U12519 (N_12519,N_10397,N_11555);
nand U12520 (N_12520,N_9565,N_10541);
or U12521 (N_12521,N_11059,N_10788);
and U12522 (N_12522,N_11874,N_10094);
or U12523 (N_12523,N_11795,N_11877);
nand U12524 (N_12524,N_9874,N_10573);
and U12525 (N_12525,N_10253,N_10776);
nor U12526 (N_12526,N_11931,N_9668);
nor U12527 (N_12527,N_10890,N_10624);
and U12528 (N_12528,N_9899,N_10229);
nor U12529 (N_12529,N_10708,N_9377);
and U12530 (N_12530,N_11126,N_11314);
nor U12531 (N_12531,N_11720,N_11483);
and U12532 (N_12532,N_11747,N_9293);
nor U12533 (N_12533,N_9024,N_10274);
nand U12534 (N_12534,N_11754,N_11093);
and U12535 (N_12535,N_10602,N_9775);
xnor U12536 (N_12536,N_11512,N_11485);
and U12537 (N_12537,N_10527,N_11936);
nor U12538 (N_12538,N_11699,N_9932);
and U12539 (N_12539,N_9036,N_11028);
and U12540 (N_12540,N_11777,N_11648);
nand U12541 (N_12541,N_11124,N_10224);
nor U12542 (N_12542,N_10053,N_11519);
or U12543 (N_12543,N_11769,N_10538);
xor U12544 (N_12544,N_9339,N_10974);
nand U12545 (N_12545,N_10716,N_11703);
nor U12546 (N_12546,N_10615,N_9518);
and U12547 (N_12547,N_11878,N_9481);
and U12548 (N_12548,N_10596,N_11723);
or U12549 (N_12549,N_9616,N_10569);
and U12550 (N_12550,N_9065,N_10611);
or U12551 (N_12551,N_9311,N_10805);
and U12552 (N_12552,N_10319,N_11262);
nor U12553 (N_12553,N_10884,N_9991);
xnor U12554 (N_12554,N_11601,N_9661);
nor U12555 (N_12555,N_11476,N_9548);
or U12556 (N_12556,N_10550,N_9779);
or U12557 (N_12557,N_11944,N_10852);
or U12558 (N_12558,N_9629,N_11246);
nor U12559 (N_12559,N_9575,N_9943);
or U12560 (N_12560,N_10687,N_10832);
and U12561 (N_12561,N_11191,N_10067);
and U12562 (N_12562,N_10426,N_9998);
nand U12563 (N_12563,N_11287,N_9852);
and U12564 (N_12564,N_10605,N_10651);
or U12565 (N_12565,N_9184,N_9071);
and U12566 (N_12566,N_9768,N_11376);
nor U12567 (N_12567,N_10880,N_10138);
nor U12568 (N_12568,N_9844,N_11380);
and U12569 (N_12569,N_9306,N_11664);
xor U12570 (N_12570,N_10630,N_10189);
nand U12571 (N_12571,N_9239,N_10748);
nand U12572 (N_12572,N_11583,N_10343);
nand U12573 (N_12573,N_9743,N_9467);
or U12574 (N_12574,N_10572,N_10937);
nor U12575 (N_12575,N_10374,N_11498);
and U12576 (N_12576,N_10565,N_10488);
or U12577 (N_12577,N_11015,N_11187);
and U12578 (N_12578,N_10889,N_9620);
nor U12579 (N_12579,N_10460,N_10600);
nor U12580 (N_12580,N_9246,N_9780);
nand U12581 (N_12581,N_11125,N_11827);
nor U12582 (N_12582,N_11785,N_11101);
nor U12583 (N_12583,N_11686,N_11891);
and U12584 (N_12584,N_11571,N_11429);
nor U12585 (N_12585,N_11839,N_10464);
or U12586 (N_12586,N_10513,N_9226);
or U12587 (N_12587,N_10697,N_10203);
nand U12588 (N_12588,N_11921,N_11600);
and U12589 (N_12589,N_9259,N_9425);
nand U12590 (N_12590,N_11065,N_10827);
xor U12591 (N_12591,N_9374,N_9247);
nor U12592 (N_12592,N_10715,N_10985);
and U12593 (N_12593,N_9624,N_9132);
nand U12594 (N_12594,N_9783,N_11967);
nand U12595 (N_12595,N_11172,N_10090);
nor U12596 (N_12596,N_10008,N_9898);
nor U12597 (N_12597,N_10515,N_10149);
nor U12598 (N_12598,N_9917,N_11970);
and U12599 (N_12599,N_11816,N_11333);
and U12600 (N_12600,N_11926,N_10404);
xor U12601 (N_12601,N_11755,N_10686);
nor U12602 (N_12602,N_10342,N_9174);
nor U12603 (N_12603,N_9681,N_10992);
xnor U12604 (N_12604,N_9434,N_11962);
or U12605 (N_12605,N_11963,N_11790);
nor U12606 (N_12606,N_11928,N_9114);
or U12607 (N_12607,N_11650,N_11079);
nor U12608 (N_12608,N_9210,N_9409);
nand U12609 (N_12609,N_10283,N_11474);
or U12610 (N_12610,N_11008,N_9813);
and U12611 (N_12611,N_11622,N_9859);
nor U12612 (N_12612,N_10147,N_10935);
nor U12613 (N_12613,N_10952,N_10164);
nand U12614 (N_12614,N_9905,N_10155);
nand U12615 (N_12615,N_11207,N_11178);
or U12616 (N_12616,N_11204,N_11150);
and U12617 (N_12617,N_11173,N_11845);
xor U12618 (N_12618,N_9638,N_10862);
xor U12619 (N_12619,N_11420,N_10929);
and U12620 (N_12620,N_11820,N_9117);
or U12621 (N_12621,N_9717,N_10743);
or U12622 (N_12622,N_9914,N_11250);
and U12623 (N_12623,N_11940,N_10191);
nand U12624 (N_12624,N_11801,N_10771);
or U12625 (N_12625,N_10999,N_10235);
or U12626 (N_12626,N_10379,N_11494);
nand U12627 (N_12627,N_10258,N_10378);
and U12628 (N_12628,N_10339,N_10114);
or U12629 (N_12629,N_11823,N_10416);
nor U12630 (N_12630,N_10013,N_11513);
or U12631 (N_12631,N_11203,N_10592);
nand U12632 (N_12632,N_11534,N_10711);
and U12633 (N_12633,N_11369,N_9671);
and U12634 (N_12634,N_11776,N_9123);
or U12635 (N_12635,N_10806,N_11045);
or U12636 (N_12636,N_10775,N_10245);
nand U12637 (N_12637,N_10587,N_10104);
or U12638 (N_12638,N_9034,N_11446);
or U12639 (N_12639,N_9165,N_9033);
or U12640 (N_12640,N_10021,N_10163);
nand U12641 (N_12641,N_9749,N_9265);
xor U12642 (N_12642,N_10330,N_11587);
nand U12643 (N_12643,N_9936,N_9402);
nor U12644 (N_12644,N_9086,N_9179);
nor U12645 (N_12645,N_9719,N_11866);
nand U12646 (N_12646,N_11450,N_10349);
nand U12647 (N_12647,N_11925,N_9438);
nor U12648 (N_12648,N_9693,N_11151);
and U12649 (N_12649,N_11054,N_9099);
nor U12650 (N_12650,N_9960,N_11454);
or U12651 (N_12651,N_11809,N_10598);
nand U12652 (N_12652,N_9237,N_11784);
and U12653 (N_12653,N_11690,N_11327);
nand U12654 (N_12654,N_11675,N_11251);
nand U12655 (N_12655,N_10778,N_11996);
nand U12656 (N_12656,N_10436,N_9814);
or U12657 (N_12657,N_11772,N_9883);
or U12658 (N_12658,N_9314,N_10850);
nor U12659 (N_12659,N_10831,N_9878);
xnor U12660 (N_12660,N_9284,N_10266);
and U12661 (N_12661,N_11618,N_9627);
nor U12662 (N_12662,N_9678,N_10012);
nor U12663 (N_12663,N_10026,N_10500);
xnor U12664 (N_12664,N_11834,N_9439);
nor U12665 (N_12665,N_11903,N_10130);
and U12666 (N_12666,N_9068,N_9995);
and U12667 (N_12667,N_10162,N_10886);
or U12668 (N_12668,N_9044,N_10802);
or U12669 (N_12669,N_10391,N_9959);
nand U12670 (N_12670,N_10578,N_9592);
nand U12671 (N_12671,N_10660,N_9950);
nor U12672 (N_12672,N_10617,N_10721);
xnor U12673 (N_12673,N_11950,N_9672);
or U12674 (N_12674,N_11465,N_10912);
xnor U12675 (N_12675,N_11470,N_10219);
nand U12676 (N_12676,N_11345,N_11215);
or U12677 (N_12677,N_9777,N_10938);
xnor U12678 (N_12678,N_10654,N_11707);
nor U12679 (N_12679,N_10882,N_9828);
and U12680 (N_12680,N_9978,N_9150);
nand U12681 (N_12681,N_10943,N_11633);
or U12682 (N_12682,N_11396,N_9388);
nor U12683 (N_12683,N_11388,N_10146);
and U12684 (N_12684,N_11523,N_11403);
nor U12685 (N_12685,N_9260,N_9682);
xnor U12686 (N_12686,N_11710,N_9465);
xnor U12687 (N_12687,N_11145,N_11424);
and U12688 (N_12688,N_10870,N_10321);
nor U12689 (N_12689,N_9185,N_10202);
nand U12690 (N_12690,N_10853,N_9767);
or U12691 (N_12691,N_9429,N_11234);
and U12692 (N_12692,N_11851,N_10448);
nand U12693 (N_12693,N_11030,N_11535);
or U12694 (N_12694,N_9333,N_11774);
nor U12695 (N_12695,N_11073,N_11560);
or U12696 (N_12696,N_10024,N_9791);
xor U12697 (N_12697,N_9188,N_10847);
or U12698 (N_12698,N_10601,N_10458);
or U12699 (N_12699,N_11579,N_11531);
nor U12700 (N_12700,N_10961,N_11349);
nor U12701 (N_12701,N_10947,N_10838);
nand U12702 (N_12702,N_11862,N_11779);
and U12703 (N_12703,N_11351,N_9865);
or U12704 (N_12704,N_11971,N_10303);
nand U12705 (N_12705,N_11289,N_10396);
nand U12706 (N_12706,N_9748,N_10386);
and U12707 (N_12707,N_9119,N_10815);
and U12708 (N_12708,N_10158,N_10220);
nor U12709 (N_12709,N_11590,N_9837);
or U12710 (N_12710,N_9302,N_9956);
and U12711 (N_12711,N_11227,N_9861);
and U12712 (N_12712,N_9077,N_10367);
or U12713 (N_12713,N_10858,N_11847);
or U12714 (N_12714,N_11761,N_10172);
nand U12715 (N_12715,N_11479,N_9168);
nor U12716 (N_12716,N_11390,N_9659);
nor U12717 (N_12717,N_11224,N_11893);
or U12718 (N_12718,N_10765,N_9772);
or U12719 (N_12719,N_11303,N_10306);
nor U12720 (N_12720,N_10874,N_9248);
nand U12721 (N_12721,N_9228,N_9568);
xnor U12722 (N_12722,N_11676,N_9325);
and U12723 (N_12723,N_9278,N_10032);
nand U12724 (N_12724,N_11230,N_10613);
and U12725 (N_12725,N_10794,N_11840);
nor U12726 (N_12726,N_11103,N_9590);
xor U12727 (N_12727,N_9358,N_11363);
or U12728 (N_12728,N_11605,N_11679);
nand U12729 (N_12729,N_9788,N_9773);
xor U12730 (N_12730,N_11998,N_10499);
nor U12731 (N_12731,N_10033,N_9315);
nor U12732 (N_12732,N_9112,N_11917);
xnor U12733 (N_12733,N_11569,N_9944);
or U12734 (N_12734,N_9337,N_9812);
and U12735 (N_12735,N_9100,N_9216);
and U12736 (N_12736,N_10264,N_10972);
nor U12737 (N_12737,N_9422,N_9200);
nand U12738 (N_12738,N_9869,N_10648);
and U12739 (N_12739,N_11733,N_11122);
nand U12740 (N_12740,N_10439,N_10480);
or U12741 (N_12741,N_11306,N_9924);
nand U12742 (N_12742,N_9417,N_9745);
nand U12743 (N_12743,N_9962,N_10497);
and U12744 (N_12744,N_10051,N_9053);
or U12745 (N_12745,N_11473,N_11395);
or U12746 (N_12746,N_11581,N_11155);
nand U12747 (N_12747,N_9359,N_9221);
nor U12748 (N_12748,N_11564,N_9449);
or U12749 (N_12749,N_10694,N_10179);
nor U12750 (N_12750,N_11121,N_11240);
or U12751 (N_12751,N_9378,N_9752);
nand U12752 (N_12752,N_9106,N_9635);
and U12753 (N_12753,N_10537,N_10477);
or U12754 (N_12754,N_11146,N_9471);
and U12755 (N_12755,N_9790,N_9965);
nand U12756 (N_12756,N_10217,N_9334);
nor U12757 (N_12757,N_9854,N_9094);
nand U12758 (N_12758,N_10704,N_11837);
nand U12759 (N_12759,N_11457,N_11545);
nor U12760 (N_12760,N_9349,N_9391);
nor U12761 (N_12761,N_11461,N_11269);
or U12762 (N_12762,N_11570,N_10891);
or U12763 (N_12763,N_10153,N_11004);
or U12764 (N_12764,N_11818,N_11012);
nand U12765 (N_12765,N_10963,N_10801);
or U12766 (N_12766,N_10420,N_10945);
nor U12767 (N_12767,N_10440,N_11911);
nor U12768 (N_12768,N_10251,N_10186);
nor U12769 (N_12769,N_9759,N_9385);
and U12770 (N_12770,N_9742,N_9398);
nand U12771 (N_12771,N_10640,N_9092);
and U12772 (N_12772,N_11659,N_10685);
nor U12773 (N_12773,N_11854,N_9554);
and U12774 (N_12774,N_9599,N_10669);
and U12775 (N_12775,N_10290,N_10839);
nor U12776 (N_12776,N_10942,N_10791);
nor U12777 (N_12777,N_11279,N_10350);
and U12778 (N_12778,N_9332,N_10482);
nor U12779 (N_12779,N_11752,N_10115);
nand U12780 (N_12780,N_10256,N_9784);
nor U12781 (N_12781,N_11144,N_11292);
or U12782 (N_12782,N_10421,N_9436);
and U12783 (N_12783,N_10210,N_11673);
nor U12784 (N_12784,N_10302,N_9448);
or U12785 (N_12785,N_11553,N_10456);
or U12786 (N_12786,N_10725,N_11236);
nor U12787 (N_12787,N_11281,N_9336);
nand U12788 (N_12788,N_10860,N_9903);
or U12789 (N_12789,N_11597,N_9104);
nand U12790 (N_12790,N_11682,N_9468);
and U12791 (N_12791,N_11313,N_11328);
or U12792 (N_12792,N_9948,N_9057);
xor U12793 (N_12793,N_11551,N_10336);
nand U12794 (N_12794,N_9986,N_10522);
nand U12795 (N_12795,N_10923,N_10100);
or U12796 (N_12796,N_10168,N_11066);
or U12797 (N_12797,N_11857,N_11083);
and U12798 (N_12798,N_9539,N_11575);
nor U12799 (N_12799,N_10875,N_11182);
nor U12800 (N_12800,N_10387,N_9387);
and U12801 (N_12801,N_10061,N_11712);
nand U12802 (N_12802,N_9608,N_9238);
and U12803 (N_12803,N_10461,N_10614);
nand U12804 (N_12804,N_10405,N_11487);
nand U12805 (N_12805,N_10354,N_10844);
or U12806 (N_12806,N_9650,N_11392);
or U12807 (N_12807,N_11604,N_10633);
nor U12808 (N_12808,N_11128,N_10593);
nand U12809 (N_12809,N_9497,N_9461);
or U12810 (N_12810,N_9240,N_10277);
nand U12811 (N_12811,N_9007,N_10174);
or U12812 (N_12812,N_11033,N_9147);
nor U12813 (N_12813,N_11401,N_10735);
nand U12814 (N_12814,N_11612,N_9256);
nand U12815 (N_12815,N_9078,N_9665);
and U12816 (N_12816,N_10446,N_10038);
xor U12817 (N_12817,N_10005,N_9963);
or U12818 (N_12818,N_10353,N_9206);
nand U12819 (N_12819,N_9908,N_9941);
or U12820 (N_12820,N_9410,N_11238);
nor U12821 (N_12821,N_9370,N_10730);
and U12822 (N_12822,N_10003,N_9093);
or U12823 (N_12823,N_10298,N_10652);
and U12824 (N_12824,N_10195,N_10714);
nor U12825 (N_12825,N_11717,N_11518);
xor U12826 (N_12826,N_10543,N_9797);
or U12827 (N_12827,N_9097,N_9056);
nor U12828 (N_12828,N_9612,N_11558);
nand U12829 (N_12829,N_10097,N_9032);
nor U12830 (N_12830,N_10304,N_11563);
or U12831 (N_12831,N_10273,N_9480);
and U12832 (N_12832,N_10742,N_9022);
and U12833 (N_12833,N_9560,N_11647);
nand U12834 (N_12834,N_10907,N_9175);
nor U12835 (N_12835,N_9866,N_10366);
xor U12836 (N_12836,N_11568,N_10635);
or U12837 (N_12837,N_11500,N_9714);
xor U12838 (N_12838,N_11915,N_11910);
nor U12839 (N_12839,N_11372,N_11814);
and U12840 (N_12840,N_9428,N_10059);
or U12841 (N_12841,N_10000,N_10236);
nor U12842 (N_12842,N_10549,N_9966);
nor U12843 (N_12843,N_9922,N_11770);
and U12844 (N_12844,N_10478,N_9732);
nor U12845 (N_12845,N_10466,N_11912);
nand U12846 (N_12846,N_9045,N_11956);
or U12847 (N_12847,N_9805,N_9460);
nor U12848 (N_12848,N_11409,N_11137);
or U12849 (N_12849,N_11449,N_11681);
and U12850 (N_12850,N_10085,N_9645);
or U12851 (N_12851,N_9102,N_11435);
nand U12852 (N_12852,N_9415,N_11094);
nand U12853 (N_12853,N_9317,N_9049);
nand U12854 (N_12854,N_11595,N_9649);
and U12855 (N_12855,N_10848,N_9756);
or U12856 (N_12856,N_9151,N_9441);
or U12857 (N_12857,N_9357,N_11280);
xnor U12858 (N_12858,N_10226,N_10450);
or U12859 (N_12859,N_9250,N_9832);
xnor U12860 (N_12860,N_11643,N_10346);
or U12861 (N_12861,N_11081,N_11199);
nand U12862 (N_12862,N_11548,N_10756);
nand U12863 (N_12863,N_9618,N_11001);
nor U12864 (N_12864,N_9591,N_9721);
and U12865 (N_12865,N_9890,N_11838);
xor U12866 (N_12866,N_10471,N_11225);
xor U12867 (N_12867,N_9916,N_10075);
or U12868 (N_12868,N_11453,N_11788);
and U12869 (N_12869,N_10113,N_10968);
nor U12870 (N_12870,N_11580,N_11080);
and U12871 (N_12871,N_11694,N_10019);
nand U12872 (N_12872,N_11653,N_10501);
xnor U12873 (N_12873,N_10201,N_9985);
xor U12874 (N_12874,N_9386,N_11935);
nor U12875 (N_12875,N_10989,N_10818);
and U12876 (N_12876,N_10677,N_11212);
xor U12877 (N_12877,N_10599,N_11089);
or U12878 (N_12878,N_11177,N_9540);
xor U12879 (N_12879,N_11257,N_11797);
or U12880 (N_12880,N_9136,N_11340);
and U12881 (N_12881,N_9892,N_11241);
and U12882 (N_12882,N_10856,N_10795);
or U12883 (N_12883,N_10863,N_9294);
or U12884 (N_12884,N_10312,N_11432);
and U12885 (N_12885,N_11393,N_11946);
or U12886 (N_12886,N_9913,N_10542);
nor U12887 (N_12887,N_11588,N_10516);
nand U12888 (N_12888,N_11586,N_9297);
nor U12889 (N_12889,N_11431,N_11591);
nor U12890 (N_12890,N_9727,N_9741);
nor U12891 (N_12891,N_11663,N_11964);
nand U12892 (N_12892,N_9648,N_9934);
or U12893 (N_12893,N_10814,N_10017);
xor U12894 (N_12894,N_10188,N_11735);
and U12895 (N_12895,N_10804,N_11621);
nand U12896 (N_12896,N_10211,N_11684);
or U12897 (N_12897,N_10639,N_10779);
or U12898 (N_12898,N_11830,N_10352);
and U12899 (N_12899,N_9804,N_11896);
nand U12900 (N_12900,N_11660,N_10493);
xnor U12901 (N_12901,N_11085,N_11934);
xor U12902 (N_12902,N_10531,N_9826);
or U12903 (N_12903,N_10141,N_9976);
nand U12904 (N_12904,N_9230,N_9118);
nand U12905 (N_12905,N_9273,N_10057);
nand U12906 (N_12906,N_10647,N_11902);
or U12907 (N_12907,N_10358,N_9330);
nor U12908 (N_12908,N_10634,N_10590);
nand U12909 (N_12909,N_9298,N_10736);
or U12910 (N_12910,N_11722,N_11484);
nand U12911 (N_12911,N_11202,N_9316);
nor U12912 (N_12912,N_10813,N_11899);
nor U12913 (N_12913,N_11695,N_11732);
or U12914 (N_12914,N_11943,N_11608);
nor U12915 (N_12915,N_10301,N_9027);
or U12916 (N_12916,N_11493,N_11898);
nor U12917 (N_12917,N_10658,N_9160);
xor U12918 (N_12918,N_9018,N_11941);
nor U12919 (N_12919,N_10232,N_11544);
nand U12920 (N_12920,N_10584,N_11428);
and U12921 (N_12921,N_11789,N_10551);
and U12922 (N_12922,N_11006,N_9793);
xor U12923 (N_12923,N_11642,N_10183);
xor U12924 (N_12924,N_11980,N_9594);
and U12925 (N_12925,N_10042,N_11055);
or U12926 (N_12926,N_9516,N_9851);
nor U12927 (N_12927,N_9277,N_9244);
or U12928 (N_12928,N_9787,N_10859);
or U12929 (N_12929,N_11958,N_10861);
xnor U12930 (N_12930,N_10595,N_10552);
xor U12931 (N_12931,N_11860,N_10533);
nor U12932 (N_12932,N_11715,N_9574);
xnor U12933 (N_12933,N_11999,N_9154);
nor U12934 (N_12934,N_9418,N_10072);
nor U12935 (N_12935,N_10740,N_10975);
and U12936 (N_12936,N_10132,N_9354);
nand U12937 (N_12937,N_11632,N_11783);
nand U12938 (N_12938,N_11875,N_11192);
or U12939 (N_12939,N_11836,N_9939);
nor U12940 (N_12940,N_10641,N_11326);
nor U12941 (N_12941,N_11852,N_9921);
nand U12942 (N_12942,N_10706,N_10228);
nand U12943 (N_12943,N_11208,N_10526);
nor U12944 (N_12944,N_11807,N_10940);
or U12945 (N_12945,N_11298,N_11913);
nand U12946 (N_12946,N_11669,N_9988);
and U12947 (N_12947,N_10070,N_10993);
nand U12948 (N_12948,N_9307,N_11399);
or U12949 (N_12949,N_11504,N_11210);
nor U12950 (N_12950,N_11288,N_10523);
nand U12951 (N_12951,N_11550,N_11441);
or U12952 (N_12952,N_10050,N_9342);
or U12953 (N_12953,N_10846,N_10389);
and U12954 (N_12954,N_9990,N_11156);
or U12955 (N_12955,N_10774,N_9328);
xor U12956 (N_12956,N_9073,N_10136);
xnor U12957 (N_12957,N_11645,N_11201);
nor U12958 (N_12958,N_11932,N_10444);
nor U12959 (N_12959,N_11729,N_10924);
xor U12960 (N_12960,N_10777,N_9456);
xor U12961 (N_12961,N_11855,N_9872);
or U12962 (N_12962,N_11331,N_10365);
nor U12963 (N_12963,N_9144,N_9020);
or U12964 (N_12964,N_10469,N_9489);
nor U12965 (N_12965,N_11338,N_11501);
or U12966 (N_12966,N_11598,N_9474);
and U12967 (N_12967,N_9488,N_11304);
xnor U12968 (N_12968,N_10833,N_10259);
and U12969 (N_12969,N_9155,N_11577);
nor U12970 (N_12970,N_9030,N_11895);
nand U12971 (N_12971,N_11270,N_9222);
nor U12972 (N_12972,N_9614,N_11927);
and U12973 (N_12973,N_9810,N_9512);
and U12974 (N_12974,N_11123,N_10780);
nand U12975 (N_12975,N_9771,N_11138);
and U12976 (N_12976,N_11670,N_9351);
nand U12977 (N_12977,N_11646,N_9268);
nor U12978 (N_12978,N_10095,N_10208);
or U12979 (N_12979,N_11742,N_9407);
nor U12980 (N_12980,N_10581,N_9432);
or U12981 (N_12981,N_9794,N_11603);
nor U12982 (N_12982,N_9224,N_9000);
and U12983 (N_12983,N_9822,N_11808);
and U12984 (N_12984,N_11418,N_11890);
nor U12985 (N_12985,N_11060,N_9857);
or U12986 (N_12986,N_10920,N_9870);
or U12987 (N_12987,N_9821,N_10628);
nor U12988 (N_12988,N_9035,N_10681);
nand U12989 (N_12989,N_10528,N_11342);
and U12990 (N_12990,N_9816,N_9341);
nand U12991 (N_12991,N_9799,N_10427);
nor U12992 (N_12992,N_10144,N_9403);
and U12993 (N_12993,N_11293,N_11773);
nor U12994 (N_12994,N_9640,N_9249);
and U12995 (N_12995,N_10338,N_11737);
and U12996 (N_12996,N_10698,N_10133);
nor U12997 (N_12997,N_10932,N_10241);
nand U12998 (N_12998,N_10407,N_10901);
and U12999 (N_12999,N_10034,N_11992);
or U13000 (N_13000,N_10490,N_10707);
and U13001 (N_13001,N_11654,N_9798);
and U13002 (N_13002,N_9849,N_10282);
and U13003 (N_13003,N_9567,N_9274);
and U13004 (N_13004,N_11526,N_9420);
or U13005 (N_13005,N_9535,N_11914);
nor U13006 (N_13006,N_9642,N_11332);
nor U13007 (N_13007,N_9399,N_10746);
xor U13008 (N_13008,N_11677,N_10684);
nor U13009 (N_13009,N_9641,N_10254);
and U13010 (N_13010,N_9371,N_9687);
nor U13011 (N_13011,N_9598,N_11050);
nor U13012 (N_13012,N_9242,N_11423);
nand U13013 (N_13013,N_9825,N_11164);
or U13014 (N_13014,N_9137,N_10849);
nand U13015 (N_13015,N_9113,N_9843);
nor U13016 (N_13016,N_10128,N_11792);
nand U13017 (N_13017,N_11947,N_11127);
nor U13018 (N_13018,N_9802,N_11832);
and U13019 (N_13019,N_9345,N_10137);
or U13020 (N_13020,N_11072,N_9309);
or U13021 (N_13021,N_9143,N_10906);
nand U13022 (N_13022,N_9338,N_9538);
nor U13023 (N_13023,N_10910,N_10372);
and U13024 (N_13024,N_9008,N_10983);
nor U13025 (N_13025,N_11803,N_10160);
nand U13026 (N_13026,N_11848,N_10322);
nand U13027 (N_13027,N_9347,N_9989);
nand U13028 (N_13028,N_11319,N_9577);
nor U13029 (N_13029,N_9735,N_9585);
and U13030 (N_13030,N_11044,N_9855);
or U13031 (N_13031,N_10384,N_11371);
nand U13032 (N_13032,N_11497,N_10415);
and U13033 (N_13033,N_10148,N_9688);
and U13034 (N_13034,N_10797,N_10289);
xnor U13035 (N_13035,N_9061,N_9920);
nor U13036 (N_13036,N_9896,N_10883);
or U13037 (N_13037,N_11680,N_9886);
nand U13038 (N_13038,N_10519,N_10430);
or U13039 (N_13039,N_9308,N_11463);
nor U13040 (N_13040,N_9764,N_9120);
nor U13041 (N_13041,N_10955,N_10392);
xnor U13042 (N_13042,N_9287,N_9815);
and U13043 (N_13043,N_10332,N_10811);
nor U13044 (N_13044,N_9884,N_11148);
nand U13045 (N_13045,N_11930,N_9047);
or U13046 (N_13046,N_11003,N_11541);
and U13047 (N_13047,N_11011,N_10769);
or U13048 (N_13048,N_11067,N_10729);
nor U13049 (N_13049,N_10842,N_9095);
nand U13050 (N_13050,N_11214,N_11350);
nand U13051 (N_13051,N_11989,N_10712);
nand U13052 (N_13052,N_9637,N_10475);
or U13053 (N_13053,N_11075,N_10145);
and U13054 (N_13054,N_11689,N_11325);
or U13055 (N_13055,N_11955,N_10823);
nand U13056 (N_13056,N_9838,N_9807);
nand U13057 (N_13057,N_9666,N_10636);
nand U13058 (N_13058,N_11165,N_9753);
nand U13059 (N_13059,N_10820,N_10468);
xor U13060 (N_13060,N_11734,N_9663);
nor U13061 (N_13061,N_11979,N_10699);
nand U13062 (N_13062,N_11638,N_11957);
nand U13063 (N_13063,N_10570,N_11198);
nor U13064 (N_13064,N_10198,N_9831);
or U13065 (N_13065,N_11687,N_11249);
or U13066 (N_13066,N_11522,N_11300);
xor U13067 (N_13067,N_9623,N_10170);
or U13068 (N_13068,N_10627,N_10525);
nand U13069 (N_13069,N_10722,N_9475);
and U13070 (N_13070,N_10991,N_10035);
nand U13071 (N_13071,N_10978,N_11540);
nand U13072 (N_13072,N_11983,N_11606);
and U13073 (N_13073,N_11565,N_11759);
nand U13074 (N_13074,N_10110,N_9023);
xnor U13075 (N_13075,N_9083,N_11344);
nor U13076 (N_13076,N_10442,N_9042);
or U13077 (N_13077,N_9647,N_10946);
and U13078 (N_13078,N_10143,N_10618);
and U13079 (N_13079,N_10548,N_10887);
nor U13080 (N_13080,N_10931,N_11871);
nor U13081 (N_13081,N_10536,N_9677);
nand U13082 (N_13082,N_11630,N_9050);
nor U13083 (N_13083,N_10710,N_9424);
and U13084 (N_13084,N_9129,N_9498);
xnor U13085 (N_13085,N_10280,N_9183);
or U13086 (N_13086,N_9431,N_10967);
or U13087 (N_13087,N_9290,N_11833);
or U13088 (N_13088,N_10546,N_10357);
nor U13089 (N_13089,N_10109,N_9466);
and U13090 (N_13090,N_11427,N_9394);
nand U13091 (N_13091,N_9867,N_11954);
xnor U13092 (N_13092,N_11120,N_11226);
nand U13093 (N_13093,N_9532,N_11562);
or U13094 (N_13094,N_9952,N_9958);
and U13095 (N_13095,N_11158,N_11299);
nor U13096 (N_13096,N_10899,N_10917);
nor U13097 (N_13097,N_9537,N_10610);
or U13098 (N_13098,N_10679,N_9509);
nor U13099 (N_13099,N_11318,N_9243);
nor U13100 (N_13100,N_10503,N_9750);
nor U13101 (N_13101,N_11367,N_11547);
and U13102 (N_13102,N_10252,N_11255);
and U13103 (N_13103,N_11511,N_10134);
or U13104 (N_13104,N_11256,N_9364);
and U13105 (N_13105,N_9186,N_10741);
nor U13106 (N_13106,N_9397,N_9817);
and U13107 (N_13107,N_11521,N_10344);
and U13108 (N_13108,N_10295,N_10755);
xnor U13109 (N_13109,N_10261,N_9457);
xnor U13110 (N_13110,N_10485,N_9833);
xnor U13111 (N_13111,N_10315,N_9545);
and U13112 (N_13112,N_11709,N_11515);
nand U13113 (N_13113,N_10031,N_11892);
and U13114 (N_13114,N_10733,N_11953);
or U13115 (N_13115,N_9075,N_9521);
nand U13116 (N_13116,N_10083,N_10218);
and U13117 (N_13117,N_11439,N_11945);
and U13118 (N_13118,N_10328,N_9726);
or U13119 (N_13119,N_10643,N_11267);
or U13120 (N_13120,N_11872,N_10954);
xor U13121 (N_13121,N_10821,N_10865);
nor U13122 (N_13122,N_11725,N_9266);
nand U13123 (N_13123,N_9344,N_9969);
or U13124 (N_13124,N_9280,N_9840);
or U13125 (N_13125,N_9972,N_10288);
or U13126 (N_13126,N_9180,N_11061);
nand U13127 (N_13127,N_10749,N_10535);
and U13128 (N_13128,N_9135,N_10693);
and U13129 (N_13129,N_11106,N_9063);
nand U13130 (N_13130,N_11781,N_11218);
nor U13131 (N_13131,N_11451,N_10911);
and U13132 (N_13132,N_9868,N_10079);
and U13133 (N_13133,N_9994,N_11185);
nand U13134 (N_13134,N_11876,N_9066);
or U13135 (N_13135,N_9079,N_10720);
nand U13136 (N_13136,N_11593,N_9761);
nor U13137 (N_13137,N_11764,N_9923);
and U13138 (N_13138,N_10753,N_11402);
or U13139 (N_13139,N_9534,N_9286);
nor U13140 (N_13140,N_10933,N_9459);
or U13141 (N_13141,N_11546,N_9152);
xnor U13142 (N_13142,N_11567,N_9904);
or U13143 (N_13143,N_11885,N_10184);
or U13144 (N_13144,N_9159,N_10689);
nand U13145 (N_13145,N_9473,N_10951);
nor U13146 (N_13146,N_9716,N_10534);
and U13147 (N_13147,N_11538,N_9289);
xor U13148 (N_13148,N_9557,N_10623);
and U13149 (N_13149,N_10949,N_11713);
and U13150 (N_13150,N_10510,N_9182);
nand U13151 (N_13151,N_10676,N_10575);
or U13152 (N_13152,N_10878,N_10425);
or U13153 (N_13153,N_9651,N_10959);
or U13154 (N_13154,N_10857,N_10656);
nand U13155 (N_13155,N_11478,N_10638);
nand U13156 (N_13156,N_9646,N_10018);
or U13157 (N_13157,N_9463,N_10877);
or U13158 (N_13158,N_11271,N_9062);
nor U13159 (N_13159,N_11102,N_10474);
and U13160 (N_13160,N_9215,N_11414);
or U13161 (N_13161,N_10696,N_9803);
nand U13162 (N_13162,N_9084,N_9811);
nor U13163 (N_13163,N_11780,N_9675);
nand U13164 (N_13164,N_10135,N_10077);
or U13165 (N_13165,N_11994,N_11095);
xor U13166 (N_13166,N_11960,N_10333);
or U13167 (N_13167,N_9353,N_10836);
nand U13168 (N_13168,N_10250,N_10375);
nand U13169 (N_13169,N_10553,N_11858);
nor U13170 (N_13170,N_10494,N_9269);
or U13171 (N_13171,N_9579,N_10369);
xnor U13172 (N_13172,N_11091,N_11264);
or U13173 (N_13173,N_10023,N_10481);
and U13174 (N_13174,N_10980,N_9800);
nor U13175 (N_13175,N_11826,N_9702);
nor U13176 (N_13176,N_10257,N_9486);
nand U13177 (N_13177,N_10316,N_10429);
nor U13178 (N_13178,N_9919,N_11539);
nor U13179 (N_13179,N_11617,N_9149);
or U13180 (N_13180,N_9170,N_10398);
xnor U13181 (N_13181,N_9502,N_11386);
nand U13182 (N_13182,N_9292,N_11793);
nand U13183 (N_13183,N_10159,N_11110);
nor U13184 (N_13184,N_10383,N_11168);
nand U13185 (N_13185,N_9705,N_10631);
nor U13186 (N_13186,N_11683,N_10998);
nand U13187 (N_13187,N_11756,N_11607);
xnor U13188 (N_13188,N_11087,N_10457);
and U13189 (N_13189,N_11475,N_9380);
nor U13190 (N_13190,N_11510,N_9524);
and U13191 (N_13191,N_9122,N_10758);
nand U13192 (N_13192,N_11667,N_9411);
and U13193 (N_13193,N_9553,N_11160);
and U13194 (N_13194,N_9970,N_11942);
or U13195 (N_13195,N_10399,N_9501);
nand U13196 (N_13196,N_9162,N_11800);
and U13197 (N_13197,N_11181,N_10556);
nor U13198 (N_13198,N_11222,N_11869);
and U13199 (N_13199,N_9774,N_11656);
or U13200 (N_13200,N_10670,N_9792);
nand U13201 (N_13201,N_10960,N_10414);
or U13202 (N_13202,N_9131,N_10453);
or U13203 (N_13203,N_10452,N_9116);
or U13204 (N_13204,N_9895,N_10313);
and U13205 (N_13205,N_11458,N_10401);
or U13206 (N_13206,N_11320,N_11097);
or U13207 (N_13207,N_11505,N_10417);
nor U13208 (N_13208,N_11398,N_10817);
or U13209 (N_13209,N_11778,N_9107);
or U13210 (N_13210,N_11961,N_11620);
xor U13211 (N_13211,N_9769,N_10297);
or U13212 (N_13212,N_9464,N_9482);
or U13213 (N_13213,N_11426,N_9296);
and U13214 (N_13214,N_9312,N_9484);
xor U13215 (N_13215,N_9219,N_10476);
nand U13216 (N_13216,N_11239,N_11169);
nand U13217 (N_13217,N_11688,N_11284);
or U13218 (N_13218,N_9711,N_9653);
or U13219 (N_13219,N_10690,N_10056);
and U13220 (N_13220,N_9472,N_10727);
and U13221 (N_13221,N_10435,N_11743);
or U13222 (N_13222,N_10566,N_11884);
nand U13223 (N_13223,N_11490,N_11486);
or U13224 (N_13224,N_10586,N_11573);
or U13225 (N_13225,N_9043,N_10793);
nand U13226 (N_13226,N_11760,N_10919);
and U13227 (N_13227,N_11969,N_10305);
nor U13228 (N_13228,N_10377,N_11116);
nand U13229 (N_13229,N_9295,N_9933);
xnor U13230 (N_13230,N_11308,N_9583);
nor U13231 (N_13231,N_11361,N_9382);
or U13232 (N_13232,N_10854,N_11464);
nor U13233 (N_13233,N_11357,N_9980);
and U13234 (N_13234,N_9809,N_11276);
and U13235 (N_13235,N_10347,N_9531);
nor U13236 (N_13236,N_10900,N_11524);
nor U13237 (N_13237,N_10037,N_10225);
nand U13238 (N_13238,N_11691,N_10888);
and U13239 (N_13239,N_9757,N_10879);
xnor U13240 (N_13240,N_11157,N_10822);
nor U13241 (N_13241,N_10751,N_10988);
nand U13242 (N_13242,N_10496,N_9754);
xor U13243 (N_13243,N_9930,N_9636);
nand U13244 (N_13244,N_9906,N_9885);
nor U13245 (N_13245,N_11196,N_9082);
or U13246 (N_13246,N_11652,N_9679);
nand U13247 (N_13247,N_9496,N_11576);
nor U13248 (N_13248,N_11064,N_9573);
nor U13249 (N_13249,N_11378,N_9169);
and U13250 (N_13250,N_11525,N_11919);
or U13251 (N_13251,N_10187,N_9673);
or U13252 (N_13252,N_9657,N_10563);
and U13253 (N_13253,N_11704,N_10688);
nor U13254 (N_13254,N_9110,N_11068);
or U13255 (N_13255,N_9413,N_11492);
nor U13256 (N_13256,N_9707,N_11077);
and U13257 (N_13257,N_9871,N_11516);
nand U13258 (N_13258,N_10521,N_11305);
nor U13259 (N_13259,N_10588,N_11035);
or U13260 (N_13260,N_9462,N_9740);
nand U13261 (N_13261,N_10509,N_10803);
nand U13262 (N_13262,N_10169,N_9600);
nor U13263 (N_13263,N_10953,N_9967);
nand U13264 (N_13264,N_9715,N_9563);
nor U13265 (N_13265,N_11724,N_10787);
and U13266 (N_13266,N_10314,N_9161);
or U13267 (N_13267,N_9167,N_10843);
nand U13268 (N_13268,N_9146,N_9442);
and U13269 (N_13269,N_9981,N_10948);
nand U13270 (N_13270,N_11828,N_9619);
and U13271 (N_13271,N_9270,N_11705);
nor U13272 (N_13272,N_9701,N_11062);
xor U13273 (N_13273,N_10340,N_11352);
or U13274 (N_13274,N_9522,N_9187);
nor U13275 (N_13275,N_10380,N_9517);
and U13276 (N_13276,N_11412,N_11017);
nor U13277 (N_13277,N_11599,N_10240);
or U13278 (N_13278,N_9048,N_11407);
or U13279 (N_13279,N_10036,N_11084);
or U13280 (N_13280,N_11757,N_10185);
or U13281 (N_13281,N_10558,N_9654);
and U13282 (N_13282,N_10166,N_11842);
nand U13283 (N_13283,N_11189,N_10199);
xnor U13284 (N_13284,N_10020,N_11582);
nor U13285 (N_13285,N_11310,N_10447);
or U13286 (N_13286,N_11437,N_11796);
xnor U13287 (N_13287,N_10323,N_9530);
or U13288 (N_13288,N_11315,N_9218);
nand U13289 (N_13289,N_11117,N_9947);
or U13290 (N_13290,N_9220,N_9940);
xnor U13291 (N_13291,N_11859,N_10650);
and U13292 (N_13292,N_10165,N_9414);
and U13293 (N_13293,N_11745,N_11990);
nand U13294 (N_13294,N_11375,N_11042);
or U13295 (N_13295,N_11018,N_9581);
or U13296 (N_13296,N_10752,N_9177);
nand U13297 (N_13297,N_11353,N_9876);
and U13298 (N_13298,N_10990,N_9997);
xor U13299 (N_13299,N_11991,N_10645);
or U13300 (N_13300,N_9982,N_9455);
nand U13301 (N_13301,N_10555,N_9847);
nand U13302 (N_13302,N_9827,N_10986);
nand U13303 (N_13303,N_11220,N_10868);
nor U13304 (N_13304,N_10577,N_10027);
or U13305 (N_13305,N_11179,N_11948);
or U13306 (N_13306,N_10483,N_10419);
or U13307 (N_13307,N_11400,N_9975);
nand U13308 (N_13308,N_10665,N_9233);
or U13309 (N_13309,N_9528,N_10267);
and U13310 (N_13310,N_11200,N_9381);
nand U13311 (N_13311,N_10894,N_11105);
xor U13312 (N_13312,N_11149,N_11397);
or U13313 (N_13313,N_10808,N_11228);
and U13314 (N_13314,N_11923,N_11377);
xnor U13315 (N_13315,N_11114,N_9596);
and U13316 (N_13316,N_10969,N_9105);
xor U13317 (N_13317,N_9140,N_11708);
nand U13318 (N_13318,N_10320,N_10325);
or U13319 (N_13319,N_9366,N_11767);
and U13320 (N_13320,N_9550,N_10238);
nand U13321 (N_13321,N_10761,N_11176);
xnor U13322 (N_13322,N_9877,N_10909);
nor U13323 (N_13323,N_10675,N_11758);
and U13324 (N_13324,N_10368,N_11171);
xnor U13325 (N_13325,N_11283,N_11311);
nand U13326 (N_13326,N_10835,N_9125);
xor U13327 (N_13327,N_9505,N_9142);
or U13328 (N_13328,N_10663,N_11448);
nand U13329 (N_13329,N_9504,N_10646);
or U13330 (N_13330,N_11822,N_11104);
or U13331 (N_13331,N_11502,N_11321);
or U13332 (N_13332,N_10719,N_10941);
nand U13333 (N_13333,N_11039,N_10180);
and U13334 (N_13334,N_11259,N_10757);
or U13335 (N_13335,N_9692,N_11235);
or U13336 (N_13336,N_10402,N_11219);
nand U13337 (N_13337,N_10962,N_9652);
nor U13338 (N_13338,N_9766,N_9335);
nor U13339 (N_13339,N_11984,N_10504);
or U13340 (N_13340,N_10629,N_10926);
or U13341 (N_13341,N_9133,N_9945);
xor U13342 (N_13342,N_11918,N_10438);
nor U13343 (N_13343,N_10869,N_11791);
or U13344 (N_13344,N_11088,N_9862);
or U13345 (N_13345,N_11082,N_10903);
nor U13346 (N_13346,N_9634,N_11460);
and U13347 (N_13347,N_9348,N_9178);
nor U13348 (N_13348,N_11846,N_10276);
nand U13349 (N_13349,N_11700,N_10125);
nor U13350 (N_13350,N_9321,N_9343);
nor U13351 (N_13351,N_9476,N_10105);
nor U13352 (N_13352,N_11561,N_11408);
xor U13353 (N_13353,N_10112,N_11810);
nand U13354 (N_13354,N_9580,N_11636);
and U13355 (N_13355,N_11099,N_9060);
and U13356 (N_13356,N_9301,N_9038);
and U13357 (N_13357,N_10173,N_10044);
xor U13358 (N_13358,N_10682,N_9011);
and U13359 (N_13359,N_11037,N_11883);
nand U13360 (N_13360,N_10082,N_9882);
and U13361 (N_13361,N_11347,N_10673);
xnor U13362 (N_13362,N_9520,N_11787);
nand U13363 (N_13363,N_9546,N_9656);
or U13364 (N_13364,N_10451,N_11503);
nor U13365 (N_13365,N_10362,N_11853);
and U13366 (N_13366,N_11763,N_9435);
nor U13367 (N_13367,N_11242,N_9639);
nand U13368 (N_13368,N_11142,N_11231);
and U13369 (N_13369,N_9469,N_11229);
nand U13370 (N_13370,N_11706,N_11096);
nand U13371 (N_13371,N_10007,N_9234);
nor U13372 (N_13372,N_10242,N_10066);
xnor U13373 (N_13373,N_11644,N_11615);
or U13374 (N_13374,N_10731,N_9621);
and U13375 (N_13375,N_10876,N_9724);
or U13376 (N_13376,N_10789,N_11263);
nor U13377 (N_13377,N_11258,N_10263);
nand U13378 (N_13378,N_11627,N_10492);
xnor U13379 (N_13379,N_10260,N_10692);
and U13380 (N_13380,N_9858,N_11184);
or U13381 (N_13381,N_11111,N_11619);
nand U13382 (N_13382,N_10724,N_9893);
nand U13383 (N_13383,N_10016,N_11692);
nor U13384 (N_13384,N_10925,N_9115);
xnor U13385 (N_13385,N_11076,N_11317);
nor U13386 (N_13386,N_9602,N_11205);
or U13387 (N_13387,N_11329,N_9604);
and U13388 (N_13388,N_9900,N_10432);
and U13389 (N_13389,N_11685,N_10728);
nor U13390 (N_13390,N_9367,N_11794);
or U13391 (N_13391,N_9617,N_11252);
nor U13392 (N_13392,N_11382,N_11900);
nand U13393 (N_13393,N_11335,N_9782);
and U13394 (N_13394,N_11614,N_10604);
nand U13395 (N_13395,N_9845,N_10517);
or U13396 (N_13396,N_10799,N_11266);
or U13397 (N_13397,N_9479,N_10667);
or U13398 (N_13398,N_9231,N_9326);
and U13399 (N_13399,N_9630,N_9846);
and U13400 (N_13400,N_10579,N_9891);
nor U13401 (N_13401,N_10472,N_10214);
nor U13402 (N_13402,N_11668,N_10355);
xor U13403 (N_13403,N_9632,N_11657);
nand U13404 (N_13404,N_10589,N_10965);
or U13405 (N_13405,N_10800,N_9427);
and U13406 (N_13406,N_10759,N_11718);
nor U13407 (N_13407,N_10086,N_11882);
xnor U13408 (N_13408,N_11109,N_9141);
and U13409 (N_13409,N_11472,N_9369);
and U13410 (N_13410,N_11730,N_9067);
nor U13411 (N_13411,N_11074,N_11275);
and U13412 (N_13412,N_11415,N_9390);
nor U13413 (N_13413,N_9021,N_10370);
nor U13414 (N_13414,N_9444,N_11908);
xnor U13415 (N_13415,N_10363,N_11360);
or U13416 (N_13416,N_11166,N_11425);
and U13417 (N_13417,N_11543,N_11139);
and U13418 (N_13418,N_10206,N_10866);
or U13419 (N_13419,N_11831,N_9703);
or U13420 (N_13420,N_9081,N_9983);
nor U13421 (N_13421,N_11232,N_10539);
or U13422 (N_13422,N_9396,N_11413);
xnor U13423 (N_13423,N_11829,N_9564);
or U13424 (N_13424,N_11938,N_9506);
or U13425 (N_13425,N_10486,N_10223);
nor U13426 (N_13426,N_10002,N_9139);
nor U13427 (N_13427,N_11233,N_9196);
or U13428 (N_13428,N_9195,N_9375);
nand U13429 (N_13429,N_10209,N_11322);
or U13430 (N_13430,N_9363,N_11740);
and U13431 (N_13431,N_10071,N_9072);
nand U13432 (N_13432,N_11141,N_10520);
nor U13433 (N_13433,N_9559,N_9551);
or U13434 (N_13434,N_10335,N_11662);
or U13435 (N_13435,N_10428,N_11071);
nand U13436 (N_13436,N_10608,N_9911);
nand U13437 (N_13437,N_10540,N_11433);
and U13438 (N_13438,N_10927,N_9368);
nand U13439 (N_13439,N_11819,N_11047);
or U13440 (N_13440,N_9426,N_11584);
or U13441 (N_13441,N_10239,N_9437);
nand U13442 (N_13442,N_11261,N_10576);
xnor U13443 (N_13443,N_10564,N_9918);
or U13444 (N_13444,N_9951,N_9644);
nor U13445 (N_13445,N_10834,N_10281);
or U13446 (N_13446,N_9003,N_10356);
and U13447 (N_13447,N_11253,N_10437);
nand U13448 (N_13448,N_10582,N_9189);
nor U13449 (N_13449,N_10977,N_10029);
nand U13450 (N_13450,N_11206,N_9194);
nor U13451 (N_13451,N_9223,N_11459);
nand U13452 (N_13452,N_11631,N_11825);
and U13453 (N_13453,N_10424,N_9181);
xnor U13454 (N_13454,N_11140,N_11405);
nand U13455 (N_13455,N_9734,N_9352);
nor U13456 (N_13456,N_9263,N_10106);
or U13457 (N_13457,N_10683,N_11370);
nor U13458 (N_13458,N_10434,N_9163);
nand U13459 (N_13459,N_10921,N_9373);
and U13460 (N_13460,N_9052,N_11530);
nor U13461 (N_13461,N_10885,N_11624);
nor U13462 (N_13462,N_11057,N_11147);
and U13463 (N_13463,N_11026,N_11162);
or U13464 (N_13464,N_11674,N_9111);
and U13465 (N_13465,N_11153,N_11907);
or U13466 (N_13466,N_9763,N_9860);
nor U13467 (N_13467,N_10081,N_9909);
and U13468 (N_13468,N_9929,N_10311);
and U13469 (N_13469,N_10873,N_10762);
xor U13470 (N_13470,N_9523,N_11324);
nand U13471 (N_13471,N_10783,N_10445);
nand U13472 (N_13472,N_9405,N_10248);
xnor U13473 (N_13473,N_10626,N_9376);
nand U13474 (N_13474,N_10770,N_11959);
and U13475 (N_13475,N_11850,N_11813);
or U13476 (N_13476,N_10441,N_9406);
or U13477 (N_13477,N_9605,N_10672);
or U13478 (N_13478,N_9842,N_10979);
and U13479 (N_13479,N_9145,N_10713);
or U13480 (N_13480,N_10996,N_11132);
or U13481 (N_13481,N_11507,N_10285);
or U13482 (N_13482,N_11136,N_9478);
or U13483 (N_13483,N_10065,N_10896);
and U13484 (N_13484,N_11496,N_9227);
xor U13485 (N_13485,N_9493,N_10664);
and U13486 (N_13486,N_9912,N_9836);
nor U13487 (N_13487,N_10030,N_11339);
nand U13488 (N_13488,N_9796,N_9320);
or U13489 (N_13489,N_11348,N_9830);
nand U13490 (N_13490,N_11366,N_9279);
nor U13491 (N_13491,N_9880,N_11815);
and U13492 (N_13492,N_9064,N_10246);
and U13493 (N_13493,N_11993,N_9907);
or U13494 (N_13494,N_10661,N_10655);
or U13495 (N_13495,N_9235,N_10612);
nand U13496 (N_13496,N_9615,N_9691);
nor U13497 (N_13497,N_9841,N_10530);
and U13498 (N_13498,N_10286,N_9031);
and U13499 (N_13499,N_10265,N_11070);
xnor U13500 (N_13500,N_10261,N_10566);
or U13501 (N_13501,N_11003,N_11931);
nand U13502 (N_13502,N_11225,N_10438);
nand U13503 (N_13503,N_11505,N_11219);
or U13504 (N_13504,N_10261,N_9703);
or U13505 (N_13505,N_11051,N_11795);
or U13506 (N_13506,N_9779,N_9132);
nor U13507 (N_13507,N_11527,N_9602);
nor U13508 (N_13508,N_10009,N_10069);
nand U13509 (N_13509,N_9758,N_9041);
or U13510 (N_13510,N_11584,N_9496);
and U13511 (N_13511,N_11268,N_9305);
nand U13512 (N_13512,N_10436,N_11550);
and U13513 (N_13513,N_10684,N_10922);
or U13514 (N_13514,N_10084,N_11042);
nor U13515 (N_13515,N_9383,N_10535);
or U13516 (N_13516,N_9516,N_11841);
nor U13517 (N_13517,N_9782,N_11780);
and U13518 (N_13518,N_10701,N_11709);
nand U13519 (N_13519,N_11824,N_10729);
nor U13520 (N_13520,N_10147,N_9791);
nor U13521 (N_13521,N_11873,N_11263);
xor U13522 (N_13522,N_10117,N_11170);
nand U13523 (N_13523,N_10059,N_10695);
nand U13524 (N_13524,N_11720,N_11934);
xnor U13525 (N_13525,N_11811,N_9140);
or U13526 (N_13526,N_10368,N_11210);
nand U13527 (N_13527,N_11674,N_11304);
xor U13528 (N_13528,N_10725,N_11784);
nor U13529 (N_13529,N_11339,N_10400);
nand U13530 (N_13530,N_9804,N_11594);
and U13531 (N_13531,N_9061,N_10707);
or U13532 (N_13532,N_9581,N_11758);
and U13533 (N_13533,N_9528,N_10072);
or U13534 (N_13534,N_10065,N_10882);
nor U13535 (N_13535,N_10765,N_10082);
nand U13536 (N_13536,N_9571,N_9489);
xor U13537 (N_13537,N_11269,N_9954);
nand U13538 (N_13538,N_10756,N_11305);
xnor U13539 (N_13539,N_9078,N_11978);
or U13540 (N_13540,N_9944,N_10035);
or U13541 (N_13541,N_9192,N_10039);
or U13542 (N_13542,N_10726,N_11106);
nor U13543 (N_13543,N_11416,N_11500);
or U13544 (N_13544,N_11515,N_9667);
nor U13545 (N_13545,N_9708,N_9408);
and U13546 (N_13546,N_11131,N_11694);
and U13547 (N_13547,N_11274,N_10019);
nand U13548 (N_13548,N_11977,N_9752);
and U13549 (N_13549,N_10204,N_11725);
nor U13550 (N_13550,N_10375,N_11562);
nor U13551 (N_13551,N_9324,N_10489);
nor U13552 (N_13552,N_10504,N_10003);
nor U13553 (N_13553,N_10264,N_10387);
xnor U13554 (N_13554,N_9905,N_10132);
and U13555 (N_13555,N_9194,N_9648);
and U13556 (N_13556,N_11606,N_9845);
and U13557 (N_13557,N_11292,N_9309);
nand U13558 (N_13558,N_9221,N_10437);
and U13559 (N_13559,N_9285,N_9250);
xnor U13560 (N_13560,N_11898,N_9048);
and U13561 (N_13561,N_10965,N_11894);
and U13562 (N_13562,N_10612,N_9072);
or U13563 (N_13563,N_9098,N_11766);
or U13564 (N_13564,N_11001,N_10641);
nand U13565 (N_13565,N_10750,N_10228);
xnor U13566 (N_13566,N_10838,N_9930);
nor U13567 (N_13567,N_9277,N_9190);
or U13568 (N_13568,N_9610,N_9370);
and U13569 (N_13569,N_11973,N_11255);
nor U13570 (N_13570,N_11445,N_9124);
xor U13571 (N_13571,N_11587,N_10325);
or U13572 (N_13572,N_11912,N_11617);
nand U13573 (N_13573,N_11908,N_9334);
nand U13574 (N_13574,N_11678,N_10415);
nand U13575 (N_13575,N_10842,N_11507);
nand U13576 (N_13576,N_10421,N_10722);
nor U13577 (N_13577,N_11297,N_9457);
nor U13578 (N_13578,N_10405,N_10411);
nand U13579 (N_13579,N_11017,N_9003);
or U13580 (N_13580,N_9325,N_10687);
and U13581 (N_13581,N_9401,N_10672);
xor U13582 (N_13582,N_11932,N_11766);
and U13583 (N_13583,N_10419,N_9184);
nor U13584 (N_13584,N_11439,N_10985);
or U13585 (N_13585,N_9584,N_10098);
nand U13586 (N_13586,N_11902,N_10574);
or U13587 (N_13587,N_9208,N_10275);
nor U13588 (N_13588,N_10125,N_9075);
and U13589 (N_13589,N_9043,N_9229);
and U13590 (N_13590,N_11208,N_11236);
nand U13591 (N_13591,N_11590,N_9984);
and U13592 (N_13592,N_10281,N_9103);
or U13593 (N_13593,N_10809,N_9144);
nor U13594 (N_13594,N_11350,N_10847);
nor U13595 (N_13595,N_9618,N_10301);
and U13596 (N_13596,N_9911,N_11419);
nand U13597 (N_13597,N_11004,N_10270);
nand U13598 (N_13598,N_10108,N_9058);
and U13599 (N_13599,N_9649,N_11984);
or U13600 (N_13600,N_11852,N_10513);
nand U13601 (N_13601,N_10887,N_9135);
nor U13602 (N_13602,N_10738,N_9780);
and U13603 (N_13603,N_9273,N_11057);
nand U13604 (N_13604,N_9096,N_10724);
nor U13605 (N_13605,N_9250,N_10986);
and U13606 (N_13606,N_11674,N_10185);
and U13607 (N_13607,N_10122,N_9088);
and U13608 (N_13608,N_10900,N_10663);
nor U13609 (N_13609,N_10351,N_11572);
nor U13610 (N_13610,N_11983,N_11921);
nand U13611 (N_13611,N_9809,N_10026);
nor U13612 (N_13612,N_9836,N_11004);
nand U13613 (N_13613,N_11444,N_10780);
or U13614 (N_13614,N_11194,N_9280);
nor U13615 (N_13615,N_9404,N_10489);
nor U13616 (N_13616,N_10265,N_10220);
and U13617 (N_13617,N_9254,N_9234);
and U13618 (N_13618,N_10353,N_10965);
or U13619 (N_13619,N_10093,N_11442);
xnor U13620 (N_13620,N_11044,N_10333);
nor U13621 (N_13621,N_11201,N_11125);
or U13622 (N_13622,N_9159,N_11294);
or U13623 (N_13623,N_11471,N_11169);
xnor U13624 (N_13624,N_10854,N_9874);
nand U13625 (N_13625,N_11234,N_9260);
or U13626 (N_13626,N_10168,N_11703);
nand U13627 (N_13627,N_10365,N_10393);
xor U13628 (N_13628,N_9362,N_10938);
nand U13629 (N_13629,N_10607,N_11176);
or U13630 (N_13630,N_11712,N_11086);
nor U13631 (N_13631,N_9667,N_10856);
or U13632 (N_13632,N_9924,N_9545);
xor U13633 (N_13633,N_11744,N_11037);
and U13634 (N_13634,N_10352,N_11230);
nand U13635 (N_13635,N_9581,N_9038);
nand U13636 (N_13636,N_10664,N_10248);
nor U13637 (N_13637,N_9114,N_9194);
nor U13638 (N_13638,N_11340,N_11942);
nand U13639 (N_13639,N_11854,N_9738);
and U13640 (N_13640,N_9346,N_11400);
or U13641 (N_13641,N_9657,N_11522);
xnor U13642 (N_13642,N_9974,N_11938);
or U13643 (N_13643,N_11788,N_11670);
and U13644 (N_13644,N_10927,N_10867);
nand U13645 (N_13645,N_9340,N_9271);
or U13646 (N_13646,N_9616,N_11222);
nand U13647 (N_13647,N_10168,N_11099);
or U13648 (N_13648,N_11719,N_11725);
and U13649 (N_13649,N_11317,N_11080);
nand U13650 (N_13650,N_10146,N_11846);
nor U13651 (N_13651,N_10515,N_9202);
and U13652 (N_13652,N_11436,N_11363);
and U13653 (N_13653,N_9611,N_11327);
and U13654 (N_13654,N_10234,N_9042);
nand U13655 (N_13655,N_11484,N_11826);
nor U13656 (N_13656,N_9591,N_9506);
nor U13657 (N_13657,N_10959,N_10080);
and U13658 (N_13658,N_9836,N_9365);
nand U13659 (N_13659,N_10599,N_9716);
and U13660 (N_13660,N_10404,N_9424);
or U13661 (N_13661,N_9507,N_9408);
nor U13662 (N_13662,N_10827,N_9997);
or U13663 (N_13663,N_9166,N_10014);
or U13664 (N_13664,N_11094,N_9462);
or U13665 (N_13665,N_9917,N_10503);
xnor U13666 (N_13666,N_10534,N_9600);
nor U13667 (N_13667,N_10501,N_10855);
nor U13668 (N_13668,N_10052,N_10314);
nand U13669 (N_13669,N_11628,N_9255);
nand U13670 (N_13670,N_10673,N_9432);
nor U13671 (N_13671,N_11453,N_9099);
nor U13672 (N_13672,N_9976,N_10162);
and U13673 (N_13673,N_10256,N_10276);
or U13674 (N_13674,N_11729,N_10647);
and U13675 (N_13675,N_10265,N_9069);
nor U13676 (N_13676,N_10054,N_11943);
nand U13677 (N_13677,N_11085,N_9666);
xor U13678 (N_13678,N_11094,N_9245);
nand U13679 (N_13679,N_10708,N_11509);
or U13680 (N_13680,N_11864,N_11330);
nand U13681 (N_13681,N_11802,N_10897);
or U13682 (N_13682,N_11479,N_10444);
nand U13683 (N_13683,N_9470,N_11494);
and U13684 (N_13684,N_9930,N_10623);
or U13685 (N_13685,N_11520,N_10329);
or U13686 (N_13686,N_10524,N_10734);
or U13687 (N_13687,N_11585,N_11962);
nand U13688 (N_13688,N_9337,N_9931);
nand U13689 (N_13689,N_9581,N_11681);
xor U13690 (N_13690,N_11450,N_9564);
or U13691 (N_13691,N_9675,N_10160);
or U13692 (N_13692,N_9180,N_10255);
nor U13693 (N_13693,N_11292,N_9244);
or U13694 (N_13694,N_11905,N_11779);
nand U13695 (N_13695,N_10833,N_10164);
xnor U13696 (N_13696,N_10225,N_10410);
nand U13697 (N_13697,N_10256,N_9117);
nand U13698 (N_13698,N_10007,N_11970);
xor U13699 (N_13699,N_9231,N_9159);
nor U13700 (N_13700,N_10542,N_9283);
and U13701 (N_13701,N_11410,N_11830);
or U13702 (N_13702,N_11117,N_9981);
nand U13703 (N_13703,N_11781,N_11682);
and U13704 (N_13704,N_9042,N_10685);
nor U13705 (N_13705,N_11862,N_10633);
nand U13706 (N_13706,N_10692,N_9942);
xnor U13707 (N_13707,N_10295,N_10649);
xnor U13708 (N_13708,N_11825,N_9592);
or U13709 (N_13709,N_9314,N_11246);
or U13710 (N_13710,N_11170,N_10132);
nand U13711 (N_13711,N_11929,N_10058);
nor U13712 (N_13712,N_10511,N_10137);
and U13713 (N_13713,N_10958,N_9278);
or U13714 (N_13714,N_10688,N_11742);
or U13715 (N_13715,N_9289,N_9456);
xnor U13716 (N_13716,N_9572,N_10196);
nor U13717 (N_13717,N_9713,N_9570);
and U13718 (N_13718,N_11631,N_9060);
nand U13719 (N_13719,N_10742,N_10856);
nor U13720 (N_13720,N_11382,N_10108);
nand U13721 (N_13721,N_10947,N_10187);
nor U13722 (N_13722,N_10761,N_9897);
and U13723 (N_13723,N_11215,N_10107);
nand U13724 (N_13724,N_9360,N_10746);
or U13725 (N_13725,N_10267,N_10776);
and U13726 (N_13726,N_10412,N_10676);
and U13727 (N_13727,N_10590,N_9771);
and U13728 (N_13728,N_10031,N_10484);
nand U13729 (N_13729,N_9805,N_10292);
or U13730 (N_13730,N_11143,N_10355);
and U13731 (N_13731,N_9399,N_9983);
nand U13732 (N_13732,N_9290,N_11536);
xor U13733 (N_13733,N_10292,N_9177);
nor U13734 (N_13734,N_11820,N_10054);
nor U13735 (N_13735,N_9008,N_10675);
and U13736 (N_13736,N_11343,N_10993);
or U13737 (N_13737,N_10444,N_9183);
nand U13738 (N_13738,N_11432,N_11798);
xnor U13739 (N_13739,N_9058,N_10601);
nand U13740 (N_13740,N_10189,N_9525);
nand U13741 (N_13741,N_10931,N_11011);
nor U13742 (N_13742,N_9127,N_10565);
nand U13743 (N_13743,N_9923,N_9529);
and U13744 (N_13744,N_11512,N_11014);
and U13745 (N_13745,N_10396,N_9197);
nor U13746 (N_13746,N_10632,N_10810);
nor U13747 (N_13747,N_10708,N_11762);
and U13748 (N_13748,N_11781,N_10512);
nor U13749 (N_13749,N_10264,N_11343);
and U13750 (N_13750,N_10872,N_9237);
nor U13751 (N_13751,N_9058,N_9123);
xnor U13752 (N_13752,N_11322,N_11125);
nand U13753 (N_13753,N_11953,N_9355);
nor U13754 (N_13754,N_11082,N_11027);
nand U13755 (N_13755,N_11579,N_9720);
nand U13756 (N_13756,N_11118,N_11054);
nor U13757 (N_13757,N_9205,N_9905);
or U13758 (N_13758,N_10254,N_9820);
nand U13759 (N_13759,N_10058,N_10524);
nand U13760 (N_13760,N_11119,N_11549);
nand U13761 (N_13761,N_10061,N_9288);
nand U13762 (N_13762,N_11091,N_9548);
nand U13763 (N_13763,N_10941,N_10335);
nor U13764 (N_13764,N_11739,N_9333);
and U13765 (N_13765,N_9465,N_10819);
nor U13766 (N_13766,N_10231,N_9883);
nand U13767 (N_13767,N_10862,N_9969);
or U13768 (N_13768,N_9013,N_9342);
or U13769 (N_13769,N_10512,N_11809);
nand U13770 (N_13770,N_11249,N_10365);
nand U13771 (N_13771,N_9199,N_9078);
nor U13772 (N_13772,N_9467,N_11440);
nor U13773 (N_13773,N_10700,N_11001);
nor U13774 (N_13774,N_9718,N_9661);
nand U13775 (N_13775,N_11704,N_10250);
or U13776 (N_13776,N_10037,N_10939);
xor U13777 (N_13777,N_11141,N_11369);
nor U13778 (N_13778,N_11352,N_9518);
nor U13779 (N_13779,N_10000,N_10802);
or U13780 (N_13780,N_11159,N_11047);
and U13781 (N_13781,N_11028,N_10248);
nand U13782 (N_13782,N_11301,N_11506);
and U13783 (N_13783,N_10388,N_11968);
and U13784 (N_13784,N_9262,N_11161);
nor U13785 (N_13785,N_11752,N_11810);
nand U13786 (N_13786,N_9900,N_11142);
and U13787 (N_13787,N_9818,N_9699);
nor U13788 (N_13788,N_11010,N_9136);
nor U13789 (N_13789,N_11328,N_9901);
nand U13790 (N_13790,N_9851,N_9591);
nor U13791 (N_13791,N_10963,N_11638);
or U13792 (N_13792,N_9109,N_10587);
nor U13793 (N_13793,N_9470,N_10988);
xor U13794 (N_13794,N_11447,N_11421);
nand U13795 (N_13795,N_9442,N_11633);
or U13796 (N_13796,N_11543,N_10000);
and U13797 (N_13797,N_11139,N_10178);
and U13798 (N_13798,N_11205,N_10867);
and U13799 (N_13799,N_9419,N_11892);
nor U13800 (N_13800,N_10483,N_11278);
or U13801 (N_13801,N_11955,N_11650);
or U13802 (N_13802,N_10843,N_10745);
nand U13803 (N_13803,N_10204,N_10945);
nor U13804 (N_13804,N_9026,N_11573);
nor U13805 (N_13805,N_11470,N_11138);
nand U13806 (N_13806,N_9806,N_9672);
and U13807 (N_13807,N_9396,N_11451);
nand U13808 (N_13808,N_9022,N_11970);
nor U13809 (N_13809,N_11686,N_11019);
nor U13810 (N_13810,N_10790,N_10066);
or U13811 (N_13811,N_10364,N_9477);
nand U13812 (N_13812,N_11905,N_11033);
or U13813 (N_13813,N_9807,N_11907);
or U13814 (N_13814,N_9343,N_9677);
nand U13815 (N_13815,N_9239,N_9007);
and U13816 (N_13816,N_9275,N_9129);
nor U13817 (N_13817,N_11034,N_11798);
and U13818 (N_13818,N_10428,N_9996);
xor U13819 (N_13819,N_10507,N_11841);
nand U13820 (N_13820,N_11894,N_11131);
xnor U13821 (N_13821,N_11696,N_11377);
nand U13822 (N_13822,N_11308,N_11500);
or U13823 (N_13823,N_10009,N_9631);
nor U13824 (N_13824,N_11045,N_10785);
nand U13825 (N_13825,N_11691,N_10379);
nand U13826 (N_13826,N_10800,N_11127);
nand U13827 (N_13827,N_9546,N_9147);
xnor U13828 (N_13828,N_10855,N_10332);
nor U13829 (N_13829,N_10698,N_10189);
xnor U13830 (N_13830,N_11625,N_9043);
nor U13831 (N_13831,N_9693,N_10308);
nand U13832 (N_13832,N_11034,N_9128);
or U13833 (N_13833,N_10081,N_10595);
nor U13834 (N_13834,N_9810,N_11898);
or U13835 (N_13835,N_10251,N_9772);
xnor U13836 (N_13836,N_11145,N_9995);
and U13837 (N_13837,N_11184,N_10890);
nor U13838 (N_13838,N_9224,N_10794);
nand U13839 (N_13839,N_11043,N_11384);
or U13840 (N_13840,N_9055,N_11605);
nand U13841 (N_13841,N_10514,N_11576);
nand U13842 (N_13842,N_10364,N_11965);
nand U13843 (N_13843,N_10906,N_11369);
and U13844 (N_13844,N_10931,N_11251);
nand U13845 (N_13845,N_11715,N_11937);
nor U13846 (N_13846,N_10766,N_10933);
and U13847 (N_13847,N_9367,N_10029);
and U13848 (N_13848,N_10301,N_11490);
nor U13849 (N_13849,N_9702,N_10846);
nor U13850 (N_13850,N_10332,N_9255);
nand U13851 (N_13851,N_9296,N_10868);
xnor U13852 (N_13852,N_10362,N_10536);
nand U13853 (N_13853,N_10385,N_9206);
nor U13854 (N_13854,N_10389,N_11883);
xor U13855 (N_13855,N_11238,N_9845);
nand U13856 (N_13856,N_10682,N_11828);
nand U13857 (N_13857,N_11711,N_10688);
nand U13858 (N_13858,N_10609,N_9731);
or U13859 (N_13859,N_9861,N_10926);
xnor U13860 (N_13860,N_10025,N_10481);
xnor U13861 (N_13861,N_9193,N_9031);
nand U13862 (N_13862,N_10266,N_10380);
xor U13863 (N_13863,N_10161,N_10157);
xnor U13864 (N_13864,N_11487,N_10422);
nand U13865 (N_13865,N_9146,N_9580);
and U13866 (N_13866,N_11573,N_11686);
nor U13867 (N_13867,N_11882,N_9062);
and U13868 (N_13868,N_10815,N_9023);
and U13869 (N_13869,N_9692,N_10689);
or U13870 (N_13870,N_10542,N_11444);
nand U13871 (N_13871,N_10552,N_9542);
xor U13872 (N_13872,N_10052,N_10158);
nor U13873 (N_13873,N_10824,N_9038);
nor U13874 (N_13874,N_10181,N_10123);
and U13875 (N_13875,N_11160,N_9291);
nor U13876 (N_13876,N_9479,N_10259);
nand U13877 (N_13877,N_10366,N_9013);
or U13878 (N_13878,N_9931,N_9761);
and U13879 (N_13879,N_9452,N_9392);
nor U13880 (N_13880,N_9494,N_10570);
nor U13881 (N_13881,N_9501,N_10027);
nand U13882 (N_13882,N_9542,N_11238);
or U13883 (N_13883,N_10936,N_10642);
nor U13884 (N_13884,N_11025,N_10310);
and U13885 (N_13885,N_10636,N_11824);
nor U13886 (N_13886,N_11162,N_9209);
nor U13887 (N_13887,N_11598,N_9382);
nand U13888 (N_13888,N_10526,N_11101);
nand U13889 (N_13889,N_11372,N_9544);
or U13890 (N_13890,N_10489,N_9866);
xnor U13891 (N_13891,N_10997,N_11651);
or U13892 (N_13892,N_11250,N_9650);
and U13893 (N_13893,N_9037,N_9055);
nor U13894 (N_13894,N_11735,N_10744);
nor U13895 (N_13895,N_10686,N_9444);
or U13896 (N_13896,N_9377,N_9252);
and U13897 (N_13897,N_9683,N_10675);
xor U13898 (N_13898,N_10203,N_11954);
and U13899 (N_13899,N_10044,N_10795);
nor U13900 (N_13900,N_11787,N_10252);
and U13901 (N_13901,N_11238,N_10233);
nand U13902 (N_13902,N_11446,N_10745);
or U13903 (N_13903,N_10859,N_10740);
nand U13904 (N_13904,N_10945,N_11528);
or U13905 (N_13905,N_10148,N_9885);
or U13906 (N_13906,N_9518,N_9295);
nand U13907 (N_13907,N_10792,N_11669);
or U13908 (N_13908,N_10941,N_9583);
nand U13909 (N_13909,N_10476,N_9124);
or U13910 (N_13910,N_10400,N_9338);
xor U13911 (N_13911,N_9740,N_10819);
and U13912 (N_13912,N_9692,N_9320);
xnor U13913 (N_13913,N_9125,N_10958);
nor U13914 (N_13914,N_11873,N_10926);
and U13915 (N_13915,N_10227,N_10970);
nor U13916 (N_13916,N_9200,N_10305);
and U13917 (N_13917,N_9375,N_9333);
nor U13918 (N_13918,N_9183,N_11506);
nor U13919 (N_13919,N_11922,N_9898);
nor U13920 (N_13920,N_9395,N_11606);
or U13921 (N_13921,N_9957,N_9263);
or U13922 (N_13922,N_9239,N_10270);
and U13923 (N_13923,N_11851,N_10788);
and U13924 (N_13924,N_9657,N_9206);
or U13925 (N_13925,N_11620,N_9380);
nand U13926 (N_13926,N_11798,N_11898);
nor U13927 (N_13927,N_9768,N_10175);
and U13928 (N_13928,N_9961,N_11045);
and U13929 (N_13929,N_9190,N_10827);
nand U13930 (N_13930,N_11283,N_10451);
and U13931 (N_13931,N_10229,N_11854);
nand U13932 (N_13932,N_9553,N_10034);
nand U13933 (N_13933,N_11412,N_10960);
or U13934 (N_13934,N_11892,N_9451);
nor U13935 (N_13935,N_9499,N_11133);
xor U13936 (N_13936,N_10486,N_11709);
and U13937 (N_13937,N_10041,N_10524);
nand U13938 (N_13938,N_10521,N_10570);
and U13939 (N_13939,N_9293,N_10069);
or U13940 (N_13940,N_11381,N_10967);
xor U13941 (N_13941,N_11421,N_9276);
xnor U13942 (N_13942,N_10305,N_11700);
nor U13943 (N_13943,N_10367,N_11555);
nor U13944 (N_13944,N_11897,N_10131);
or U13945 (N_13945,N_10158,N_11103);
and U13946 (N_13946,N_11021,N_11840);
and U13947 (N_13947,N_11709,N_11231);
or U13948 (N_13948,N_9251,N_10936);
xor U13949 (N_13949,N_10702,N_9501);
nor U13950 (N_13950,N_10459,N_11015);
nor U13951 (N_13951,N_9344,N_11887);
xor U13952 (N_13952,N_9585,N_10983);
or U13953 (N_13953,N_10604,N_11531);
xor U13954 (N_13954,N_9614,N_11132);
or U13955 (N_13955,N_11698,N_11072);
nor U13956 (N_13956,N_11594,N_9077);
xnor U13957 (N_13957,N_11024,N_10137);
nand U13958 (N_13958,N_10651,N_10557);
and U13959 (N_13959,N_9953,N_10232);
and U13960 (N_13960,N_11910,N_9489);
nand U13961 (N_13961,N_11740,N_10950);
or U13962 (N_13962,N_9840,N_9966);
or U13963 (N_13963,N_9772,N_10534);
or U13964 (N_13964,N_10596,N_10982);
nor U13965 (N_13965,N_9153,N_11271);
nor U13966 (N_13966,N_10778,N_10014);
nor U13967 (N_13967,N_9726,N_11163);
nor U13968 (N_13968,N_10408,N_10513);
and U13969 (N_13969,N_10314,N_11419);
or U13970 (N_13970,N_11487,N_10641);
or U13971 (N_13971,N_9836,N_11092);
nand U13972 (N_13972,N_10690,N_10048);
nor U13973 (N_13973,N_10102,N_9272);
xor U13974 (N_13974,N_10016,N_11223);
xor U13975 (N_13975,N_11208,N_10515);
or U13976 (N_13976,N_9034,N_9432);
and U13977 (N_13977,N_9182,N_11421);
or U13978 (N_13978,N_10299,N_10808);
nor U13979 (N_13979,N_11763,N_11533);
or U13980 (N_13980,N_10661,N_10093);
nor U13981 (N_13981,N_10441,N_11154);
or U13982 (N_13982,N_10444,N_10882);
nor U13983 (N_13983,N_11202,N_10358);
and U13984 (N_13984,N_11510,N_11298);
nor U13985 (N_13985,N_9070,N_10665);
and U13986 (N_13986,N_11687,N_9276);
and U13987 (N_13987,N_11995,N_11096);
nand U13988 (N_13988,N_9005,N_11477);
or U13989 (N_13989,N_11793,N_9745);
or U13990 (N_13990,N_9243,N_9637);
nand U13991 (N_13991,N_9082,N_10155);
or U13992 (N_13992,N_10363,N_9631);
or U13993 (N_13993,N_10206,N_11444);
or U13994 (N_13994,N_11214,N_11029);
nand U13995 (N_13995,N_9814,N_9590);
nor U13996 (N_13996,N_11835,N_11160);
xnor U13997 (N_13997,N_10040,N_11317);
nand U13998 (N_13998,N_11366,N_9981);
nand U13999 (N_13999,N_11280,N_10057);
nand U14000 (N_14000,N_9327,N_9729);
xnor U14001 (N_14001,N_11622,N_11222);
nor U14002 (N_14002,N_9439,N_9788);
or U14003 (N_14003,N_10671,N_10262);
nand U14004 (N_14004,N_10452,N_11208);
nand U14005 (N_14005,N_9883,N_10449);
and U14006 (N_14006,N_11191,N_10539);
and U14007 (N_14007,N_10425,N_10247);
nor U14008 (N_14008,N_11336,N_10221);
or U14009 (N_14009,N_9416,N_10287);
or U14010 (N_14010,N_11315,N_9671);
nand U14011 (N_14011,N_9389,N_10809);
and U14012 (N_14012,N_10111,N_9778);
nand U14013 (N_14013,N_10703,N_10698);
xnor U14014 (N_14014,N_9369,N_9568);
nand U14015 (N_14015,N_11558,N_9502);
or U14016 (N_14016,N_11382,N_10011);
and U14017 (N_14017,N_11369,N_10213);
nor U14018 (N_14018,N_9854,N_10011);
nor U14019 (N_14019,N_9155,N_9658);
and U14020 (N_14020,N_11814,N_11236);
nand U14021 (N_14021,N_10323,N_11908);
nor U14022 (N_14022,N_9291,N_10768);
nand U14023 (N_14023,N_11888,N_11722);
or U14024 (N_14024,N_9253,N_11748);
nor U14025 (N_14025,N_11916,N_11396);
nor U14026 (N_14026,N_10161,N_9726);
or U14027 (N_14027,N_9330,N_11741);
and U14028 (N_14028,N_9523,N_9153);
or U14029 (N_14029,N_10195,N_10317);
nand U14030 (N_14030,N_11709,N_10571);
nor U14031 (N_14031,N_10765,N_9946);
or U14032 (N_14032,N_10997,N_10002);
nand U14033 (N_14033,N_10760,N_9891);
nor U14034 (N_14034,N_10136,N_11016);
nor U14035 (N_14035,N_10530,N_11338);
and U14036 (N_14036,N_10605,N_10307);
nor U14037 (N_14037,N_9669,N_10496);
and U14038 (N_14038,N_11142,N_11330);
or U14039 (N_14039,N_11566,N_11908);
nor U14040 (N_14040,N_9783,N_10849);
or U14041 (N_14041,N_9566,N_10122);
nor U14042 (N_14042,N_10462,N_10142);
nand U14043 (N_14043,N_9993,N_10745);
and U14044 (N_14044,N_9680,N_11833);
nand U14045 (N_14045,N_9477,N_9302);
nor U14046 (N_14046,N_9516,N_11578);
nor U14047 (N_14047,N_11118,N_11587);
nor U14048 (N_14048,N_10411,N_10317);
and U14049 (N_14049,N_10756,N_9627);
or U14050 (N_14050,N_11297,N_11906);
nor U14051 (N_14051,N_10581,N_10061);
nor U14052 (N_14052,N_10526,N_9019);
nand U14053 (N_14053,N_10973,N_10225);
nor U14054 (N_14054,N_11590,N_11399);
or U14055 (N_14055,N_11348,N_9102);
nand U14056 (N_14056,N_9614,N_9357);
and U14057 (N_14057,N_9562,N_10850);
nand U14058 (N_14058,N_9045,N_10916);
or U14059 (N_14059,N_10535,N_11554);
and U14060 (N_14060,N_9710,N_9770);
nand U14061 (N_14061,N_10047,N_9089);
nor U14062 (N_14062,N_11088,N_9107);
xnor U14063 (N_14063,N_10255,N_10347);
nand U14064 (N_14064,N_11797,N_9284);
nor U14065 (N_14065,N_9740,N_10045);
nand U14066 (N_14066,N_11385,N_9688);
or U14067 (N_14067,N_9770,N_11542);
nand U14068 (N_14068,N_9158,N_9153);
nor U14069 (N_14069,N_10068,N_10895);
or U14070 (N_14070,N_10136,N_11374);
or U14071 (N_14071,N_9974,N_11762);
nor U14072 (N_14072,N_10802,N_10070);
nand U14073 (N_14073,N_10488,N_9889);
or U14074 (N_14074,N_11535,N_10305);
and U14075 (N_14075,N_11103,N_9599);
and U14076 (N_14076,N_9738,N_11946);
and U14077 (N_14077,N_9147,N_10850);
or U14078 (N_14078,N_11312,N_11363);
xnor U14079 (N_14079,N_10071,N_11533);
and U14080 (N_14080,N_11777,N_11086);
and U14081 (N_14081,N_11332,N_10919);
and U14082 (N_14082,N_11164,N_10350);
nor U14083 (N_14083,N_11135,N_11055);
and U14084 (N_14084,N_11924,N_9228);
and U14085 (N_14085,N_11418,N_11752);
nor U14086 (N_14086,N_9923,N_10200);
nor U14087 (N_14087,N_11687,N_9885);
and U14088 (N_14088,N_11640,N_10912);
nor U14089 (N_14089,N_9960,N_9166);
nor U14090 (N_14090,N_9806,N_10397);
and U14091 (N_14091,N_10106,N_9116);
and U14092 (N_14092,N_10516,N_10595);
nor U14093 (N_14093,N_11479,N_9546);
nand U14094 (N_14094,N_10011,N_9749);
nor U14095 (N_14095,N_11964,N_11597);
and U14096 (N_14096,N_10035,N_10203);
nand U14097 (N_14097,N_10402,N_11465);
nand U14098 (N_14098,N_9062,N_10311);
nand U14099 (N_14099,N_9330,N_11715);
and U14100 (N_14100,N_10360,N_11708);
nor U14101 (N_14101,N_9559,N_9900);
and U14102 (N_14102,N_10320,N_10729);
nand U14103 (N_14103,N_10748,N_10300);
nand U14104 (N_14104,N_10564,N_9442);
and U14105 (N_14105,N_9753,N_10405);
nand U14106 (N_14106,N_10696,N_10198);
nand U14107 (N_14107,N_10230,N_10987);
or U14108 (N_14108,N_10483,N_10200);
and U14109 (N_14109,N_11335,N_10902);
and U14110 (N_14110,N_9101,N_11463);
and U14111 (N_14111,N_9336,N_10361);
nor U14112 (N_14112,N_10992,N_9838);
nand U14113 (N_14113,N_9586,N_9191);
nor U14114 (N_14114,N_11685,N_11929);
nor U14115 (N_14115,N_10153,N_9653);
or U14116 (N_14116,N_10824,N_9665);
nor U14117 (N_14117,N_10132,N_11830);
or U14118 (N_14118,N_9913,N_11722);
xor U14119 (N_14119,N_11891,N_10572);
or U14120 (N_14120,N_11277,N_10089);
nand U14121 (N_14121,N_10527,N_11242);
nor U14122 (N_14122,N_10822,N_9229);
or U14123 (N_14123,N_11222,N_10704);
xnor U14124 (N_14124,N_10844,N_9146);
xor U14125 (N_14125,N_11620,N_10689);
nor U14126 (N_14126,N_11990,N_11934);
nand U14127 (N_14127,N_10443,N_11559);
or U14128 (N_14128,N_11720,N_10759);
or U14129 (N_14129,N_9130,N_10957);
or U14130 (N_14130,N_11886,N_11942);
nand U14131 (N_14131,N_10303,N_11132);
and U14132 (N_14132,N_9201,N_9700);
xnor U14133 (N_14133,N_11257,N_9078);
nor U14134 (N_14134,N_11927,N_9573);
nor U14135 (N_14135,N_10511,N_9699);
and U14136 (N_14136,N_10752,N_9408);
nor U14137 (N_14137,N_10812,N_11271);
nor U14138 (N_14138,N_11733,N_9165);
or U14139 (N_14139,N_11208,N_10545);
or U14140 (N_14140,N_10707,N_10224);
nor U14141 (N_14141,N_9316,N_9048);
nand U14142 (N_14142,N_11458,N_10813);
nand U14143 (N_14143,N_11480,N_10151);
nor U14144 (N_14144,N_11011,N_10721);
and U14145 (N_14145,N_11632,N_10731);
nand U14146 (N_14146,N_11620,N_10087);
or U14147 (N_14147,N_10730,N_11566);
and U14148 (N_14148,N_9192,N_9227);
nor U14149 (N_14149,N_11588,N_10092);
xor U14150 (N_14150,N_9205,N_11934);
and U14151 (N_14151,N_10930,N_11170);
nand U14152 (N_14152,N_9417,N_11016);
nand U14153 (N_14153,N_9036,N_9459);
or U14154 (N_14154,N_11555,N_10044);
and U14155 (N_14155,N_11656,N_9521);
or U14156 (N_14156,N_11597,N_10643);
xnor U14157 (N_14157,N_10466,N_11641);
nor U14158 (N_14158,N_9927,N_9095);
or U14159 (N_14159,N_11945,N_10428);
and U14160 (N_14160,N_10894,N_10087);
xor U14161 (N_14161,N_10854,N_11125);
nor U14162 (N_14162,N_10923,N_9022);
or U14163 (N_14163,N_10067,N_11056);
nand U14164 (N_14164,N_10822,N_11898);
nor U14165 (N_14165,N_11591,N_11898);
xor U14166 (N_14166,N_9836,N_9702);
nand U14167 (N_14167,N_9635,N_9823);
and U14168 (N_14168,N_9901,N_10912);
nor U14169 (N_14169,N_11493,N_10709);
nor U14170 (N_14170,N_11486,N_9892);
and U14171 (N_14171,N_11843,N_10751);
xnor U14172 (N_14172,N_9804,N_10201);
nor U14173 (N_14173,N_11201,N_10634);
nor U14174 (N_14174,N_10527,N_10116);
and U14175 (N_14175,N_9379,N_9933);
xor U14176 (N_14176,N_9255,N_10357);
or U14177 (N_14177,N_10789,N_11259);
and U14178 (N_14178,N_10503,N_10849);
nor U14179 (N_14179,N_9256,N_9468);
nand U14180 (N_14180,N_9957,N_9247);
xnor U14181 (N_14181,N_9862,N_9027);
or U14182 (N_14182,N_9228,N_11780);
nand U14183 (N_14183,N_11107,N_11659);
or U14184 (N_14184,N_11128,N_11629);
or U14185 (N_14185,N_10567,N_9432);
or U14186 (N_14186,N_10913,N_10515);
xnor U14187 (N_14187,N_11984,N_10010);
xnor U14188 (N_14188,N_9069,N_9192);
xor U14189 (N_14189,N_11592,N_10127);
nand U14190 (N_14190,N_10753,N_9367);
or U14191 (N_14191,N_9002,N_10024);
xor U14192 (N_14192,N_10625,N_9121);
nand U14193 (N_14193,N_9547,N_11716);
or U14194 (N_14194,N_11693,N_11010);
nand U14195 (N_14195,N_10220,N_9023);
nand U14196 (N_14196,N_11836,N_10333);
or U14197 (N_14197,N_11260,N_11565);
nor U14198 (N_14198,N_11449,N_10439);
and U14199 (N_14199,N_11278,N_11343);
nand U14200 (N_14200,N_10126,N_10496);
nand U14201 (N_14201,N_10604,N_9754);
xnor U14202 (N_14202,N_9156,N_9649);
nor U14203 (N_14203,N_9598,N_10388);
nor U14204 (N_14204,N_9145,N_11422);
nand U14205 (N_14205,N_9394,N_11610);
and U14206 (N_14206,N_10211,N_11782);
or U14207 (N_14207,N_9727,N_9905);
nand U14208 (N_14208,N_10045,N_10778);
nor U14209 (N_14209,N_9235,N_10717);
or U14210 (N_14210,N_10314,N_10853);
nor U14211 (N_14211,N_11208,N_10048);
or U14212 (N_14212,N_10184,N_9765);
or U14213 (N_14213,N_10914,N_10828);
and U14214 (N_14214,N_10988,N_10285);
nand U14215 (N_14215,N_11062,N_11287);
nand U14216 (N_14216,N_9194,N_11765);
nand U14217 (N_14217,N_11657,N_10773);
nor U14218 (N_14218,N_11735,N_11407);
nor U14219 (N_14219,N_11407,N_9838);
xnor U14220 (N_14220,N_9350,N_10832);
nand U14221 (N_14221,N_11762,N_11434);
and U14222 (N_14222,N_9287,N_9397);
xor U14223 (N_14223,N_11618,N_10089);
or U14224 (N_14224,N_10710,N_11755);
or U14225 (N_14225,N_9388,N_9376);
and U14226 (N_14226,N_11076,N_10373);
xor U14227 (N_14227,N_9676,N_9247);
nor U14228 (N_14228,N_11352,N_11148);
nand U14229 (N_14229,N_9124,N_10958);
or U14230 (N_14230,N_10490,N_11835);
and U14231 (N_14231,N_10553,N_9723);
xnor U14232 (N_14232,N_11961,N_11301);
and U14233 (N_14233,N_11524,N_9896);
or U14234 (N_14234,N_11485,N_10559);
or U14235 (N_14235,N_10342,N_11610);
or U14236 (N_14236,N_11668,N_11754);
and U14237 (N_14237,N_11649,N_11757);
and U14238 (N_14238,N_11200,N_11866);
nor U14239 (N_14239,N_9135,N_9516);
or U14240 (N_14240,N_11285,N_9502);
and U14241 (N_14241,N_11256,N_9738);
nand U14242 (N_14242,N_11406,N_11448);
nand U14243 (N_14243,N_9206,N_10559);
nand U14244 (N_14244,N_9070,N_11485);
nor U14245 (N_14245,N_10904,N_11199);
nor U14246 (N_14246,N_11459,N_10890);
and U14247 (N_14247,N_11115,N_9449);
and U14248 (N_14248,N_9102,N_10893);
or U14249 (N_14249,N_9391,N_9553);
xor U14250 (N_14250,N_9601,N_10678);
and U14251 (N_14251,N_9434,N_9111);
nor U14252 (N_14252,N_11615,N_11452);
nor U14253 (N_14253,N_11924,N_9961);
or U14254 (N_14254,N_11733,N_10015);
or U14255 (N_14255,N_10359,N_9944);
and U14256 (N_14256,N_11574,N_9404);
nand U14257 (N_14257,N_10405,N_9247);
nand U14258 (N_14258,N_11981,N_9902);
and U14259 (N_14259,N_9231,N_11608);
or U14260 (N_14260,N_9976,N_10979);
nor U14261 (N_14261,N_11428,N_11773);
nand U14262 (N_14262,N_10329,N_11321);
nand U14263 (N_14263,N_9785,N_10383);
nand U14264 (N_14264,N_9183,N_10059);
or U14265 (N_14265,N_9879,N_11851);
xor U14266 (N_14266,N_11167,N_9774);
nor U14267 (N_14267,N_10948,N_9068);
or U14268 (N_14268,N_9006,N_11650);
nand U14269 (N_14269,N_9568,N_10056);
nor U14270 (N_14270,N_9950,N_11531);
or U14271 (N_14271,N_9802,N_10086);
nor U14272 (N_14272,N_10204,N_11327);
or U14273 (N_14273,N_11374,N_9580);
nor U14274 (N_14274,N_11151,N_11072);
nand U14275 (N_14275,N_10439,N_11720);
or U14276 (N_14276,N_9522,N_9054);
or U14277 (N_14277,N_11090,N_11543);
nor U14278 (N_14278,N_10312,N_9306);
nand U14279 (N_14279,N_11102,N_11910);
or U14280 (N_14280,N_9477,N_10164);
nor U14281 (N_14281,N_9343,N_10791);
or U14282 (N_14282,N_11915,N_9867);
or U14283 (N_14283,N_9899,N_10521);
nand U14284 (N_14284,N_10161,N_10962);
xnor U14285 (N_14285,N_9683,N_10084);
or U14286 (N_14286,N_9705,N_10412);
or U14287 (N_14287,N_10415,N_9380);
nand U14288 (N_14288,N_9825,N_11786);
or U14289 (N_14289,N_9284,N_9297);
and U14290 (N_14290,N_9379,N_9666);
xnor U14291 (N_14291,N_9888,N_9767);
or U14292 (N_14292,N_10548,N_10122);
and U14293 (N_14293,N_9444,N_10333);
or U14294 (N_14294,N_9711,N_10232);
or U14295 (N_14295,N_10536,N_9972);
nand U14296 (N_14296,N_11637,N_10091);
and U14297 (N_14297,N_10168,N_9658);
and U14298 (N_14298,N_11967,N_11543);
nand U14299 (N_14299,N_9952,N_10104);
or U14300 (N_14300,N_9175,N_11526);
nor U14301 (N_14301,N_9781,N_9745);
nand U14302 (N_14302,N_9518,N_10826);
nand U14303 (N_14303,N_9699,N_9323);
nand U14304 (N_14304,N_11831,N_10256);
or U14305 (N_14305,N_11515,N_11356);
nor U14306 (N_14306,N_11563,N_9822);
or U14307 (N_14307,N_10526,N_9520);
and U14308 (N_14308,N_11880,N_9277);
or U14309 (N_14309,N_11022,N_10669);
nand U14310 (N_14310,N_9996,N_10897);
or U14311 (N_14311,N_9995,N_11927);
or U14312 (N_14312,N_9284,N_11821);
xnor U14313 (N_14313,N_9782,N_10448);
nand U14314 (N_14314,N_10778,N_10477);
xor U14315 (N_14315,N_9982,N_11466);
nor U14316 (N_14316,N_10277,N_11784);
and U14317 (N_14317,N_11660,N_9122);
nor U14318 (N_14318,N_11660,N_9135);
nand U14319 (N_14319,N_10477,N_11994);
nor U14320 (N_14320,N_11339,N_11529);
and U14321 (N_14321,N_11800,N_10948);
nand U14322 (N_14322,N_10556,N_10125);
nand U14323 (N_14323,N_9860,N_10476);
nor U14324 (N_14324,N_9659,N_10625);
nand U14325 (N_14325,N_9189,N_11395);
nand U14326 (N_14326,N_11958,N_10005);
xor U14327 (N_14327,N_11304,N_10237);
and U14328 (N_14328,N_10555,N_11726);
and U14329 (N_14329,N_10085,N_11765);
or U14330 (N_14330,N_11625,N_9024);
or U14331 (N_14331,N_10413,N_11237);
nand U14332 (N_14332,N_11106,N_9658);
nand U14333 (N_14333,N_11282,N_10885);
nor U14334 (N_14334,N_9119,N_11424);
nor U14335 (N_14335,N_9534,N_10013);
nand U14336 (N_14336,N_10673,N_11513);
nand U14337 (N_14337,N_9905,N_10365);
xor U14338 (N_14338,N_9776,N_10538);
nand U14339 (N_14339,N_11446,N_10947);
nand U14340 (N_14340,N_11122,N_10773);
and U14341 (N_14341,N_11947,N_10368);
nand U14342 (N_14342,N_9038,N_11425);
and U14343 (N_14343,N_10777,N_11599);
xor U14344 (N_14344,N_9060,N_11151);
and U14345 (N_14345,N_11552,N_10507);
xor U14346 (N_14346,N_10696,N_11485);
nor U14347 (N_14347,N_11133,N_11621);
and U14348 (N_14348,N_11798,N_11040);
or U14349 (N_14349,N_9531,N_11007);
and U14350 (N_14350,N_9686,N_11338);
or U14351 (N_14351,N_9893,N_11959);
nor U14352 (N_14352,N_11245,N_10570);
or U14353 (N_14353,N_9487,N_10453);
or U14354 (N_14354,N_9958,N_9020);
and U14355 (N_14355,N_11747,N_11242);
nor U14356 (N_14356,N_11141,N_11616);
and U14357 (N_14357,N_9617,N_11269);
xor U14358 (N_14358,N_9747,N_11493);
or U14359 (N_14359,N_10022,N_9708);
and U14360 (N_14360,N_9113,N_9643);
nand U14361 (N_14361,N_11036,N_10912);
nor U14362 (N_14362,N_9896,N_10306);
or U14363 (N_14363,N_11253,N_9692);
or U14364 (N_14364,N_9813,N_11196);
nor U14365 (N_14365,N_10399,N_10629);
and U14366 (N_14366,N_11711,N_9790);
nor U14367 (N_14367,N_9296,N_11926);
nor U14368 (N_14368,N_9058,N_11225);
and U14369 (N_14369,N_10263,N_11347);
or U14370 (N_14370,N_11212,N_11148);
nand U14371 (N_14371,N_9022,N_11926);
xor U14372 (N_14372,N_11163,N_11862);
nand U14373 (N_14373,N_11356,N_11062);
nor U14374 (N_14374,N_11293,N_9525);
and U14375 (N_14375,N_10962,N_10089);
nand U14376 (N_14376,N_11398,N_10977);
and U14377 (N_14377,N_11722,N_10763);
xor U14378 (N_14378,N_11520,N_9831);
or U14379 (N_14379,N_9978,N_10520);
nor U14380 (N_14380,N_9651,N_11284);
or U14381 (N_14381,N_11053,N_9835);
nor U14382 (N_14382,N_9539,N_11680);
nor U14383 (N_14383,N_10756,N_10925);
nand U14384 (N_14384,N_9531,N_11400);
nor U14385 (N_14385,N_9448,N_11101);
and U14386 (N_14386,N_11784,N_11666);
nor U14387 (N_14387,N_11744,N_11969);
and U14388 (N_14388,N_10351,N_9039);
or U14389 (N_14389,N_10284,N_11235);
nand U14390 (N_14390,N_11861,N_10859);
xor U14391 (N_14391,N_9700,N_11841);
and U14392 (N_14392,N_10579,N_9543);
or U14393 (N_14393,N_11261,N_9436);
or U14394 (N_14394,N_11334,N_9773);
and U14395 (N_14395,N_11202,N_9450);
nand U14396 (N_14396,N_10806,N_10415);
and U14397 (N_14397,N_11308,N_9689);
nand U14398 (N_14398,N_9466,N_11098);
or U14399 (N_14399,N_9772,N_10669);
and U14400 (N_14400,N_10170,N_10829);
nor U14401 (N_14401,N_9777,N_10251);
and U14402 (N_14402,N_10145,N_10963);
or U14403 (N_14403,N_11785,N_11612);
nand U14404 (N_14404,N_11271,N_11009);
and U14405 (N_14405,N_9555,N_10701);
xnor U14406 (N_14406,N_10601,N_10564);
and U14407 (N_14407,N_9125,N_10323);
and U14408 (N_14408,N_10825,N_11940);
nand U14409 (N_14409,N_9404,N_11683);
or U14410 (N_14410,N_10307,N_10035);
nand U14411 (N_14411,N_10404,N_11075);
nand U14412 (N_14412,N_10349,N_11828);
and U14413 (N_14413,N_11295,N_10248);
or U14414 (N_14414,N_10433,N_11358);
nor U14415 (N_14415,N_10664,N_9159);
xor U14416 (N_14416,N_11551,N_10982);
nor U14417 (N_14417,N_9912,N_9027);
or U14418 (N_14418,N_10486,N_10131);
nand U14419 (N_14419,N_9577,N_10534);
nor U14420 (N_14420,N_10358,N_11914);
and U14421 (N_14421,N_10328,N_9411);
and U14422 (N_14422,N_10954,N_9118);
and U14423 (N_14423,N_11271,N_11689);
and U14424 (N_14424,N_9408,N_10936);
or U14425 (N_14425,N_10115,N_11603);
nand U14426 (N_14426,N_10437,N_10267);
or U14427 (N_14427,N_9650,N_11621);
nand U14428 (N_14428,N_11255,N_11388);
nor U14429 (N_14429,N_10369,N_11974);
or U14430 (N_14430,N_10570,N_11663);
nor U14431 (N_14431,N_11544,N_9130);
and U14432 (N_14432,N_11848,N_9543);
or U14433 (N_14433,N_10978,N_10589);
nand U14434 (N_14434,N_10335,N_9675);
or U14435 (N_14435,N_11902,N_10368);
and U14436 (N_14436,N_10849,N_10213);
or U14437 (N_14437,N_9557,N_9595);
or U14438 (N_14438,N_10440,N_11890);
xor U14439 (N_14439,N_10078,N_10580);
and U14440 (N_14440,N_10418,N_10247);
nand U14441 (N_14441,N_9477,N_10399);
or U14442 (N_14442,N_10518,N_11130);
xor U14443 (N_14443,N_9658,N_10923);
and U14444 (N_14444,N_11455,N_11329);
xnor U14445 (N_14445,N_9138,N_11338);
or U14446 (N_14446,N_9061,N_9327);
and U14447 (N_14447,N_10264,N_9998);
or U14448 (N_14448,N_11454,N_9345);
nor U14449 (N_14449,N_11079,N_9195);
nor U14450 (N_14450,N_9415,N_9526);
or U14451 (N_14451,N_11553,N_9866);
and U14452 (N_14452,N_10742,N_9770);
and U14453 (N_14453,N_11745,N_9173);
nand U14454 (N_14454,N_10205,N_10793);
xnor U14455 (N_14455,N_10540,N_9395);
or U14456 (N_14456,N_9224,N_11019);
nor U14457 (N_14457,N_10440,N_9598);
or U14458 (N_14458,N_11158,N_9996);
nor U14459 (N_14459,N_9349,N_9961);
nand U14460 (N_14460,N_10847,N_11182);
nand U14461 (N_14461,N_9115,N_11168);
or U14462 (N_14462,N_10661,N_9914);
or U14463 (N_14463,N_9012,N_11156);
nand U14464 (N_14464,N_9363,N_10046);
or U14465 (N_14465,N_9507,N_9708);
nand U14466 (N_14466,N_11153,N_9216);
or U14467 (N_14467,N_10249,N_10180);
or U14468 (N_14468,N_9600,N_10859);
and U14469 (N_14469,N_9262,N_10444);
nor U14470 (N_14470,N_11560,N_9916);
and U14471 (N_14471,N_11498,N_11781);
or U14472 (N_14472,N_10245,N_10784);
or U14473 (N_14473,N_10700,N_11865);
xnor U14474 (N_14474,N_10016,N_10914);
or U14475 (N_14475,N_11573,N_9276);
and U14476 (N_14476,N_9850,N_9676);
nor U14477 (N_14477,N_11547,N_11182);
nand U14478 (N_14478,N_11866,N_9193);
nor U14479 (N_14479,N_11912,N_11062);
nor U14480 (N_14480,N_10733,N_9563);
nand U14481 (N_14481,N_11407,N_9609);
nand U14482 (N_14482,N_9225,N_9403);
and U14483 (N_14483,N_11346,N_9095);
nand U14484 (N_14484,N_11818,N_10937);
nand U14485 (N_14485,N_10259,N_9624);
or U14486 (N_14486,N_11007,N_11614);
or U14487 (N_14487,N_9533,N_11591);
nand U14488 (N_14488,N_11199,N_10180);
xnor U14489 (N_14489,N_9912,N_9299);
nand U14490 (N_14490,N_9024,N_10742);
nand U14491 (N_14491,N_11455,N_10601);
or U14492 (N_14492,N_10595,N_11572);
and U14493 (N_14493,N_10823,N_10687);
nor U14494 (N_14494,N_9795,N_10916);
or U14495 (N_14495,N_9643,N_10641);
nor U14496 (N_14496,N_10295,N_11301);
or U14497 (N_14497,N_9872,N_11393);
nand U14498 (N_14498,N_11317,N_11430);
nand U14499 (N_14499,N_11114,N_11381);
nor U14500 (N_14500,N_9036,N_11947);
nor U14501 (N_14501,N_9486,N_11031);
or U14502 (N_14502,N_11818,N_9945);
nor U14503 (N_14503,N_10195,N_10405);
or U14504 (N_14504,N_9811,N_9114);
and U14505 (N_14505,N_9695,N_9635);
and U14506 (N_14506,N_9846,N_11748);
nand U14507 (N_14507,N_9530,N_10816);
or U14508 (N_14508,N_9630,N_10642);
and U14509 (N_14509,N_9048,N_10850);
or U14510 (N_14510,N_9270,N_9128);
nand U14511 (N_14511,N_11123,N_9445);
or U14512 (N_14512,N_9746,N_9691);
nor U14513 (N_14513,N_10725,N_9939);
nor U14514 (N_14514,N_10876,N_10511);
and U14515 (N_14515,N_9962,N_10883);
and U14516 (N_14516,N_10136,N_9140);
nand U14517 (N_14517,N_11682,N_10602);
or U14518 (N_14518,N_10607,N_10804);
nand U14519 (N_14519,N_10988,N_9185);
and U14520 (N_14520,N_11367,N_9658);
or U14521 (N_14521,N_11689,N_9786);
and U14522 (N_14522,N_11785,N_10948);
or U14523 (N_14523,N_10151,N_10217);
or U14524 (N_14524,N_9755,N_11772);
nor U14525 (N_14525,N_9088,N_10306);
or U14526 (N_14526,N_10585,N_9453);
nand U14527 (N_14527,N_10494,N_10084);
nand U14528 (N_14528,N_10648,N_10480);
nand U14529 (N_14529,N_9850,N_9884);
nor U14530 (N_14530,N_10002,N_10312);
and U14531 (N_14531,N_9625,N_9003);
and U14532 (N_14532,N_10376,N_11210);
nand U14533 (N_14533,N_10861,N_9022);
and U14534 (N_14534,N_11635,N_11424);
and U14535 (N_14535,N_11743,N_11887);
nor U14536 (N_14536,N_11166,N_10367);
nor U14537 (N_14537,N_10874,N_9831);
or U14538 (N_14538,N_11070,N_11497);
xnor U14539 (N_14539,N_9179,N_9285);
or U14540 (N_14540,N_11329,N_11527);
xnor U14541 (N_14541,N_11618,N_11041);
nor U14542 (N_14542,N_9579,N_10471);
or U14543 (N_14543,N_10396,N_9637);
or U14544 (N_14544,N_9557,N_10368);
nor U14545 (N_14545,N_11577,N_10296);
nand U14546 (N_14546,N_10340,N_9202);
and U14547 (N_14547,N_9589,N_9788);
and U14548 (N_14548,N_11322,N_11079);
or U14549 (N_14549,N_9752,N_11708);
or U14550 (N_14550,N_10043,N_9499);
nor U14551 (N_14551,N_10700,N_9391);
nor U14552 (N_14552,N_9942,N_11000);
nor U14553 (N_14553,N_10149,N_9325);
nand U14554 (N_14554,N_10039,N_10936);
xor U14555 (N_14555,N_10879,N_10392);
nor U14556 (N_14556,N_10529,N_11575);
xnor U14557 (N_14557,N_9219,N_10224);
or U14558 (N_14558,N_9598,N_9101);
and U14559 (N_14559,N_10064,N_11519);
nor U14560 (N_14560,N_10165,N_11116);
and U14561 (N_14561,N_9807,N_11333);
and U14562 (N_14562,N_9849,N_10417);
and U14563 (N_14563,N_11946,N_10735);
nor U14564 (N_14564,N_9402,N_11294);
or U14565 (N_14565,N_10001,N_9115);
and U14566 (N_14566,N_10990,N_10159);
and U14567 (N_14567,N_11106,N_10742);
xnor U14568 (N_14568,N_10969,N_9598);
xor U14569 (N_14569,N_9218,N_10028);
nand U14570 (N_14570,N_11837,N_10399);
nor U14571 (N_14571,N_9651,N_9722);
or U14572 (N_14572,N_10010,N_10116);
nand U14573 (N_14573,N_11251,N_9983);
xor U14574 (N_14574,N_11948,N_9507);
and U14575 (N_14575,N_11908,N_9118);
or U14576 (N_14576,N_10311,N_10595);
nor U14577 (N_14577,N_10952,N_11568);
nand U14578 (N_14578,N_10880,N_9572);
nand U14579 (N_14579,N_9256,N_10062);
nor U14580 (N_14580,N_9837,N_10277);
or U14581 (N_14581,N_10431,N_11723);
nor U14582 (N_14582,N_9511,N_9238);
nor U14583 (N_14583,N_10068,N_11895);
nor U14584 (N_14584,N_9220,N_9992);
or U14585 (N_14585,N_9909,N_10423);
or U14586 (N_14586,N_9934,N_10501);
nor U14587 (N_14587,N_11154,N_9995);
or U14588 (N_14588,N_9748,N_11783);
nor U14589 (N_14589,N_11206,N_11081);
nor U14590 (N_14590,N_10090,N_11036);
and U14591 (N_14591,N_9300,N_9614);
nand U14592 (N_14592,N_11179,N_11908);
or U14593 (N_14593,N_11174,N_11085);
and U14594 (N_14594,N_9443,N_11489);
and U14595 (N_14595,N_10363,N_11050);
xor U14596 (N_14596,N_9905,N_10323);
and U14597 (N_14597,N_9476,N_11723);
or U14598 (N_14598,N_10944,N_10976);
and U14599 (N_14599,N_11050,N_11414);
nor U14600 (N_14600,N_9613,N_10014);
or U14601 (N_14601,N_9580,N_10088);
nor U14602 (N_14602,N_10289,N_9180);
and U14603 (N_14603,N_9552,N_11402);
or U14604 (N_14604,N_10003,N_9234);
and U14605 (N_14605,N_11540,N_9605);
nand U14606 (N_14606,N_10200,N_11289);
xor U14607 (N_14607,N_9422,N_11949);
nand U14608 (N_14608,N_11310,N_11860);
or U14609 (N_14609,N_9785,N_10800);
nand U14610 (N_14610,N_10402,N_9925);
and U14611 (N_14611,N_9066,N_11577);
nand U14612 (N_14612,N_10274,N_9828);
nor U14613 (N_14613,N_9617,N_10737);
or U14614 (N_14614,N_10299,N_9398);
nand U14615 (N_14615,N_11976,N_11591);
and U14616 (N_14616,N_10587,N_9304);
nor U14617 (N_14617,N_11316,N_11640);
nand U14618 (N_14618,N_10973,N_11849);
nand U14619 (N_14619,N_9739,N_11966);
and U14620 (N_14620,N_11572,N_9977);
xnor U14621 (N_14621,N_9899,N_11697);
xor U14622 (N_14622,N_11715,N_9295);
or U14623 (N_14623,N_9843,N_9205);
or U14624 (N_14624,N_10700,N_9322);
and U14625 (N_14625,N_10585,N_10474);
or U14626 (N_14626,N_9453,N_9038);
or U14627 (N_14627,N_11844,N_11169);
and U14628 (N_14628,N_10067,N_11993);
or U14629 (N_14629,N_9978,N_10662);
nor U14630 (N_14630,N_10102,N_10632);
or U14631 (N_14631,N_11849,N_11698);
nor U14632 (N_14632,N_10257,N_10837);
nand U14633 (N_14633,N_11612,N_9179);
and U14634 (N_14634,N_11036,N_10150);
nor U14635 (N_14635,N_9692,N_11577);
and U14636 (N_14636,N_10103,N_10763);
nand U14637 (N_14637,N_9141,N_11450);
xor U14638 (N_14638,N_11997,N_11679);
nor U14639 (N_14639,N_10907,N_10059);
or U14640 (N_14640,N_9528,N_9930);
or U14641 (N_14641,N_11949,N_11648);
nor U14642 (N_14642,N_9523,N_9683);
nand U14643 (N_14643,N_10654,N_11702);
or U14644 (N_14644,N_10779,N_10789);
and U14645 (N_14645,N_10756,N_11116);
and U14646 (N_14646,N_10586,N_9417);
nand U14647 (N_14647,N_10988,N_9013);
or U14648 (N_14648,N_10988,N_10596);
and U14649 (N_14649,N_10223,N_11349);
and U14650 (N_14650,N_11390,N_9194);
nand U14651 (N_14651,N_9873,N_9621);
and U14652 (N_14652,N_10219,N_11093);
nand U14653 (N_14653,N_9691,N_9864);
or U14654 (N_14654,N_11213,N_10651);
nand U14655 (N_14655,N_11092,N_11379);
and U14656 (N_14656,N_9063,N_11431);
nand U14657 (N_14657,N_11615,N_11514);
nand U14658 (N_14658,N_10001,N_11345);
and U14659 (N_14659,N_10225,N_10363);
or U14660 (N_14660,N_10985,N_11857);
xnor U14661 (N_14661,N_10654,N_11581);
nor U14662 (N_14662,N_11093,N_11544);
or U14663 (N_14663,N_10384,N_9116);
nor U14664 (N_14664,N_10618,N_9033);
xor U14665 (N_14665,N_9843,N_11346);
or U14666 (N_14666,N_11091,N_9665);
nand U14667 (N_14667,N_9346,N_9984);
and U14668 (N_14668,N_9839,N_10351);
or U14669 (N_14669,N_9383,N_11194);
or U14670 (N_14670,N_9610,N_11763);
nor U14671 (N_14671,N_10479,N_11728);
xnor U14672 (N_14672,N_9422,N_11725);
and U14673 (N_14673,N_10418,N_11009);
nor U14674 (N_14674,N_9882,N_9750);
nand U14675 (N_14675,N_10191,N_9489);
or U14676 (N_14676,N_9741,N_10096);
nand U14677 (N_14677,N_10787,N_11740);
xor U14678 (N_14678,N_11693,N_11966);
nand U14679 (N_14679,N_11246,N_9587);
and U14680 (N_14680,N_11721,N_10668);
nor U14681 (N_14681,N_10177,N_9823);
or U14682 (N_14682,N_10531,N_9184);
and U14683 (N_14683,N_11981,N_9176);
or U14684 (N_14684,N_10880,N_10475);
xnor U14685 (N_14685,N_9165,N_9315);
and U14686 (N_14686,N_10551,N_10675);
and U14687 (N_14687,N_10534,N_9340);
and U14688 (N_14688,N_11780,N_11885);
nand U14689 (N_14689,N_9658,N_10339);
or U14690 (N_14690,N_10176,N_11698);
and U14691 (N_14691,N_10891,N_10744);
nand U14692 (N_14692,N_9190,N_11750);
and U14693 (N_14693,N_11412,N_11176);
or U14694 (N_14694,N_11092,N_9217);
nand U14695 (N_14695,N_10296,N_9125);
nor U14696 (N_14696,N_9182,N_9110);
nor U14697 (N_14697,N_9267,N_10387);
nand U14698 (N_14698,N_10010,N_9736);
nand U14699 (N_14699,N_11511,N_11409);
and U14700 (N_14700,N_9825,N_10053);
nor U14701 (N_14701,N_11367,N_9074);
nor U14702 (N_14702,N_11787,N_10596);
nor U14703 (N_14703,N_9732,N_11601);
or U14704 (N_14704,N_9814,N_9522);
nor U14705 (N_14705,N_11009,N_11354);
or U14706 (N_14706,N_10024,N_10383);
nand U14707 (N_14707,N_11004,N_11945);
and U14708 (N_14708,N_11987,N_10166);
nor U14709 (N_14709,N_11700,N_11364);
nor U14710 (N_14710,N_9977,N_11379);
nand U14711 (N_14711,N_11356,N_10890);
nor U14712 (N_14712,N_10829,N_11133);
nand U14713 (N_14713,N_11837,N_10631);
nor U14714 (N_14714,N_11238,N_11094);
nand U14715 (N_14715,N_11500,N_9890);
and U14716 (N_14716,N_9253,N_11855);
and U14717 (N_14717,N_11597,N_9054);
or U14718 (N_14718,N_11664,N_10303);
nor U14719 (N_14719,N_10033,N_10979);
nor U14720 (N_14720,N_10777,N_9972);
nand U14721 (N_14721,N_9449,N_9286);
nand U14722 (N_14722,N_9505,N_9808);
and U14723 (N_14723,N_10751,N_9436);
nor U14724 (N_14724,N_10117,N_11409);
or U14725 (N_14725,N_10073,N_11540);
xnor U14726 (N_14726,N_11458,N_9303);
and U14727 (N_14727,N_10810,N_11570);
nor U14728 (N_14728,N_10979,N_9986);
or U14729 (N_14729,N_11606,N_10512);
nor U14730 (N_14730,N_9680,N_10795);
or U14731 (N_14731,N_9707,N_10036);
xnor U14732 (N_14732,N_10149,N_11549);
nor U14733 (N_14733,N_10195,N_10703);
nor U14734 (N_14734,N_11767,N_11609);
or U14735 (N_14735,N_9240,N_9417);
nand U14736 (N_14736,N_10516,N_11826);
nand U14737 (N_14737,N_9062,N_11398);
nand U14738 (N_14738,N_11971,N_10291);
nor U14739 (N_14739,N_10240,N_10223);
nor U14740 (N_14740,N_9637,N_11258);
and U14741 (N_14741,N_11091,N_9961);
nand U14742 (N_14742,N_11035,N_11585);
nand U14743 (N_14743,N_10853,N_11803);
or U14744 (N_14744,N_10193,N_10351);
and U14745 (N_14745,N_10492,N_9782);
and U14746 (N_14746,N_11490,N_10960);
or U14747 (N_14747,N_10167,N_10019);
or U14748 (N_14748,N_10071,N_10529);
or U14749 (N_14749,N_10094,N_10630);
and U14750 (N_14750,N_9661,N_11803);
nand U14751 (N_14751,N_9236,N_11570);
xor U14752 (N_14752,N_9783,N_9900);
or U14753 (N_14753,N_10395,N_10773);
and U14754 (N_14754,N_11510,N_9739);
xnor U14755 (N_14755,N_9445,N_9203);
or U14756 (N_14756,N_11227,N_11864);
or U14757 (N_14757,N_10073,N_10211);
xor U14758 (N_14758,N_9768,N_9920);
or U14759 (N_14759,N_10616,N_9956);
nand U14760 (N_14760,N_11272,N_10892);
or U14761 (N_14761,N_9381,N_10536);
and U14762 (N_14762,N_10587,N_9059);
and U14763 (N_14763,N_9404,N_11427);
nor U14764 (N_14764,N_9865,N_9576);
nand U14765 (N_14765,N_11009,N_10932);
or U14766 (N_14766,N_9958,N_11314);
or U14767 (N_14767,N_11756,N_11244);
or U14768 (N_14768,N_10079,N_9639);
and U14769 (N_14769,N_11457,N_11256);
or U14770 (N_14770,N_11357,N_11044);
nand U14771 (N_14771,N_10958,N_9969);
nand U14772 (N_14772,N_9586,N_11555);
nor U14773 (N_14773,N_10097,N_10912);
nor U14774 (N_14774,N_10480,N_11697);
nor U14775 (N_14775,N_11123,N_11934);
or U14776 (N_14776,N_11188,N_9269);
and U14777 (N_14777,N_10936,N_9870);
and U14778 (N_14778,N_11916,N_9339);
xor U14779 (N_14779,N_11371,N_10812);
nand U14780 (N_14780,N_11685,N_10308);
xor U14781 (N_14781,N_11708,N_11729);
nand U14782 (N_14782,N_11433,N_9755);
or U14783 (N_14783,N_9427,N_10066);
nand U14784 (N_14784,N_10087,N_11062);
nor U14785 (N_14785,N_11562,N_10807);
and U14786 (N_14786,N_10937,N_11821);
nand U14787 (N_14787,N_10059,N_9209);
or U14788 (N_14788,N_9879,N_9432);
or U14789 (N_14789,N_11953,N_10906);
or U14790 (N_14790,N_11616,N_10853);
and U14791 (N_14791,N_11963,N_10743);
or U14792 (N_14792,N_9165,N_10750);
nor U14793 (N_14793,N_11958,N_10880);
or U14794 (N_14794,N_11120,N_11718);
nand U14795 (N_14795,N_10649,N_11006);
xnor U14796 (N_14796,N_9369,N_9298);
and U14797 (N_14797,N_11431,N_11906);
and U14798 (N_14798,N_10092,N_9843);
or U14799 (N_14799,N_9532,N_11598);
and U14800 (N_14800,N_10824,N_10351);
or U14801 (N_14801,N_10540,N_9632);
and U14802 (N_14802,N_10317,N_10712);
and U14803 (N_14803,N_11521,N_11926);
nand U14804 (N_14804,N_10154,N_11085);
nor U14805 (N_14805,N_9465,N_10658);
xor U14806 (N_14806,N_10343,N_11934);
nand U14807 (N_14807,N_9381,N_9937);
and U14808 (N_14808,N_9641,N_10328);
nor U14809 (N_14809,N_11167,N_9478);
nand U14810 (N_14810,N_11761,N_10918);
nand U14811 (N_14811,N_11791,N_10897);
and U14812 (N_14812,N_11471,N_10046);
xnor U14813 (N_14813,N_10549,N_9415);
nor U14814 (N_14814,N_9612,N_10094);
xor U14815 (N_14815,N_11795,N_11957);
or U14816 (N_14816,N_10955,N_9240);
nor U14817 (N_14817,N_10395,N_11388);
nand U14818 (N_14818,N_9868,N_11667);
nand U14819 (N_14819,N_9769,N_10671);
or U14820 (N_14820,N_9409,N_11327);
or U14821 (N_14821,N_10678,N_9326);
or U14822 (N_14822,N_10314,N_9864);
or U14823 (N_14823,N_10037,N_10560);
or U14824 (N_14824,N_11432,N_9600);
nor U14825 (N_14825,N_9654,N_9731);
nand U14826 (N_14826,N_11786,N_9010);
or U14827 (N_14827,N_9631,N_10590);
and U14828 (N_14828,N_9539,N_10428);
nor U14829 (N_14829,N_9478,N_9618);
or U14830 (N_14830,N_10701,N_11842);
nand U14831 (N_14831,N_10939,N_10933);
and U14832 (N_14832,N_9435,N_11658);
or U14833 (N_14833,N_9363,N_9262);
and U14834 (N_14834,N_10159,N_9213);
nand U14835 (N_14835,N_9730,N_10545);
xor U14836 (N_14836,N_10028,N_9326);
and U14837 (N_14837,N_11562,N_11425);
and U14838 (N_14838,N_9276,N_11023);
and U14839 (N_14839,N_11705,N_10573);
xnor U14840 (N_14840,N_9468,N_9555);
or U14841 (N_14841,N_9628,N_10388);
or U14842 (N_14842,N_9653,N_10635);
nand U14843 (N_14843,N_9458,N_9572);
and U14844 (N_14844,N_9232,N_9602);
nand U14845 (N_14845,N_11690,N_11979);
or U14846 (N_14846,N_11699,N_11323);
nand U14847 (N_14847,N_11008,N_10072);
nand U14848 (N_14848,N_11942,N_9633);
and U14849 (N_14849,N_11688,N_11602);
or U14850 (N_14850,N_9523,N_9456);
or U14851 (N_14851,N_10659,N_9804);
and U14852 (N_14852,N_10889,N_11619);
or U14853 (N_14853,N_10586,N_10619);
nor U14854 (N_14854,N_11929,N_9031);
nor U14855 (N_14855,N_10445,N_11236);
and U14856 (N_14856,N_10641,N_10734);
nor U14857 (N_14857,N_11803,N_10429);
nor U14858 (N_14858,N_10588,N_11115);
or U14859 (N_14859,N_11651,N_9651);
nor U14860 (N_14860,N_11133,N_9172);
nand U14861 (N_14861,N_10783,N_9540);
xnor U14862 (N_14862,N_10123,N_9785);
and U14863 (N_14863,N_10755,N_9431);
or U14864 (N_14864,N_9266,N_10933);
nand U14865 (N_14865,N_11493,N_11230);
nor U14866 (N_14866,N_11392,N_10612);
nand U14867 (N_14867,N_9411,N_11599);
nor U14868 (N_14868,N_9415,N_9411);
nor U14869 (N_14869,N_10123,N_11081);
or U14870 (N_14870,N_11776,N_10208);
xor U14871 (N_14871,N_10724,N_10094);
and U14872 (N_14872,N_11410,N_11389);
or U14873 (N_14873,N_11992,N_10994);
nand U14874 (N_14874,N_9382,N_9820);
and U14875 (N_14875,N_9066,N_9609);
nand U14876 (N_14876,N_9531,N_9340);
or U14877 (N_14877,N_9961,N_9089);
and U14878 (N_14878,N_9717,N_9827);
or U14879 (N_14879,N_11183,N_11742);
or U14880 (N_14880,N_10666,N_10140);
or U14881 (N_14881,N_9077,N_11324);
nand U14882 (N_14882,N_11959,N_11681);
nor U14883 (N_14883,N_9268,N_9320);
or U14884 (N_14884,N_11664,N_9572);
xnor U14885 (N_14885,N_11620,N_11042);
or U14886 (N_14886,N_11284,N_10900);
xor U14887 (N_14887,N_9805,N_10148);
and U14888 (N_14888,N_10271,N_11666);
and U14889 (N_14889,N_9217,N_11889);
and U14890 (N_14890,N_10059,N_11825);
nand U14891 (N_14891,N_10179,N_11187);
or U14892 (N_14892,N_11131,N_9479);
or U14893 (N_14893,N_10831,N_11306);
nand U14894 (N_14894,N_10285,N_9975);
xor U14895 (N_14895,N_9512,N_10499);
nor U14896 (N_14896,N_11978,N_9403);
and U14897 (N_14897,N_10794,N_11484);
and U14898 (N_14898,N_11762,N_9708);
nand U14899 (N_14899,N_9010,N_10509);
or U14900 (N_14900,N_10391,N_10078);
nor U14901 (N_14901,N_10084,N_10419);
and U14902 (N_14902,N_11537,N_9991);
xnor U14903 (N_14903,N_11376,N_9407);
nor U14904 (N_14904,N_9510,N_9384);
nand U14905 (N_14905,N_11873,N_10840);
or U14906 (N_14906,N_9464,N_10728);
or U14907 (N_14907,N_11370,N_10689);
or U14908 (N_14908,N_10974,N_10929);
or U14909 (N_14909,N_11500,N_10942);
nor U14910 (N_14910,N_10108,N_11224);
or U14911 (N_14911,N_11405,N_11097);
and U14912 (N_14912,N_9050,N_10885);
and U14913 (N_14913,N_10438,N_11357);
or U14914 (N_14914,N_9134,N_9782);
nor U14915 (N_14915,N_9640,N_11776);
and U14916 (N_14916,N_11556,N_9130);
or U14917 (N_14917,N_11075,N_9739);
xor U14918 (N_14918,N_9135,N_11695);
or U14919 (N_14919,N_9401,N_10193);
xor U14920 (N_14920,N_10158,N_9732);
xor U14921 (N_14921,N_11763,N_9219);
nand U14922 (N_14922,N_10927,N_9306);
and U14923 (N_14923,N_10741,N_9559);
nand U14924 (N_14924,N_11043,N_9324);
nor U14925 (N_14925,N_11566,N_10803);
or U14926 (N_14926,N_11958,N_9574);
xnor U14927 (N_14927,N_11723,N_11229);
xnor U14928 (N_14928,N_9044,N_10014);
nand U14929 (N_14929,N_10053,N_11284);
xnor U14930 (N_14930,N_11555,N_9454);
xnor U14931 (N_14931,N_9286,N_11916);
nor U14932 (N_14932,N_10066,N_11125);
nand U14933 (N_14933,N_9098,N_9311);
or U14934 (N_14934,N_9666,N_10354);
nand U14935 (N_14935,N_10256,N_9572);
nand U14936 (N_14936,N_11549,N_10700);
nand U14937 (N_14937,N_11362,N_10211);
nand U14938 (N_14938,N_9253,N_9368);
nor U14939 (N_14939,N_10028,N_9509);
and U14940 (N_14940,N_9424,N_9635);
xor U14941 (N_14941,N_11055,N_9153);
nand U14942 (N_14942,N_11912,N_11625);
nand U14943 (N_14943,N_10372,N_11011);
xnor U14944 (N_14944,N_11500,N_11838);
nand U14945 (N_14945,N_10975,N_11030);
and U14946 (N_14946,N_11866,N_10047);
nor U14947 (N_14947,N_10058,N_10860);
or U14948 (N_14948,N_11980,N_10058);
or U14949 (N_14949,N_9616,N_9960);
or U14950 (N_14950,N_10224,N_11041);
and U14951 (N_14951,N_9348,N_10918);
nand U14952 (N_14952,N_11165,N_9689);
or U14953 (N_14953,N_9223,N_9899);
xor U14954 (N_14954,N_10512,N_9607);
and U14955 (N_14955,N_11807,N_9940);
or U14956 (N_14956,N_9354,N_10123);
and U14957 (N_14957,N_9192,N_9336);
nand U14958 (N_14958,N_10914,N_9182);
and U14959 (N_14959,N_11744,N_9116);
or U14960 (N_14960,N_9211,N_10688);
or U14961 (N_14961,N_11417,N_11789);
xnor U14962 (N_14962,N_10283,N_10484);
nor U14963 (N_14963,N_11898,N_11076);
or U14964 (N_14964,N_11170,N_10467);
nand U14965 (N_14965,N_10012,N_11920);
nand U14966 (N_14966,N_11838,N_10276);
nand U14967 (N_14967,N_11393,N_10423);
or U14968 (N_14968,N_10510,N_9434);
nand U14969 (N_14969,N_11217,N_11583);
or U14970 (N_14970,N_11839,N_11915);
or U14971 (N_14971,N_11356,N_10547);
or U14972 (N_14972,N_11598,N_9062);
nor U14973 (N_14973,N_10018,N_10749);
nor U14974 (N_14974,N_10568,N_9750);
nor U14975 (N_14975,N_9654,N_10588);
and U14976 (N_14976,N_10930,N_10166);
and U14977 (N_14977,N_11274,N_10666);
nand U14978 (N_14978,N_11107,N_11041);
or U14979 (N_14979,N_9026,N_11643);
nand U14980 (N_14980,N_9540,N_11605);
or U14981 (N_14981,N_10742,N_9633);
or U14982 (N_14982,N_9521,N_10392);
nand U14983 (N_14983,N_10408,N_10052);
and U14984 (N_14984,N_11381,N_9249);
nand U14985 (N_14985,N_11210,N_11858);
nor U14986 (N_14986,N_10171,N_9820);
xnor U14987 (N_14987,N_11734,N_9949);
nor U14988 (N_14988,N_10155,N_9275);
nor U14989 (N_14989,N_10132,N_10619);
xor U14990 (N_14990,N_10597,N_9988);
and U14991 (N_14991,N_11679,N_11643);
xor U14992 (N_14992,N_11109,N_10240);
nor U14993 (N_14993,N_9007,N_10292);
nand U14994 (N_14994,N_9811,N_10478);
xor U14995 (N_14995,N_9161,N_9071);
nand U14996 (N_14996,N_11743,N_11704);
or U14997 (N_14997,N_10435,N_11375);
and U14998 (N_14998,N_10155,N_10801);
or U14999 (N_14999,N_10026,N_9720);
and UO_0 (O_0,N_14604,N_14268);
and UO_1 (O_1,N_14500,N_13372);
and UO_2 (O_2,N_12631,N_13619);
and UO_3 (O_3,N_12037,N_12031);
xor UO_4 (O_4,N_12465,N_13587);
and UO_5 (O_5,N_13633,N_14985);
nand UO_6 (O_6,N_13919,N_14719);
or UO_7 (O_7,N_14889,N_12416);
nand UO_8 (O_8,N_13858,N_14409);
nand UO_9 (O_9,N_14063,N_12119);
and UO_10 (O_10,N_14159,N_14521);
and UO_11 (O_11,N_12346,N_13037);
and UO_12 (O_12,N_14216,N_14878);
nor UO_13 (O_13,N_14304,N_12920);
and UO_14 (O_14,N_12514,N_14145);
nand UO_15 (O_15,N_12134,N_12055);
and UO_16 (O_16,N_12138,N_13747);
or UO_17 (O_17,N_14323,N_13398);
nand UO_18 (O_18,N_13833,N_14242);
or UO_19 (O_19,N_12802,N_12110);
xor UO_20 (O_20,N_13639,N_13750);
xnor UO_21 (O_21,N_13048,N_13681);
nor UO_22 (O_22,N_12361,N_12438);
xnor UO_23 (O_23,N_12641,N_13455);
or UO_24 (O_24,N_12670,N_12358);
nand UO_25 (O_25,N_12863,N_12790);
and UO_26 (O_26,N_14493,N_14096);
nor UO_27 (O_27,N_12902,N_14948);
or UO_28 (O_28,N_14142,N_12196);
or UO_29 (O_29,N_14205,N_13056);
and UO_30 (O_30,N_14025,N_13964);
nor UO_31 (O_31,N_13551,N_13796);
and UO_32 (O_32,N_12407,N_13780);
and UO_33 (O_33,N_12314,N_14415);
and UO_34 (O_34,N_14263,N_13617);
or UO_35 (O_35,N_12972,N_14672);
nor UO_36 (O_36,N_12447,N_13898);
and UO_37 (O_37,N_13189,N_12728);
and UO_38 (O_38,N_12461,N_12370);
and UO_39 (O_39,N_13277,N_14586);
and UO_40 (O_40,N_14450,N_13343);
nor UO_41 (O_41,N_14937,N_13176);
and UO_42 (O_42,N_13351,N_14964);
nor UO_43 (O_43,N_14193,N_14869);
nand UO_44 (O_44,N_12477,N_13443);
and UO_45 (O_45,N_13230,N_14087);
nor UO_46 (O_46,N_13640,N_13427);
nor UO_47 (O_47,N_13506,N_14720);
nor UO_48 (O_48,N_14446,N_12486);
nor UO_49 (O_49,N_13549,N_14747);
or UO_50 (O_50,N_12455,N_13144);
nand UO_51 (O_51,N_14234,N_12418);
and UO_52 (O_52,N_13843,N_13799);
and UO_53 (O_53,N_13305,N_14297);
or UO_54 (O_54,N_14452,N_14749);
nor UO_55 (O_55,N_12924,N_13872);
or UO_56 (O_56,N_14210,N_12703);
or UO_57 (O_57,N_12056,N_14111);
and UO_58 (O_58,N_13870,N_12483);
and UO_59 (O_59,N_13622,N_13771);
and UO_60 (O_60,N_14480,N_14845);
and UO_61 (O_61,N_14814,N_13378);
and UO_62 (O_62,N_14295,N_12843);
nor UO_63 (O_63,N_14546,N_14932);
or UO_64 (O_64,N_13560,N_12371);
or UO_65 (O_65,N_13415,N_13270);
nand UO_66 (O_66,N_12946,N_13987);
nand UO_67 (O_67,N_12608,N_12600);
nor UO_68 (O_68,N_14613,N_12554);
nor UO_69 (O_69,N_12998,N_13059);
and UO_70 (O_70,N_14091,N_12649);
nand UO_71 (O_71,N_13786,N_13995);
and UO_72 (O_72,N_13460,N_12406);
xor UO_73 (O_73,N_12300,N_12783);
and UO_74 (O_74,N_12984,N_14543);
nand UO_75 (O_75,N_14614,N_12223);
and UO_76 (O_76,N_14565,N_14013);
nand UO_77 (O_77,N_14507,N_14092);
xor UO_78 (O_78,N_13761,N_14868);
nor UO_79 (O_79,N_14661,N_14300);
nor UO_80 (O_80,N_14527,N_12965);
and UO_81 (O_81,N_12642,N_12870);
or UO_82 (O_82,N_12986,N_14978);
or UO_83 (O_83,N_14417,N_14523);
and UO_84 (O_84,N_13654,N_13718);
and UO_85 (O_85,N_14942,N_13288);
nor UO_86 (O_86,N_12501,N_14681);
nand UO_87 (O_87,N_12516,N_14305);
nor UO_88 (O_88,N_14360,N_14346);
or UO_89 (O_89,N_13135,N_14541);
nor UO_90 (O_90,N_13051,N_14405);
or UO_91 (O_91,N_14775,N_13271);
nor UO_92 (O_92,N_13468,N_14718);
nand UO_93 (O_93,N_13697,N_14441);
or UO_94 (O_94,N_13969,N_14260);
nor UO_95 (O_95,N_12817,N_12759);
or UO_96 (O_96,N_12357,N_12680);
nand UO_97 (O_97,N_14435,N_12372);
nor UO_98 (O_98,N_14572,N_12154);
nand UO_99 (O_99,N_14605,N_13322);
nor UO_100 (O_100,N_12704,N_14017);
or UO_101 (O_101,N_13211,N_13340);
and UO_102 (O_102,N_12212,N_12456);
and UO_103 (O_103,N_14075,N_14684);
or UO_104 (O_104,N_12498,N_13347);
and UO_105 (O_105,N_13708,N_12412);
and UO_106 (O_106,N_13118,N_12927);
and UO_107 (O_107,N_12257,N_14161);
nor UO_108 (O_108,N_12356,N_14199);
nor UO_109 (O_109,N_13132,N_13483);
and UO_110 (O_110,N_13970,N_12235);
or UO_111 (O_111,N_12127,N_12743);
xor UO_112 (O_112,N_13156,N_13294);
nor UO_113 (O_113,N_12682,N_12744);
nand UO_114 (O_114,N_14174,N_13912);
nand UO_115 (O_115,N_12240,N_13044);
nand UO_116 (O_116,N_14739,N_14080);
or UO_117 (O_117,N_12029,N_13553);
nor UO_118 (O_118,N_13717,N_13744);
or UO_119 (O_119,N_13104,N_14921);
nor UO_120 (O_120,N_14428,N_12145);
nand UO_121 (O_121,N_14813,N_12316);
nor UO_122 (O_122,N_13171,N_12512);
and UO_123 (O_123,N_13451,N_12643);
or UO_124 (O_124,N_14781,N_14952);
and UO_125 (O_125,N_13143,N_12878);
or UO_126 (O_126,N_13857,N_14959);
nand UO_127 (O_127,N_13349,N_12312);
xnor UO_128 (O_128,N_12260,N_14862);
or UO_129 (O_129,N_12667,N_12030);
nor UO_130 (O_130,N_14812,N_14197);
nand UO_131 (O_131,N_13173,N_12176);
and UO_132 (O_132,N_13660,N_12933);
nor UO_133 (O_133,N_13330,N_13107);
nand UO_134 (O_134,N_13971,N_14352);
nand UO_135 (O_135,N_14476,N_14120);
nor UO_136 (O_136,N_14946,N_14423);
or UO_137 (O_137,N_13213,N_12915);
xor UO_138 (O_138,N_14916,N_13784);
xnor UO_139 (O_139,N_12202,N_13810);
nor UO_140 (O_140,N_12849,N_14461);
nand UO_141 (O_141,N_12094,N_14807);
or UO_142 (O_142,N_13689,N_13982);
nor UO_143 (O_143,N_14036,N_12228);
nor UO_144 (O_144,N_14686,N_12846);
or UO_145 (O_145,N_13653,N_14756);
or UO_146 (O_146,N_14420,N_14855);
and UO_147 (O_147,N_14628,N_13975);
nor UO_148 (O_148,N_13325,N_12873);
nor UO_149 (O_149,N_12023,N_14490);
or UO_150 (O_150,N_13223,N_13576);
or UO_151 (O_151,N_12135,N_13000);
nor UO_152 (O_152,N_13986,N_14930);
or UO_153 (O_153,N_12190,N_12085);
nand UO_154 (O_154,N_14588,N_13563);
nor UO_155 (O_155,N_12877,N_13245);
nand UO_156 (O_156,N_12114,N_14341);
or UO_157 (O_157,N_12285,N_14678);
and UO_158 (O_158,N_13848,N_13863);
nand UO_159 (O_159,N_13400,N_13880);
or UO_160 (O_160,N_13019,N_14540);
and UO_161 (O_161,N_13678,N_12570);
and UO_162 (O_162,N_14357,N_14047);
and UO_163 (O_163,N_14806,N_14129);
or UO_164 (O_164,N_14859,N_14671);
and UO_165 (O_165,N_12875,N_13184);
nand UO_166 (O_166,N_14679,N_14503);
and UO_167 (O_167,N_14645,N_14574);
nor UO_168 (O_168,N_13268,N_13536);
nor UO_169 (O_169,N_14625,N_12695);
nor UO_170 (O_170,N_14282,N_13357);
nor UO_171 (O_171,N_14976,N_12754);
and UO_172 (O_172,N_13824,N_13578);
and UO_173 (O_173,N_14848,N_12651);
or UO_174 (O_174,N_12468,N_13169);
nand UO_175 (O_175,N_13258,N_14416);
nand UO_176 (O_176,N_12921,N_14984);
xor UO_177 (O_177,N_14289,N_13494);
nand UO_178 (O_178,N_12320,N_14750);
xor UO_179 (O_179,N_14391,N_12018);
xor UO_180 (O_180,N_12130,N_14024);
and UO_181 (O_181,N_14861,N_14912);
nor UO_182 (O_182,N_14832,N_14641);
nand UO_183 (O_183,N_13229,N_12237);
and UO_184 (O_184,N_12241,N_14674);
and UO_185 (O_185,N_14436,N_12658);
or UO_186 (O_186,N_13055,N_12051);
or UO_187 (O_187,N_12277,N_14113);
nand UO_188 (O_188,N_12052,N_12479);
nand UO_189 (O_189,N_12059,N_13826);
nor UO_190 (O_190,N_12671,N_12463);
nand UO_191 (O_191,N_14669,N_13785);
nand UO_192 (O_192,N_14783,N_12497);
nand UO_193 (O_193,N_14876,N_12839);
xnor UO_194 (O_194,N_12229,N_13136);
nand UO_195 (O_195,N_13374,N_12753);
and UO_196 (O_196,N_13170,N_12601);
nand UO_197 (O_197,N_14421,N_13484);
or UO_198 (O_198,N_13387,N_12307);
and UO_199 (O_199,N_13803,N_13196);
xnor UO_200 (O_200,N_12340,N_13428);
and UO_201 (O_201,N_13083,N_12204);
nor UO_202 (O_202,N_14284,N_12916);
nor UO_203 (O_203,N_12719,N_12978);
nand UO_204 (O_204,N_13839,N_14779);
or UO_205 (O_205,N_12354,N_14817);
xnor UO_206 (O_206,N_12113,N_14518);
and UO_207 (O_207,N_13666,N_13525);
nand UO_208 (O_208,N_14240,N_13462);
xnor UO_209 (O_209,N_12171,N_14164);
and UO_210 (O_210,N_14255,N_13187);
nor UO_211 (O_211,N_13237,N_12015);
nor UO_212 (O_212,N_13557,N_13940);
nand UO_213 (O_213,N_13147,N_14067);
nor UO_214 (O_214,N_13746,N_13221);
nor UO_215 (O_215,N_13172,N_13518);
nor UO_216 (O_216,N_12609,N_14808);
nand UO_217 (O_217,N_13495,N_12689);
nor UO_218 (O_218,N_14156,N_12521);
and UO_219 (O_219,N_12803,N_14973);
or UO_220 (O_220,N_14874,N_14371);
nor UO_221 (O_221,N_12355,N_14902);
or UO_222 (O_222,N_13045,N_12768);
xnor UO_223 (O_223,N_12861,N_14955);
and UO_224 (O_224,N_13657,N_12390);
nand UO_225 (O_225,N_14636,N_13238);
nor UO_226 (O_226,N_14922,N_14189);
or UO_227 (O_227,N_12112,N_13847);
nand UO_228 (O_228,N_12931,N_14597);
nor UO_229 (O_229,N_12076,N_13269);
nor UO_230 (O_230,N_12188,N_13684);
nand UO_231 (O_231,N_14451,N_14584);
or UO_232 (O_232,N_12304,N_13099);
xnor UO_233 (O_233,N_13508,N_13683);
nand UO_234 (O_234,N_12969,N_13737);
nand UO_235 (O_235,N_14851,N_14481);
and UO_236 (O_236,N_13155,N_14603);
nor UO_237 (O_237,N_12540,N_14175);
and UO_238 (O_238,N_12505,N_12777);
nand UO_239 (O_239,N_13859,N_13797);
and UO_240 (O_240,N_14342,N_14000);
nand UO_241 (O_241,N_13485,N_13084);
or UO_242 (O_242,N_12904,N_13119);
nor UO_243 (O_243,N_12057,N_12940);
or UO_244 (O_244,N_12218,N_13758);
nor UO_245 (O_245,N_13868,N_13405);
nand UO_246 (O_246,N_12611,N_14638);
nand UO_247 (O_247,N_12518,N_13193);
and UO_248 (O_248,N_13822,N_12458);
nor UO_249 (O_249,N_13649,N_13539);
nor UO_250 (O_250,N_14012,N_13113);
and UO_251 (O_251,N_13738,N_12276);
and UO_252 (O_252,N_14600,N_12795);
nand UO_253 (O_253,N_13191,N_14666);
nand UO_254 (O_254,N_14691,N_14362);
xnor UO_255 (O_255,N_13130,N_14366);
nor UO_256 (O_256,N_13958,N_14022);
or UO_257 (O_257,N_12879,N_13673);
nand UO_258 (O_258,N_14810,N_12733);
nand UO_259 (O_259,N_14953,N_12441);
nand UO_260 (O_260,N_13634,N_13150);
nand UO_261 (O_261,N_13441,N_12367);
nor UO_262 (O_262,N_13556,N_12131);
and UO_263 (O_263,N_13167,N_14052);
nor UO_264 (O_264,N_13032,N_14350);
nor UO_265 (O_265,N_12886,N_14270);
nor UO_266 (O_266,N_14777,N_13181);
nand UO_267 (O_267,N_14760,N_13984);
or UO_268 (O_268,N_13205,N_12003);
nand UO_269 (O_269,N_14787,N_12216);
or UO_270 (O_270,N_12149,N_12325);
or UO_271 (O_271,N_13475,N_12097);
xnor UO_272 (O_272,N_14738,N_14339);
and UO_273 (O_273,N_12413,N_14183);
nand UO_274 (O_274,N_13890,N_14979);
nor UO_275 (O_275,N_13403,N_14786);
nor UO_276 (O_276,N_14630,N_13517);
or UO_277 (O_277,N_14867,N_12368);
and UO_278 (O_278,N_14085,N_12928);
and UO_279 (O_279,N_13088,N_12061);
and UO_280 (O_280,N_14384,N_14517);
nand UO_281 (O_281,N_14338,N_14103);
nand UO_282 (O_282,N_13179,N_12645);
or UO_283 (O_283,N_13310,N_14485);
and UO_284 (O_284,N_13770,N_12930);
or UO_285 (O_285,N_14078,N_12952);
and UO_286 (O_286,N_14139,N_13935);
nor UO_287 (O_287,N_12360,N_13909);
or UO_288 (O_288,N_14892,N_14020);
xnor UO_289 (O_289,N_14019,N_13470);
nor UO_290 (O_290,N_13510,N_13605);
nor UO_291 (O_291,N_12905,N_12382);
nand UO_292 (O_292,N_12823,N_12289);
or UO_293 (O_293,N_12583,N_13411);
or UO_294 (O_294,N_12122,N_12079);
nor UO_295 (O_295,N_13532,N_13162);
and UO_296 (O_296,N_12250,N_13543);
nand UO_297 (O_297,N_14722,N_12578);
or UO_298 (O_298,N_13389,N_12353);
and UO_299 (O_299,N_14727,N_13233);
nand UO_300 (O_300,N_13243,N_13203);
nor UO_301 (O_301,N_14533,N_12948);
and UO_302 (O_302,N_14884,N_14254);
nand UO_303 (O_303,N_13390,N_13137);
nor UO_304 (O_304,N_12396,N_12071);
nand UO_305 (O_305,N_13953,N_14336);
and UO_306 (O_306,N_14796,N_14150);
or UO_307 (O_307,N_13877,N_14181);
and UO_308 (O_308,N_14689,N_14321);
nand UO_309 (O_309,N_12837,N_12748);
nor UO_310 (O_310,N_12901,N_12894);
or UO_311 (O_311,N_14549,N_13655);
nor UO_312 (O_312,N_14650,N_14140);
nand UO_313 (O_313,N_12747,N_14232);
nor UO_314 (O_314,N_12811,N_12892);
or UO_315 (O_315,N_14007,N_12951);
and UO_316 (O_316,N_12797,N_14882);
and UO_317 (O_317,N_14797,N_14870);
nor UO_318 (O_318,N_12476,N_12918);
nor UO_319 (O_319,N_13377,N_12462);
and UO_320 (O_320,N_14782,N_13814);
and UO_321 (O_321,N_12472,N_14881);
and UO_322 (O_322,N_12214,N_13108);
or UO_323 (O_323,N_13776,N_13600);
nand UO_324 (O_324,N_13727,N_14028);
nor UO_325 (O_325,N_12482,N_13914);
nor UO_326 (O_326,N_13365,N_12552);
or UO_327 (O_327,N_12793,N_12936);
nand UO_328 (O_328,N_12193,N_13285);
and UO_329 (O_329,N_13337,N_12457);
and UO_330 (O_330,N_14179,N_14196);
or UO_331 (O_331,N_13345,N_12246);
and UO_332 (O_332,N_14514,N_14457);
and UO_333 (O_333,N_13125,N_12133);
or UO_334 (O_334,N_14149,N_12439);
or UO_335 (O_335,N_12267,N_12684);
or UO_336 (O_336,N_12323,N_14839);
nor UO_337 (O_337,N_14466,N_13142);
xor UO_338 (O_338,N_12393,N_12640);
and UO_339 (O_339,N_12213,N_14261);
or UO_340 (O_340,N_13547,N_12943);
and UO_341 (O_341,N_14626,N_14072);
nand UO_342 (O_342,N_13936,N_12781);
nand UO_343 (O_343,N_13450,N_13110);
nor UO_344 (O_344,N_12115,N_14909);
nor UO_345 (O_345,N_14692,N_12180);
nand UO_346 (O_346,N_14525,N_13835);
nand UO_347 (O_347,N_12153,N_14236);
nor UO_348 (O_348,N_12173,N_13049);
and UO_349 (O_349,N_14045,N_14492);
xor UO_350 (O_350,N_13502,N_13180);
nor UO_351 (O_351,N_12077,N_14235);
or UO_352 (O_352,N_14475,N_14348);
and UO_353 (O_353,N_13577,N_14253);
xnor UO_354 (O_354,N_14846,N_12495);
nand UO_355 (O_355,N_12132,N_13446);
xnor UO_356 (O_356,N_13628,N_12709);
and UO_357 (O_357,N_13458,N_12401);
and UO_358 (O_358,N_12408,N_12542);
and UO_359 (O_359,N_14136,N_14194);
nand UO_360 (O_360,N_12819,N_14702);
nand UO_361 (O_361,N_12047,N_13231);
and UO_362 (O_362,N_14455,N_14137);
xnor UO_363 (O_363,N_13082,N_12278);
or UO_364 (O_364,N_12100,N_12523);
or UO_365 (O_365,N_13053,N_12624);
xnor UO_366 (O_366,N_12508,N_12898);
or UO_367 (O_367,N_12923,N_12900);
and UO_368 (O_368,N_12021,N_13063);
or UO_369 (O_369,N_13741,N_12752);
and UO_370 (O_370,N_12857,N_14315);
or UO_371 (O_371,N_13615,N_14146);
nor UO_372 (O_372,N_13457,N_14050);
nor UO_373 (O_373,N_14040,N_12243);
nand UO_374 (O_374,N_14249,N_13621);
nor UO_375 (O_375,N_14975,N_13667);
and UO_376 (O_376,N_14033,N_12812);
nor UO_377 (O_377,N_12387,N_14863);
nor UO_378 (O_378,N_13081,N_13521);
and UO_379 (O_379,N_13094,N_14230);
nor UO_380 (O_380,N_13210,N_12226);
or UO_381 (O_381,N_12705,N_14991);
nor UO_382 (O_382,N_14429,N_12259);
nor UO_383 (O_383,N_14318,N_13816);
and UO_384 (O_384,N_13514,N_14322);
nand UO_385 (O_385,N_14073,N_12347);
or UO_386 (O_386,N_14035,N_12075);
or UO_387 (O_387,N_12063,N_14169);
and UO_388 (O_388,N_12268,N_13572);
nand UO_389 (O_389,N_13244,N_13293);
nand UO_390 (O_390,N_12862,N_13735);
or UO_391 (O_391,N_13627,N_12379);
nand UO_392 (O_392,N_14333,N_13752);
and UO_393 (O_393,N_13896,N_14898);
or UO_394 (O_394,N_12573,N_14667);
or UO_395 (O_395,N_14785,N_12872);
nor UO_396 (O_396,N_14585,N_13190);
or UO_397 (O_397,N_12326,N_14462);
or UO_398 (O_398,N_13149,N_12840);
nand UO_399 (O_399,N_13381,N_13906);
nor UO_400 (O_400,N_14377,N_12349);
and UO_401 (O_401,N_12517,N_13492);
or UO_402 (O_402,N_14372,N_14180);
nand UO_403 (O_403,N_13146,N_13674);
nand UO_404 (O_404,N_14997,N_14723);
or UO_405 (O_405,N_14653,N_12263);
or UO_406 (O_406,N_12017,N_14619);
and UO_407 (O_407,N_12687,N_12977);
nor UO_408 (O_408,N_12546,N_13275);
or UO_409 (O_409,N_12919,N_12222);
nor UO_410 (O_410,N_14502,N_12702);
and UO_411 (O_411,N_12086,N_14850);
and UO_412 (O_412,N_13946,N_14097);
and UO_413 (O_413,N_13069,N_13897);
nor UO_414 (O_414,N_13215,N_13421);
or UO_415 (O_415,N_13070,N_12646);
or UO_416 (O_416,N_12588,N_14893);
and UO_417 (O_417,N_12120,N_13817);
or UO_418 (O_418,N_14109,N_14313);
nand UO_419 (O_419,N_13908,N_12502);
and UO_420 (O_420,N_13943,N_13703);
and UO_421 (O_421,N_13133,N_14567);
xnor UO_422 (O_422,N_12853,N_13864);
and UO_423 (O_423,N_14849,N_12869);
nand UO_424 (O_424,N_12039,N_14202);
or UO_425 (O_425,N_14539,N_13422);
and UO_426 (O_426,N_12062,N_13003);
nand UO_427 (O_427,N_13429,N_14675);
nor UO_428 (O_428,N_12435,N_12348);
and UO_429 (O_429,N_14456,N_12524);
or UO_430 (O_430,N_12992,N_12065);
nand UO_431 (O_431,N_13910,N_12906);
or UO_432 (O_432,N_13361,N_12825);
nor UO_433 (O_433,N_12958,N_13881);
or UO_434 (O_434,N_12659,N_14144);
or UO_435 (O_435,N_13740,N_14376);
nand UO_436 (O_436,N_14066,N_12746);
xor UO_437 (O_437,N_14755,N_14542);
nand UO_438 (O_438,N_12574,N_12708);
nand UO_439 (O_439,N_14030,N_13922);
or UO_440 (O_440,N_12549,N_13823);
nor UO_441 (O_441,N_12652,N_14079);
or UO_442 (O_442,N_13961,N_14612);
and UO_443 (O_443,N_12816,N_12108);
and UO_444 (O_444,N_12548,N_13360);
nand UO_445 (O_445,N_13076,N_14238);
nand UO_446 (O_446,N_14206,N_13933);
nor UO_447 (O_447,N_12740,N_14399);
nand UO_448 (O_448,N_12553,N_14448);
nand UO_449 (O_449,N_12866,N_14733);
nand UO_450 (O_450,N_14920,N_13074);
nor UO_451 (O_451,N_12026,N_13296);
and UO_452 (O_452,N_12706,N_14116);
or UO_453 (O_453,N_14647,N_12230);
and UO_454 (O_454,N_14355,N_14496);
and UO_455 (O_455,N_12907,N_13795);
or UO_456 (O_456,N_14617,N_13197);
and UO_457 (O_457,N_14117,N_14660);
or UO_458 (O_458,N_12162,N_12507);
nor UO_459 (O_459,N_14334,N_12398);
nand UO_460 (O_460,N_14463,N_12238);
nor UO_461 (O_461,N_13339,N_13808);
nand UO_462 (O_462,N_12850,N_14217);
xor UO_463 (O_463,N_13449,N_14375);
and UO_464 (O_464,N_14611,N_13208);
or UO_465 (O_465,N_12504,N_12206);
nand UO_466 (O_466,N_12432,N_12625);
nand UO_467 (O_467,N_12765,N_13713);
xor UO_468 (O_468,N_12774,N_13867);
and UO_469 (O_469,N_13767,N_13777);
and UO_470 (O_470,N_12297,N_14425);
or UO_471 (O_471,N_14730,N_14044);
nand UO_472 (O_472,N_12858,N_12815);
nor UO_473 (O_473,N_13386,N_14852);
or UO_474 (O_474,N_13109,N_12178);
nor UO_475 (O_475,N_12156,N_13299);
and UO_476 (O_476,N_14530,N_12606);
and UO_477 (O_477,N_13853,N_14601);
or UO_478 (O_478,N_14726,N_14225);
xor UO_479 (O_479,N_13954,N_12810);
or UO_480 (O_480,N_12536,N_12440);
nor UO_481 (O_481,N_13077,N_12442);
nor UO_482 (O_482,N_12818,N_12696);
nor UO_483 (O_483,N_13103,N_14472);
or UO_484 (O_484,N_13555,N_14830);
and UO_485 (O_485,N_12917,N_13592);
and UO_486 (O_486,N_14844,N_13827);
or UO_487 (O_487,N_12555,N_13682);
nand UO_488 (O_488,N_12616,N_14105);
xnor UO_489 (O_489,N_14519,N_12644);
nor UO_490 (O_490,N_14986,N_13601);
or UO_491 (O_491,N_14776,N_12587);
or UO_492 (O_492,N_14590,N_13175);
or UO_493 (O_493,N_12896,N_13650);
nor UO_494 (O_494,N_14491,N_14387);
and UO_495 (O_495,N_14792,N_14167);
xnor UO_496 (O_496,N_12532,N_13298);
and UO_497 (O_497,N_13590,N_13126);
nor UO_498 (O_498,N_12828,N_12718);
and UO_499 (O_499,N_14215,N_13743);
nand UO_500 (O_500,N_14568,N_13043);
and UO_501 (O_501,N_12184,N_13200);
nand UO_502 (O_502,N_14014,N_13008);
nand UO_503 (O_503,N_13161,N_14258);
nand UO_504 (O_504,N_12591,N_14061);
and UO_505 (O_505,N_14992,N_12690);
nand UO_506 (O_506,N_13861,N_13062);
or UO_507 (O_507,N_13716,N_12205);
or UO_508 (O_508,N_12650,N_12473);
and UO_509 (O_509,N_13134,N_14413);
nor UO_510 (O_510,N_13302,N_14888);
xor UO_511 (O_511,N_14246,N_12107);
or UO_512 (O_512,N_13410,N_14126);
nor UO_513 (O_513,N_12043,N_12851);
nand UO_514 (O_514,N_13105,N_14556);
nand UO_515 (O_515,N_14563,N_13932);
nand UO_516 (O_516,N_14509,N_14743);
and UO_517 (O_517,N_12426,N_14482);
nor UO_518 (O_518,N_14634,N_12807);
and UO_519 (O_519,N_14969,N_13570);
or UO_520 (O_520,N_12451,N_14635);
and UO_521 (O_521,N_12602,N_13362);
nand UO_522 (O_522,N_12050,N_14903);
and UO_523 (O_523,N_12264,N_12971);
nand UO_524 (O_524,N_14982,N_12123);
nor UO_525 (O_525,N_14245,N_14108);
nor UO_526 (O_526,N_12410,N_13967);
and UO_527 (O_527,N_12720,N_12046);
and UO_528 (O_528,N_13905,N_12090);
or UO_529 (O_529,N_14478,N_13895);
nand UO_530 (O_530,N_13774,N_13720);
nor UO_531 (O_531,N_13901,N_12950);
nor UO_532 (O_532,N_12957,N_13145);
nor UO_533 (O_533,N_13039,N_13091);
nor UO_534 (O_534,N_13680,N_12932);
nand UO_535 (O_535,N_13670,N_14981);
xnor UO_536 (O_536,N_13529,N_13513);
or UO_537 (O_537,N_12848,N_12707);
and UO_538 (O_538,N_14303,N_14799);
and UO_539 (O_539,N_14655,N_14835);
and UO_540 (O_540,N_13790,N_12064);
nor UO_541 (O_541,N_13809,N_12493);
or UO_542 (O_542,N_13005,N_14398);
and UO_543 (O_543,N_13756,N_12199);
and UO_544 (O_544,N_13439,N_12185);
nor UO_545 (O_545,N_12799,N_13481);
and UO_546 (O_546,N_12912,N_12760);
nor UO_547 (O_547,N_12494,N_14594);
nor UO_548 (O_548,N_12420,N_13260);
nand UO_549 (O_549,N_12730,N_14957);
nand UO_550 (O_550,N_13616,N_14919);
nand UO_551 (O_551,N_14276,N_12419);
or UO_552 (O_552,N_13073,N_12800);
and UO_553 (O_553,N_12448,N_12727);
nor UO_554 (O_554,N_13687,N_14358);
or UO_555 (O_555,N_12531,N_14373);
or UO_556 (O_556,N_12701,N_14860);
or UO_557 (O_557,N_14737,N_12403);
nor UO_558 (O_558,N_13035,N_14840);
nor UO_559 (O_559,N_12639,N_12281);
and UO_560 (O_560,N_12247,N_14731);
nor UO_561 (O_561,N_14359,N_14370);
xnor UO_562 (O_562,N_14171,N_12195);
nor UO_563 (O_563,N_13028,N_13938);
or UO_564 (O_564,N_12234,N_12510);
and UO_565 (O_565,N_12543,N_14654);
and UO_566 (O_566,N_13876,N_13391);
nand UO_567 (O_567,N_13384,N_14569);
or UO_568 (O_568,N_12648,N_12256);
xnor UO_569 (O_569,N_14272,N_13962);
xor UO_570 (O_570,N_13596,N_13524);
or UO_571 (O_571,N_13583,N_14005);
xnor UO_572 (O_572,N_12835,N_14700);
and UO_573 (O_573,N_14790,N_14228);
nor UO_574 (O_574,N_14771,N_14018);
nor UO_575 (O_575,N_12344,N_13806);
and UO_576 (O_576,N_12874,N_14823);
or UO_577 (O_577,N_13437,N_13937);
nand UO_578 (O_578,N_13732,N_14904);
and UO_579 (O_579,N_14032,N_12201);
nand UO_580 (O_580,N_12738,N_14999);
or UO_581 (O_581,N_13544,N_14742);
nand UO_582 (O_582,N_13128,N_14656);
or UO_583 (O_583,N_12359,N_13779);
xor UO_584 (O_584,N_14071,N_14250);
nor UO_585 (O_585,N_12035,N_12559);
or UO_586 (O_586,N_13818,N_14214);
nor UO_587 (O_587,N_14389,N_12485);
nand UO_588 (O_588,N_12069,N_14487);
nor UO_589 (O_589,N_12073,N_12425);
nand UO_590 (O_590,N_12617,N_14595);
or UO_591 (O_591,N_13382,N_13204);
nand UO_592 (O_592,N_14060,N_14621);
nand UO_593 (O_593,N_13501,N_12296);
nor UO_594 (O_594,N_13012,N_12144);
or UO_595 (O_595,N_13001,N_14770);
nor UO_596 (O_596,N_12391,N_12245);
or UO_597 (O_597,N_12189,N_12980);
nor UO_598 (O_598,N_14573,N_12556);
nand UO_599 (O_599,N_13885,N_12306);
nor UO_600 (O_600,N_13139,N_12762);
and UO_601 (O_601,N_12963,N_13546);
xnor UO_602 (O_602,N_13342,N_14598);
or UO_603 (O_603,N_12737,N_14841);
or UO_604 (O_604,N_14100,N_14374);
and UO_605 (O_605,N_13272,N_12530);
nand UO_606 (O_606,N_12566,N_14735);
xor UO_607 (O_607,N_12944,N_14728);
and UO_608 (O_608,N_14538,N_13246);
xor UO_609 (O_609,N_12383,N_13388);
and UO_610 (O_610,N_13955,N_14699);
and UO_611 (O_611,N_12421,N_14314);
and UO_612 (O_612,N_13247,N_12852);
and UO_613 (O_613,N_13218,N_12890);
nand UO_614 (O_614,N_13527,N_14696);
nor UO_615 (O_615,N_14177,N_13503);
nand UO_616 (O_616,N_13760,N_14163);
or UO_617 (O_617,N_12968,N_13804);
xnor UO_618 (O_618,N_12166,N_14074);
and UO_619 (O_619,N_13913,N_12253);
nor UO_620 (O_620,N_13127,N_14512);
and UO_621 (O_621,N_12067,N_13907);
or UO_622 (O_622,N_13304,N_14037);
or UO_623 (O_623,N_14331,N_14778);
nor UO_624 (O_624,N_13652,N_12098);
and UO_625 (O_625,N_14537,N_14524);
nor UO_626 (O_626,N_13722,N_12750);
or UO_627 (O_627,N_13614,N_13412);
or UO_628 (O_628,N_12088,N_12544);
nand UO_629 (O_629,N_12632,N_12389);
and UO_630 (O_630,N_14883,N_13250);
nand UO_631 (O_631,N_13566,N_12280);
nand UO_632 (O_632,N_12509,N_14578);
nand UO_633 (O_633,N_13631,N_14836);
xnor UO_634 (O_634,N_14763,N_12036);
and UO_635 (O_635,N_12937,N_14433);
and UO_636 (O_636,N_12970,N_12124);
nand UO_637 (O_637,N_14422,N_14062);
nand UO_638 (O_638,N_14320,N_13526);
or UO_639 (O_639,N_12395,N_13471);
nor UO_640 (O_640,N_14712,N_13846);
and UO_641 (O_641,N_12339,N_13297);
or UO_642 (O_642,N_13821,N_14688);
nor UO_643 (O_643,N_14768,N_14887);
and UO_644 (O_644,N_14293,N_12249);
or UO_645 (O_645,N_13591,N_12830);
xnor UO_646 (O_646,N_14048,N_13033);
nor UO_647 (O_647,N_13749,N_12568);
nand UO_648 (O_648,N_12329,N_14141);
nand UO_649 (O_649,N_14651,N_13862);
or UO_650 (O_650,N_14833,N_12778);
and UO_651 (O_651,N_14744,N_14950);
or UO_652 (O_652,N_12048,N_13992);
and UO_653 (O_653,N_12922,N_13368);
nand UO_654 (O_654,N_13493,N_14155);
nor UO_655 (O_655,N_12791,N_12342);
nor UO_656 (O_656,N_14148,N_12788);
or UO_657 (O_657,N_13994,N_14351);
and UO_658 (O_658,N_12732,N_12688);
or UO_659 (O_659,N_12460,N_12585);
xnor UO_660 (O_660,N_14941,N_12716);
or UO_661 (O_661,N_13768,N_12910);
and UO_662 (O_662,N_13224,N_13844);
nand UO_663 (O_663,N_13178,N_14685);
and UO_664 (O_664,N_13057,N_12677);
xnor UO_665 (O_665,N_14762,N_14286);
and UO_666 (O_666,N_13497,N_12480);
and UO_667 (O_667,N_14344,N_13561);
nand UO_668 (O_668,N_12629,N_12964);
nand UO_669 (O_669,N_12563,N_14998);
nand UO_670 (O_670,N_12712,N_12002);
or UO_671 (O_671,N_12192,N_12225);
nor UO_672 (O_672,N_14243,N_14827);
or UO_673 (O_673,N_14658,N_12129);
nor UO_674 (O_674,N_12891,N_12673);
nor UO_675 (O_675,N_13997,N_14853);
nor UO_676 (O_676,N_14327,N_12302);
nand UO_677 (O_677,N_14464,N_13482);
nor UO_678 (O_678,N_13990,N_12041);
and UO_679 (O_679,N_14977,N_12157);
xnor UO_680 (O_680,N_14198,N_14774);
and UO_681 (O_681,N_13278,N_12895);
nor UO_682 (O_682,N_13637,N_12464);
xor UO_683 (O_683,N_13726,N_12564);
or UO_684 (O_684,N_13900,N_14908);
nor UO_685 (O_685,N_13973,N_13663);
or UO_686 (O_686,N_14528,N_13217);
or UO_687 (O_687,N_13939,N_12224);
nand UO_688 (O_688,N_14460,N_14695);
nand UO_689 (O_689,N_12560,N_13788);
or UO_690 (O_690,N_13255,N_12148);
nand UO_691 (O_691,N_12722,N_12411);
or UO_692 (O_692,N_13168,N_13542);
xnor UO_693 (O_693,N_14011,N_13991);
and UO_694 (O_694,N_12829,N_12976);
nand UO_695 (O_695,N_12386,N_12773);
or UO_696 (O_696,N_12884,N_14864);
or UO_697 (O_697,N_13284,N_14767);
nor UO_698 (O_698,N_13324,N_14925);
and UO_699 (O_699,N_12273,N_12911);
nand UO_700 (O_700,N_14165,N_12522);
and UO_701 (O_701,N_14115,N_12146);
xor UO_702 (O_702,N_12938,N_14683);
or UO_703 (O_703,N_13509,N_12763);
nand UO_704 (O_704,N_12429,N_14520);
nor UO_705 (O_705,N_14309,N_13957);
nor UO_706 (O_706,N_14239,N_13963);
nor UO_707 (O_707,N_13463,N_13425);
nand UO_708 (O_708,N_14504,N_12538);
nor UO_709 (O_709,N_14274,N_14772);
and UO_710 (O_710,N_13899,N_12197);
and UO_711 (O_711,N_13887,N_14042);
and UO_712 (O_712,N_14039,N_13263);
nor UO_713 (O_713,N_12111,N_12500);
nand UO_714 (O_714,N_12595,N_14620);
nor UO_715 (O_715,N_12529,N_14547);
xnor UO_716 (O_716,N_13367,N_12001);
nand UO_717 (O_717,N_13267,N_12973);
nor UO_718 (O_718,N_12613,N_13079);
nor UO_719 (O_719,N_14642,N_13625);
and UO_720 (O_720,N_12045,N_12596);
nor UO_721 (O_721,N_14328,N_14132);
or UO_722 (O_722,N_12116,N_13329);
or UO_723 (O_723,N_13778,N_12697);
nand UO_724 (O_724,N_13589,N_13461);
nor UO_725 (O_725,N_12779,N_14897);
nand UO_726 (O_726,N_13865,N_13280);
nand UO_727 (O_727,N_12775,N_12191);
nor UO_728 (O_728,N_13723,N_14789);
and UO_729 (O_729,N_12313,N_14418);
or UO_730 (O_730,N_14343,N_12939);
or UO_731 (O_731,N_14203,N_13157);
nand UO_732 (O_732,N_12981,N_12335);
nand UO_733 (O_733,N_12203,N_13420);
nor UO_734 (O_734,N_12317,N_14086);
or UO_735 (O_735,N_13878,N_14185);
and UO_736 (O_736,N_12985,N_13159);
nand UO_737 (O_737,N_13308,N_14191);
nor UO_738 (O_738,N_13281,N_13414);
and UO_739 (O_739,N_13941,N_14515);
nor UO_740 (O_740,N_13336,N_14879);
and UO_741 (O_741,N_14160,N_14332);
nor UO_742 (O_742,N_12422,N_12060);
or UO_743 (O_743,N_12633,N_12859);
nand UO_744 (O_744,N_14974,N_14842);
nand UO_745 (O_745,N_14968,N_14473);
and UO_746 (O_746,N_13516,N_12598);
and UO_747 (O_747,N_13626,N_13522);
nor UO_748 (O_748,N_12366,N_14128);
nor UO_749 (O_749,N_13927,N_13891);
or UO_750 (O_750,N_13866,N_12266);
and UO_751 (O_751,N_12832,N_12251);
or UO_752 (O_752,N_14412,N_13602);
nand UO_753 (O_753,N_14560,N_12836);
xnor UO_754 (O_754,N_12693,N_12581);
nand UO_755 (O_755,N_13464,N_12236);
nor UO_756 (O_756,N_13911,N_14577);
and UO_757 (O_757,N_13315,N_12083);
nor UO_758 (O_758,N_12376,N_12995);
and UO_759 (O_759,N_12089,N_12334);
and UO_760 (O_760,N_14673,N_13773);
or UO_761 (O_761,N_12488,N_12745);
and UO_762 (O_762,N_14938,N_13849);
nor UO_763 (O_763,N_13840,N_12780);
and UO_764 (O_764,N_14280,N_13801);
or UO_765 (O_765,N_13448,N_14102);
xnor UO_766 (O_766,N_14469,N_14736);
nand UO_767 (O_767,N_12751,N_12742);
nand UO_768 (O_768,N_14427,N_14361);
nor UO_769 (O_769,N_12215,N_13445);
nor UO_770 (O_770,N_14459,N_13309);
nand UO_771 (O_771,N_12013,N_13392);
and UO_772 (O_772,N_13724,N_13307);
nand UO_773 (O_773,N_14665,N_13884);
or UO_774 (O_774,N_12956,N_14449);
or UO_775 (O_775,N_14084,N_13668);
or UO_776 (O_776,N_14965,N_14392);
or UO_777 (O_777,N_14394,N_12322);
or UO_778 (O_778,N_14388,N_14773);
and UO_779 (O_779,N_14501,N_12945);
or UO_780 (O_780,N_13515,N_12343);
or UO_781 (O_781,N_13292,N_14529);
xnor UO_782 (O_782,N_12373,N_12489);
and UO_783 (O_783,N_12279,N_14345);
and UO_784 (O_784,N_13220,N_13854);
nand UO_785 (O_785,N_14758,N_14368);
xnor UO_786 (O_786,N_14551,N_14820);
and UO_787 (O_787,N_13535,N_12935);
nor UO_788 (O_788,N_14337,N_14290);
nor UO_789 (O_789,N_13504,N_12729);
nand UO_790 (O_790,N_13394,N_13571);
and UO_791 (O_791,N_12806,N_14488);
nor UO_792 (O_792,N_13020,N_13782);
or UO_793 (O_793,N_13794,N_14178);
xor UO_794 (O_794,N_12860,N_14531);
or UO_795 (O_795,N_13588,N_14058);
or UO_796 (O_796,N_13375,N_12764);
nor UO_797 (O_797,N_14707,N_14277);
or UO_798 (O_798,N_13301,N_14380);
nand UO_799 (O_799,N_13869,N_13537);
and UO_800 (O_800,N_14367,N_12526);
xnor UO_801 (O_801,N_14710,N_13282);
or UO_802 (O_802,N_14690,N_13883);
or UO_803 (O_803,N_13174,N_13498);
or UO_804 (O_804,N_14550,N_13279);
or UO_805 (O_805,N_14815,N_14499);
nand UO_806 (O_806,N_14581,N_12929);
and UO_807 (O_807,N_12513,N_12614);
and UO_808 (O_808,N_13072,N_13067);
nor UO_809 (O_809,N_14195,N_13642);
nor UO_810 (O_810,N_12635,N_13015);
nand UO_811 (O_811,N_12987,N_13447);
or UO_812 (O_812,N_12337,N_13274);
or UO_813 (O_813,N_14935,N_12838);
nand UO_814 (O_814,N_12292,N_14143);
nor UO_815 (O_815,N_13265,N_12656);
nand UO_816 (O_816,N_12864,N_13273);
and UO_817 (O_817,N_14222,N_14135);
and UO_818 (O_818,N_13212,N_12409);
xnor UO_819 (O_819,N_14054,N_12770);
nor UO_820 (O_820,N_12481,N_12139);
nand UO_821 (O_821,N_13915,N_14281);
nand UO_822 (O_822,N_14907,N_12262);
and UO_823 (O_823,N_14340,N_13798);
xnor UO_824 (O_824,N_13488,N_13418);
nor UO_825 (O_825,N_14308,N_14798);
nor UO_826 (O_826,N_12310,N_13636);
nand UO_827 (O_827,N_14765,N_14800);
or UO_828 (O_828,N_14670,N_13597);
nor UO_829 (O_829,N_13585,N_14431);
and UO_830 (O_830,N_13759,N_13541);
and UO_831 (O_831,N_13089,N_14107);
and UO_832 (O_832,N_13234,N_13228);
and UO_833 (O_833,N_12181,N_14353);
or UO_834 (O_834,N_13712,N_13606);
nor UO_835 (O_835,N_13831,N_12081);
nor UO_836 (O_836,N_12179,N_12433);
or UO_837 (O_837,N_14508,N_12888);
and UO_838 (O_838,N_13754,N_12321);
and UO_839 (O_839,N_13860,N_14479);
or UO_840 (O_840,N_14880,N_13344);
and UO_841 (O_841,N_14704,N_12772);
and UO_842 (O_842,N_14292,N_14218);
nand UO_843 (O_843,N_12674,N_14716);
nand UO_844 (O_844,N_14426,N_13734);
and UO_845 (O_845,N_12845,N_12630);
nand UO_846 (O_846,N_13974,N_13071);
nor UO_847 (O_847,N_12503,N_13248);
and UO_848 (O_848,N_14947,N_13328);
xnor UO_849 (O_849,N_14555,N_13165);
nand UO_850 (O_850,N_12612,N_14363);
or UO_851 (O_851,N_12242,N_13295);
xor UO_852 (O_852,N_13610,N_12437);
and UO_853 (O_853,N_14223,N_13192);
and UO_854 (O_854,N_13487,N_14390);
or UO_855 (O_855,N_12140,N_14023);
nand UO_856 (O_856,N_14831,N_12217);
and UO_857 (O_857,N_13453,N_13417);
nor UO_858 (O_858,N_14319,N_12767);
and UO_859 (O_859,N_14629,N_13007);
xor UO_860 (O_860,N_14306,N_12074);
nor UO_861 (O_861,N_12686,N_12006);
nor UO_862 (O_862,N_14029,N_13473);
nand UO_863 (O_863,N_12662,N_13286);
or UO_864 (O_864,N_13916,N_13219);
nand UO_865 (O_865,N_14609,N_12996);
nor UO_866 (O_866,N_13772,N_12805);
nor UO_867 (O_867,N_14856,N_12994);
nor UO_868 (O_868,N_12125,N_14262);
or UO_869 (O_869,N_13356,N_14648);
or UO_870 (O_870,N_14534,N_12385);
or UO_871 (O_871,N_13027,N_14640);
and UO_872 (O_872,N_12669,N_12593);
xor UO_873 (O_873,N_12883,N_13499);
nand UO_874 (O_874,N_12311,N_14041);
and UO_875 (O_875,N_14652,N_14990);
or UO_876 (O_876,N_13316,N_14386);
nand UO_877 (O_877,N_14378,N_14335);
or UO_878 (O_878,N_12095,N_13253);
or UO_879 (O_879,N_12654,N_13163);
and UO_880 (O_880,N_12865,N_12681);
xor UO_881 (O_881,N_14312,N_12636);
or UO_882 (O_882,N_12796,N_14006);
nand UO_883 (O_883,N_14070,N_14622);
nand UO_884 (O_884,N_13751,N_13721);
nor UO_885 (O_885,N_14721,N_14349);
and UO_886 (O_886,N_12597,N_14204);
or UO_887 (O_887,N_13892,N_13755);
nand UO_888 (O_888,N_13528,N_14381);
nand UO_889 (O_889,N_13327,N_13677);
nand UO_890 (O_890,N_14470,N_13120);
nand UO_891 (O_891,N_12299,N_13988);
xor UO_892 (O_892,N_14837,N_14051);
nor UO_893 (O_893,N_13511,N_12626);
nand UO_894 (O_894,N_12966,N_13407);
and UO_895 (O_895,N_13651,N_13534);
nand UO_896 (O_896,N_12525,N_14872);
or UO_897 (O_897,N_13141,N_12159);
nor UO_898 (O_898,N_13252,N_12492);
or UO_899 (O_899,N_14419,N_14406);
or UO_900 (O_900,N_14766,N_12787);
and UO_901 (O_901,N_12913,N_14090);
and UO_902 (O_902,N_14483,N_14127);
xnor UO_903 (O_903,N_13584,N_14151);
nand UO_904 (O_904,N_12121,N_14708);
xnor UO_905 (O_905,N_13856,N_13875);
xnor UO_906 (O_906,N_14330,N_12628);
and UO_907 (O_907,N_14447,N_14121);
or UO_908 (O_908,N_14123,N_14212);
or UO_909 (O_909,N_13021,N_14962);
or UO_910 (O_910,N_13952,N_12757);
nor UO_911 (O_911,N_14602,N_12983);
and UO_912 (O_912,N_13688,N_13138);
nor UO_913 (O_913,N_13519,N_12084);
and UO_914 (O_914,N_14592,N_13569);
or UO_915 (O_915,N_14004,N_12925);
nand UO_916 (O_916,N_12871,N_14677);
or UO_917 (O_917,N_13106,N_13432);
nand UO_918 (O_918,N_13235,N_12012);
or UO_919 (O_919,N_12103,N_14201);
or UO_920 (O_920,N_13512,N_13216);
nor UO_921 (O_921,N_12897,N_13256);
and UO_922 (O_922,N_14983,N_12967);
nand UO_923 (O_923,N_14497,N_13520);
nor UO_924 (O_924,N_14031,N_12714);
and UO_925 (O_925,N_13568,N_14873);
xor UO_926 (O_926,N_12049,N_14076);
or UO_927 (O_927,N_13701,N_12586);
xor UO_928 (O_928,N_14987,N_14112);
xnor UO_929 (O_929,N_14285,N_13396);
nor UO_930 (O_930,N_12988,N_14996);
or UO_931 (O_931,N_13690,N_13820);
nor UO_932 (O_932,N_14558,N_12676);
nand UO_933 (O_933,N_12506,N_13757);
or UO_934 (O_934,N_14188,N_13659);
nor UO_935 (O_935,N_14561,N_12567);
and UO_936 (O_936,N_12305,N_14208);
nor UO_937 (O_937,N_12515,N_14053);
nor UO_938 (O_938,N_12019,N_13882);
xnor UO_939 (O_939,N_12561,N_12618);
nor UO_940 (O_940,N_14307,N_14026);
or UO_941 (O_941,N_13624,N_13629);
and UO_942 (O_942,N_12827,N_13424);
and UO_943 (O_943,N_12953,N_12731);
and UO_944 (O_944,N_12170,N_14928);
nand UO_945 (O_945,N_13114,N_14082);
xnor UO_946 (O_946,N_13486,N_13929);
nor UO_947 (O_947,N_13662,N_14899);
and UO_948 (O_948,N_14988,N_12534);
nor UO_949 (O_949,N_13573,N_13580);
nor UO_950 (O_950,N_14877,N_14251);
and UO_951 (O_951,N_12248,N_14933);
and UO_952 (O_952,N_13956,N_13841);
nor UO_953 (O_953,N_12137,N_14659);
nand UO_954 (O_954,N_13131,N_13748);
and UO_955 (O_955,N_12054,N_14838);
nand UO_956 (O_956,N_13635,N_12975);
or UO_957 (O_957,N_14278,N_13733);
nand UO_958 (O_958,N_13671,N_13006);
xor UO_959 (O_959,N_14963,N_12982);
nor UO_960 (O_960,N_13719,N_14632);
nand UO_961 (O_961,N_13183,N_13036);
nor UO_962 (O_962,N_14379,N_14168);
nor UO_963 (O_963,N_13034,N_12165);
nand UO_964 (O_964,N_12068,N_14559);
and UO_965 (O_965,N_14811,N_13641);
nor UO_966 (O_966,N_12698,N_14544);
and UO_967 (O_967,N_13710,N_13704);
or UO_968 (O_968,N_12599,N_14077);
or UO_969 (O_969,N_13151,N_12352);
nand UO_970 (O_970,N_14383,N_14929);
xnor UO_971 (O_971,N_12692,N_14676);
and UO_972 (O_972,N_12327,N_14697);
nand UO_973 (O_973,N_14553,N_13152);
or UO_974 (O_974,N_13829,N_12666);
nand UO_975 (O_975,N_12961,N_12539);
or UO_976 (O_976,N_14923,N_12168);
nand UO_977 (O_977,N_14526,N_13825);
nor UO_978 (O_978,N_13314,N_13010);
and UO_979 (O_979,N_13608,N_14414);
or UO_980 (O_980,N_14471,N_12847);
or UO_981 (O_981,N_14458,N_12594);
or UO_982 (O_982,N_12102,N_13871);
and UO_983 (O_983,N_12634,N_14438);
and UO_984 (O_984,N_13017,N_12721);
or UO_985 (O_985,N_14094,N_14580);
nor UO_986 (O_986,N_14532,N_14795);
and UO_987 (O_987,N_12661,N_14442);
and UO_988 (O_988,N_12428,N_14570);
or UO_989 (O_989,N_12183,N_14494);
nand UO_990 (O_990,N_13186,N_12274);
nand UO_991 (O_991,N_13993,N_12694);
or UO_992 (O_992,N_12155,N_12298);
or UO_993 (O_993,N_14275,N_14316);
nor UO_994 (O_994,N_14101,N_13593);
or UO_995 (O_995,N_14068,N_12293);
or UO_996 (O_996,N_13431,N_12683);
nand UO_997 (O_997,N_12724,N_14453);
and UO_998 (O_998,N_13438,N_12283);
and UO_999 (O_999,N_13575,N_13085);
or UO_1000 (O_1000,N_12926,N_12459);
nand UO_1001 (O_1001,N_14926,N_12009);
nor UO_1002 (O_1002,N_13241,N_13052);
or UO_1003 (O_1003,N_12855,N_14637);
nand UO_1004 (O_1004,N_14663,N_14021);
or UO_1005 (O_1005,N_12186,N_13550);
and UO_1006 (O_1006,N_13917,N_12619);
nand UO_1007 (O_1007,N_13338,N_13401);
nand UO_1008 (O_1008,N_13061,N_14994);
xor UO_1009 (O_1009,N_13346,N_14283);
nand UO_1010 (O_1010,N_13266,N_12960);
nor UO_1011 (O_1011,N_13489,N_12194);
xnor UO_1012 (O_1012,N_12315,N_14248);
nor UO_1013 (O_1013,N_12092,N_13287);
nor UO_1014 (O_1014,N_13623,N_13254);
and UO_1015 (O_1015,N_12882,N_13728);
and UO_1016 (O_1016,N_14972,N_13018);
nor UO_1017 (O_1017,N_14484,N_14081);
nor UO_1018 (O_1018,N_12484,N_13259);
nor UO_1019 (O_1019,N_13249,N_14010);
and UO_1020 (O_1020,N_13582,N_13323);
nand UO_1021 (O_1021,N_14894,N_13586);
or UO_1022 (O_1022,N_13011,N_13364);
or UO_1023 (O_1023,N_14701,N_13004);
or UO_1024 (O_1024,N_12275,N_14657);
nor UO_1025 (O_1025,N_13842,N_14209);
and UO_1026 (O_1026,N_13977,N_12258);
nand UO_1027 (O_1027,N_13332,N_13334);
and UO_1028 (O_1028,N_12160,N_12499);
or UO_1029 (O_1029,N_13080,N_12290);
and UO_1030 (O_1030,N_13466,N_12603);
nor UO_1031 (O_1031,N_13198,N_13115);
nor UO_1032 (O_1032,N_13177,N_12637);
nand UO_1033 (O_1033,N_13373,N_12804);
or UO_1034 (O_1034,N_13185,N_12331);
nand UO_1035 (O_1035,N_12627,N_14124);
or UO_1036 (O_1036,N_14751,N_13802);
or UO_1037 (O_1037,N_13402,N_14562);
nand UO_1038 (O_1038,N_13594,N_14034);
nand UO_1039 (O_1039,N_13350,N_14954);
xnor UO_1040 (O_1040,N_14847,N_14917);
and UO_1041 (O_1041,N_12908,N_14369);
nand UO_1042 (O_1042,N_13202,N_14891);
and UO_1043 (O_1043,N_14172,N_14265);
nor UO_1044 (O_1044,N_14825,N_12533);
nand UO_1045 (O_1045,N_14411,N_14264);
nor UO_1046 (O_1046,N_12161,N_14966);
and UO_1047 (O_1047,N_14187,N_12399);
and UO_1048 (O_1048,N_12550,N_13996);
nor UO_1049 (O_1049,N_12377,N_12685);
nor UO_1050 (O_1050,N_12990,N_12545);
or UO_1051 (O_1051,N_12109,N_14008);
or UO_1052 (O_1052,N_13698,N_12101);
or UO_1053 (O_1053,N_14582,N_14454);
nor UO_1054 (O_1054,N_14513,N_12415);
and UO_1055 (O_1055,N_12219,N_13983);
nand UO_1056 (O_1056,N_13630,N_14713);
nand UO_1057 (O_1057,N_13959,N_14949);
nor UO_1058 (O_1058,N_14410,N_12319);
xor UO_1059 (O_1059,N_12381,N_13706);
nand UO_1060 (O_1060,N_12117,N_12182);
and UO_1061 (O_1061,N_12024,N_13811);
and UO_1062 (O_1062,N_13852,N_13765);
nor UO_1063 (O_1063,N_12657,N_14644);
and UO_1064 (O_1064,N_12786,N_13472);
nor UO_1065 (O_1065,N_13567,N_13739);
or UO_1066 (O_1066,N_14046,N_14002);
or UO_1067 (O_1067,N_13320,N_12106);
nor UO_1068 (O_1068,N_13800,N_12841);
nand UO_1069 (O_1069,N_14649,N_14131);
and UO_1070 (O_1070,N_13934,N_14714);
nand UO_1071 (O_1071,N_14804,N_12328);
xor UO_1072 (O_1072,N_12496,N_12660);
or UO_1073 (O_1073,N_13715,N_13423);
nor UO_1074 (O_1074,N_12384,N_13469);
xor UO_1075 (O_1075,N_14971,N_13507);
nand UO_1076 (O_1076,N_13545,N_13972);
nor UO_1077 (O_1077,N_13819,N_12338);
or UO_1078 (O_1078,N_12078,N_12607);
and UO_1079 (O_1079,N_14114,N_12087);
xor UO_1080 (O_1080,N_12776,N_14104);
nor UO_1081 (O_1081,N_13025,N_14769);
nor UO_1082 (O_1082,N_12717,N_12834);
xor UO_1083 (O_1083,N_13122,N_13679);
xor UO_1084 (O_1084,N_13505,N_12715);
nor UO_1085 (O_1085,N_12769,N_12962);
or UO_1086 (O_1086,N_12147,N_13333);
nor UO_1087 (O_1087,N_13574,N_13923);
or UO_1088 (O_1088,N_13928,N_13014);
xor UO_1089 (O_1089,N_14819,N_14147);
or UO_1090 (O_1090,N_13949,N_13645);
nor UO_1091 (O_1091,N_14596,N_12239);
and UO_1092 (O_1092,N_14043,N_14694);
xor UO_1093 (O_1093,N_12301,N_12082);
or UO_1094 (O_1094,N_14324,N_12151);
and UO_1095 (O_1095,N_13251,N_13321);
and UO_1096 (O_1096,N_12392,N_13707);
or UO_1097 (O_1097,N_13257,N_12887);
nor UO_1098 (O_1098,N_12020,N_12749);
or UO_1099 (O_1099,N_13098,N_12979);
nor UO_1100 (O_1100,N_14382,N_14809);
xnor UO_1101 (O_1101,N_12167,N_12755);
nor UO_1102 (O_1102,N_13393,N_13355);
nand UO_1103 (O_1103,N_13564,N_12941);
or UO_1104 (O_1104,N_13124,N_14803);
nor UO_1105 (O_1105,N_14166,N_13658);
nor UO_1106 (O_1106,N_12034,N_13024);
or UO_1107 (O_1107,N_13419,N_14298);
nand UO_1108 (O_1108,N_14993,N_12726);
and UO_1109 (O_1109,N_13791,N_14056);
nand UO_1110 (O_1110,N_12000,N_12211);
xor UO_1111 (O_1111,N_14003,N_13369);
xor UO_1112 (O_1112,N_14843,N_13101);
nand UO_1113 (O_1113,N_12070,N_14259);
or UO_1114 (O_1114,N_13413,N_12589);
nor UO_1115 (O_1115,N_14397,N_12295);
or UO_1116 (O_1116,N_13480,N_13533);
and UO_1117 (O_1117,N_14816,N_12005);
nor UO_1118 (O_1118,N_13792,N_13989);
nand UO_1119 (O_1119,N_13066,N_14711);
nor UO_1120 (O_1120,N_14705,N_14896);
and UO_1121 (O_1121,N_12363,N_14385);
or UO_1122 (O_1122,N_12443,N_14828);
nand UO_1123 (O_1123,N_14583,N_14118);
nor UO_1124 (O_1124,N_13787,N_13406);
and UO_1125 (O_1125,N_14294,N_14591);
xor UO_1126 (O_1126,N_14354,N_12997);
and UO_1127 (O_1127,N_12375,N_12822);
nand UO_1128 (O_1128,N_12177,N_14400);
or UO_1129 (O_1129,N_14498,N_12672);
or UO_1130 (O_1130,N_12404,N_14271);
nand UO_1131 (O_1131,N_14200,N_13612);
nand UO_1132 (O_1132,N_13926,N_14257);
xor UO_1133 (O_1133,N_13930,N_13467);
nor UO_1134 (O_1134,N_12380,N_12809);
or UO_1135 (O_1135,N_12288,N_13558);
or UO_1136 (O_1136,N_13980,N_13086);
xnor UO_1137 (O_1137,N_13359,N_14119);
nor UO_1138 (O_1138,N_13598,N_13199);
nand UO_1139 (O_1139,N_12675,N_14211);
or UO_1140 (O_1140,N_13888,N_13764);
xnor UO_1141 (O_1141,N_13538,N_14049);
or UO_1142 (O_1142,N_14122,N_12332);
and UO_1143 (O_1143,N_13479,N_12011);
and UO_1144 (O_1144,N_12318,N_13646);
or UO_1145 (O_1145,N_12040,N_14913);
or UO_1146 (O_1146,N_14858,N_14310);
and UO_1147 (O_1147,N_13478,N_13319);
nand UO_1148 (O_1148,N_14724,N_12949);
or UO_1149 (O_1149,N_12066,N_12725);
or UO_1150 (O_1150,N_13775,N_14302);
nor UO_1151 (O_1151,N_12333,N_14157);
xnor UO_1152 (O_1152,N_12833,N_12400);
xor UO_1153 (O_1153,N_13290,N_12402);
and UO_1154 (O_1154,N_14901,N_13830);
and UO_1155 (O_1155,N_13552,N_14516);
or UO_1156 (O_1156,N_13097,N_13695);
xor UO_1157 (O_1157,N_14432,N_12033);
xnor UO_1158 (O_1158,N_12454,N_13813);
nand UO_1159 (O_1159,N_12826,N_12038);
xnor UO_1160 (O_1160,N_12664,N_12736);
nand UO_1161 (O_1161,N_13300,N_13491);
nor UO_1162 (O_1162,N_12362,N_14098);
and UO_1163 (O_1163,N_13700,N_13026);
or UO_1164 (O_1164,N_14233,N_12475);
and UO_1165 (O_1165,N_13607,N_13158);
or UO_1166 (O_1166,N_12220,N_12576);
and UO_1167 (O_1167,N_13879,N_13685);
nand UO_1168 (O_1168,N_12104,N_13609);
or UO_1169 (O_1169,N_13948,N_12284);
nor UO_1170 (O_1170,N_14317,N_13944);
nor UO_1171 (O_1171,N_13058,N_14401);
or UO_1172 (O_1172,N_14668,N_14761);
and UO_1173 (O_1173,N_14886,N_13604);
nand UO_1174 (O_1174,N_12814,N_14593);
nand UO_1175 (O_1175,N_13579,N_13490);
or UO_1176 (O_1176,N_12663,N_12208);
nand UO_1177 (O_1177,N_12711,N_13087);
nor UO_1178 (O_1178,N_12934,N_13530);
nand UO_1179 (O_1179,N_13664,N_14911);
xor UO_1180 (O_1180,N_14443,N_13893);
nor UO_1181 (O_1181,N_13894,N_14445);
nand UO_1182 (O_1182,N_13054,N_13311);
nor UO_1183 (O_1183,N_12854,N_13153);
or UO_1184 (O_1184,N_13194,N_12231);
nand UO_1185 (O_1185,N_12453,N_14329);
and UO_1186 (O_1186,N_12261,N_14162);
nor UO_1187 (O_1187,N_13023,N_12233);
or UO_1188 (O_1188,N_12255,N_14956);
nand UO_1189 (O_1189,N_14545,N_14535);
xor UO_1190 (O_1190,N_13030,N_12388);
or UO_1191 (O_1191,N_12282,N_12324);
or UO_1192 (O_1192,N_14746,N_14133);
nor UO_1193 (O_1193,N_14465,N_12893);
or UO_1194 (O_1194,N_14444,N_12294);
xnor UO_1195 (O_1195,N_13276,N_12444);
or UO_1196 (O_1196,N_14753,N_14821);
and UO_1197 (O_1197,N_14055,N_14326);
or UO_1198 (O_1198,N_12174,N_12575);
and UO_1199 (O_1199,N_12655,N_13404);
nand UO_1200 (O_1200,N_13548,N_13408);
or UO_1201 (O_1201,N_13924,N_12899);
nand UO_1202 (O_1202,N_12378,N_12571);
or UO_1203 (O_1203,N_12942,N_13611);
and UO_1204 (O_1204,N_12016,N_13562);
xor UO_1205 (O_1205,N_12198,N_14607);
nor UO_1206 (O_1206,N_12615,N_14505);
and UO_1207 (O_1207,N_14757,N_13121);
and UO_1208 (O_1208,N_14474,N_12232);
and UO_1209 (O_1209,N_13903,N_14407);
and UO_1210 (O_1210,N_12881,N_13188);
nor UO_1211 (O_1211,N_13440,N_13236);
nor UO_1212 (O_1212,N_12158,N_13354);
nand UO_1213 (O_1213,N_14924,N_14213);
and UO_1214 (O_1214,N_13766,N_13376);
nand UO_1215 (O_1215,N_14106,N_13709);
nand UO_1216 (O_1216,N_12028,N_14511);
and UO_1217 (O_1217,N_13978,N_13696);
nand UO_1218 (O_1218,N_12042,N_13353);
xor UO_1219 (O_1219,N_13815,N_13164);
nor UO_1220 (O_1220,N_12187,N_12647);
or UO_1221 (O_1221,N_13416,N_12254);
nand UO_1222 (O_1222,N_12820,N_12999);
and UO_1223 (O_1223,N_12470,N_13326);
nor UO_1224 (O_1224,N_12678,N_12350);
or UO_1225 (O_1225,N_12735,N_13060);
and UO_1226 (O_1226,N_13009,N_14631);
nand UO_1227 (O_1227,N_12579,N_13022);
and UO_1228 (O_1228,N_14154,N_12801);
xor UO_1229 (O_1229,N_13783,N_12519);
nand UO_1230 (O_1230,N_14754,N_14794);
and UO_1231 (O_1231,N_12007,N_14015);
nor UO_1232 (O_1232,N_13554,N_13214);
nor UO_1233 (O_1233,N_12209,N_14914);
nor UO_1234 (O_1234,N_13632,N_12252);
and UO_1235 (O_1235,N_13540,N_14299);
and UO_1236 (O_1236,N_14229,N_14961);
nor UO_1237 (O_1237,N_12782,N_13047);
or UO_1238 (O_1238,N_14970,N_13476);
or UO_1239 (O_1239,N_13599,N_13559);
xnor UO_1240 (O_1240,N_14725,N_14662);
nor UO_1241 (O_1241,N_14610,N_14495);
nand UO_1242 (O_1242,N_14424,N_12771);
nand UO_1243 (O_1243,N_12424,N_14805);
or UO_1244 (O_1244,N_14226,N_13154);
nor UO_1245 (O_1245,N_13676,N_13838);
nor UO_1246 (O_1246,N_12541,N_14095);
and UO_1247 (O_1247,N_12008,N_14057);
and UO_1248 (O_1248,N_13046,N_14664);
nand UO_1249 (O_1249,N_13742,N_14548);
and UO_1250 (O_1250,N_13725,N_13729);
nand UO_1251 (O_1251,N_13855,N_14279);
nor UO_1252 (O_1252,N_13904,N_14267);
or UO_1253 (O_1253,N_13283,N_14715);
nand UO_1254 (O_1254,N_13638,N_13500);
nand UO_1255 (O_1255,N_14967,N_13886);
nand UO_1256 (O_1256,N_13366,N_14939);
nor UO_1257 (O_1257,N_12143,N_12452);
nand UO_1258 (O_1258,N_12487,N_12032);
and UO_1259 (O_1259,N_14606,N_14089);
and UO_1260 (O_1260,N_14301,N_13850);
or UO_1261 (O_1261,N_13711,N_14729);
nand UO_1262 (O_1262,N_14687,N_12562);
or UO_1263 (O_1263,N_13945,N_12590);
nor UO_1264 (O_1264,N_12336,N_14296);
nor UO_1265 (O_1265,N_14943,N_13102);
or UO_1266 (O_1266,N_12128,N_13041);
nor UO_1267 (O_1267,N_12699,N_13303);
nand UO_1268 (O_1268,N_14780,N_12269);
and UO_1269 (O_1269,N_14069,N_12053);
nor UO_1270 (O_1270,N_14951,N_12200);
or UO_1271 (O_1271,N_13182,N_12844);
nand UO_1272 (O_1272,N_12959,N_12027);
nor UO_1273 (O_1273,N_12303,N_12954);
or UO_1274 (O_1274,N_13064,N_13117);
nand UO_1275 (O_1275,N_12175,N_13042);
nand UO_1276 (O_1276,N_14554,N_12478);
nor UO_1277 (O_1277,N_14477,N_13123);
nand UO_1278 (O_1278,N_13807,N_14138);
nand UO_1279 (O_1279,N_14170,N_14576);
nor UO_1280 (O_1280,N_13812,N_12580);
or UO_1281 (O_1281,N_13832,N_13675);
nand UO_1282 (O_1282,N_12947,N_14125);
or UO_1283 (O_1283,N_14989,N_13341);
nand UO_1284 (O_1284,N_12798,N_14311);
nor UO_1285 (O_1285,N_13762,N_14099);
nand UO_1286 (O_1286,N_12734,N_14356);
or UO_1287 (O_1287,N_14639,N_14936);
xnor UO_1288 (O_1288,N_12427,N_14709);
nand UO_1289 (O_1289,N_13496,N_12784);
and UO_1290 (O_1290,N_14347,N_12592);
nor UO_1291 (O_1291,N_12118,N_13789);
nor UO_1292 (O_1292,N_13383,N_12345);
nand UO_1293 (O_1293,N_12004,N_12172);
nand UO_1294 (O_1294,N_12287,N_13313);
nor UO_1295 (O_1295,N_12405,N_12813);
or UO_1296 (O_1296,N_13581,N_13647);
and UO_1297 (O_1297,N_12136,N_12291);
nand UO_1298 (O_1298,N_13613,N_13371);
xnor UO_1299 (O_1299,N_14906,N_13459);
and UO_1300 (O_1300,N_12831,N_13444);
nand UO_1301 (O_1301,N_13648,N_12914);
nand UO_1302 (O_1302,N_14269,N_12856);
nor UO_1303 (O_1303,N_13565,N_14396);
or UO_1304 (O_1304,N_14182,N_14866);
xnor UO_1305 (O_1305,N_14288,N_13031);
nor UO_1306 (O_1306,N_12169,N_13950);
nand UO_1307 (O_1307,N_14915,N_13692);
and UO_1308 (O_1308,N_14633,N_14958);
or UO_1309 (O_1309,N_14027,N_13318);
and UO_1310 (O_1310,N_13227,N_13686);
nand UO_1311 (O_1311,N_12265,N_13452);
nor UO_1312 (O_1312,N_13793,N_12364);
or UO_1313 (O_1313,N_12096,N_12842);
xor UO_1314 (O_1314,N_14910,N_13985);
xor UO_1315 (O_1315,N_14486,N_14557);
nand UO_1316 (O_1316,N_14408,N_12126);
and UO_1317 (O_1317,N_12638,N_14393);
or UO_1318 (O_1318,N_12351,N_13465);
or UO_1319 (O_1319,N_13331,N_14152);
or UO_1320 (O_1320,N_12080,N_12141);
and UO_1321 (O_1321,N_13523,N_12414);
xor UO_1322 (O_1322,N_14434,N_13845);
and UO_1323 (O_1323,N_13029,N_13603);
or UO_1324 (O_1324,N_12221,N_13745);
xnor UO_1325 (O_1325,N_14134,N_13395);
or UO_1326 (O_1326,N_14693,N_14186);
or UO_1327 (O_1327,N_13918,N_12397);
nor UO_1328 (O_1328,N_12766,N_12739);
or UO_1329 (O_1329,N_14818,N_13620);
nand UO_1330 (O_1330,N_14706,N_12621);
nor UO_1331 (O_1331,N_13370,N_12010);
or UO_1332 (O_1332,N_13038,N_14717);
xnor UO_1333 (O_1333,N_13998,N_13264);
nor UO_1334 (O_1334,N_13921,N_14291);
nand UO_1335 (O_1335,N_13753,N_14759);
or UO_1336 (O_1336,N_14088,N_13456);
nor UO_1337 (O_1337,N_13531,N_12142);
nand UO_1338 (O_1338,N_13195,N_14745);
nor UO_1339 (O_1339,N_12467,N_13399);
and UO_1340 (O_1340,N_12794,N_12511);
nand UO_1341 (O_1341,N_13222,N_12374);
nand UO_1342 (O_1342,N_14207,N_12547);
and UO_1343 (O_1343,N_14918,N_14065);
nand UO_1344 (O_1344,N_14552,N_14110);
xor UO_1345 (O_1345,N_14252,N_12824);
nor UO_1346 (O_1346,N_13951,N_13040);
nand UO_1347 (O_1347,N_13976,N_12527);
nand UO_1348 (O_1348,N_12244,N_12903);
nand UO_1349 (O_1349,N_13979,N_12105);
and UO_1350 (O_1350,N_14905,N_12551);
nor UO_1351 (O_1351,N_13409,N_12474);
and UO_1352 (O_1352,N_12569,N_14934);
nor UO_1353 (O_1353,N_14227,N_14623);
or UO_1354 (O_1354,N_12785,N_13016);
or UO_1355 (O_1355,N_12789,N_12207);
or UO_1356 (O_1356,N_12365,N_14575);
nor UO_1357 (O_1357,N_12025,N_13262);
nor UO_1358 (O_1358,N_14564,N_13699);
nor UO_1359 (O_1359,N_14571,N_13050);
or UO_1360 (O_1360,N_14682,N_13874);
nor UO_1361 (O_1361,N_13665,N_14589);
and UO_1362 (O_1362,N_13306,N_12099);
xor UO_1363 (O_1363,N_13380,N_13352);
and UO_1364 (O_1364,N_12668,N_13442);
and UO_1365 (O_1365,N_14219,N_13261);
nand UO_1366 (O_1366,N_12163,N_12286);
xor UO_1367 (O_1367,N_13999,N_13289);
nor UO_1368 (O_1368,N_14247,N_12436);
and UO_1369 (O_1369,N_13643,N_13966);
and UO_1370 (O_1370,N_12394,N_12710);
nand UO_1371 (O_1371,N_12955,N_13769);
xor UO_1372 (O_1372,N_13931,N_12821);
and UO_1373 (O_1373,N_13965,N_14857);
and UO_1374 (O_1374,N_12535,N_14158);
and UO_1375 (O_1375,N_13434,N_12491);
nor UO_1376 (O_1376,N_14791,N_13837);
nand UO_1377 (O_1377,N_12423,N_14618);
or UO_1378 (O_1378,N_13902,N_12974);
xor UO_1379 (O_1379,N_14364,N_12466);
and UO_1380 (O_1380,N_13226,N_12093);
and UO_1381 (O_1381,N_14430,N_12991);
and UO_1382 (O_1382,N_12309,N_12210);
or UO_1383 (O_1383,N_14184,N_14643);
or UO_1384 (O_1384,N_14822,N_14900);
nor UO_1385 (O_1385,N_14064,N_13096);
xor UO_1386 (O_1386,N_12610,N_13730);
nand UO_1387 (O_1387,N_14960,N_13166);
or UO_1388 (O_1388,N_12885,N_12623);
nand UO_1389 (O_1389,N_14467,N_14536);
and UO_1390 (O_1390,N_14793,N_12572);
and UO_1391 (O_1391,N_13805,N_14522);
and UO_1392 (O_1392,N_12756,N_14752);
nand UO_1393 (O_1393,N_14748,N_14365);
and UO_1394 (O_1394,N_13714,N_14784);
or UO_1395 (O_1395,N_13065,N_12445);
and UO_1396 (O_1396,N_14834,N_13669);
or UO_1397 (O_1397,N_13691,N_12758);
nand UO_1398 (O_1398,N_14680,N_13112);
or UO_1399 (O_1399,N_14940,N_14788);
nand UO_1400 (O_1400,N_12909,N_13981);
and UO_1401 (O_1401,N_13232,N_14566);
xnor UO_1402 (O_1402,N_12577,N_14931);
and UO_1403 (O_1403,N_12792,N_13335);
nand UO_1404 (O_1404,N_13093,N_13656);
nand UO_1405 (O_1405,N_13209,N_14616);
and UO_1406 (O_1406,N_13111,N_13242);
and UO_1407 (O_1407,N_14826,N_14403);
nand UO_1408 (O_1408,N_13358,N_12152);
and UO_1409 (O_1409,N_12868,N_12620);
and UO_1410 (O_1410,N_13925,N_14579);
or UO_1411 (O_1411,N_14980,N_12528);
or UO_1412 (O_1412,N_14927,N_14871);
and UO_1413 (O_1413,N_14945,N_14287);
nor UO_1414 (O_1414,N_14153,N_13889);
nor UO_1415 (O_1415,N_13090,N_13454);
nor UO_1416 (O_1416,N_12557,N_12431);
xor UO_1417 (O_1417,N_14895,N_14801);
xnor UO_1418 (O_1418,N_12604,N_12490);
nand UO_1419 (O_1419,N_14615,N_13672);
or UO_1420 (O_1420,N_14256,N_12471);
nand UO_1421 (O_1421,N_13836,N_14220);
nor UO_1422 (O_1422,N_13436,N_14093);
nor UO_1423 (O_1423,N_14439,N_13312);
or UO_1424 (O_1424,N_14001,N_12665);
or UO_1425 (O_1425,N_12014,N_13968);
nand UO_1426 (O_1426,N_12272,N_14875);
nand UO_1427 (O_1427,N_12741,N_13095);
or UO_1428 (O_1428,N_14489,N_14395);
or UO_1429 (O_1429,N_13201,N_13348);
nand UO_1430 (O_1430,N_12889,N_14854);
or UO_1431 (O_1431,N_12876,N_12989);
nand UO_1432 (O_1432,N_14740,N_14890);
and UO_1433 (O_1433,N_12808,N_12723);
or UO_1434 (O_1434,N_12520,N_13207);
nor UO_1435 (O_1435,N_14599,N_13873);
nor UO_1436 (O_1436,N_12653,N_12700);
nor UO_1437 (O_1437,N_13474,N_14130);
nor UO_1438 (O_1438,N_12430,N_14009);
or UO_1439 (O_1439,N_13129,N_13291);
nor UO_1440 (O_1440,N_12691,N_12271);
nand UO_1441 (O_1441,N_14732,N_14192);
nor UO_1442 (O_1442,N_12622,N_12605);
nor UO_1443 (O_1443,N_14802,N_14404);
and UO_1444 (O_1444,N_14325,N_13092);
nand UO_1445 (O_1445,N_14059,N_13644);
and UO_1446 (O_1446,N_12679,N_12713);
or UO_1447 (O_1447,N_13225,N_12044);
xnor UO_1448 (O_1448,N_12867,N_12446);
nand UO_1449 (O_1449,N_12582,N_14944);
xnor UO_1450 (O_1450,N_13100,N_13595);
nor UO_1451 (O_1451,N_14829,N_14587);
and UO_1452 (O_1452,N_12450,N_14190);
and UO_1453 (O_1453,N_14885,N_12880);
and UO_1454 (O_1454,N_12072,N_13140);
or UO_1455 (O_1455,N_13828,N_13702);
or UO_1456 (O_1456,N_13477,N_12434);
or UO_1457 (O_1457,N_14646,N_13240);
nor UO_1458 (O_1458,N_12558,N_13435);
xnor UO_1459 (O_1459,N_12469,N_13160);
or UO_1460 (O_1460,N_13947,N_12164);
or UO_1461 (O_1461,N_12091,N_14224);
nor UO_1462 (O_1462,N_14016,N_13763);
or UO_1463 (O_1463,N_13834,N_13781);
and UO_1464 (O_1464,N_12449,N_13693);
nand UO_1465 (O_1465,N_13206,N_14506);
xnor UO_1466 (O_1466,N_13430,N_12341);
and UO_1467 (O_1467,N_14038,N_14734);
or UO_1468 (O_1468,N_13385,N_12417);
nand UO_1469 (O_1469,N_14402,N_14083);
or UO_1470 (O_1470,N_13705,N_13148);
and UO_1471 (O_1471,N_14241,N_13618);
nand UO_1472 (O_1472,N_13731,N_13433);
or UO_1473 (O_1473,N_14173,N_13920);
nor UO_1474 (O_1474,N_13116,N_14437);
and UO_1475 (O_1475,N_12993,N_14703);
xor UO_1476 (O_1476,N_13942,N_14764);
xor UO_1477 (O_1477,N_14266,N_13078);
nor UO_1478 (O_1478,N_14176,N_13661);
nand UO_1479 (O_1479,N_13317,N_14624);
nor UO_1480 (O_1480,N_13851,N_12308);
xor UO_1481 (O_1481,N_14865,N_14608);
nor UO_1482 (O_1482,N_14741,N_14237);
xor UO_1483 (O_1483,N_13426,N_12022);
nand UO_1484 (O_1484,N_14273,N_12058);
and UO_1485 (O_1485,N_14510,N_12761);
xor UO_1486 (O_1486,N_13960,N_12150);
and UO_1487 (O_1487,N_14468,N_12565);
nor UO_1488 (O_1488,N_14995,N_13397);
xnor UO_1489 (O_1489,N_13379,N_12330);
xnor UO_1490 (O_1490,N_13363,N_13068);
or UO_1491 (O_1491,N_14627,N_12227);
nor UO_1492 (O_1492,N_13694,N_14221);
xor UO_1493 (O_1493,N_13239,N_12369);
nor UO_1494 (O_1494,N_14824,N_14440);
and UO_1495 (O_1495,N_12270,N_12537);
nand UO_1496 (O_1496,N_14231,N_14244);
or UO_1497 (O_1497,N_12584,N_13075);
and UO_1498 (O_1498,N_13002,N_13013);
nand UO_1499 (O_1499,N_13736,N_14698);
nand UO_1500 (O_1500,N_14708,N_13344);
nor UO_1501 (O_1501,N_12697,N_12361);
and UO_1502 (O_1502,N_13662,N_12152);
nand UO_1503 (O_1503,N_12790,N_13898);
nor UO_1504 (O_1504,N_12194,N_13645);
or UO_1505 (O_1505,N_14744,N_12944);
and UO_1506 (O_1506,N_13239,N_13848);
nand UO_1507 (O_1507,N_12744,N_14569);
nand UO_1508 (O_1508,N_12675,N_14030);
or UO_1509 (O_1509,N_14685,N_13205);
nand UO_1510 (O_1510,N_12662,N_14054);
and UO_1511 (O_1511,N_14394,N_13478);
nand UO_1512 (O_1512,N_12032,N_12455);
xor UO_1513 (O_1513,N_14096,N_12628);
nor UO_1514 (O_1514,N_14388,N_14868);
or UO_1515 (O_1515,N_13127,N_13460);
nor UO_1516 (O_1516,N_13151,N_14359);
and UO_1517 (O_1517,N_12860,N_12201);
and UO_1518 (O_1518,N_13882,N_13469);
and UO_1519 (O_1519,N_12208,N_14744);
nor UO_1520 (O_1520,N_14256,N_13309);
nand UO_1521 (O_1521,N_13626,N_12942);
or UO_1522 (O_1522,N_14673,N_12789);
or UO_1523 (O_1523,N_13717,N_13318);
and UO_1524 (O_1524,N_13947,N_12935);
and UO_1525 (O_1525,N_14405,N_14875);
and UO_1526 (O_1526,N_14257,N_12231);
xnor UO_1527 (O_1527,N_13247,N_13318);
xnor UO_1528 (O_1528,N_14663,N_13955);
and UO_1529 (O_1529,N_14027,N_13092);
and UO_1530 (O_1530,N_12230,N_12428);
xnor UO_1531 (O_1531,N_13233,N_14690);
xnor UO_1532 (O_1532,N_12139,N_14767);
nand UO_1533 (O_1533,N_12506,N_13615);
or UO_1534 (O_1534,N_14978,N_12785);
xnor UO_1535 (O_1535,N_14418,N_13650);
or UO_1536 (O_1536,N_14956,N_12452);
or UO_1537 (O_1537,N_14498,N_14013);
nand UO_1538 (O_1538,N_14059,N_12464);
or UO_1539 (O_1539,N_12489,N_12776);
nor UO_1540 (O_1540,N_13613,N_13907);
or UO_1541 (O_1541,N_14943,N_13580);
or UO_1542 (O_1542,N_12421,N_12811);
and UO_1543 (O_1543,N_14714,N_14865);
and UO_1544 (O_1544,N_12876,N_12943);
nand UO_1545 (O_1545,N_14478,N_12945);
nor UO_1546 (O_1546,N_12691,N_14363);
and UO_1547 (O_1547,N_14743,N_14011);
nor UO_1548 (O_1548,N_12031,N_12999);
or UO_1549 (O_1549,N_14889,N_13020);
nand UO_1550 (O_1550,N_13816,N_12364);
nor UO_1551 (O_1551,N_12661,N_13649);
nand UO_1552 (O_1552,N_14726,N_14292);
nor UO_1553 (O_1553,N_12542,N_14965);
nor UO_1554 (O_1554,N_12828,N_12285);
and UO_1555 (O_1555,N_12778,N_13920);
and UO_1556 (O_1556,N_14138,N_14112);
nor UO_1557 (O_1557,N_12200,N_12994);
nand UO_1558 (O_1558,N_13174,N_13948);
nand UO_1559 (O_1559,N_14300,N_14266);
nand UO_1560 (O_1560,N_14132,N_12402);
nand UO_1561 (O_1561,N_13646,N_13865);
nand UO_1562 (O_1562,N_13760,N_12810);
nand UO_1563 (O_1563,N_14491,N_13319);
and UO_1564 (O_1564,N_12796,N_13649);
or UO_1565 (O_1565,N_12465,N_12410);
nor UO_1566 (O_1566,N_13239,N_14894);
and UO_1567 (O_1567,N_13019,N_12921);
nor UO_1568 (O_1568,N_13617,N_12784);
and UO_1569 (O_1569,N_13938,N_14871);
xnor UO_1570 (O_1570,N_14507,N_13121);
and UO_1571 (O_1571,N_14076,N_13495);
or UO_1572 (O_1572,N_13014,N_13204);
nor UO_1573 (O_1573,N_14708,N_12615);
or UO_1574 (O_1574,N_13846,N_12984);
nor UO_1575 (O_1575,N_13475,N_14231);
and UO_1576 (O_1576,N_14046,N_12846);
xor UO_1577 (O_1577,N_14420,N_12320);
xor UO_1578 (O_1578,N_13659,N_12752);
nor UO_1579 (O_1579,N_12969,N_12085);
xnor UO_1580 (O_1580,N_13627,N_14675);
nor UO_1581 (O_1581,N_13276,N_14155);
or UO_1582 (O_1582,N_13114,N_13070);
nand UO_1583 (O_1583,N_14393,N_12243);
nand UO_1584 (O_1584,N_12852,N_12377);
nand UO_1585 (O_1585,N_13997,N_12776);
and UO_1586 (O_1586,N_14072,N_14669);
nor UO_1587 (O_1587,N_14802,N_12117);
nor UO_1588 (O_1588,N_13538,N_12202);
or UO_1589 (O_1589,N_12058,N_13983);
or UO_1590 (O_1590,N_14175,N_14425);
nor UO_1591 (O_1591,N_14214,N_12248);
nand UO_1592 (O_1592,N_14102,N_12258);
nor UO_1593 (O_1593,N_14774,N_13441);
xor UO_1594 (O_1594,N_14581,N_13207);
nand UO_1595 (O_1595,N_14630,N_14121);
or UO_1596 (O_1596,N_12742,N_13300);
or UO_1597 (O_1597,N_12120,N_12992);
and UO_1598 (O_1598,N_14378,N_13626);
nor UO_1599 (O_1599,N_13703,N_12744);
and UO_1600 (O_1600,N_12924,N_13158);
nand UO_1601 (O_1601,N_14008,N_13760);
xor UO_1602 (O_1602,N_14740,N_12082);
nor UO_1603 (O_1603,N_14470,N_14731);
and UO_1604 (O_1604,N_12893,N_12718);
nor UO_1605 (O_1605,N_12845,N_14429);
or UO_1606 (O_1606,N_12101,N_12523);
or UO_1607 (O_1607,N_14063,N_14715);
nand UO_1608 (O_1608,N_14063,N_12874);
nand UO_1609 (O_1609,N_14621,N_14031);
nand UO_1610 (O_1610,N_12560,N_14466);
nor UO_1611 (O_1611,N_12985,N_13572);
and UO_1612 (O_1612,N_13334,N_12861);
or UO_1613 (O_1613,N_12028,N_14585);
or UO_1614 (O_1614,N_13929,N_14011);
nand UO_1615 (O_1615,N_13942,N_14035);
or UO_1616 (O_1616,N_14770,N_14533);
and UO_1617 (O_1617,N_13697,N_13342);
nor UO_1618 (O_1618,N_12253,N_12158);
and UO_1619 (O_1619,N_14644,N_12496);
xnor UO_1620 (O_1620,N_14486,N_13749);
and UO_1621 (O_1621,N_12341,N_12217);
nand UO_1622 (O_1622,N_12157,N_14237);
and UO_1623 (O_1623,N_12519,N_14102);
nand UO_1624 (O_1624,N_12808,N_14012);
nor UO_1625 (O_1625,N_12791,N_12702);
or UO_1626 (O_1626,N_14768,N_14713);
or UO_1627 (O_1627,N_14302,N_14205);
nand UO_1628 (O_1628,N_12067,N_14881);
and UO_1629 (O_1629,N_13129,N_13642);
or UO_1630 (O_1630,N_14219,N_12907);
xor UO_1631 (O_1631,N_14991,N_13034);
xnor UO_1632 (O_1632,N_14610,N_13251);
and UO_1633 (O_1633,N_14594,N_14983);
nand UO_1634 (O_1634,N_14610,N_13949);
nor UO_1635 (O_1635,N_13046,N_12122);
and UO_1636 (O_1636,N_14259,N_12762);
and UO_1637 (O_1637,N_13812,N_14151);
and UO_1638 (O_1638,N_12487,N_14629);
and UO_1639 (O_1639,N_14383,N_12647);
nand UO_1640 (O_1640,N_12208,N_14649);
nor UO_1641 (O_1641,N_13946,N_12608);
nand UO_1642 (O_1642,N_13290,N_13195);
nand UO_1643 (O_1643,N_13410,N_12642);
and UO_1644 (O_1644,N_12013,N_14405);
nor UO_1645 (O_1645,N_12009,N_14492);
or UO_1646 (O_1646,N_12596,N_12689);
nor UO_1647 (O_1647,N_12544,N_12086);
nor UO_1648 (O_1648,N_12017,N_14426);
nand UO_1649 (O_1649,N_13374,N_13390);
nor UO_1650 (O_1650,N_13535,N_12085);
nor UO_1651 (O_1651,N_12926,N_13739);
or UO_1652 (O_1652,N_12041,N_14362);
and UO_1653 (O_1653,N_13605,N_12920);
nand UO_1654 (O_1654,N_12016,N_14775);
nor UO_1655 (O_1655,N_13853,N_12798);
and UO_1656 (O_1656,N_14535,N_12408);
and UO_1657 (O_1657,N_13201,N_13635);
xor UO_1658 (O_1658,N_14502,N_12756);
nand UO_1659 (O_1659,N_14184,N_14132);
nor UO_1660 (O_1660,N_13628,N_14683);
nor UO_1661 (O_1661,N_13483,N_12911);
and UO_1662 (O_1662,N_14347,N_14557);
nand UO_1663 (O_1663,N_14105,N_13517);
nor UO_1664 (O_1664,N_14663,N_12221);
and UO_1665 (O_1665,N_12771,N_13268);
xor UO_1666 (O_1666,N_14242,N_14008);
and UO_1667 (O_1667,N_13193,N_12861);
nor UO_1668 (O_1668,N_13858,N_12110);
or UO_1669 (O_1669,N_14241,N_12473);
or UO_1670 (O_1670,N_14016,N_14097);
nor UO_1671 (O_1671,N_12167,N_13029);
and UO_1672 (O_1672,N_13894,N_12474);
nand UO_1673 (O_1673,N_14416,N_13940);
nor UO_1674 (O_1674,N_13884,N_14027);
nor UO_1675 (O_1675,N_13253,N_13708);
nand UO_1676 (O_1676,N_14246,N_13526);
xor UO_1677 (O_1677,N_12449,N_13316);
nand UO_1678 (O_1678,N_14394,N_13367);
nor UO_1679 (O_1679,N_12280,N_13016);
nor UO_1680 (O_1680,N_13735,N_14105);
and UO_1681 (O_1681,N_12242,N_12357);
nand UO_1682 (O_1682,N_12504,N_12384);
and UO_1683 (O_1683,N_13292,N_14675);
and UO_1684 (O_1684,N_14931,N_14581);
or UO_1685 (O_1685,N_13620,N_14157);
and UO_1686 (O_1686,N_13704,N_12746);
nand UO_1687 (O_1687,N_14344,N_13416);
or UO_1688 (O_1688,N_14363,N_12539);
and UO_1689 (O_1689,N_13490,N_13868);
nor UO_1690 (O_1690,N_13438,N_13853);
and UO_1691 (O_1691,N_12717,N_14162);
nor UO_1692 (O_1692,N_12550,N_13780);
nand UO_1693 (O_1693,N_14072,N_12193);
nor UO_1694 (O_1694,N_13563,N_14555);
or UO_1695 (O_1695,N_14460,N_12384);
or UO_1696 (O_1696,N_14541,N_12393);
nand UO_1697 (O_1697,N_12376,N_13343);
or UO_1698 (O_1698,N_14328,N_13791);
or UO_1699 (O_1699,N_13361,N_12385);
nand UO_1700 (O_1700,N_12116,N_13012);
and UO_1701 (O_1701,N_12647,N_14888);
or UO_1702 (O_1702,N_13911,N_13358);
and UO_1703 (O_1703,N_14035,N_13719);
nand UO_1704 (O_1704,N_12593,N_13462);
nand UO_1705 (O_1705,N_14925,N_14873);
and UO_1706 (O_1706,N_14915,N_13935);
nand UO_1707 (O_1707,N_13698,N_14540);
nand UO_1708 (O_1708,N_13888,N_13399);
and UO_1709 (O_1709,N_13696,N_12149);
and UO_1710 (O_1710,N_14621,N_13464);
or UO_1711 (O_1711,N_12897,N_14786);
xnor UO_1712 (O_1712,N_13597,N_13138);
and UO_1713 (O_1713,N_12565,N_14268);
nor UO_1714 (O_1714,N_13003,N_14002);
and UO_1715 (O_1715,N_14042,N_14191);
nand UO_1716 (O_1716,N_12845,N_14268);
and UO_1717 (O_1717,N_14381,N_13307);
or UO_1718 (O_1718,N_12271,N_13662);
or UO_1719 (O_1719,N_12820,N_12547);
or UO_1720 (O_1720,N_14531,N_13613);
and UO_1721 (O_1721,N_12627,N_14255);
xnor UO_1722 (O_1722,N_13150,N_12377);
nand UO_1723 (O_1723,N_12769,N_13456);
nor UO_1724 (O_1724,N_12846,N_13357);
nor UO_1725 (O_1725,N_13397,N_13051);
nor UO_1726 (O_1726,N_13629,N_13854);
or UO_1727 (O_1727,N_12208,N_14950);
or UO_1728 (O_1728,N_13223,N_14389);
and UO_1729 (O_1729,N_14091,N_12568);
or UO_1730 (O_1730,N_13161,N_12433);
and UO_1731 (O_1731,N_13711,N_12293);
nand UO_1732 (O_1732,N_14573,N_14823);
nand UO_1733 (O_1733,N_13899,N_14513);
and UO_1734 (O_1734,N_14676,N_13162);
and UO_1735 (O_1735,N_14897,N_14542);
and UO_1736 (O_1736,N_13626,N_13321);
nor UO_1737 (O_1737,N_12288,N_14783);
or UO_1738 (O_1738,N_13927,N_14013);
nor UO_1739 (O_1739,N_12350,N_13545);
nor UO_1740 (O_1740,N_14121,N_12133);
nand UO_1741 (O_1741,N_14721,N_14723);
and UO_1742 (O_1742,N_14904,N_12965);
or UO_1743 (O_1743,N_12000,N_12311);
xnor UO_1744 (O_1744,N_12944,N_12440);
and UO_1745 (O_1745,N_13939,N_14450);
nand UO_1746 (O_1746,N_14389,N_13593);
nor UO_1747 (O_1747,N_14236,N_13951);
and UO_1748 (O_1748,N_14893,N_14627);
nor UO_1749 (O_1749,N_14693,N_12405);
nor UO_1750 (O_1750,N_12016,N_13865);
nor UO_1751 (O_1751,N_14791,N_12949);
nand UO_1752 (O_1752,N_14946,N_13939);
and UO_1753 (O_1753,N_12913,N_14053);
or UO_1754 (O_1754,N_14605,N_14884);
xnor UO_1755 (O_1755,N_14555,N_14572);
and UO_1756 (O_1756,N_12411,N_13118);
xnor UO_1757 (O_1757,N_13636,N_12155);
or UO_1758 (O_1758,N_14594,N_14513);
nand UO_1759 (O_1759,N_13047,N_12724);
nor UO_1760 (O_1760,N_12019,N_14987);
nor UO_1761 (O_1761,N_12202,N_12600);
and UO_1762 (O_1762,N_13672,N_13310);
nor UO_1763 (O_1763,N_14179,N_14773);
xor UO_1764 (O_1764,N_14522,N_13183);
or UO_1765 (O_1765,N_13555,N_14235);
nand UO_1766 (O_1766,N_14013,N_14698);
nor UO_1767 (O_1767,N_12667,N_13606);
nand UO_1768 (O_1768,N_13198,N_14445);
nand UO_1769 (O_1769,N_12563,N_14968);
and UO_1770 (O_1770,N_14357,N_12968);
nand UO_1771 (O_1771,N_12845,N_14242);
or UO_1772 (O_1772,N_13043,N_12942);
nor UO_1773 (O_1773,N_14155,N_12702);
nand UO_1774 (O_1774,N_14452,N_14943);
or UO_1775 (O_1775,N_12007,N_14161);
or UO_1776 (O_1776,N_14331,N_14582);
xor UO_1777 (O_1777,N_12066,N_13976);
nor UO_1778 (O_1778,N_14570,N_12064);
xor UO_1779 (O_1779,N_12508,N_14245);
or UO_1780 (O_1780,N_12935,N_14790);
xnor UO_1781 (O_1781,N_12511,N_12690);
nand UO_1782 (O_1782,N_13516,N_12114);
xor UO_1783 (O_1783,N_12137,N_12209);
nand UO_1784 (O_1784,N_14911,N_13027);
nor UO_1785 (O_1785,N_14184,N_12702);
xnor UO_1786 (O_1786,N_14463,N_12990);
nor UO_1787 (O_1787,N_14482,N_12287);
nand UO_1788 (O_1788,N_14914,N_14833);
nor UO_1789 (O_1789,N_12600,N_14415);
or UO_1790 (O_1790,N_13717,N_14640);
nand UO_1791 (O_1791,N_14501,N_12968);
xor UO_1792 (O_1792,N_12421,N_12526);
nor UO_1793 (O_1793,N_14767,N_13396);
or UO_1794 (O_1794,N_12685,N_14122);
nor UO_1795 (O_1795,N_14962,N_13486);
nand UO_1796 (O_1796,N_13706,N_13199);
nor UO_1797 (O_1797,N_14246,N_14104);
or UO_1798 (O_1798,N_13295,N_14193);
nor UO_1799 (O_1799,N_13310,N_14406);
nand UO_1800 (O_1800,N_14186,N_14671);
and UO_1801 (O_1801,N_14240,N_14926);
nand UO_1802 (O_1802,N_14289,N_12991);
xor UO_1803 (O_1803,N_14210,N_14955);
or UO_1804 (O_1804,N_13299,N_12277);
nor UO_1805 (O_1805,N_14786,N_13156);
and UO_1806 (O_1806,N_14137,N_12221);
nand UO_1807 (O_1807,N_12842,N_13250);
nand UO_1808 (O_1808,N_12004,N_12667);
xor UO_1809 (O_1809,N_14404,N_14174);
nand UO_1810 (O_1810,N_12208,N_14216);
nor UO_1811 (O_1811,N_13177,N_12493);
or UO_1812 (O_1812,N_14401,N_14693);
xnor UO_1813 (O_1813,N_13175,N_13082);
nand UO_1814 (O_1814,N_13265,N_13012);
xor UO_1815 (O_1815,N_14923,N_14714);
nand UO_1816 (O_1816,N_14220,N_13937);
nor UO_1817 (O_1817,N_13814,N_13548);
nor UO_1818 (O_1818,N_13243,N_12841);
or UO_1819 (O_1819,N_14116,N_14663);
nor UO_1820 (O_1820,N_13118,N_14326);
or UO_1821 (O_1821,N_13915,N_13972);
nor UO_1822 (O_1822,N_12958,N_13201);
nor UO_1823 (O_1823,N_14735,N_12077);
nand UO_1824 (O_1824,N_13965,N_13729);
nand UO_1825 (O_1825,N_13193,N_12136);
nor UO_1826 (O_1826,N_13334,N_12739);
or UO_1827 (O_1827,N_12154,N_13968);
nor UO_1828 (O_1828,N_14572,N_12390);
or UO_1829 (O_1829,N_12803,N_12258);
nand UO_1830 (O_1830,N_14762,N_13337);
xnor UO_1831 (O_1831,N_13642,N_14508);
nor UO_1832 (O_1832,N_13207,N_12730);
and UO_1833 (O_1833,N_12681,N_12649);
or UO_1834 (O_1834,N_12043,N_12432);
nand UO_1835 (O_1835,N_13453,N_14738);
nor UO_1836 (O_1836,N_12891,N_12452);
nand UO_1837 (O_1837,N_13096,N_14461);
nor UO_1838 (O_1838,N_14705,N_14554);
nand UO_1839 (O_1839,N_13078,N_12009);
and UO_1840 (O_1840,N_13878,N_12052);
nor UO_1841 (O_1841,N_14526,N_14644);
or UO_1842 (O_1842,N_13869,N_12577);
nor UO_1843 (O_1843,N_14295,N_13938);
nand UO_1844 (O_1844,N_12242,N_13912);
nand UO_1845 (O_1845,N_13866,N_12029);
xnor UO_1846 (O_1846,N_13061,N_12362);
and UO_1847 (O_1847,N_14442,N_12840);
or UO_1848 (O_1848,N_12793,N_13403);
nand UO_1849 (O_1849,N_12149,N_12203);
and UO_1850 (O_1850,N_14372,N_14311);
nor UO_1851 (O_1851,N_12316,N_12310);
or UO_1852 (O_1852,N_12585,N_14249);
and UO_1853 (O_1853,N_13612,N_13551);
nand UO_1854 (O_1854,N_14815,N_13771);
nor UO_1855 (O_1855,N_14543,N_14930);
nor UO_1856 (O_1856,N_14990,N_14126);
and UO_1857 (O_1857,N_14665,N_14716);
nand UO_1858 (O_1858,N_12014,N_12001);
xor UO_1859 (O_1859,N_14746,N_13276);
or UO_1860 (O_1860,N_13680,N_12522);
and UO_1861 (O_1861,N_13974,N_12791);
and UO_1862 (O_1862,N_12952,N_14981);
and UO_1863 (O_1863,N_14543,N_13877);
xor UO_1864 (O_1864,N_13247,N_12030);
nand UO_1865 (O_1865,N_14379,N_12795);
nor UO_1866 (O_1866,N_12724,N_12241);
nand UO_1867 (O_1867,N_14654,N_14671);
or UO_1868 (O_1868,N_14463,N_12128);
nand UO_1869 (O_1869,N_13968,N_14751);
nor UO_1870 (O_1870,N_14179,N_14385);
xnor UO_1871 (O_1871,N_13398,N_14981);
xnor UO_1872 (O_1872,N_14795,N_14057);
or UO_1873 (O_1873,N_12757,N_12946);
nor UO_1874 (O_1874,N_12242,N_12571);
nor UO_1875 (O_1875,N_12665,N_13117);
nor UO_1876 (O_1876,N_14057,N_12418);
and UO_1877 (O_1877,N_12677,N_12310);
xor UO_1878 (O_1878,N_12329,N_12218);
nand UO_1879 (O_1879,N_12578,N_13681);
nand UO_1880 (O_1880,N_12661,N_12422);
nand UO_1881 (O_1881,N_14104,N_12122);
nand UO_1882 (O_1882,N_13709,N_14705);
and UO_1883 (O_1883,N_12305,N_14623);
and UO_1884 (O_1884,N_14924,N_14332);
and UO_1885 (O_1885,N_14758,N_12839);
and UO_1886 (O_1886,N_14877,N_14925);
nor UO_1887 (O_1887,N_12552,N_13844);
or UO_1888 (O_1888,N_14809,N_13060);
and UO_1889 (O_1889,N_14378,N_13434);
nor UO_1890 (O_1890,N_14170,N_13453);
and UO_1891 (O_1891,N_13729,N_13245);
nand UO_1892 (O_1892,N_13522,N_14887);
nand UO_1893 (O_1893,N_12871,N_14067);
nand UO_1894 (O_1894,N_14063,N_12349);
nor UO_1895 (O_1895,N_13853,N_14397);
nand UO_1896 (O_1896,N_14512,N_14724);
and UO_1897 (O_1897,N_14664,N_13759);
and UO_1898 (O_1898,N_14684,N_13748);
or UO_1899 (O_1899,N_12470,N_12632);
or UO_1900 (O_1900,N_13452,N_14193);
or UO_1901 (O_1901,N_12761,N_13504);
or UO_1902 (O_1902,N_13346,N_12217);
nor UO_1903 (O_1903,N_14878,N_13630);
and UO_1904 (O_1904,N_14725,N_12292);
nand UO_1905 (O_1905,N_12671,N_14733);
nand UO_1906 (O_1906,N_12371,N_13927);
or UO_1907 (O_1907,N_14786,N_14171);
nand UO_1908 (O_1908,N_13760,N_13939);
or UO_1909 (O_1909,N_14099,N_14600);
or UO_1910 (O_1910,N_12471,N_12245);
xnor UO_1911 (O_1911,N_12477,N_13882);
nor UO_1912 (O_1912,N_12181,N_13501);
nor UO_1913 (O_1913,N_12429,N_14519);
or UO_1914 (O_1914,N_14942,N_12171);
nor UO_1915 (O_1915,N_12870,N_14279);
or UO_1916 (O_1916,N_13362,N_14756);
or UO_1917 (O_1917,N_12019,N_14261);
xnor UO_1918 (O_1918,N_13455,N_12759);
nor UO_1919 (O_1919,N_12325,N_12767);
or UO_1920 (O_1920,N_12311,N_14985);
or UO_1921 (O_1921,N_12762,N_14278);
nor UO_1922 (O_1922,N_14916,N_13204);
nand UO_1923 (O_1923,N_12374,N_13257);
or UO_1924 (O_1924,N_14255,N_12996);
and UO_1925 (O_1925,N_12701,N_13757);
nor UO_1926 (O_1926,N_14719,N_12792);
nor UO_1927 (O_1927,N_13604,N_12068);
nor UO_1928 (O_1928,N_14710,N_14885);
or UO_1929 (O_1929,N_12109,N_13957);
nand UO_1930 (O_1930,N_13667,N_12841);
or UO_1931 (O_1931,N_12649,N_12411);
nor UO_1932 (O_1932,N_14806,N_14034);
or UO_1933 (O_1933,N_12762,N_12654);
or UO_1934 (O_1934,N_13297,N_12806);
nor UO_1935 (O_1935,N_13195,N_12556);
and UO_1936 (O_1936,N_12334,N_13380);
or UO_1937 (O_1937,N_13688,N_14194);
and UO_1938 (O_1938,N_12181,N_14877);
and UO_1939 (O_1939,N_14553,N_14853);
and UO_1940 (O_1940,N_12378,N_13069);
nor UO_1941 (O_1941,N_14971,N_13161);
or UO_1942 (O_1942,N_14284,N_14240);
or UO_1943 (O_1943,N_12617,N_13097);
nor UO_1944 (O_1944,N_14473,N_14530);
and UO_1945 (O_1945,N_12508,N_13265);
xor UO_1946 (O_1946,N_13443,N_14674);
nor UO_1947 (O_1947,N_12367,N_12045);
and UO_1948 (O_1948,N_12154,N_14764);
and UO_1949 (O_1949,N_12852,N_13547);
and UO_1950 (O_1950,N_13893,N_12801);
nor UO_1951 (O_1951,N_13190,N_14895);
and UO_1952 (O_1952,N_13565,N_14828);
nor UO_1953 (O_1953,N_14238,N_12359);
nor UO_1954 (O_1954,N_13263,N_12502);
or UO_1955 (O_1955,N_14417,N_14642);
nand UO_1956 (O_1956,N_14837,N_14947);
or UO_1957 (O_1957,N_12655,N_14896);
and UO_1958 (O_1958,N_13299,N_12448);
or UO_1959 (O_1959,N_12205,N_12147);
nand UO_1960 (O_1960,N_12455,N_12776);
nand UO_1961 (O_1961,N_13421,N_14274);
and UO_1962 (O_1962,N_14659,N_13893);
nand UO_1963 (O_1963,N_14853,N_12318);
or UO_1964 (O_1964,N_12666,N_14345);
or UO_1965 (O_1965,N_13577,N_13798);
or UO_1966 (O_1966,N_13149,N_13544);
or UO_1967 (O_1967,N_14827,N_14742);
nor UO_1968 (O_1968,N_14235,N_12614);
or UO_1969 (O_1969,N_13834,N_12593);
and UO_1970 (O_1970,N_14857,N_12015);
and UO_1971 (O_1971,N_13334,N_14258);
and UO_1972 (O_1972,N_14582,N_12149);
and UO_1973 (O_1973,N_12815,N_13667);
nand UO_1974 (O_1974,N_12079,N_12017);
and UO_1975 (O_1975,N_14986,N_12580);
and UO_1976 (O_1976,N_13595,N_12771);
and UO_1977 (O_1977,N_14427,N_12620);
nand UO_1978 (O_1978,N_13083,N_12077);
nor UO_1979 (O_1979,N_14386,N_12627);
or UO_1980 (O_1980,N_12966,N_13914);
nor UO_1981 (O_1981,N_12103,N_12459);
nor UO_1982 (O_1982,N_12832,N_13419);
and UO_1983 (O_1983,N_14888,N_12776);
or UO_1984 (O_1984,N_12020,N_12442);
and UO_1985 (O_1985,N_14071,N_13763);
and UO_1986 (O_1986,N_14058,N_12188);
nor UO_1987 (O_1987,N_14618,N_13414);
nand UO_1988 (O_1988,N_13035,N_14061);
or UO_1989 (O_1989,N_13939,N_13380);
nor UO_1990 (O_1990,N_14096,N_12428);
nand UO_1991 (O_1991,N_12436,N_14947);
and UO_1992 (O_1992,N_13431,N_13171);
nor UO_1993 (O_1993,N_12113,N_13161);
or UO_1994 (O_1994,N_12408,N_14903);
nand UO_1995 (O_1995,N_12279,N_13065);
and UO_1996 (O_1996,N_13064,N_14639);
or UO_1997 (O_1997,N_13280,N_12707);
nor UO_1998 (O_1998,N_12156,N_12678);
and UO_1999 (O_1999,N_14276,N_12967);
endmodule