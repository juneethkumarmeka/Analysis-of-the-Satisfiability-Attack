module basic_2500_25000_3000_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_872,In_860);
xor U1 (N_1,In_2149,In_679);
or U2 (N_2,In_1171,In_1853);
xor U3 (N_3,In_931,In_77);
nor U4 (N_4,In_1566,In_1406);
or U5 (N_5,In_2489,In_792);
nand U6 (N_6,In_1060,In_1900);
nor U7 (N_7,In_1573,In_2417);
or U8 (N_8,In_2407,In_342);
nand U9 (N_9,In_2441,In_81);
and U10 (N_10,In_983,In_51);
nor U11 (N_11,In_1798,In_423);
nor U12 (N_12,In_63,In_1950);
or U13 (N_13,In_958,In_208);
or U14 (N_14,In_743,In_1311);
or U15 (N_15,In_2446,In_583);
xor U16 (N_16,In_1731,In_1021);
xnor U17 (N_17,In_432,In_2207);
nor U18 (N_18,In_950,In_998);
and U19 (N_19,In_1807,In_2364);
xor U20 (N_20,In_2223,In_869);
and U21 (N_21,In_1939,In_1961);
nor U22 (N_22,In_1527,In_2112);
nand U23 (N_23,In_692,In_1804);
or U24 (N_24,In_1735,In_121);
or U25 (N_25,In_1622,In_2444);
or U26 (N_26,In_766,In_1334);
nand U27 (N_27,In_1193,In_1351);
or U28 (N_28,In_1941,In_458);
and U29 (N_29,In_153,In_443);
nand U30 (N_30,In_1500,In_191);
and U31 (N_31,In_532,In_176);
or U32 (N_32,In_1958,In_408);
or U33 (N_33,In_1817,In_1238);
and U34 (N_34,In_363,In_1671);
nand U35 (N_35,In_1448,In_1197);
xnor U36 (N_36,In_1858,In_2042);
nand U37 (N_37,In_2408,In_1106);
xnor U38 (N_38,In_635,In_1675);
or U39 (N_39,In_435,In_2015);
nor U40 (N_40,In_317,In_638);
nand U41 (N_41,In_225,In_670);
and U42 (N_42,In_899,In_1755);
xor U43 (N_43,In_2063,In_2142);
nand U44 (N_44,In_2495,In_1584);
nand U45 (N_45,In_86,In_298);
nor U46 (N_46,In_1885,In_337);
and U47 (N_47,In_1149,In_1418);
and U48 (N_48,In_976,In_1157);
and U49 (N_49,In_2006,In_2272);
nand U50 (N_50,In_555,In_1367);
and U51 (N_51,In_207,In_2114);
xnor U52 (N_52,In_1013,In_46);
nand U53 (N_53,In_1844,In_1672);
or U54 (N_54,In_1983,In_1813);
xnor U55 (N_55,In_2439,In_358);
xor U56 (N_56,In_1727,In_1923);
or U57 (N_57,In_1342,In_2175);
and U58 (N_58,In_2254,In_2422);
nor U59 (N_59,In_1,In_29);
nor U60 (N_60,In_346,In_1525);
xor U61 (N_61,In_463,In_1370);
and U62 (N_62,In_951,In_185);
nor U63 (N_63,In_101,In_372);
or U64 (N_64,In_988,In_1291);
nand U65 (N_65,In_1806,In_857);
or U66 (N_66,In_634,In_406);
nor U67 (N_67,In_1452,In_464);
nand U68 (N_68,In_1666,In_152);
nand U69 (N_69,In_791,In_780);
and U70 (N_70,In_130,In_851);
nor U71 (N_71,In_1563,In_498);
or U72 (N_72,In_1933,In_2125);
xor U73 (N_73,In_1786,In_1619);
nor U74 (N_74,In_420,In_1594);
nand U75 (N_75,In_1078,In_833);
and U76 (N_76,In_1092,In_2371);
and U77 (N_77,In_771,In_1372);
and U78 (N_78,In_182,In_1456);
and U79 (N_79,In_1582,In_466);
or U80 (N_80,In_2413,In_345);
and U81 (N_81,In_1419,In_90);
xnor U82 (N_82,In_1907,In_1832);
xnor U83 (N_83,In_1232,In_1679);
xnor U84 (N_84,In_1052,In_37);
xor U85 (N_85,In_737,In_1898);
or U86 (N_86,In_278,In_841);
and U87 (N_87,In_48,In_687);
and U88 (N_88,In_2454,In_1026);
nor U89 (N_89,In_1000,In_897);
and U90 (N_90,In_2206,In_2294);
and U91 (N_91,In_1315,In_883);
and U92 (N_92,In_132,In_485);
and U93 (N_93,In_91,In_1951);
or U94 (N_94,In_401,In_1842);
or U95 (N_95,In_1760,In_1324);
nand U96 (N_96,In_2434,In_1240);
and U97 (N_97,In_184,In_1914);
nand U98 (N_98,In_2067,In_1880);
nor U99 (N_99,In_2470,In_2193);
nor U100 (N_100,In_217,In_285);
xor U101 (N_101,In_172,In_2350);
and U102 (N_102,In_539,In_1191);
nor U103 (N_103,In_399,In_531);
xor U104 (N_104,In_1765,In_1190);
nand U105 (N_105,In_1940,In_740);
nand U106 (N_106,In_202,In_1520);
xnor U107 (N_107,In_965,In_1710);
or U108 (N_108,In_331,In_1720);
or U109 (N_109,In_327,In_2004);
xnor U110 (N_110,In_2411,In_350);
and U111 (N_111,In_255,In_144);
nand U112 (N_112,In_2136,In_992);
or U113 (N_113,In_215,In_667);
nand U114 (N_114,In_1131,In_440);
or U115 (N_115,In_2382,In_666);
nand U116 (N_116,In_1423,In_1398);
and U117 (N_117,In_1467,In_525);
and U118 (N_118,In_122,In_1553);
or U119 (N_119,In_1850,In_753);
and U120 (N_120,In_1641,In_307);
and U121 (N_121,In_123,In_1773);
and U122 (N_122,In_1975,In_112);
nor U123 (N_123,In_1705,In_2076);
or U124 (N_124,In_1373,In_199);
nand U125 (N_125,In_2440,In_2260);
nor U126 (N_126,In_2266,In_158);
xor U127 (N_127,In_1690,In_419);
nand U128 (N_128,In_1970,In_2462);
and U129 (N_129,In_304,In_287);
and U130 (N_130,In_1884,In_703);
nor U131 (N_131,In_368,In_714);
xnor U132 (N_132,In_1667,In_1175);
xnor U133 (N_133,In_716,In_1460);
and U134 (N_134,In_2017,In_603);
or U135 (N_135,In_561,In_696);
xnor U136 (N_136,In_460,In_1123);
and U137 (N_137,In_1437,In_2262);
or U138 (N_138,In_492,In_529);
xnor U139 (N_139,In_2134,In_1545);
xnor U140 (N_140,In_2152,In_1200);
or U141 (N_141,In_2154,In_1924);
nand U142 (N_142,In_236,In_1287);
or U143 (N_143,In_2397,In_2164);
nor U144 (N_144,In_930,In_943);
and U145 (N_145,In_1080,In_1736);
nand U146 (N_146,In_1426,In_2459);
xnor U147 (N_147,In_1475,In_516);
xnor U148 (N_148,In_1103,In_1852);
xnor U149 (N_149,In_827,In_1715);
or U150 (N_150,In_1177,In_302);
or U151 (N_151,In_767,In_2079);
or U152 (N_152,In_1361,In_247);
and U153 (N_153,In_545,In_418);
xor U154 (N_154,In_542,In_816);
and U155 (N_155,In_654,In_248);
nand U156 (N_156,In_1082,In_709);
nand U157 (N_157,In_1102,In_607);
nand U158 (N_158,In_1024,In_1045);
xor U159 (N_159,In_1274,In_1857);
and U160 (N_160,In_1308,In_396);
xor U161 (N_161,In_1255,In_1020);
and U162 (N_162,In_888,In_1101);
and U163 (N_163,In_818,In_2131);
xnor U164 (N_164,In_2068,In_2346);
nand U165 (N_165,In_1586,In_486);
or U166 (N_166,In_2200,In_1038);
nor U167 (N_167,In_711,In_1389);
or U168 (N_168,In_1574,In_2299);
xnor U169 (N_169,In_1336,In_1058);
and U170 (N_170,In_2121,In_397);
or U171 (N_171,In_2003,In_413);
nand U172 (N_172,In_328,In_633);
xor U173 (N_173,In_40,In_839);
or U174 (N_174,In_1495,In_2415);
or U175 (N_175,In_2248,In_1347);
and U176 (N_176,In_237,In_1963);
nor U177 (N_177,In_1658,In_2107);
nor U178 (N_178,In_1906,In_656);
or U179 (N_179,In_871,In_1911);
and U180 (N_180,In_2265,In_415);
xor U181 (N_181,In_2324,In_1791);
xor U182 (N_182,In_1615,In_447);
nand U183 (N_183,In_1415,In_273);
nand U184 (N_184,In_1323,In_1638);
or U185 (N_185,In_365,In_54);
xor U186 (N_186,In_1579,In_610);
nor U187 (N_187,In_102,In_22);
nor U188 (N_188,In_1986,In_741);
nor U189 (N_189,In_1879,In_1381);
and U190 (N_190,In_837,In_2332);
nor U191 (N_191,In_1051,In_470);
or U192 (N_192,In_2330,In_1814);
or U193 (N_193,In_2051,In_918);
or U194 (N_194,In_2080,In_1386);
xor U195 (N_195,In_1778,In_1442);
nand U196 (N_196,In_1141,In_2030);
xnor U197 (N_197,In_1547,In_1449);
nand U198 (N_198,In_1805,In_659);
or U199 (N_199,In_1833,In_1698);
nor U200 (N_200,In_1492,In_1481);
or U201 (N_201,In_1083,In_1030);
and U202 (N_202,In_763,In_1624);
nand U203 (N_203,In_619,In_186);
or U204 (N_204,In_524,In_2116);
nor U205 (N_205,In_1830,In_626);
nand U206 (N_206,In_1823,In_1496);
nor U207 (N_207,In_230,In_1144);
xnor U208 (N_208,In_1510,In_836);
nand U209 (N_209,In_734,In_1075);
xor U210 (N_210,In_1212,In_842);
xor U211 (N_211,In_873,In_884);
xor U212 (N_212,In_1578,In_523);
xnor U213 (N_213,In_866,In_2102);
xnor U214 (N_214,In_1790,In_1338);
nor U215 (N_215,In_1189,In_1077);
nor U216 (N_216,In_280,In_921);
or U217 (N_217,In_1304,In_2420);
xnor U218 (N_218,In_2348,In_1081);
xnor U219 (N_219,In_1378,In_1726);
nand U220 (N_220,In_2232,In_2428);
nand U221 (N_221,In_2479,In_919);
nand U222 (N_222,In_1974,In_675);
xnor U223 (N_223,In_1743,In_658);
and U224 (N_224,In_2442,In_2061);
xnor U225 (N_225,In_1922,In_246);
nor U226 (N_226,In_822,In_1241);
or U227 (N_227,In_23,In_1507);
nor U228 (N_228,In_2176,In_50);
nor U229 (N_229,In_800,In_1623);
or U230 (N_230,In_575,In_2409);
or U231 (N_231,In_2401,In_1952);
and U232 (N_232,In_731,In_1919);
nand U233 (N_233,In_1503,In_394);
xnor U234 (N_234,In_2233,In_128);
and U235 (N_235,In_1214,In_162);
or U236 (N_236,In_2386,In_2481);
nor U237 (N_237,In_2438,In_2424);
xor U238 (N_238,In_1027,In_1136);
or U239 (N_239,In_1668,In_2383);
or U240 (N_240,In_2072,In_1905);
xor U241 (N_241,In_430,In_966);
nand U242 (N_242,In_2201,In_1712);
nand U243 (N_243,In_2421,In_349);
and U244 (N_244,In_266,In_326);
nand U245 (N_245,In_1376,In_2240);
or U246 (N_246,In_2243,In_563);
and U247 (N_247,In_1938,In_2000);
nor U248 (N_248,In_1687,In_2054);
and U249 (N_249,In_2419,In_863);
or U250 (N_250,In_2297,In_522);
nor U251 (N_251,In_621,In_1816);
nand U252 (N_252,In_2029,In_233);
xnor U253 (N_253,In_1549,In_2037);
nor U254 (N_254,In_1607,In_1569);
nor U255 (N_255,In_1462,In_2141);
xor U256 (N_256,In_2021,In_935);
and U257 (N_257,In_499,In_12);
xor U258 (N_258,In_438,In_2331);
nor U259 (N_259,In_1133,In_1697);
nor U260 (N_260,In_39,In_2282);
or U261 (N_261,In_1180,In_2216);
nand U262 (N_262,In_2322,In_171);
nor U263 (N_263,In_682,In_794);
and U264 (N_264,In_1886,In_1368);
nor U265 (N_265,In_457,In_1068);
xnor U266 (N_266,In_469,In_125);
or U267 (N_267,In_650,In_437);
and U268 (N_268,In_214,In_807);
nand U269 (N_269,In_1856,In_712);
or U270 (N_270,In_671,In_1352);
nand U271 (N_271,In_1427,In_288);
nand U272 (N_272,In_1395,In_1004);
nand U273 (N_273,In_513,In_209);
or U274 (N_274,In_2335,In_1978);
nor U275 (N_275,In_1680,In_1770);
xnor U276 (N_276,In_954,In_1965);
or U277 (N_277,In_1776,In_1132);
nand U278 (N_278,In_1673,In_790);
or U279 (N_279,In_1236,In_1223);
xnor U280 (N_280,In_473,In_1440);
or U281 (N_281,In_721,In_1069);
nand U282 (N_282,In_1616,In_1454);
nand U283 (N_283,In_749,In_1931);
nor U284 (N_284,In_204,In_2052);
or U285 (N_285,In_19,In_197);
or U286 (N_286,In_1966,In_425);
or U287 (N_287,In_136,In_1100);
or U288 (N_288,In_1916,In_1247);
xnor U289 (N_289,In_1725,In_526);
nor U290 (N_290,In_572,In_1526);
xor U291 (N_291,In_1788,In_1815);
and U292 (N_292,In_2448,In_3);
xnor U293 (N_293,In_1413,In_1262);
xnor U294 (N_294,In_681,In_2097);
nand U295 (N_295,In_1493,In_964);
nand U296 (N_296,In_2115,In_110);
nor U297 (N_297,In_616,In_1650);
nand U298 (N_298,In_2086,In_2416);
nand U299 (N_299,In_2089,In_1016);
xnor U300 (N_300,In_926,In_1126);
and U301 (N_301,In_1565,In_375);
nor U302 (N_302,In_2473,In_722);
xor U303 (N_303,In_109,In_1178);
or U304 (N_304,In_643,In_874);
nor U305 (N_305,In_1895,In_1837);
xor U306 (N_306,In_10,In_284);
nor U307 (N_307,In_165,In_2098);
and U308 (N_308,In_1618,In_1359);
and U309 (N_309,In_632,In_1990);
or U310 (N_310,In_174,In_95);
xnor U311 (N_311,In_2437,In_1882);
or U312 (N_312,In_953,In_16);
xnor U313 (N_313,In_330,In_79);
xor U314 (N_314,In_1337,In_2393);
nor U315 (N_315,In_1548,In_2226);
nand U316 (N_316,In_1003,In_1992);
or U317 (N_317,In_75,In_2083);
and U318 (N_318,In_1903,In_2179);
or U319 (N_319,In_2339,In_2399);
or U320 (N_320,In_2341,In_2038);
nor U321 (N_321,In_1766,In_187);
and U322 (N_322,In_496,In_343);
and U323 (N_323,In_1560,In_891);
nor U324 (N_324,In_1872,In_798);
xor U325 (N_325,In_520,In_1756);
xor U326 (N_326,In_892,In_489);
xnor U327 (N_327,In_454,In_35);
or U328 (N_328,In_1982,In_894);
or U329 (N_329,In_1320,In_757);
nand U330 (N_330,In_713,In_1384);
and U331 (N_331,In_1487,In_2129);
or U332 (N_332,In_2047,In_85);
nand U333 (N_333,In_1195,In_488);
nor U334 (N_334,In_2120,In_2135);
xnor U335 (N_335,In_2103,In_221);
nor U336 (N_336,In_1758,In_427);
nor U337 (N_337,In_547,In_1581);
and U338 (N_338,In_1264,In_2188);
nor U339 (N_339,In_1237,In_1501);
xor U340 (N_340,In_2453,In_1301);
nand U341 (N_341,In_571,In_2334);
nor U342 (N_342,In_1310,In_1637);
nand U343 (N_343,In_2106,In_1944);
or U344 (N_344,In_625,In_242);
and U345 (N_345,In_831,In_502);
xor U346 (N_346,In_710,In_1403);
nor U347 (N_347,In_1828,In_1119);
nor U348 (N_348,In_213,In_927);
nor U349 (N_349,In_678,In_517);
and U350 (N_350,In_2212,In_1523);
nand U351 (N_351,In_809,In_1404);
or U352 (N_352,In_846,In_1993);
or U353 (N_353,In_360,In_1091);
nand U354 (N_354,In_2259,In_1929);
nor U355 (N_355,In_505,In_459);
xor U356 (N_356,In_2325,In_1011);
xor U357 (N_357,In_1685,In_2363);
or U358 (N_358,In_2249,In_404);
xor U359 (N_359,In_824,In_87);
nand U360 (N_360,In_1847,In_728);
xnor U361 (N_361,In_1151,In_1893);
or U362 (N_362,In_1818,In_584);
or U363 (N_363,In_503,In_937);
or U364 (N_364,In_108,In_674);
xnor U365 (N_365,In_2251,In_7);
nor U366 (N_366,In_1665,In_1401);
or U367 (N_367,In_2264,In_2155);
nor U368 (N_368,In_407,In_1709);
nor U369 (N_369,In_1216,In_2392);
nand U370 (N_370,In_1250,In_2447);
and U371 (N_371,In_1787,In_1009);
xor U372 (N_372,In_2192,In_2485);
xor U373 (N_373,In_1887,In_2309);
or U374 (N_374,In_1782,In_758);
nor U375 (N_375,In_1994,In_777);
xnor U376 (N_376,In_2379,In_1261);
nand U377 (N_377,In_2190,In_647);
and U378 (N_378,In_1112,In_1087);
nor U379 (N_379,In_985,In_1670);
or U380 (N_380,In_979,In_1686);
xnor U381 (N_381,In_2242,In_1445);
xor U382 (N_382,In_1848,In_557);
nand U383 (N_383,In_868,In_854);
and U384 (N_384,In_989,In_835);
and U385 (N_385,In_2234,In_1774);
xor U386 (N_386,In_2291,In_701);
xnor U387 (N_387,In_968,In_2024);
and U388 (N_388,In_88,In_1985);
nand U389 (N_389,In_795,In_1346);
or U390 (N_390,In_1589,In_1871);
xnor U391 (N_391,In_668,In_1265);
nand U392 (N_392,In_1278,In_482);
nor U393 (N_393,In_693,In_2443);
nor U394 (N_394,In_944,In_1194);
or U395 (N_395,In_49,In_506);
nand U396 (N_396,In_1821,In_1646);
nand U397 (N_397,In_1256,In_746);
nand U398 (N_398,In_1964,In_356);
and U399 (N_399,In_2238,In_240);
and U400 (N_400,In_1533,In_1785);
nor U401 (N_401,In_1438,In_1235);
nor U402 (N_402,In_1831,In_2378);
xnor U403 (N_403,In_243,In_1161);
nand U404 (N_404,In_803,In_289);
nand U405 (N_405,In_120,In_388);
nor U406 (N_406,In_2261,In_393);
nor U407 (N_407,In_1738,In_760);
nand U408 (N_408,In_1170,In_2214);
nand U409 (N_409,In_1228,In_694);
nor U410 (N_410,In_198,In_2170);
or U411 (N_411,In_1797,In_1834);
or U412 (N_412,In_323,In_1097);
nand U413 (N_413,In_880,In_817);
nand U414 (N_414,In_861,In_1312);
nand U415 (N_415,In_1629,In_2314);
and U416 (N_416,In_476,In_62);
and U417 (N_417,In_774,In_1459);
xor U418 (N_418,In_471,In_259);
and U419 (N_419,In_1991,In_1407);
and U420 (N_420,In_1322,In_1281);
xor U421 (N_421,In_550,In_2405);
xnor U422 (N_422,In_1105,In_1759);
or U423 (N_423,In_468,In_959);
nand U424 (N_424,In_957,In_2498);
xor U425 (N_425,In_751,In_1450);
nand U426 (N_426,In_73,In_380);
nand U427 (N_427,In_1702,In_2491);
and U428 (N_428,In_453,In_2285);
nand U429 (N_429,In_684,In_1913);
or U430 (N_430,In_422,In_1962);
nor U431 (N_431,In_2113,In_2287);
xor U432 (N_432,In_131,In_2457);
nand U433 (N_433,In_84,In_1321);
or U434 (N_434,In_223,In_1851);
and U435 (N_435,In_2053,In_1657);
nand U436 (N_436,In_412,In_2445);
and U437 (N_437,In_400,In_664);
nand U438 (N_438,In_1683,In_739);
xnor U439 (N_439,In_612,In_1703);
nor U440 (N_440,In_878,In_773);
nand U441 (N_441,In_2384,In_986);
and U442 (N_442,In_2169,In_1762);
xor U443 (N_443,In_2403,In_843);
or U444 (N_444,In_2245,In_613);
nor U445 (N_445,In_456,In_1339);
xnor U446 (N_446,In_995,In_2349);
xor U447 (N_447,In_1267,In_2369);
and U448 (N_448,In_1639,In_697);
nor U449 (N_449,In_1570,In_723);
nor U450 (N_450,In_1692,In_1752);
or U451 (N_451,In_2119,In_1143);
nor U452 (N_452,In_1433,In_922);
xor U453 (N_453,In_1543,In_2108);
xnor U454 (N_454,In_1122,In_47);
xor U455 (N_455,In_1681,In_2241);
nor U456 (N_456,In_590,In_2090);
nor U457 (N_457,In_1789,In_1676);
and U458 (N_458,In_1904,In_885);
and U459 (N_459,In_219,In_410);
xnor U460 (N_460,In_2497,In_1971);
nand U461 (N_461,In_662,In_821);
xor U462 (N_462,In_2163,In_1253);
nand U463 (N_463,In_1414,In_1019);
nor U464 (N_464,In_1358,In_2064);
or U465 (N_465,In_2123,In_1208);
xnor U466 (N_466,In_494,In_352);
or U467 (N_467,In_805,In_752);
xor U468 (N_468,In_942,In_1239);
nor U469 (N_469,In_170,In_1432);
nand U470 (N_470,In_1822,In_1585);
xor U471 (N_471,In_535,In_1204);
nand U472 (N_472,In_1572,In_1561);
nor U473 (N_473,In_1173,In_1059);
nand U474 (N_474,In_759,In_1096);
or U475 (N_475,In_778,In_1063);
xor U476 (N_476,In_1205,In_1443);
nor U477 (N_477,In_1271,In_1206);
and U478 (N_478,In_2026,In_727);
or U479 (N_479,In_1217,In_1120);
and U480 (N_480,In_377,In_367);
xnor U481 (N_481,In_936,In_1869);
nand U482 (N_482,In_1592,In_2209);
nor U483 (N_483,In_996,In_1568);
nor U484 (N_484,In_1099,In_113);
or U485 (N_485,In_1155,In_2157);
or U486 (N_486,In_484,In_2019);
nand U487 (N_487,In_452,In_2084);
or U488 (N_488,In_1098,In_1768);
nor U489 (N_489,In_1660,In_2333);
and U490 (N_490,In_374,In_181);
and U491 (N_491,In_1722,In_245);
xnor U492 (N_492,In_2329,In_2307);
or U493 (N_493,In_1458,In_2255);
nand U494 (N_494,In_137,In_2048);
xor U495 (N_495,In_2186,In_1953);
xnor U496 (N_496,In_1135,In_411);
nand U497 (N_497,In_1263,In_2423);
xnor U498 (N_498,In_2452,In_1380);
nand U499 (N_499,In_810,In_455);
nand U500 (N_500,In_1695,In_1156);
xor U501 (N_501,In_1588,In_1138);
xnor U502 (N_502,In_501,In_2496);
or U503 (N_503,In_1444,In_275);
nor U504 (N_504,In_1942,In_1041);
and U505 (N_505,In_689,In_1272);
xor U506 (N_506,In_1465,In_705);
nand U507 (N_507,In_2321,In_1227);
and U508 (N_508,In_2343,In_1128);
nor U509 (N_509,In_26,In_1335);
xor U510 (N_510,In_858,In_2326);
or U511 (N_511,In_1486,In_840);
and U512 (N_512,In_655,In_834);
xor U513 (N_513,In_2044,In_2191);
xnor U514 (N_514,In_1434,In_96);
xor U515 (N_515,In_2099,In_2146);
nand U516 (N_516,In_2060,In_421);
and U517 (N_517,In_1775,In_1392);
xor U518 (N_518,In_1514,In_1046);
nor U519 (N_519,In_2027,In_1891);
or U520 (N_520,In_639,In_1184);
and U521 (N_521,In_450,In_1357);
or U522 (N_522,In_2269,In_537);
xor U523 (N_523,In_386,In_663);
nor U524 (N_524,In_446,In_1583);
or U525 (N_525,In_228,In_799);
or U526 (N_526,In_972,In_1167);
and U527 (N_527,In_1628,In_1137);
or U528 (N_528,In_882,In_934);
nand U529 (N_529,In_2088,In_2130);
nand U530 (N_530,In_1150,In_89);
xor U531 (N_531,In_38,In_1488);
nand U532 (N_532,In_1436,In_1967);
nor U533 (N_533,In_1899,In_923);
and U534 (N_534,In_1305,In_1073);
and U535 (N_535,In_71,In_2323);
or U536 (N_536,In_1973,In_251);
xor U537 (N_537,In_1843,In_1251);
xnor U538 (N_538,In_1896,In_1693);
xnor U539 (N_539,In_2073,In_1248);
or U540 (N_540,In_2124,In_672);
or U541 (N_541,In_61,In_776);
nand U542 (N_542,In_416,In_754);
and U543 (N_543,In_2217,In_373);
nand U544 (N_544,In_353,In_2337);
and U545 (N_545,In_956,In_559);
and U546 (N_546,In_1793,In_1751);
nand U547 (N_547,In_1332,In_146);
or U548 (N_548,In_683,In_2189);
nand U549 (N_549,In_2278,In_1769);
xor U550 (N_550,In_2410,In_478);
nand U551 (N_551,In_235,In_2300);
and U552 (N_552,In_1348,In_297);
nand U553 (N_553,In_2014,In_1820);
nor U554 (N_554,In_1863,In_1421);
nor U555 (N_555,In_1127,In_1980);
and U556 (N_556,In_383,In_1551);
xor U557 (N_557,In_2071,In_2150);
nor U558 (N_558,In_581,In_566);
and U559 (N_559,In_1412,In_629);
nor U560 (N_560,In_1331,In_2365);
or U561 (N_561,In_585,In_1541);
nor U562 (N_562,In_67,In_1417);
nand U563 (N_563,In_1613,In_2182);
or U564 (N_564,In_1478,In_1435);
or U565 (N_565,In_2059,In_1382);
nor U566 (N_566,In_2177,In_997);
nor U567 (N_567,In_1375,In_551);
or U568 (N_568,In_2195,In_653);
or U569 (N_569,In_1186,In_828);
xnor U570 (N_570,In_1270,In_354);
xnor U571 (N_571,In_45,In_1374);
xor U572 (N_572,In_444,In_2388);
or U573 (N_573,In_945,In_139);
xnor U574 (N_574,In_1654,In_474);
or U575 (N_575,In_2055,In_180);
xnor U576 (N_576,In_2045,In_1397);
and U577 (N_577,In_2020,In_1729);
xor U578 (N_578,In_309,In_1015);
nand U579 (N_579,In_1688,In_2174);
or U580 (N_580,In_903,In_1620);
and U581 (N_581,In_1279,In_1659);
nand U582 (N_582,In_1405,In_1152);
nand U583 (N_583,In_1745,In_1949);
nor U584 (N_584,In_1095,In_2199);
xnor U585 (N_585,In_1918,In_1656);
nor U586 (N_586,In_1108,In_462);
and U587 (N_587,In_2425,In_2069);
xor U588 (N_588,In_138,In_1093);
nor U589 (N_589,In_1306,In_1148);
xor U590 (N_590,In_2185,In_2256);
nand U591 (N_591,In_1391,In_1839);
nor U592 (N_592,In_1341,In_82);
nand U593 (N_593,In_1694,In_1499);
xnor U594 (N_594,In_1612,In_796);
and U595 (N_595,In_212,In_433);
or U596 (N_596,In_1065,In_481);
xnor U597 (N_597,In_1537,In_801);
nor U598 (N_598,In_564,In_2327);
xor U599 (N_599,In_1411,In_2284);
nor U600 (N_600,In_2077,In_1511);
xor U601 (N_601,In_1948,In_1608);
nor U602 (N_602,In_1145,In_2008);
nand U603 (N_603,In_1984,In_205);
and U604 (N_604,In_907,In_2040);
or U605 (N_605,In_177,In_2373);
and U606 (N_606,In_60,In_414);
nand U607 (N_607,In_2357,In_933);
or U608 (N_608,In_1064,In_2168);
or U609 (N_609,In_1183,In_1877);
nor U610 (N_610,In_1439,In_1734);
and U611 (N_611,In_265,In_2078);
xor U612 (N_612,In_491,In_1244);
nand U613 (N_613,In_306,In_898);
xnor U614 (N_614,In_1811,In_33);
nor U615 (N_615,In_434,In_2075);
nor U616 (N_616,In_1633,In_912);
xnor U617 (N_617,In_43,In_1981);
nor U618 (N_618,In_1366,In_1874);
xor U619 (N_619,In_1614,In_1490);
or U620 (N_620,In_1809,In_1649);
nor U621 (N_621,In_1610,In_2283);
xnor U622 (N_622,In_2062,In_1598);
and U623 (N_623,In_2181,In_1536);
xor U624 (N_624,In_646,In_1689);
nor U625 (N_625,In_98,In_1606);
or U626 (N_626,In_870,In_890);
nor U627 (N_627,In_249,In_622);
nand U628 (N_628,In_1353,In_2474);
or U629 (N_629,In_1243,In_2305);
or U630 (N_630,In_1640,In_2375);
or U631 (N_631,In_2400,In_475);
nand U632 (N_632,In_2050,In_97);
or U633 (N_633,In_2429,In_1048);
and U634 (N_634,In_2057,In_2165);
nor U635 (N_635,In_2340,In_2158);
xnor U636 (N_636,In_381,In_2279);
nand U637 (N_637,In_733,In_718);
nand U638 (N_638,In_614,In_1054);
nor U639 (N_639,In_258,In_829);
or U640 (N_640,In_134,In_2087);
or U641 (N_641,In_2390,In_2093);
xnor U642 (N_642,In_1972,In_917);
and U643 (N_643,In_1626,In_104);
nand U644 (N_644,In_2304,In_881);
and U645 (N_645,In_8,In_1977);
nor U646 (N_646,In_2302,In_320);
xor U647 (N_647,In_2056,In_941);
nand U648 (N_648,In_527,In_2235);
nand U649 (N_649,In_2301,In_2144);
nand U650 (N_650,In_2412,In_2065);
and U651 (N_651,In_1748,In_224);
nor U652 (N_652,In_511,In_465);
and U653 (N_653,In_479,In_984);
or U654 (N_654,In_1288,In_348);
or U655 (N_655,In_1841,In_1512);
or U656 (N_656,In_14,In_1268);
or U657 (N_657,In_804,In_1314);
and U658 (N_658,In_1684,In_745);
xor U659 (N_659,In_1846,In_975);
nand U660 (N_660,In_426,In_147);
and U661 (N_661,In_1280,In_1169);
nand U662 (N_662,In_6,In_1316);
nor U663 (N_663,In_2482,In_847);
and U664 (N_664,In_2451,In_1036);
or U665 (N_665,In_1721,In_334);
or U666 (N_666,In_387,In_591);
or U667 (N_667,In_442,In_1464);
and U668 (N_668,In_519,In_11);
nor U669 (N_669,In_1231,In_2085);
nor U670 (N_670,In_1825,In_850);
or U671 (N_671,In_2338,In_156);
nor U672 (N_672,In_630,In_2140);
xnor U673 (N_673,In_1201,In_1043);
nand U674 (N_674,In_1480,In_1164);
or U675 (N_675,In_1528,In_1181);
nor U676 (N_676,In_877,In_2172);
xnor U677 (N_677,In_1746,In_9);
and U678 (N_678,In_1057,In_1915);
or U679 (N_679,In_2171,In_1234);
nor U680 (N_680,In_124,In_553);
or U681 (N_681,In_2387,In_1242);
xor U682 (N_682,In_1025,In_1783);
or U683 (N_683,In_1664,In_364);
nor U684 (N_684,In_1908,In_405);
and U685 (N_685,In_887,In_895);
nor U686 (N_686,In_2253,In_1158);
nand U687 (N_687,In_1559,In_1163);
nor U688 (N_688,In_1218,In_1544);
xnor U689 (N_689,In_1047,In_1110);
nor U690 (N_690,In_1071,In_1303);
or U691 (N_691,In_1757,In_2456);
nor U692 (N_692,In_362,In_391);
nand U693 (N_693,In_1707,In_1580);
and U694 (N_694,In_2160,In_715);
xnor U695 (N_695,In_2023,In_1935);
nand U696 (N_696,In_148,In_1801);
nor U697 (N_697,In_750,In_627);
or U698 (N_698,In_1090,In_1636);
nor U699 (N_699,In_2466,In_154);
or U700 (N_700,In_1796,In_2345);
nor U701 (N_701,In_602,In_2257);
nand U702 (N_702,In_1955,In_2303);
nand U703 (N_703,In_963,In_1601);
nand U704 (N_704,In_1425,In_1394);
nor U705 (N_705,In_1957,In_806);
or U706 (N_706,In_1595,In_1873);
xor U707 (N_707,In_578,In_1635);
nor U708 (N_708,In_2270,In_651);
nor U709 (N_709,In_1883,In_973);
or U710 (N_710,In_1309,In_1014);
xnor U711 (N_711,In_900,In_1210);
nor U712 (N_712,In_2230,In_1954);
nor U713 (N_713,In_1576,In_521);
nand U714 (N_714,In_548,In_2109);
and U715 (N_715,In_779,In_2128);
nand U716 (N_716,In_232,In_142);
and U717 (N_717,In_786,In_1540);
nand U718 (N_718,In_637,In_644);
nand U719 (N_719,In_2035,In_1111);
or U720 (N_720,In_2458,In_577);
and U721 (N_721,In_149,In_2012);
and U722 (N_722,In_889,In_141);
nor U723 (N_723,In_1468,In_949);
and U724 (N_724,In_814,In_313);
xnor U725 (N_725,In_269,In_1764);
or U726 (N_726,In_955,In_294);
nor U727 (N_727,In_241,In_2127);
nor U728 (N_728,In_133,In_385);
nand U729 (N_729,In_1491,In_2194);
xor U730 (N_730,In_1469,In_1661);
nand U731 (N_731,In_719,In_1655);
and U732 (N_732,In_500,In_1067);
or U733 (N_733,In_1719,In_1130);
nand U734 (N_734,In_852,In_1897);
and U735 (N_735,In_1596,In_250);
xnor U736 (N_736,In_770,In_1424);
xor U737 (N_737,In_1276,In_1730);
and U738 (N_738,In_1408,In_1836);
and U739 (N_739,In_2263,In_2319);
and U740 (N_740,In_1179,In_1864);
xnor U741 (N_741,In_1711,In_299);
nor U742 (N_742,In_640,In_1724);
xnor U743 (N_743,In_1917,In_1865);
xor U744 (N_744,In_315,In_179);
nor U745 (N_745,In_2041,In_339);
xor U746 (N_746,In_1682,In_1162);
nor U747 (N_747,In_665,In_1430);
and U748 (N_748,In_117,In_2362);
and U749 (N_749,In_1088,In_1538);
xor U750 (N_750,In_2376,In_1153);
nand U751 (N_751,In_2215,In_764);
or U752 (N_752,In_660,In_1835);
nand U753 (N_753,In_832,In_1387);
xor U754 (N_754,In_2025,In_2227);
or U755 (N_755,In_164,In_1154);
nand U756 (N_756,In_256,In_1989);
or U757 (N_757,In_1741,In_56);
nand U758 (N_758,In_64,In_1747);
xor U759 (N_759,In_1621,In_2361);
or U760 (N_760,In_1737,In_1653);
and U761 (N_761,In_1266,In_310);
or U762 (N_762,In_2471,In_1627);
nor U763 (N_763,In_1032,In_1333);
or U764 (N_764,In_2208,In_558);
or U765 (N_765,In_724,In_1364);
nor U766 (N_766,In_560,In_267);
nor U767 (N_767,In_1325,In_1187);
xnor U768 (N_768,In_282,In_744);
nand U769 (N_769,In_1987,In_1945);
nor U770 (N_770,In_2081,In_2427);
nand U771 (N_771,In_2290,In_409);
or U772 (N_772,In_2032,In_1630);
and U773 (N_773,In_1479,In_1005);
xnor U774 (N_774,In_1894,In_1300);
or U775 (N_775,In_2092,In_2306);
xnor U776 (N_776,In_1763,In_855);
nand U777 (N_777,In_2460,In_784);
xnor U778 (N_778,In_1085,In_2139);
nand U779 (N_779,In_2036,In_2281);
xnor U780 (N_780,In_1166,In_335);
nand U781 (N_781,In_1504,In_556);
nand U782 (N_782,In_1554,In_69);
xor U783 (N_783,In_826,In_735);
xnor U784 (N_784,In_1319,In_1182);
nand U785 (N_785,In_2132,In_1498);
or U786 (N_786,In_1470,In_1860);
xnor U787 (N_787,In_2033,In_2344);
nor U788 (N_788,In_2398,In_190);
xnor U789 (N_789,In_1192,In_515);
nor U790 (N_790,In_1477,In_20);
xor U791 (N_791,In_823,In_2198);
and U792 (N_792,In_1593,In_2389);
or U793 (N_793,In_729,In_1866);
and U794 (N_794,In_1890,In_642);
nor U795 (N_795,In_1211,In_536);
or U796 (N_796,In_902,In_732);
and U797 (N_797,In_107,In_318);
nor U798 (N_798,In_1799,In_1508);
and U799 (N_799,In_595,In_1859);
or U800 (N_800,In_1410,In_1428);
or U801 (N_801,In_999,In_908);
nand U802 (N_802,In_78,In_1780);
xor U803 (N_803,In_982,In_1371);
nor U804 (N_804,In_1845,In_1976);
and U805 (N_805,In_17,In_2368);
nor U806 (N_806,In_2465,In_2353);
xnor U807 (N_807,In_845,In_322);
nor U808 (N_808,In_2431,In_2385);
or U809 (N_809,In_1299,In_1517);
xor U810 (N_810,In_1889,In_1455);
nand U811 (N_811,In_72,In_1349);
nand U812 (N_812,In_1617,In_332);
or U813 (N_813,In_24,In_1562);
xor U814 (N_814,In_2111,In_417);
or U815 (N_815,In_606,In_756);
and U816 (N_816,In_914,In_592);
or U817 (N_817,In_305,In_338);
nor U818 (N_818,In_604,In_126);
or U819 (N_819,In_1084,In_1516);
nor U820 (N_820,In_730,In_636);
xnor U821 (N_821,In_582,In_2);
nor U822 (N_822,In_1076,In_2483);
xnor U823 (N_823,In_2316,In_1326);
xnor U824 (N_824,In_1006,In_815);
and U825 (N_825,In_1509,In_1207);
nand U826 (N_826,In_2280,In_41);
nor U827 (N_827,In_196,In_1892);
xor U828 (N_828,In_159,In_301);
nor U829 (N_829,In_333,In_403);
xnor U830 (N_830,In_2433,In_1055);
and U831 (N_831,In_155,In_586);
and U832 (N_832,In_166,In_978);
nand U833 (N_833,In_676,In_210);
or U834 (N_834,In_234,In_1591);
xor U835 (N_835,In_2178,In_1979);
or U836 (N_836,In_1956,In_1925);
and U837 (N_837,In_2156,In_962);
xor U838 (N_838,In_52,In_649);
xor U839 (N_839,In_1476,In_1605);
xnor U840 (N_840,In_2289,In_2468);
and U841 (N_841,In_2404,In_1061);
and U842 (N_842,In_105,In_2184);
nor U843 (N_843,In_2058,In_472);
and U844 (N_844,In_1328,In_21);
or U845 (N_845,In_1772,In_761);
nand U846 (N_846,In_2315,In_1546);
or U847 (N_847,In_1302,In_2166);
or U848 (N_848,In_1031,In_1202);
and U849 (N_849,In_769,In_83);
nor U850 (N_850,In_229,In_2475);
nand U851 (N_851,In_2202,In_2418);
nor U852 (N_852,In_2358,In_2039);
and U853 (N_853,In_1224,In_319);
xor U854 (N_854,In_276,In_2347);
nor U855 (N_855,In_1564,In_2370);
and U856 (N_856,In_2359,In_762);
xnor U857 (N_857,In_2492,In_1779);
or U858 (N_858,In_2043,In_1313);
and U859 (N_859,In_1447,In_283);
and U860 (N_860,In_512,In_1691);
nor U861 (N_861,In_1739,In_2173);
nor U862 (N_862,In_347,In_119);
nand U863 (N_863,In_2082,In_961);
or U864 (N_864,In_2224,In_15);
or U865 (N_865,In_1350,In_573);
or U866 (N_866,In_991,In_589);
nand U867 (N_867,In_428,In_600);
nand U868 (N_868,In_1446,In_1577);
or U869 (N_869,In_1113,In_439);
and U870 (N_870,In_1713,In_1222);
or U871 (N_871,In_1840,In_1039);
nand U872 (N_872,In_1733,In_1539);
xnor U873 (N_873,In_311,In_1296);
or U874 (N_874,In_295,In_596);
nand U875 (N_875,In_2484,In_1385);
nor U876 (N_876,In_1862,In_2449);
and U877 (N_877,In_797,In_344);
nor U878 (N_878,In_2426,In_366);
or U879 (N_879,In_748,In_947);
and U880 (N_880,In_1909,In_2351);
xor U881 (N_881,In_2046,In_441);
and U882 (N_882,In_2213,In_2472);
or U883 (N_883,In_608,In_1484);
or U884 (N_884,In_80,In_875);
and U885 (N_885,In_669,In_1800);
and U886 (N_886,In_1632,In_1714);
or U887 (N_887,In_1888,In_92);
nor U888 (N_888,In_169,In_544);
nand U889 (N_889,In_106,In_969);
nor U890 (N_890,In_395,In_2196);
xnor U891 (N_891,In_1959,In_1466);
and U892 (N_892,In_994,In_2395);
nand U893 (N_893,In_2487,In_1472);
nor U894 (N_894,In_68,In_2486);
nor U895 (N_895,In_1285,In_1937);
nand U896 (N_896,In_300,In_1829);
and U897 (N_897,In_1631,In_1604);
or U898 (N_898,In_493,In_720);
nor U899 (N_899,In_1515,In_2274);
or U900 (N_900,In_308,In_1643);
or U901 (N_901,In_429,In_987);
or U902 (N_902,In_1901,In_534);
or U903 (N_903,In_2145,In_260);
nor U904 (N_904,In_1485,In_93);
xnor U905 (N_905,In_30,In_1042);
or U906 (N_906,In_2286,In_896);
nand U907 (N_907,In_1165,In_59);
and U908 (N_908,In_392,In_76);
xor U909 (N_909,In_2239,In_389);
or U910 (N_910,In_820,In_2317);
or U911 (N_911,In_787,In_2211);
nor U912 (N_912,In_702,In_1920);
nand U913 (N_913,In_788,In_867);
and U914 (N_914,In_2180,In_1997);
and U915 (N_915,In_967,In_1482);
or U916 (N_916,In_18,In_2009);
nand U917 (N_917,In_1483,In_1116);
xnor U918 (N_918,In_115,In_1086);
nand U919 (N_919,In_1229,In_1744);
xnor U920 (N_920,In_993,In_1552);
xnor U921 (N_921,In_830,In_1587);
xor U922 (N_922,In_862,In_783);
nor U923 (N_923,In_1260,In_1400);
or U924 (N_924,In_1089,In_1934);
or U925 (N_925,In_708,In_1988);
and U926 (N_926,In_1362,In_1603);
nand U927 (N_927,In_402,In_768);
nor U928 (N_928,In_2018,In_1740);
nor U929 (N_929,In_1176,In_1219);
nor U930 (N_930,In_925,In_325);
nand U931 (N_931,In_853,In_1599);
nand U932 (N_932,In_1704,In_222);
nand U933 (N_933,In_58,In_1356);
or U934 (N_934,In_2477,In_1927);
nor U935 (N_935,In_1118,In_2028);
nor U936 (N_936,In_974,In_183);
nand U937 (N_937,In_1531,In_1803);
nand U938 (N_938,In_2402,In_1209);
nor U939 (N_939,In_201,In_1226);
nand U940 (N_940,In_2187,In_1812);
xor U941 (N_941,In_1114,In_2311);
nand U942 (N_942,In_1700,In_971);
and U943 (N_943,In_495,In_775);
xnor U944 (N_944,In_948,In_1420);
nor U945 (N_945,In_1327,In_707);
and U946 (N_946,In_576,In_1104);
and U947 (N_947,In_371,In_2074);
nand U948 (N_948,In_538,In_487);
and U949 (N_949,In_257,In_1040);
nand U950 (N_950,In_1094,In_272);
nor U951 (N_951,In_5,In_699);
nor U952 (N_952,In_1012,In_2013);
nand U953 (N_953,In_1029,In_74);
or U954 (N_954,In_226,In_1028);
nand U955 (N_955,In_1597,In_2016);
xor U956 (N_956,In_624,In_281);
nor U957 (N_957,In_2318,In_1557);
nand U958 (N_958,In_1074,In_2377);
nand U959 (N_959,In_252,In_1461);
nand U960 (N_960,In_316,In_1708);
xnor U961 (N_961,In_2360,In_129);
and U962 (N_962,In_2374,In_1451);
xor U963 (N_963,In_1867,In_605);
xor U964 (N_964,In_1878,In_1124);
and U965 (N_965,In_1388,In_270);
nor U966 (N_966,In_436,In_268);
xor U967 (N_967,In_2246,In_2096);
nand U968 (N_968,In_1363,In_911);
nor U969 (N_969,In_178,In_203);
nand U970 (N_970,In_1473,In_2228);
nand U971 (N_971,In_567,In_2394);
nor U972 (N_972,In_1996,In_2220);
xnor U973 (N_973,In_2354,In_765);
or U974 (N_974,In_27,In_554);
nand U975 (N_975,In_1471,In_916);
nor U976 (N_976,In_657,In_1340);
or U977 (N_977,In_1474,In_940);
and U978 (N_978,In_1292,In_2137);
and U979 (N_979,In_274,In_562);
or U980 (N_980,In_648,In_264);
nand U981 (N_981,In_1298,In_1379);
and U982 (N_982,In_593,In_789);
or U983 (N_983,In_424,In_254);
or U984 (N_984,In_1505,In_1960);
nor U985 (N_985,In_929,In_1645);
nand U986 (N_986,In_2237,In_477);
and U987 (N_987,In_2104,In_1307);
and U988 (N_988,In_483,In_569);
and U989 (N_989,In_704,In_864);
or U990 (N_990,In_1521,In_1609);
xnor U991 (N_991,In_1932,In_497);
nor U992 (N_992,In_1761,In_2310);
nand U993 (N_993,In_116,In_1188);
nor U994 (N_994,In_1056,In_1611);
xor U995 (N_995,In_1567,In_1289);
and U996 (N_996,In_1018,In_540);
xor U997 (N_997,In_2276,In_2143);
nand U998 (N_998,In_1220,In_2478);
xor U999 (N_999,In_238,In_1518);
xor U1000 (N_1000,In_227,In_1494);
nand U1001 (N_1001,In_1838,In_726);
or U1002 (N_1002,In_695,In_66);
and U1003 (N_1003,In_2001,In_1795);
nand U1004 (N_1004,In_1017,In_2271);
or U1005 (N_1005,In_594,In_290);
or U1006 (N_1006,In_2499,In_140);
and U1007 (N_1007,In_2414,In_1794);
or U1008 (N_1008,In_189,In_1728);
or U1009 (N_1009,In_1530,In_2122);
or U1010 (N_1010,In_915,In_893);
or U1011 (N_1011,In_2221,In_449);
or U1012 (N_1012,In_239,In_886);
or U1013 (N_1013,In_188,In_145);
nand U1014 (N_1014,In_1294,In_685);
or U1015 (N_1015,In_2153,In_574);
or U1016 (N_1016,In_1277,In_2258);
or U1017 (N_1017,In_467,In_2005);
or U1018 (N_1018,In_271,In_1969);
or U1019 (N_1019,In_1172,In_1855);
nand U1020 (N_1020,In_1140,In_340);
xnor U1021 (N_1021,In_1079,In_2244);
or U1022 (N_1022,In_1431,In_1213);
nand U1023 (N_1023,In_587,In_598);
nand U1024 (N_1024,In_1767,In_844);
nor U1025 (N_1025,In_1429,In_876);
nand U1026 (N_1026,In_793,In_1926);
nor U1027 (N_1027,In_928,In_65);
and U1028 (N_1028,In_2210,In_384);
and U1029 (N_1029,In_261,In_1995);
xnor U1030 (N_1030,In_1254,In_1196);
xor U1031 (N_1031,In_2252,In_1022);
nor U1032 (N_1032,In_167,In_1273);
and U1033 (N_1033,In_528,In_909);
or U1034 (N_1034,In_1524,In_661);
and U1035 (N_1035,In_2328,In_747);
or U1036 (N_1036,In_725,In_211);
xor U1037 (N_1037,In_2372,In_1875);
or U1038 (N_1038,In_218,In_94);
or U1039 (N_1039,In_1648,In_781);
and U1040 (N_1040,In_220,In_151);
nor U1041 (N_1041,In_329,In_1678);
and U1042 (N_1042,In_2273,In_2022);
and U1043 (N_1043,In_31,In_1810);
nand U1044 (N_1044,In_2476,In_2148);
nor U1045 (N_1045,In_277,In_1513);
xor U1046 (N_1046,In_565,In_293);
nor U1047 (N_1047,In_1225,In_1930);
nand U1048 (N_1048,In_645,In_691);
nand U1049 (N_1049,In_1522,In_1802);
nand U1050 (N_1050,In_1861,In_579);
nand U1051 (N_1051,In_1257,In_42);
xor U1052 (N_1052,In_324,In_2292);
nor U1053 (N_1053,In_1125,In_127);
or U1054 (N_1054,In_2490,In_2367);
nor U1055 (N_1055,In_1674,In_1535);
nand U1056 (N_1056,In_382,In_286);
xnor U1057 (N_1057,In_1117,In_1007);
nand U1058 (N_1058,In_970,In_785);
nand U1059 (N_1059,In_231,In_2204);
or U1060 (N_1060,In_1781,In_1868);
or U1061 (N_1061,In_28,In_292);
and U1062 (N_1062,In_262,In_2288);
nand U1063 (N_1063,In_1902,In_1928);
xor U1064 (N_1064,In_631,In_2267);
nand U1065 (N_1065,In_1701,In_2101);
xnor U1066 (N_1066,In_879,In_1044);
nand U1067 (N_1067,In_1037,In_808);
nor U1068 (N_1068,In_1753,In_706);
nor U1069 (N_1069,In_2203,In_615);
or U1070 (N_1070,In_623,In_359);
xnor U1071 (N_1071,In_2147,In_312);
xor U1072 (N_1072,In_192,In_1002);
xnor U1073 (N_1073,In_157,In_2275);
nor U1074 (N_1074,In_1998,In_2031);
and U1075 (N_1075,In_398,In_1297);
and U1076 (N_1076,In_32,In_1390);
nand U1077 (N_1077,In_849,In_1035);
or U1078 (N_1078,In_193,In_36);
and U1079 (N_1079,In_1558,In_1230);
or U1080 (N_1080,In_1634,In_599);
nor U1081 (N_1081,In_1034,In_336);
xnor U1082 (N_1082,In_1999,In_2250);
nor U1083 (N_1083,In_1870,In_580);
xor U1084 (N_1084,In_2219,In_1529);
and U1085 (N_1085,In_1160,In_2197);
and U1086 (N_1086,In_2034,In_111);
nand U1087 (N_1087,In_2091,In_431);
and U1088 (N_1088,In_2455,In_1147);
nor U1089 (N_1089,In_2049,In_2406);
nor U1090 (N_1090,In_2095,In_1377);
xnor U1091 (N_1091,In_1383,In_1246);
xor U1092 (N_1092,In_357,In_1506);
xnor U1093 (N_1093,In_1718,In_838);
nand U1094 (N_1094,In_938,In_1198);
nand U1095 (N_1095,In_1876,In_1399);
and U1096 (N_1096,In_1159,In_1463);
or U1097 (N_1097,In_848,In_461);
xor U1098 (N_1098,In_2308,In_2162);
nand U1099 (N_1099,In_4,In_1947);
nand U1100 (N_1100,In_1912,In_351);
and U1101 (N_1101,In_1534,In_2320);
or U1102 (N_1102,In_2094,In_1749);
and U1103 (N_1103,In_44,In_1532);
and U1104 (N_1104,In_620,In_2432);
nand U1105 (N_1105,In_2205,In_1854);
nand U1106 (N_1106,In_1826,In_1139);
nor U1107 (N_1107,In_2293,In_2494);
nand U1108 (N_1108,In_717,In_2117);
and U1109 (N_1109,In_609,In_480);
nor U1110 (N_1110,In_1771,In_2159);
nand U1111 (N_1111,In_611,In_1600);
nor U1112 (N_1112,In_379,In_946);
nor U1113 (N_1113,In_2268,In_1663);
or U1114 (N_1114,In_1109,In_2225);
and U1115 (N_1115,In_990,In_1345);
and U1116 (N_1116,In_2277,In_200);
or U1117 (N_1117,In_825,In_1146);
nor U1118 (N_1118,In_1519,In_291);
and U1119 (N_1119,In_1318,In_2296);
or U1120 (N_1120,In_952,In_1001);
or U1121 (N_1121,In_530,In_1669);
and U1122 (N_1122,In_1275,In_2110);
and U1123 (N_1123,In_163,In_150);
nor U1124 (N_1124,In_1115,In_2105);
nand U1125 (N_1125,In_2467,In_686);
and U1126 (N_1126,In_303,In_1142);
nand U1127 (N_1127,In_568,In_1033);
or U1128 (N_1128,In_932,In_1221);
nand U1129 (N_1129,In_906,In_1290);
and U1130 (N_1130,In_369,In_2342);
and U1131 (N_1131,In_57,In_1295);
nand U1132 (N_1132,In_341,In_905);
xor U1133 (N_1133,In_1716,In_296);
nor U1134 (N_1134,In_1777,In_2430);
and U1135 (N_1135,In_2469,In_370);
nor U1136 (N_1136,In_2010,In_2222);
or U1137 (N_1137,In_2167,In_1355);
nand U1138 (N_1138,In_55,In_448);
nand U1139 (N_1139,In_53,In_0);
and U1140 (N_1140,In_641,In_2118);
or U1141 (N_1141,In_2355,In_1317);
nand U1142 (N_1142,In_135,In_1010);
and U1143 (N_1143,In_279,In_1819);
nor U1144 (N_1144,In_175,In_698);
or U1145 (N_1145,In_1072,In_1943);
nor U1146 (N_1146,In_1644,In_103);
nor U1147 (N_1147,In_1750,In_2366);
or U1148 (N_1148,In_1849,In_738);
or U1149 (N_1149,In_2463,In_2161);
or U1150 (N_1150,In_100,In_1107);
or U1151 (N_1151,In_1354,In_1754);
xor U1152 (N_1152,In_1129,In_736);
nand U1153 (N_1153,In_504,In_2100);
nor U1154 (N_1154,In_910,In_1881);
nand U1155 (N_1155,In_2183,In_1199);
nor U1156 (N_1156,In_1457,In_2218);
or U1157 (N_1157,In_1827,In_541);
xnor U1158 (N_1158,In_99,In_2133);
or U1159 (N_1159,In_1824,In_913);
or U1160 (N_1160,In_772,In_904);
nor U1161 (N_1161,In_1784,In_2070);
and U1162 (N_1162,In_1696,In_2011);
xor U1163 (N_1163,In_2450,In_2313);
or U1164 (N_1164,In_1259,In_194);
nand U1165 (N_1165,In_445,In_1416);
and U1166 (N_1166,In_1732,In_34);
nand U1167 (N_1167,In_451,In_1215);
nand U1168 (N_1168,In_570,In_1717);
xnor U1169 (N_1169,In_1283,In_1402);
or U1170 (N_1170,In_673,In_206);
nor U1171 (N_1171,In_509,In_510);
or U1172 (N_1172,In_1168,In_1441);
nand U1173 (N_1173,In_617,In_2138);
nand U1174 (N_1174,In_508,In_314);
nor U1175 (N_1175,In_543,In_490);
xnor U1176 (N_1176,In_1662,In_253);
or U1177 (N_1177,In_195,In_618);
xor U1178 (N_1178,In_1651,In_1706);
and U1179 (N_1179,In_25,In_161);
nor U1180 (N_1180,In_680,In_1699);
or U1181 (N_1181,In_782,In_552);
and U1182 (N_1182,In_263,In_1393);
or U1183 (N_1183,In_1008,In_755);
nor U1184 (N_1184,In_390,In_355);
nor U1185 (N_1185,In_2312,In_1344);
xor U1186 (N_1186,In_819,In_2391);
nor U1187 (N_1187,In_1489,In_1396);
or U1188 (N_1188,In_1023,In_1542);
and U1189 (N_1189,In_2126,In_700);
nor U1190 (N_1190,In_813,In_321);
nand U1191 (N_1191,In_1066,In_1049);
or U1192 (N_1192,In_1742,In_518);
or U1193 (N_1193,In_1121,In_677);
or U1194 (N_1194,In_1556,In_114);
nand U1195 (N_1195,In_376,In_652);
nor U1196 (N_1196,In_2480,In_2229);
nor U1197 (N_1197,In_1946,In_597);
nand U1198 (N_1198,In_920,In_549);
or U1199 (N_1199,In_2336,In_546);
and U1200 (N_1200,In_601,In_1453);
nor U1201 (N_1201,In_1555,In_812);
xnor U1202 (N_1202,In_1571,In_2435);
or U1203 (N_1203,In_1723,In_143);
or U1204 (N_1204,In_533,In_2381);
nand U1205 (N_1205,In_2488,In_2295);
nor U1206 (N_1206,In_1497,In_1808);
nor U1207 (N_1207,In_977,In_2066);
nor U1208 (N_1208,In_1625,In_2236);
nand U1209 (N_1209,In_2461,In_1249);
or U1210 (N_1210,In_1062,In_811);
nor U1211 (N_1211,In_1968,In_1329);
nor U1212 (N_1212,In_1258,In_628);
or U1213 (N_1213,In_924,In_168);
nand U1214 (N_1214,In_1910,In_1252);
nand U1215 (N_1215,In_1365,In_688);
nand U1216 (N_1216,In_1936,In_2380);
nand U1217 (N_1217,In_1369,In_901);
and U1218 (N_1218,In_1203,In_690);
or U1219 (N_1219,In_514,In_2002);
nand U1220 (N_1220,In_1647,In_118);
xor U1221 (N_1221,In_1053,In_2436);
and U1222 (N_1222,In_1284,In_2356);
nand U1223 (N_1223,In_856,In_2464);
nand U1224 (N_1224,In_1286,In_960);
and U1225 (N_1225,In_1792,In_1233);
xnor U1226 (N_1226,In_2247,In_939);
nand U1227 (N_1227,In_1550,In_742);
and U1228 (N_1228,In_2151,In_2007);
or U1229 (N_1229,In_160,In_1343);
nor U1230 (N_1230,In_2352,In_1360);
and U1231 (N_1231,In_1174,In_244);
nand U1232 (N_1232,In_1677,In_1422);
nor U1233 (N_1233,In_859,In_2231);
xnor U1234 (N_1234,In_1575,In_981);
nand U1235 (N_1235,In_1134,In_1185);
xor U1236 (N_1236,In_1921,In_70);
or U1237 (N_1237,In_1282,In_1330);
and U1238 (N_1238,In_378,In_1245);
or U1239 (N_1239,In_865,In_1269);
xor U1240 (N_1240,In_173,In_588);
nand U1241 (N_1241,In_13,In_361);
nor U1242 (N_1242,In_802,In_2396);
nor U1243 (N_1243,In_1293,In_507);
nand U1244 (N_1244,In_216,In_1590);
nand U1245 (N_1245,In_1502,In_2298);
and U1246 (N_1246,In_980,In_1602);
nor U1247 (N_1247,In_1642,In_1409);
nor U1248 (N_1248,In_1050,In_1070);
or U1249 (N_1249,In_2493,In_1652);
nor U1250 (N_1250,In_617,In_293);
or U1251 (N_1251,In_2176,In_276);
nand U1252 (N_1252,In_254,In_164);
or U1253 (N_1253,In_850,In_1363);
xnor U1254 (N_1254,In_16,In_288);
nand U1255 (N_1255,In_1415,In_586);
xor U1256 (N_1256,In_981,In_1428);
or U1257 (N_1257,In_526,In_34);
nand U1258 (N_1258,In_1372,In_868);
xor U1259 (N_1259,In_1414,In_757);
nor U1260 (N_1260,In_179,In_2369);
nand U1261 (N_1261,In_2383,In_1728);
or U1262 (N_1262,In_373,In_1867);
nand U1263 (N_1263,In_1406,In_1);
nand U1264 (N_1264,In_199,In_1907);
xor U1265 (N_1265,In_2135,In_512);
and U1266 (N_1266,In_1891,In_1422);
nand U1267 (N_1267,In_1682,In_1650);
and U1268 (N_1268,In_1849,In_468);
nand U1269 (N_1269,In_333,In_2402);
and U1270 (N_1270,In_2346,In_1111);
nand U1271 (N_1271,In_1266,In_309);
nor U1272 (N_1272,In_882,In_1548);
and U1273 (N_1273,In_752,In_2101);
xor U1274 (N_1274,In_1715,In_1572);
nor U1275 (N_1275,In_1157,In_1373);
and U1276 (N_1276,In_2457,In_211);
xor U1277 (N_1277,In_212,In_1511);
xor U1278 (N_1278,In_266,In_805);
xor U1279 (N_1279,In_463,In_2378);
nor U1280 (N_1280,In_2037,In_571);
nor U1281 (N_1281,In_1506,In_1833);
or U1282 (N_1282,In_112,In_491);
nor U1283 (N_1283,In_51,In_128);
or U1284 (N_1284,In_1000,In_770);
xnor U1285 (N_1285,In_2318,In_1767);
xnor U1286 (N_1286,In_2338,In_1561);
or U1287 (N_1287,In_1004,In_1850);
or U1288 (N_1288,In_142,In_2137);
and U1289 (N_1289,In_1627,In_773);
xor U1290 (N_1290,In_598,In_1667);
and U1291 (N_1291,In_8,In_372);
or U1292 (N_1292,In_558,In_2048);
xnor U1293 (N_1293,In_877,In_958);
and U1294 (N_1294,In_2378,In_1905);
nor U1295 (N_1295,In_542,In_2154);
nand U1296 (N_1296,In_1916,In_1645);
nand U1297 (N_1297,In_960,In_1445);
nand U1298 (N_1298,In_920,In_1473);
nor U1299 (N_1299,In_2260,In_2471);
nand U1300 (N_1300,In_1040,In_1892);
nor U1301 (N_1301,In_124,In_753);
and U1302 (N_1302,In_1209,In_581);
xnor U1303 (N_1303,In_338,In_782);
nand U1304 (N_1304,In_1992,In_1619);
xnor U1305 (N_1305,In_1844,In_1406);
xor U1306 (N_1306,In_1904,In_1829);
or U1307 (N_1307,In_1070,In_1560);
or U1308 (N_1308,In_2232,In_624);
or U1309 (N_1309,In_321,In_1513);
nor U1310 (N_1310,In_1348,In_1676);
xor U1311 (N_1311,In_1709,In_2145);
nor U1312 (N_1312,In_494,In_2189);
nand U1313 (N_1313,In_1951,In_1542);
and U1314 (N_1314,In_1764,In_609);
nor U1315 (N_1315,In_742,In_1431);
nor U1316 (N_1316,In_644,In_1808);
xnor U1317 (N_1317,In_240,In_2478);
nand U1318 (N_1318,In_183,In_601);
nor U1319 (N_1319,In_411,In_1189);
or U1320 (N_1320,In_867,In_1145);
nor U1321 (N_1321,In_1883,In_1824);
nor U1322 (N_1322,In_314,In_318);
xnor U1323 (N_1323,In_1409,In_443);
nor U1324 (N_1324,In_989,In_484);
and U1325 (N_1325,In_139,In_566);
xnor U1326 (N_1326,In_963,In_2232);
xor U1327 (N_1327,In_27,In_21);
xnor U1328 (N_1328,In_448,In_2018);
or U1329 (N_1329,In_1131,In_93);
nor U1330 (N_1330,In_1004,In_2014);
and U1331 (N_1331,In_2397,In_1034);
or U1332 (N_1332,In_336,In_452);
xnor U1333 (N_1333,In_2131,In_596);
nor U1334 (N_1334,In_584,In_1322);
and U1335 (N_1335,In_2280,In_854);
and U1336 (N_1336,In_1239,In_2192);
nand U1337 (N_1337,In_1527,In_1817);
nand U1338 (N_1338,In_2325,In_2157);
nand U1339 (N_1339,In_749,In_514);
nor U1340 (N_1340,In_1537,In_27);
and U1341 (N_1341,In_684,In_376);
and U1342 (N_1342,In_710,In_249);
or U1343 (N_1343,In_1124,In_236);
or U1344 (N_1344,In_1716,In_1577);
xor U1345 (N_1345,In_827,In_616);
nand U1346 (N_1346,In_2028,In_1359);
or U1347 (N_1347,In_1057,In_1121);
and U1348 (N_1348,In_328,In_2068);
nand U1349 (N_1349,In_1937,In_1777);
or U1350 (N_1350,In_1438,In_1034);
nor U1351 (N_1351,In_1930,In_766);
and U1352 (N_1352,In_1068,In_802);
and U1353 (N_1353,In_537,In_1424);
or U1354 (N_1354,In_113,In_2325);
nor U1355 (N_1355,In_363,In_265);
or U1356 (N_1356,In_417,In_2232);
nor U1357 (N_1357,In_1854,In_1037);
and U1358 (N_1358,In_2133,In_246);
nand U1359 (N_1359,In_973,In_1893);
or U1360 (N_1360,In_228,In_734);
nand U1361 (N_1361,In_1575,In_1237);
nor U1362 (N_1362,In_1131,In_763);
nand U1363 (N_1363,In_1195,In_2091);
xor U1364 (N_1364,In_1382,In_925);
nand U1365 (N_1365,In_2352,In_1070);
and U1366 (N_1366,In_2233,In_134);
nand U1367 (N_1367,In_1331,In_1375);
xnor U1368 (N_1368,In_2167,In_2168);
and U1369 (N_1369,In_1573,In_2455);
nor U1370 (N_1370,In_1502,In_908);
or U1371 (N_1371,In_1926,In_1939);
and U1372 (N_1372,In_1662,In_163);
nand U1373 (N_1373,In_655,In_1808);
and U1374 (N_1374,In_1084,In_1775);
nor U1375 (N_1375,In_1360,In_223);
nand U1376 (N_1376,In_52,In_1970);
nor U1377 (N_1377,In_446,In_2495);
nand U1378 (N_1378,In_2116,In_634);
or U1379 (N_1379,In_2139,In_2370);
and U1380 (N_1380,In_1126,In_1632);
and U1381 (N_1381,In_1048,In_1898);
nor U1382 (N_1382,In_852,In_1772);
xor U1383 (N_1383,In_90,In_1573);
and U1384 (N_1384,In_637,In_1813);
and U1385 (N_1385,In_1764,In_296);
nor U1386 (N_1386,In_1674,In_232);
and U1387 (N_1387,In_1622,In_2288);
nor U1388 (N_1388,In_1269,In_1081);
nor U1389 (N_1389,In_919,In_907);
or U1390 (N_1390,In_1549,In_14);
or U1391 (N_1391,In_998,In_1470);
nand U1392 (N_1392,In_463,In_831);
nand U1393 (N_1393,In_2288,In_46);
and U1394 (N_1394,In_417,In_1431);
xor U1395 (N_1395,In_1930,In_525);
and U1396 (N_1396,In_2175,In_970);
nand U1397 (N_1397,In_1287,In_643);
xnor U1398 (N_1398,In_2270,In_87);
nor U1399 (N_1399,In_747,In_1571);
xnor U1400 (N_1400,In_1182,In_2450);
and U1401 (N_1401,In_14,In_1813);
nor U1402 (N_1402,In_1858,In_1396);
or U1403 (N_1403,In_1393,In_420);
and U1404 (N_1404,In_1064,In_791);
or U1405 (N_1405,In_759,In_2095);
nand U1406 (N_1406,In_273,In_1209);
and U1407 (N_1407,In_1752,In_2326);
nand U1408 (N_1408,In_377,In_859);
nor U1409 (N_1409,In_823,In_2457);
or U1410 (N_1410,In_1760,In_389);
or U1411 (N_1411,In_160,In_2140);
and U1412 (N_1412,In_1351,In_1139);
or U1413 (N_1413,In_1662,In_468);
or U1414 (N_1414,In_1416,In_508);
and U1415 (N_1415,In_413,In_2008);
or U1416 (N_1416,In_2163,In_1376);
xnor U1417 (N_1417,In_1854,In_1182);
nand U1418 (N_1418,In_84,In_101);
nor U1419 (N_1419,In_1414,In_2041);
and U1420 (N_1420,In_2222,In_455);
xor U1421 (N_1421,In_2078,In_33);
or U1422 (N_1422,In_57,In_268);
or U1423 (N_1423,In_1349,In_1842);
and U1424 (N_1424,In_98,In_829);
nor U1425 (N_1425,In_1445,In_1060);
xnor U1426 (N_1426,In_1627,In_2429);
and U1427 (N_1427,In_1143,In_1814);
and U1428 (N_1428,In_1599,In_660);
xnor U1429 (N_1429,In_181,In_2104);
or U1430 (N_1430,In_619,In_940);
xor U1431 (N_1431,In_739,In_829);
or U1432 (N_1432,In_453,In_2040);
or U1433 (N_1433,In_1934,In_2484);
or U1434 (N_1434,In_877,In_801);
and U1435 (N_1435,In_196,In_235);
xor U1436 (N_1436,In_2389,In_2308);
nor U1437 (N_1437,In_1140,In_1566);
xnor U1438 (N_1438,In_131,In_233);
or U1439 (N_1439,In_572,In_1783);
nor U1440 (N_1440,In_803,In_1023);
or U1441 (N_1441,In_2152,In_2468);
nor U1442 (N_1442,In_157,In_298);
xnor U1443 (N_1443,In_144,In_2358);
or U1444 (N_1444,In_6,In_1041);
and U1445 (N_1445,In_981,In_1412);
and U1446 (N_1446,In_353,In_171);
or U1447 (N_1447,In_887,In_1780);
and U1448 (N_1448,In_1400,In_1645);
and U1449 (N_1449,In_217,In_1406);
and U1450 (N_1450,In_947,In_2416);
or U1451 (N_1451,In_365,In_1601);
xor U1452 (N_1452,In_1754,In_870);
nor U1453 (N_1453,In_377,In_2292);
nor U1454 (N_1454,In_870,In_2209);
nand U1455 (N_1455,In_1951,In_1394);
and U1456 (N_1456,In_1660,In_2471);
nor U1457 (N_1457,In_986,In_1931);
xor U1458 (N_1458,In_1412,In_1655);
and U1459 (N_1459,In_2385,In_834);
xor U1460 (N_1460,In_2081,In_685);
and U1461 (N_1461,In_969,In_2119);
nor U1462 (N_1462,In_1451,In_972);
xnor U1463 (N_1463,In_612,In_2142);
xor U1464 (N_1464,In_2499,In_989);
xnor U1465 (N_1465,In_1624,In_476);
nor U1466 (N_1466,In_2410,In_2019);
xnor U1467 (N_1467,In_960,In_2031);
xnor U1468 (N_1468,In_1215,In_498);
and U1469 (N_1469,In_1060,In_144);
nand U1470 (N_1470,In_465,In_743);
or U1471 (N_1471,In_384,In_1601);
nor U1472 (N_1472,In_1394,In_51);
nand U1473 (N_1473,In_1188,In_1507);
nand U1474 (N_1474,In_421,In_1948);
xnor U1475 (N_1475,In_442,In_912);
nor U1476 (N_1476,In_1773,In_1453);
xnor U1477 (N_1477,In_329,In_1554);
and U1478 (N_1478,In_2411,In_1396);
nor U1479 (N_1479,In_1372,In_1196);
or U1480 (N_1480,In_162,In_1505);
xor U1481 (N_1481,In_37,In_1016);
or U1482 (N_1482,In_834,In_2291);
nand U1483 (N_1483,In_1936,In_261);
xor U1484 (N_1484,In_1643,In_337);
xnor U1485 (N_1485,In_1069,In_1692);
nor U1486 (N_1486,In_1311,In_1235);
or U1487 (N_1487,In_2250,In_2157);
or U1488 (N_1488,In_290,In_1603);
and U1489 (N_1489,In_1190,In_1885);
nand U1490 (N_1490,In_744,In_1674);
xor U1491 (N_1491,In_875,In_2228);
and U1492 (N_1492,In_442,In_1526);
nand U1493 (N_1493,In_966,In_784);
nor U1494 (N_1494,In_379,In_1389);
xor U1495 (N_1495,In_2088,In_642);
or U1496 (N_1496,In_1354,In_1161);
nor U1497 (N_1497,In_125,In_2477);
nor U1498 (N_1498,In_2,In_2426);
and U1499 (N_1499,In_2343,In_914);
nand U1500 (N_1500,In_66,In_750);
and U1501 (N_1501,In_989,In_526);
and U1502 (N_1502,In_2282,In_207);
xor U1503 (N_1503,In_242,In_1229);
xor U1504 (N_1504,In_1069,In_503);
xor U1505 (N_1505,In_2351,In_198);
nor U1506 (N_1506,In_1611,In_1229);
or U1507 (N_1507,In_1361,In_2212);
or U1508 (N_1508,In_1694,In_1835);
nor U1509 (N_1509,In_1561,In_2406);
or U1510 (N_1510,In_906,In_837);
nand U1511 (N_1511,In_1030,In_1090);
nor U1512 (N_1512,In_378,In_628);
xnor U1513 (N_1513,In_1995,In_1033);
and U1514 (N_1514,In_121,In_897);
nor U1515 (N_1515,In_19,In_489);
and U1516 (N_1516,In_1841,In_1224);
nand U1517 (N_1517,In_1353,In_1158);
and U1518 (N_1518,In_1929,In_5);
xor U1519 (N_1519,In_2458,In_1921);
or U1520 (N_1520,In_211,In_1710);
nor U1521 (N_1521,In_1587,In_1872);
or U1522 (N_1522,In_2039,In_521);
nand U1523 (N_1523,In_503,In_513);
xnor U1524 (N_1524,In_422,In_1761);
xor U1525 (N_1525,In_321,In_1774);
nor U1526 (N_1526,In_1663,In_404);
nor U1527 (N_1527,In_2148,In_545);
nor U1528 (N_1528,In_398,In_133);
nand U1529 (N_1529,In_948,In_424);
or U1530 (N_1530,In_2170,In_1907);
or U1531 (N_1531,In_2476,In_86);
or U1532 (N_1532,In_526,In_758);
nand U1533 (N_1533,In_1319,In_2198);
or U1534 (N_1534,In_427,In_1766);
and U1535 (N_1535,In_2453,In_640);
and U1536 (N_1536,In_2365,In_819);
or U1537 (N_1537,In_248,In_2252);
nand U1538 (N_1538,In_1191,In_1259);
or U1539 (N_1539,In_539,In_1399);
and U1540 (N_1540,In_2392,In_752);
and U1541 (N_1541,In_1510,In_1211);
nor U1542 (N_1542,In_1403,In_1099);
or U1543 (N_1543,In_1186,In_1458);
or U1544 (N_1544,In_688,In_1568);
or U1545 (N_1545,In_554,In_2123);
and U1546 (N_1546,In_2187,In_1654);
and U1547 (N_1547,In_367,In_1157);
xnor U1548 (N_1548,In_928,In_2117);
nand U1549 (N_1549,In_1044,In_1924);
and U1550 (N_1550,In_1864,In_1424);
and U1551 (N_1551,In_2153,In_1068);
xnor U1552 (N_1552,In_1668,In_1783);
nand U1553 (N_1553,In_65,In_317);
xnor U1554 (N_1554,In_1959,In_896);
nor U1555 (N_1555,In_1881,In_1577);
nand U1556 (N_1556,In_859,In_2482);
nand U1557 (N_1557,In_888,In_2342);
or U1558 (N_1558,In_1424,In_2428);
and U1559 (N_1559,In_1752,In_2319);
or U1560 (N_1560,In_993,In_1491);
xor U1561 (N_1561,In_2314,In_1016);
xor U1562 (N_1562,In_625,In_1518);
xor U1563 (N_1563,In_1146,In_1918);
xor U1564 (N_1564,In_1405,In_406);
and U1565 (N_1565,In_2057,In_225);
nand U1566 (N_1566,In_578,In_75);
nor U1567 (N_1567,In_2073,In_770);
or U1568 (N_1568,In_454,In_1768);
or U1569 (N_1569,In_2186,In_368);
or U1570 (N_1570,In_1558,In_1609);
and U1571 (N_1571,In_1509,In_1);
xor U1572 (N_1572,In_130,In_1570);
nand U1573 (N_1573,In_2377,In_1292);
or U1574 (N_1574,In_1918,In_410);
nand U1575 (N_1575,In_2022,In_981);
xor U1576 (N_1576,In_1266,In_1038);
nor U1577 (N_1577,In_1373,In_2472);
xnor U1578 (N_1578,In_1558,In_168);
and U1579 (N_1579,In_170,In_812);
nand U1580 (N_1580,In_1711,In_60);
xor U1581 (N_1581,In_659,In_2364);
and U1582 (N_1582,In_2232,In_2446);
xnor U1583 (N_1583,In_677,In_2379);
nand U1584 (N_1584,In_1421,In_1933);
xor U1585 (N_1585,In_2418,In_199);
and U1586 (N_1586,In_1117,In_2046);
nand U1587 (N_1587,In_630,In_1582);
nand U1588 (N_1588,In_917,In_1483);
or U1589 (N_1589,In_484,In_2180);
or U1590 (N_1590,In_1677,In_669);
or U1591 (N_1591,In_38,In_1135);
xnor U1592 (N_1592,In_735,In_1200);
or U1593 (N_1593,In_2409,In_1100);
nand U1594 (N_1594,In_1299,In_2296);
xor U1595 (N_1595,In_1922,In_1967);
xor U1596 (N_1596,In_1662,In_1890);
and U1597 (N_1597,In_1043,In_1141);
nor U1598 (N_1598,In_2475,In_2093);
or U1599 (N_1599,In_938,In_1982);
or U1600 (N_1600,In_382,In_2000);
nand U1601 (N_1601,In_1685,In_2390);
nand U1602 (N_1602,In_1087,In_2419);
nand U1603 (N_1603,In_382,In_701);
nand U1604 (N_1604,In_1272,In_1821);
nor U1605 (N_1605,In_1726,In_2063);
nor U1606 (N_1606,In_781,In_554);
nor U1607 (N_1607,In_1275,In_407);
nand U1608 (N_1608,In_530,In_155);
nand U1609 (N_1609,In_465,In_329);
nand U1610 (N_1610,In_1800,In_195);
nor U1611 (N_1611,In_1644,In_2283);
nor U1612 (N_1612,In_2444,In_1651);
or U1613 (N_1613,In_1213,In_675);
xor U1614 (N_1614,In_2268,In_19);
and U1615 (N_1615,In_1632,In_1568);
xor U1616 (N_1616,In_1067,In_1786);
nor U1617 (N_1617,In_2210,In_2137);
nor U1618 (N_1618,In_670,In_799);
nand U1619 (N_1619,In_1749,In_380);
and U1620 (N_1620,In_1510,In_1514);
and U1621 (N_1621,In_1972,In_1265);
xor U1622 (N_1622,In_1495,In_1363);
nor U1623 (N_1623,In_1688,In_4);
and U1624 (N_1624,In_2451,In_2414);
nor U1625 (N_1625,In_1802,In_1730);
xnor U1626 (N_1626,In_1986,In_1548);
nor U1627 (N_1627,In_1378,In_708);
nand U1628 (N_1628,In_995,In_126);
nand U1629 (N_1629,In_2137,In_814);
or U1630 (N_1630,In_2035,In_108);
nand U1631 (N_1631,In_1088,In_566);
nand U1632 (N_1632,In_827,In_1595);
and U1633 (N_1633,In_861,In_1946);
and U1634 (N_1634,In_1574,In_1512);
xnor U1635 (N_1635,In_1067,In_1470);
xnor U1636 (N_1636,In_1189,In_327);
nor U1637 (N_1637,In_921,In_26);
nor U1638 (N_1638,In_1077,In_983);
xnor U1639 (N_1639,In_1536,In_1551);
nand U1640 (N_1640,In_1873,In_584);
and U1641 (N_1641,In_2417,In_1253);
nand U1642 (N_1642,In_332,In_552);
nand U1643 (N_1643,In_1072,In_1355);
xnor U1644 (N_1644,In_1413,In_1470);
nor U1645 (N_1645,In_1612,In_2312);
nor U1646 (N_1646,In_1598,In_158);
nand U1647 (N_1647,In_540,In_358);
nor U1648 (N_1648,In_1617,In_65);
xnor U1649 (N_1649,In_655,In_1274);
nand U1650 (N_1650,In_2471,In_709);
nor U1651 (N_1651,In_1933,In_588);
nand U1652 (N_1652,In_659,In_377);
or U1653 (N_1653,In_2277,In_1653);
xor U1654 (N_1654,In_1731,In_314);
or U1655 (N_1655,In_639,In_1503);
nand U1656 (N_1656,In_1198,In_1778);
or U1657 (N_1657,In_431,In_2344);
nand U1658 (N_1658,In_1778,In_1544);
nor U1659 (N_1659,In_1603,In_1875);
or U1660 (N_1660,In_1122,In_374);
and U1661 (N_1661,In_170,In_2119);
nand U1662 (N_1662,In_1414,In_2209);
or U1663 (N_1663,In_1806,In_1390);
or U1664 (N_1664,In_2178,In_714);
xor U1665 (N_1665,In_1000,In_426);
nor U1666 (N_1666,In_1790,In_6);
xnor U1667 (N_1667,In_1570,In_1730);
nand U1668 (N_1668,In_2330,In_2267);
nor U1669 (N_1669,In_99,In_292);
nor U1670 (N_1670,In_749,In_1976);
and U1671 (N_1671,In_2055,In_2066);
nor U1672 (N_1672,In_2387,In_747);
nor U1673 (N_1673,In_1320,In_1350);
and U1674 (N_1674,In_295,In_422);
nand U1675 (N_1675,In_652,In_774);
nor U1676 (N_1676,In_2067,In_2440);
nor U1677 (N_1677,In_1027,In_2254);
and U1678 (N_1678,In_851,In_175);
nor U1679 (N_1679,In_1105,In_2127);
nor U1680 (N_1680,In_1725,In_1066);
nor U1681 (N_1681,In_1362,In_1221);
nor U1682 (N_1682,In_107,In_72);
nand U1683 (N_1683,In_1511,In_1353);
nand U1684 (N_1684,In_1541,In_922);
xor U1685 (N_1685,In_1772,In_1071);
nand U1686 (N_1686,In_695,In_2428);
and U1687 (N_1687,In_1912,In_1886);
and U1688 (N_1688,In_363,In_463);
nand U1689 (N_1689,In_74,In_1325);
nor U1690 (N_1690,In_108,In_1610);
nor U1691 (N_1691,In_1843,In_2423);
nor U1692 (N_1692,In_1558,In_1930);
and U1693 (N_1693,In_1518,In_952);
and U1694 (N_1694,In_17,In_1549);
xor U1695 (N_1695,In_348,In_1113);
or U1696 (N_1696,In_1852,In_2057);
and U1697 (N_1697,In_368,In_1455);
xnor U1698 (N_1698,In_1780,In_68);
or U1699 (N_1699,In_880,In_2404);
nor U1700 (N_1700,In_1655,In_517);
xnor U1701 (N_1701,In_2496,In_2298);
or U1702 (N_1702,In_556,In_1264);
nand U1703 (N_1703,In_2118,In_257);
nand U1704 (N_1704,In_622,In_1051);
and U1705 (N_1705,In_2075,In_945);
nand U1706 (N_1706,In_1568,In_1859);
xnor U1707 (N_1707,In_2454,In_2233);
xnor U1708 (N_1708,In_755,In_1222);
nor U1709 (N_1709,In_592,In_1502);
nand U1710 (N_1710,In_2434,In_210);
or U1711 (N_1711,In_73,In_2443);
and U1712 (N_1712,In_520,In_875);
nor U1713 (N_1713,In_1499,In_819);
or U1714 (N_1714,In_2187,In_821);
xnor U1715 (N_1715,In_1343,In_1106);
and U1716 (N_1716,In_1409,In_1297);
nand U1717 (N_1717,In_1659,In_2121);
xor U1718 (N_1718,In_1274,In_1669);
nand U1719 (N_1719,In_1288,In_2329);
or U1720 (N_1720,In_1543,In_982);
nor U1721 (N_1721,In_1871,In_2229);
nand U1722 (N_1722,In_1561,In_2357);
xor U1723 (N_1723,In_1642,In_1654);
nor U1724 (N_1724,In_2479,In_1614);
xor U1725 (N_1725,In_1881,In_1451);
and U1726 (N_1726,In_2179,In_27);
xnor U1727 (N_1727,In_666,In_1612);
and U1728 (N_1728,In_807,In_1351);
and U1729 (N_1729,In_1768,In_1895);
xnor U1730 (N_1730,In_650,In_1601);
and U1731 (N_1731,In_1784,In_700);
nor U1732 (N_1732,In_165,In_677);
xor U1733 (N_1733,In_1747,In_1870);
or U1734 (N_1734,In_113,In_2348);
nand U1735 (N_1735,In_1521,In_1454);
or U1736 (N_1736,In_849,In_137);
nand U1737 (N_1737,In_1664,In_2055);
and U1738 (N_1738,In_892,In_1475);
and U1739 (N_1739,In_343,In_2450);
xnor U1740 (N_1740,In_265,In_101);
or U1741 (N_1741,In_1769,In_228);
and U1742 (N_1742,In_1978,In_1338);
nor U1743 (N_1743,In_329,In_470);
nor U1744 (N_1744,In_1336,In_1199);
xnor U1745 (N_1745,In_1876,In_561);
nand U1746 (N_1746,In_1039,In_923);
nor U1747 (N_1747,In_2498,In_2425);
nand U1748 (N_1748,In_919,In_1440);
or U1749 (N_1749,In_2120,In_1634);
nand U1750 (N_1750,In_1818,In_461);
xnor U1751 (N_1751,In_684,In_1974);
nand U1752 (N_1752,In_1017,In_1150);
xor U1753 (N_1753,In_1499,In_1869);
and U1754 (N_1754,In_1810,In_1434);
or U1755 (N_1755,In_1677,In_1663);
and U1756 (N_1756,In_1706,In_599);
nand U1757 (N_1757,In_475,In_2475);
nor U1758 (N_1758,In_1073,In_2266);
nor U1759 (N_1759,In_1088,In_633);
and U1760 (N_1760,In_1010,In_2462);
xor U1761 (N_1761,In_1361,In_107);
and U1762 (N_1762,In_660,In_2298);
nand U1763 (N_1763,In_1984,In_1086);
nand U1764 (N_1764,In_315,In_1980);
nor U1765 (N_1765,In_2412,In_1284);
or U1766 (N_1766,In_1012,In_991);
xnor U1767 (N_1767,In_46,In_301);
or U1768 (N_1768,In_1536,In_269);
xnor U1769 (N_1769,In_2459,In_710);
and U1770 (N_1770,In_1905,In_2025);
xnor U1771 (N_1771,In_96,In_1465);
and U1772 (N_1772,In_539,In_407);
nor U1773 (N_1773,In_1939,In_938);
and U1774 (N_1774,In_2235,In_1281);
nand U1775 (N_1775,In_958,In_2141);
and U1776 (N_1776,In_2248,In_2433);
and U1777 (N_1777,In_1984,In_2447);
and U1778 (N_1778,In_208,In_2206);
xor U1779 (N_1779,In_347,In_433);
nand U1780 (N_1780,In_1525,In_766);
or U1781 (N_1781,In_158,In_1299);
or U1782 (N_1782,In_678,In_1952);
nor U1783 (N_1783,In_739,In_897);
or U1784 (N_1784,In_2237,In_1674);
or U1785 (N_1785,In_441,In_1020);
nor U1786 (N_1786,In_1154,In_2155);
nor U1787 (N_1787,In_1363,In_2458);
nor U1788 (N_1788,In_1928,In_782);
nor U1789 (N_1789,In_123,In_1860);
xor U1790 (N_1790,In_2438,In_379);
xor U1791 (N_1791,In_1390,In_1509);
nor U1792 (N_1792,In_2344,In_890);
xnor U1793 (N_1793,In_937,In_1017);
nor U1794 (N_1794,In_2359,In_584);
nor U1795 (N_1795,In_1251,In_988);
nor U1796 (N_1796,In_1856,In_197);
nor U1797 (N_1797,In_1868,In_1992);
xor U1798 (N_1798,In_1507,In_1139);
xnor U1799 (N_1799,In_1936,In_979);
or U1800 (N_1800,In_953,In_1950);
nand U1801 (N_1801,In_2056,In_1343);
or U1802 (N_1802,In_1098,In_1785);
or U1803 (N_1803,In_924,In_299);
xor U1804 (N_1804,In_132,In_2403);
xor U1805 (N_1805,In_812,In_2200);
xnor U1806 (N_1806,In_867,In_431);
or U1807 (N_1807,In_465,In_1131);
and U1808 (N_1808,In_998,In_2483);
xor U1809 (N_1809,In_790,In_1439);
nor U1810 (N_1810,In_1837,In_465);
xnor U1811 (N_1811,In_1868,In_863);
or U1812 (N_1812,In_642,In_1566);
xor U1813 (N_1813,In_581,In_2049);
and U1814 (N_1814,In_937,In_477);
nor U1815 (N_1815,In_2399,In_1320);
or U1816 (N_1816,In_2325,In_1750);
nand U1817 (N_1817,In_1087,In_2398);
xnor U1818 (N_1818,In_2235,In_1963);
and U1819 (N_1819,In_1030,In_2045);
xnor U1820 (N_1820,In_1298,In_51);
xor U1821 (N_1821,In_833,In_949);
and U1822 (N_1822,In_2025,In_2445);
and U1823 (N_1823,In_428,In_663);
nand U1824 (N_1824,In_505,In_1086);
xor U1825 (N_1825,In_2408,In_225);
nand U1826 (N_1826,In_925,In_190);
nor U1827 (N_1827,In_1232,In_185);
nand U1828 (N_1828,In_1244,In_1605);
nor U1829 (N_1829,In_393,In_1986);
or U1830 (N_1830,In_1719,In_892);
and U1831 (N_1831,In_728,In_818);
nand U1832 (N_1832,In_2199,In_936);
xnor U1833 (N_1833,In_80,In_40);
and U1834 (N_1834,In_367,In_410);
nand U1835 (N_1835,In_1055,In_814);
nand U1836 (N_1836,In_609,In_1790);
nor U1837 (N_1837,In_2493,In_18);
nor U1838 (N_1838,In_906,In_2166);
nor U1839 (N_1839,In_1557,In_573);
nand U1840 (N_1840,In_501,In_386);
nor U1841 (N_1841,In_667,In_1721);
xor U1842 (N_1842,In_862,In_2025);
nand U1843 (N_1843,In_1591,In_2155);
nor U1844 (N_1844,In_788,In_329);
or U1845 (N_1845,In_2272,In_1993);
nor U1846 (N_1846,In_878,In_212);
nand U1847 (N_1847,In_1120,In_319);
or U1848 (N_1848,In_2007,In_1354);
nand U1849 (N_1849,In_1621,In_1897);
nand U1850 (N_1850,In_609,In_85);
nand U1851 (N_1851,In_172,In_2268);
nand U1852 (N_1852,In_1513,In_1381);
nor U1853 (N_1853,In_6,In_217);
and U1854 (N_1854,In_1970,In_819);
xor U1855 (N_1855,In_2398,In_704);
nor U1856 (N_1856,In_864,In_1877);
xnor U1857 (N_1857,In_94,In_2337);
xnor U1858 (N_1858,In_2142,In_1019);
xor U1859 (N_1859,In_1069,In_1673);
nor U1860 (N_1860,In_1843,In_901);
nand U1861 (N_1861,In_637,In_2107);
nand U1862 (N_1862,In_1233,In_2016);
nand U1863 (N_1863,In_1420,In_781);
or U1864 (N_1864,In_1372,In_881);
xnor U1865 (N_1865,In_1393,In_1442);
and U1866 (N_1866,In_726,In_1950);
or U1867 (N_1867,In_1845,In_1871);
nand U1868 (N_1868,In_484,In_1357);
nor U1869 (N_1869,In_785,In_1749);
and U1870 (N_1870,In_788,In_643);
nand U1871 (N_1871,In_2133,In_1268);
nand U1872 (N_1872,In_2494,In_849);
or U1873 (N_1873,In_2189,In_2445);
xor U1874 (N_1874,In_1346,In_902);
and U1875 (N_1875,In_1611,In_2041);
and U1876 (N_1876,In_2490,In_2204);
or U1877 (N_1877,In_869,In_822);
or U1878 (N_1878,In_1776,In_41);
nand U1879 (N_1879,In_41,In_2157);
xnor U1880 (N_1880,In_2107,In_2325);
nand U1881 (N_1881,In_721,In_1740);
xor U1882 (N_1882,In_2380,In_1950);
xor U1883 (N_1883,In_79,In_1289);
and U1884 (N_1884,In_12,In_1939);
nor U1885 (N_1885,In_656,In_1249);
xnor U1886 (N_1886,In_1024,In_450);
nor U1887 (N_1887,In_2311,In_2289);
and U1888 (N_1888,In_505,In_2323);
and U1889 (N_1889,In_1952,In_1867);
and U1890 (N_1890,In_802,In_2091);
xor U1891 (N_1891,In_304,In_1050);
xnor U1892 (N_1892,In_264,In_2121);
nand U1893 (N_1893,In_1961,In_2177);
nor U1894 (N_1894,In_1171,In_803);
xor U1895 (N_1895,In_277,In_1748);
and U1896 (N_1896,In_1572,In_912);
xor U1897 (N_1897,In_1157,In_1678);
and U1898 (N_1898,In_1651,In_223);
xnor U1899 (N_1899,In_1065,In_868);
or U1900 (N_1900,In_1916,In_1992);
xor U1901 (N_1901,In_252,In_2480);
nor U1902 (N_1902,In_1308,In_1432);
nand U1903 (N_1903,In_1136,In_322);
nor U1904 (N_1904,In_1013,In_432);
or U1905 (N_1905,In_2303,In_2184);
or U1906 (N_1906,In_818,In_607);
nor U1907 (N_1907,In_85,In_421);
xor U1908 (N_1908,In_304,In_2001);
nand U1909 (N_1909,In_567,In_709);
nand U1910 (N_1910,In_2410,In_45);
nand U1911 (N_1911,In_57,In_1323);
or U1912 (N_1912,In_1534,In_2026);
or U1913 (N_1913,In_656,In_2344);
and U1914 (N_1914,In_1954,In_2231);
nor U1915 (N_1915,In_1505,In_1181);
and U1916 (N_1916,In_2060,In_2136);
or U1917 (N_1917,In_1564,In_2006);
xor U1918 (N_1918,In_1230,In_995);
and U1919 (N_1919,In_503,In_1951);
and U1920 (N_1920,In_1192,In_2441);
nor U1921 (N_1921,In_1431,In_1314);
nand U1922 (N_1922,In_1940,In_1891);
and U1923 (N_1923,In_916,In_1335);
or U1924 (N_1924,In_1935,In_1008);
nor U1925 (N_1925,In_1172,In_1144);
and U1926 (N_1926,In_1519,In_1974);
and U1927 (N_1927,In_1604,In_2048);
xor U1928 (N_1928,In_518,In_675);
nor U1929 (N_1929,In_56,In_1038);
and U1930 (N_1930,In_245,In_221);
nand U1931 (N_1931,In_181,In_1769);
nand U1932 (N_1932,In_90,In_1399);
xor U1933 (N_1933,In_513,In_2325);
and U1934 (N_1934,In_603,In_1571);
nor U1935 (N_1935,In_1706,In_192);
xor U1936 (N_1936,In_912,In_1899);
nand U1937 (N_1937,In_340,In_531);
xor U1938 (N_1938,In_285,In_274);
nor U1939 (N_1939,In_180,In_2330);
nor U1940 (N_1940,In_708,In_743);
xor U1941 (N_1941,In_1194,In_1435);
nor U1942 (N_1942,In_1165,In_1545);
nand U1943 (N_1943,In_2378,In_1659);
or U1944 (N_1944,In_1071,In_1989);
and U1945 (N_1945,In_287,In_2143);
nor U1946 (N_1946,In_322,In_860);
nand U1947 (N_1947,In_1348,In_768);
or U1948 (N_1948,In_2403,In_2341);
nor U1949 (N_1949,In_611,In_420);
nor U1950 (N_1950,In_1800,In_809);
nand U1951 (N_1951,In_1263,In_679);
and U1952 (N_1952,In_1742,In_1447);
or U1953 (N_1953,In_36,In_1463);
xor U1954 (N_1954,In_194,In_2304);
and U1955 (N_1955,In_1435,In_2060);
nor U1956 (N_1956,In_1038,In_2330);
and U1957 (N_1957,In_971,In_1481);
and U1958 (N_1958,In_683,In_1850);
nor U1959 (N_1959,In_99,In_1833);
xor U1960 (N_1960,In_1294,In_389);
xor U1961 (N_1961,In_260,In_506);
nand U1962 (N_1962,In_1321,In_2401);
and U1963 (N_1963,In_1091,In_2480);
nand U1964 (N_1964,In_2275,In_2301);
nand U1965 (N_1965,In_1435,In_1674);
or U1966 (N_1966,In_511,In_1548);
and U1967 (N_1967,In_453,In_1387);
nor U1968 (N_1968,In_232,In_476);
and U1969 (N_1969,In_839,In_2461);
xor U1970 (N_1970,In_45,In_130);
xnor U1971 (N_1971,In_2349,In_570);
or U1972 (N_1972,In_357,In_906);
xnor U1973 (N_1973,In_1272,In_2021);
or U1974 (N_1974,In_982,In_1468);
and U1975 (N_1975,In_1676,In_1546);
xnor U1976 (N_1976,In_2092,In_965);
nor U1977 (N_1977,In_2427,In_1395);
nor U1978 (N_1978,In_2174,In_1172);
or U1979 (N_1979,In_2320,In_2331);
or U1980 (N_1980,In_2029,In_1816);
nand U1981 (N_1981,In_804,In_1386);
or U1982 (N_1982,In_981,In_857);
or U1983 (N_1983,In_716,In_2066);
xnor U1984 (N_1984,In_1604,In_79);
and U1985 (N_1985,In_1415,In_855);
nand U1986 (N_1986,In_1954,In_1386);
xnor U1987 (N_1987,In_2157,In_1305);
and U1988 (N_1988,In_249,In_433);
and U1989 (N_1989,In_430,In_480);
and U1990 (N_1990,In_172,In_878);
and U1991 (N_1991,In_1887,In_2300);
or U1992 (N_1992,In_1969,In_1475);
or U1993 (N_1993,In_278,In_1643);
xnor U1994 (N_1994,In_1407,In_997);
and U1995 (N_1995,In_1985,In_2069);
or U1996 (N_1996,In_2111,In_2106);
nand U1997 (N_1997,In_744,In_2419);
or U1998 (N_1998,In_2118,In_2119);
xor U1999 (N_1999,In_84,In_1703);
nor U2000 (N_2000,In_619,In_1380);
nand U2001 (N_2001,In_2012,In_1798);
or U2002 (N_2002,In_339,In_500);
nand U2003 (N_2003,In_557,In_1658);
and U2004 (N_2004,In_171,In_172);
xnor U2005 (N_2005,In_1416,In_1967);
xor U2006 (N_2006,In_1240,In_423);
nand U2007 (N_2007,In_259,In_30);
xnor U2008 (N_2008,In_961,In_1989);
and U2009 (N_2009,In_2283,In_1778);
xnor U2010 (N_2010,In_506,In_228);
or U2011 (N_2011,In_1575,In_220);
xor U2012 (N_2012,In_2417,In_1079);
and U2013 (N_2013,In_2006,In_204);
nor U2014 (N_2014,In_21,In_1187);
or U2015 (N_2015,In_1467,In_1308);
nor U2016 (N_2016,In_1999,In_826);
nand U2017 (N_2017,In_2366,In_840);
nor U2018 (N_2018,In_30,In_436);
and U2019 (N_2019,In_445,In_1859);
nand U2020 (N_2020,In_361,In_180);
nand U2021 (N_2021,In_1077,In_1635);
nand U2022 (N_2022,In_2054,In_64);
nor U2023 (N_2023,In_1357,In_1384);
xor U2024 (N_2024,In_1711,In_2297);
xor U2025 (N_2025,In_1769,In_1019);
nand U2026 (N_2026,In_1837,In_1003);
and U2027 (N_2027,In_1904,In_2147);
and U2028 (N_2028,In_1739,In_684);
or U2029 (N_2029,In_515,In_2430);
and U2030 (N_2030,In_1297,In_1249);
and U2031 (N_2031,In_1261,In_748);
nand U2032 (N_2032,In_861,In_1693);
or U2033 (N_2033,In_857,In_61);
and U2034 (N_2034,In_814,In_691);
and U2035 (N_2035,In_1363,In_2265);
nand U2036 (N_2036,In_1218,In_921);
or U2037 (N_2037,In_1638,In_897);
nor U2038 (N_2038,In_2269,In_2176);
and U2039 (N_2039,In_925,In_2367);
or U2040 (N_2040,In_9,In_1651);
xor U2041 (N_2041,In_369,In_195);
nand U2042 (N_2042,In_1800,In_1910);
or U2043 (N_2043,In_1319,In_973);
or U2044 (N_2044,In_423,In_2041);
xor U2045 (N_2045,In_1389,In_22);
xor U2046 (N_2046,In_710,In_1878);
xor U2047 (N_2047,In_1855,In_2332);
or U2048 (N_2048,In_273,In_2166);
and U2049 (N_2049,In_1714,In_2260);
and U2050 (N_2050,In_1516,In_115);
and U2051 (N_2051,In_729,In_2007);
nand U2052 (N_2052,In_622,In_2315);
and U2053 (N_2053,In_969,In_1982);
xor U2054 (N_2054,In_1246,In_406);
xnor U2055 (N_2055,In_1025,In_2163);
nor U2056 (N_2056,In_706,In_452);
xor U2057 (N_2057,In_2247,In_425);
nand U2058 (N_2058,In_2267,In_2346);
nand U2059 (N_2059,In_1728,In_526);
nor U2060 (N_2060,In_768,In_165);
nand U2061 (N_2061,In_397,In_358);
or U2062 (N_2062,In_1251,In_1555);
and U2063 (N_2063,In_159,In_1912);
xor U2064 (N_2064,In_264,In_1658);
nor U2065 (N_2065,In_1406,In_2420);
nand U2066 (N_2066,In_1323,In_873);
nand U2067 (N_2067,In_46,In_2221);
or U2068 (N_2068,In_1238,In_1003);
nand U2069 (N_2069,In_2429,In_534);
nor U2070 (N_2070,In_2306,In_480);
xor U2071 (N_2071,In_2024,In_772);
or U2072 (N_2072,In_2286,In_428);
xnor U2073 (N_2073,In_810,In_2233);
or U2074 (N_2074,In_1781,In_2479);
nand U2075 (N_2075,In_1018,In_2344);
xor U2076 (N_2076,In_1886,In_658);
or U2077 (N_2077,In_1538,In_404);
nand U2078 (N_2078,In_1774,In_1723);
xor U2079 (N_2079,In_212,In_1029);
and U2080 (N_2080,In_1140,In_979);
and U2081 (N_2081,In_839,In_2468);
or U2082 (N_2082,In_1977,In_1662);
or U2083 (N_2083,In_73,In_667);
nor U2084 (N_2084,In_2083,In_1487);
and U2085 (N_2085,In_1936,In_649);
nand U2086 (N_2086,In_2186,In_1901);
xnor U2087 (N_2087,In_1788,In_2190);
nor U2088 (N_2088,In_2190,In_1757);
xnor U2089 (N_2089,In_1032,In_2389);
nand U2090 (N_2090,In_1595,In_1449);
nor U2091 (N_2091,In_1410,In_448);
nor U2092 (N_2092,In_465,In_392);
and U2093 (N_2093,In_2219,In_1078);
or U2094 (N_2094,In_1164,In_174);
or U2095 (N_2095,In_327,In_986);
or U2096 (N_2096,In_1811,In_828);
xor U2097 (N_2097,In_696,In_1657);
and U2098 (N_2098,In_1909,In_675);
nand U2099 (N_2099,In_837,In_2356);
nor U2100 (N_2100,In_1987,In_1567);
nor U2101 (N_2101,In_1934,In_288);
nand U2102 (N_2102,In_1073,In_2218);
xnor U2103 (N_2103,In_881,In_787);
xnor U2104 (N_2104,In_2031,In_1286);
nor U2105 (N_2105,In_2217,In_921);
nor U2106 (N_2106,In_1553,In_1625);
xnor U2107 (N_2107,In_1051,In_1400);
xor U2108 (N_2108,In_1816,In_409);
nor U2109 (N_2109,In_2290,In_1980);
xor U2110 (N_2110,In_625,In_1342);
nor U2111 (N_2111,In_2448,In_2169);
nor U2112 (N_2112,In_1989,In_1937);
and U2113 (N_2113,In_248,In_1535);
or U2114 (N_2114,In_2497,In_287);
or U2115 (N_2115,In_2108,In_1985);
nand U2116 (N_2116,In_859,In_2467);
nand U2117 (N_2117,In_329,In_241);
or U2118 (N_2118,In_1494,In_1455);
xnor U2119 (N_2119,In_297,In_1449);
nor U2120 (N_2120,In_2176,In_4);
xor U2121 (N_2121,In_1939,In_2039);
nand U2122 (N_2122,In_2162,In_1618);
or U2123 (N_2123,In_527,In_1925);
or U2124 (N_2124,In_547,In_2346);
nor U2125 (N_2125,In_53,In_2029);
nor U2126 (N_2126,In_2215,In_918);
and U2127 (N_2127,In_1174,In_360);
nor U2128 (N_2128,In_830,In_166);
xnor U2129 (N_2129,In_21,In_1304);
nor U2130 (N_2130,In_2349,In_2295);
or U2131 (N_2131,In_1091,In_649);
and U2132 (N_2132,In_2198,In_362);
nand U2133 (N_2133,In_1379,In_2250);
or U2134 (N_2134,In_1329,In_1478);
and U2135 (N_2135,In_1314,In_1575);
and U2136 (N_2136,In_728,In_2408);
nor U2137 (N_2137,In_996,In_2475);
nand U2138 (N_2138,In_2016,In_1272);
xor U2139 (N_2139,In_356,In_1728);
or U2140 (N_2140,In_2298,In_212);
nand U2141 (N_2141,In_1474,In_2272);
nor U2142 (N_2142,In_1750,In_1336);
or U2143 (N_2143,In_733,In_851);
nor U2144 (N_2144,In_1046,In_1753);
or U2145 (N_2145,In_2305,In_713);
nor U2146 (N_2146,In_708,In_2368);
or U2147 (N_2147,In_501,In_933);
nor U2148 (N_2148,In_129,In_73);
and U2149 (N_2149,In_342,In_1579);
nand U2150 (N_2150,In_1256,In_544);
nand U2151 (N_2151,In_1464,In_830);
or U2152 (N_2152,In_1268,In_223);
or U2153 (N_2153,In_111,In_364);
nor U2154 (N_2154,In_1203,In_1748);
and U2155 (N_2155,In_526,In_1390);
xor U2156 (N_2156,In_502,In_1952);
nand U2157 (N_2157,In_2096,In_1518);
nor U2158 (N_2158,In_2020,In_556);
and U2159 (N_2159,In_1120,In_1573);
and U2160 (N_2160,In_2299,In_195);
xor U2161 (N_2161,In_769,In_1903);
nand U2162 (N_2162,In_2154,In_1463);
or U2163 (N_2163,In_1200,In_588);
or U2164 (N_2164,In_72,In_874);
nor U2165 (N_2165,In_340,In_898);
and U2166 (N_2166,In_2257,In_355);
nand U2167 (N_2167,In_1219,In_1813);
xnor U2168 (N_2168,In_555,In_1403);
nor U2169 (N_2169,In_2439,In_1111);
xor U2170 (N_2170,In_854,In_2480);
nor U2171 (N_2171,In_438,In_813);
nor U2172 (N_2172,In_1432,In_1965);
nor U2173 (N_2173,In_2438,In_582);
nand U2174 (N_2174,In_2076,In_2024);
and U2175 (N_2175,In_977,In_2299);
or U2176 (N_2176,In_1247,In_570);
and U2177 (N_2177,In_250,In_1925);
nor U2178 (N_2178,In_1558,In_1451);
nor U2179 (N_2179,In_1625,In_1788);
nor U2180 (N_2180,In_930,In_1233);
or U2181 (N_2181,In_1083,In_97);
nor U2182 (N_2182,In_1410,In_1308);
and U2183 (N_2183,In_1115,In_550);
xnor U2184 (N_2184,In_267,In_750);
nor U2185 (N_2185,In_1239,In_1620);
xor U2186 (N_2186,In_216,In_137);
nor U2187 (N_2187,In_1451,In_1680);
xnor U2188 (N_2188,In_729,In_2052);
nand U2189 (N_2189,In_2405,In_1780);
nor U2190 (N_2190,In_668,In_345);
or U2191 (N_2191,In_1410,In_1400);
nor U2192 (N_2192,In_1452,In_1764);
xor U2193 (N_2193,In_567,In_2036);
or U2194 (N_2194,In_2257,In_1351);
nand U2195 (N_2195,In_1710,In_525);
nand U2196 (N_2196,In_1152,In_1204);
nor U2197 (N_2197,In_234,In_1614);
and U2198 (N_2198,In_585,In_1056);
and U2199 (N_2199,In_2262,In_2014);
or U2200 (N_2200,In_437,In_463);
nand U2201 (N_2201,In_1944,In_1542);
nand U2202 (N_2202,In_2029,In_1350);
nor U2203 (N_2203,In_2219,In_581);
nor U2204 (N_2204,In_1973,In_203);
or U2205 (N_2205,In_1642,In_247);
nand U2206 (N_2206,In_1604,In_952);
or U2207 (N_2207,In_372,In_1915);
nand U2208 (N_2208,In_863,In_421);
nor U2209 (N_2209,In_2476,In_1102);
nand U2210 (N_2210,In_2360,In_736);
or U2211 (N_2211,In_1731,In_2010);
or U2212 (N_2212,In_1037,In_1510);
and U2213 (N_2213,In_1442,In_1882);
and U2214 (N_2214,In_1192,In_1581);
xor U2215 (N_2215,In_270,In_1972);
and U2216 (N_2216,In_797,In_679);
and U2217 (N_2217,In_635,In_157);
xor U2218 (N_2218,In_1639,In_845);
nand U2219 (N_2219,In_1864,In_1127);
nand U2220 (N_2220,In_1264,In_348);
nand U2221 (N_2221,In_1705,In_1936);
or U2222 (N_2222,In_293,In_274);
nor U2223 (N_2223,In_1809,In_1111);
nand U2224 (N_2224,In_1477,In_1108);
or U2225 (N_2225,In_170,In_1468);
or U2226 (N_2226,In_2419,In_631);
or U2227 (N_2227,In_1473,In_950);
and U2228 (N_2228,In_2358,In_1701);
nor U2229 (N_2229,In_1148,In_339);
nor U2230 (N_2230,In_1704,In_1099);
nor U2231 (N_2231,In_2074,In_367);
nand U2232 (N_2232,In_101,In_2224);
or U2233 (N_2233,In_899,In_1761);
nor U2234 (N_2234,In_368,In_1758);
xor U2235 (N_2235,In_1546,In_1479);
nand U2236 (N_2236,In_54,In_811);
or U2237 (N_2237,In_1111,In_722);
nand U2238 (N_2238,In_520,In_312);
nor U2239 (N_2239,In_1000,In_534);
or U2240 (N_2240,In_999,In_72);
nand U2241 (N_2241,In_1666,In_349);
nor U2242 (N_2242,In_2486,In_302);
nor U2243 (N_2243,In_340,In_1681);
nand U2244 (N_2244,In_1844,In_720);
xnor U2245 (N_2245,In_1018,In_2322);
and U2246 (N_2246,In_259,In_1838);
nand U2247 (N_2247,In_405,In_37);
or U2248 (N_2248,In_114,In_1775);
xnor U2249 (N_2249,In_44,In_2049);
nand U2250 (N_2250,In_629,In_1619);
or U2251 (N_2251,In_1162,In_1499);
nor U2252 (N_2252,In_83,In_974);
and U2253 (N_2253,In_149,In_972);
nor U2254 (N_2254,In_18,In_767);
or U2255 (N_2255,In_2392,In_1663);
xnor U2256 (N_2256,In_233,In_1303);
nor U2257 (N_2257,In_2336,In_569);
xor U2258 (N_2258,In_571,In_667);
or U2259 (N_2259,In_275,In_1264);
xnor U2260 (N_2260,In_2475,In_555);
or U2261 (N_2261,In_1695,In_367);
xor U2262 (N_2262,In_1246,In_1133);
nor U2263 (N_2263,In_1452,In_630);
nand U2264 (N_2264,In_1127,In_1988);
or U2265 (N_2265,In_2111,In_53);
nor U2266 (N_2266,In_1143,In_1985);
and U2267 (N_2267,In_39,In_907);
and U2268 (N_2268,In_936,In_1317);
and U2269 (N_2269,In_1913,In_1878);
or U2270 (N_2270,In_1435,In_1428);
or U2271 (N_2271,In_261,In_390);
and U2272 (N_2272,In_1208,In_1555);
and U2273 (N_2273,In_2034,In_1718);
and U2274 (N_2274,In_1171,In_699);
or U2275 (N_2275,In_106,In_2017);
or U2276 (N_2276,In_112,In_1783);
nand U2277 (N_2277,In_22,In_1959);
and U2278 (N_2278,In_2125,In_2034);
or U2279 (N_2279,In_922,In_456);
and U2280 (N_2280,In_1276,In_1694);
nor U2281 (N_2281,In_1018,In_1096);
or U2282 (N_2282,In_1449,In_1548);
or U2283 (N_2283,In_1977,In_388);
nor U2284 (N_2284,In_960,In_863);
and U2285 (N_2285,In_1613,In_1670);
xnor U2286 (N_2286,In_1628,In_2118);
nor U2287 (N_2287,In_1462,In_2193);
nor U2288 (N_2288,In_1481,In_1101);
and U2289 (N_2289,In_1666,In_878);
xnor U2290 (N_2290,In_282,In_47);
or U2291 (N_2291,In_1687,In_1054);
and U2292 (N_2292,In_2071,In_2258);
nand U2293 (N_2293,In_553,In_1567);
xnor U2294 (N_2294,In_606,In_1895);
or U2295 (N_2295,In_1332,In_584);
and U2296 (N_2296,In_1843,In_2281);
or U2297 (N_2297,In_2316,In_1023);
nor U2298 (N_2298,In_1542,In_2111);
xnor U2299 (N_2299,In_176,In_1107);
or U2300 (N_2300,In_837,In_923);
and U2301 (N_2301,In_1481,In_974);
nor U2302 (N_2302,In_1049,In_2014);
xnor U2303 (N_2303,In_920,In_573);
xnor U2304 (N_2304,In_1207,In_554);
and U2305 (N_2305,In_2306,In_548);
xor U2306 (N_2306,In_2180,In_2164);
xnor U2307 (N_2307,In_1286,In_865);
nand U2308 (N_2308,In_1717,In_1882);
nor U2309 (N_2309,In_1808,In_962);
or U2310 (N_2310,In_1488,In_2063);
and U2311 (N_2311,In_2175,In_1180);
nor U2312 (N_2312,In_127,In_680);
xnor U2313 (N_2313,In_854,In_1636);
or U2314 (N_2314,In_2038,In_1838);
and U2315 (N_2315,In_921,In_391);
nor U2316 (N_2316,In_2150,In_449);
and U2317 (N_2317,In_1268,In_827);
xnor U2318 (N_2318,In_1555,In_1183);
or U2319 (N_2319,In_1903,In_492);
xnor U2320 (N_2320,In_2105,In_2216);
or U2321 (N_2321,In_1279,In_1741);
nor U2322 (N_2322,In_855,In_359);
nand U2323 (N_2323,In_1209,In_1595);
or U2324 (N_2324,In_2220,In_1747);
nor U2325 (N_2325,In_1946,In_37);
xor U2326 (N_2326,In_523,In_1157);
and U2327 (N_2327,In_863,In_961);
and U2328 (N_2328,In_968,In_338);
and U2329 (N_2329,In_157,In_804);
and U2330 (N_2330,In_2333,In_1867);
and U2331 (N_2331,In_2052,In_12);
or U2332 (N_2332,In_146,In_1696);
nor U2333 (N_2333,In_2413,In_1986);
or U2334 (N_2334,In_2081,In_188);
or U2335 (N_2335,In_1801,In_1710);
xnor U2336 (N_2336,In_1785,In_553);
and U2337 (N_2337,In_1427,In_2388);
nor U2338 (N_2338,In_1910,In_1904);
or U2339 (N_2339,In_403,In_14);
nor U2340 (N_2340,In_600,In_895);
nand U2341 (N_2341,In_732,In_2);
nor U2342 (N_2342,In_211,In_1541);
xnor U2343 (N_2343,In_290,In_160);
xnor U2344 (N_2344,In_1650,In_172);
nor U2345 (N_2345,In_437,In_1389);
nor U2346 (N_2346,In_1640,In_1483);
xnor U2347 (N_2347,In_1074,In_396);
nand U2348 (N_2348,In_986,In_1814);
xnor U2349 (N_2349,In_1186,In_802);
xor U2350 (N_2350,In_2189,In_0);
nor U2351 (N_2351,In_2104,In_1576);
xnor U2352 (N_2352,In_803,In_1947);
nand U2353 (N_2353,In_1417,In_1744);
or U2354 (N_2354,In_2367,In_597);
nor U2355 (N_2355,In_1708,In_25);
or U2356 (N_2356,In_2495,In_524);
nand U2357 (N_2357,In_1518,In_2262);
and U2358 (N_2358,In_1348,In_2189);
and U2359 (N_2359,In_1570,In_570);
nand U2360 (N_2360,In_1687,In_1276);
or U2361 (N_2361,In_47,In_1806);
nor U2362 (N_2362,In_1144,In_801);
nor U2363 (N_2363,In_984,In_2319);
or U2364 (N_2364,In_1577,In_541);
nand U2365 (N_2365,In_2083,In_1786);
xor U2366 (N_2366,In_1785,In_1489);
xor U2367 (N_2367,In_519,In_2195);
nor U2368 (N_2368,In_2312,In_615);
nor U2369 (N_2369,In_344,In_1820);
xnor U2370 (N_2370,In_1982,In_707);
xnor U2371 (N_2371,In_2350,In_746);
and U2372 (N_2372,In_272,In_375);
and U2373 (N_2373,In_1440,In_265);
xor U2374 (N_2374,In_1827,In_415);
and U2375 (N_2375,In_1901,In_1782);
nand U2376 (N_2376,In_1216,In_996);
and U2377 (N_2377,In_28,In_2032);
and U2378 (N_2378,In_1836,In_297);
nor U2379 (N_2379,In_2096,In_1753);
and U2380 (N_2380,In_430,In_2470);
xor U2381 (N_2381,In_192,In_2203);
and U2382 (N_2382,In_2139,In_1472);
xnor U2383 (N_2383,In_818,In_691);
or U2384 (N_2384,In_746,In_1231);
and U2385 (N_2385,In_171,In_1939);
or U2386 (N_2386,In_1283,In_461);
and U2387 (N_2387,In_1209,In_629);
nand U2388 (N_2388,In_1114,In_2375);
nor U2389 (N_2389,In_476,In_1617);
nor U2390 (N_2390,In_1949,In_86);
nand U2391 (N_2391,In_711,In_2292);
or U2392 (N_2392,In_658,In_1051);
and U2393 (N_2393,In_423,In_1171);
nand U2394 (N_2394,In_108,In_2365);
nor U2395 (N_2395,In_1945,In_1230);
or U2396 (N_2396,In_944,In_839);
xor U2397 (N_2397,In_1826,In_1713);
nand U2398 (N_2398,In_1761,In_1407);
or U2399 (N_2399,In_1508,In_729);
or U2400 (N_2400,In_2246,In_195);
xor U2401 (N_2401,In_2283,In_1922);
nand U2402 (N_2402,In_2263,In_722);
nand U2403 (N_2403,In_1004,In_1412);
or U2404 (N_2404,In_1366,In_1651);
nor U2405 (N_2405,In_1024,In_1256);
nand U2406 (N_2406,In_777,In_1806);
nand U2407 (N_2407,In_2105,In_1778);
xnor U2408 (N_2408,In_2045,In_1638);
xnor U2409 (N_2409,In_1920,In_824);
nor U2410 (N_2410,In_2394,In_1451);
nor U2411 (N_2411,In_1313,In_1140);
nor U2412 (N_2412,In_4,In_1933);
or U2413 (N_2413,In_360,In_940);
xor U2414 (N_2414,In_405,In_1869);
xor U2415 (N_2415,In_2111,In_27);
and U2416 (N_2416,In_701,In_1702);
xnor U2417 (N_2417,In_778,In_664);
and U2418 (N_2418,In_1351,In_265);
or U2419 (N_2419,In_1244,In_1514);
or U2420 (N_2420,In_1228,In_337);
nor U2421 (N_2421,In_1704,In_2124);
xnor U2422 (N_2422,In_1997,In_1061);
and U2423 (N_2423,In_2162,In_731);
or U2424 (N_2424,In_541,In_1939);
and U2425 (N_2425,In_2012,In_341);
nor U2426 (N_2426,In_296,In_2460);
nand U2427 (N_2427,In_1561,In_2137);
nor U2428 (N_2428,In_1757,In_133);
and U2429 (N_2429,In_2161,In_1028);
or U2430 (N_2430,In_289,In_110);
and U2431 (N_2431,In_1752,In_649);
nand U2432 (N_2432,In_1555,In_1244);
and U2433 (N_2433,In_17,In_217);
or U2434 (N_2434,In_2140,In_1565);
and U2435 (N_2435,In_1570,In_1537);
nor U2436 (N_2436,In_2057,In_2376);
nor U2437 (N_2437,In_669,In_555);
nor U2438 (N_2438,In_372,In_1001);
nand U2439 (N_2439,In_1168,In_2468);
nor U2440 (N_2440,In_791,In_732);
nand U2441 (N_2441,In_2098,In_2233);
or U2442 (N_2442,In_2417,In_280);
nand U2443 (N_2443,In_229,In_248);
nand U2444 (N_2444,In_26,In_1988);
nor U2445 (N_2445,In_674,In_935);
nor U2446 (N_2446,In_2287,In_1293);
nand U2447 (N_2447,In_1208,In_1295);
nor U2448 (N_2448,In_1414,In_347);
or U2449 (N_2449,In_1417,In_1872);
or U2450 (N_2450,In_2094,In_1580);
xnor U2451 (N_2451,In_756,In_380);
or U2452 (N_2452,In_2188,In_2254);
xnor U2453 (N_2453,In_1921,In_2138);
xor U2454 (N_2454,In_1126,In_1367);
nor U2455 (N_2455,In_318,In_2078);
and U2456 (N_2456,In_1875,In_1606);
or U2457 (N_2457,In_2473,In_1287);
nor U2458 (N_2458,In_242,In_1707);
nand U2459 (N_2459,In_494,In_1624);
xor U2460 (N_2460,In_1489,In_88);
or U2461 (N_2461,In_959,In_2390);
or U2462 (N_2462,In_2090,In_686);
and U2463 (N_2463,In_2476,In_2350);
nor U2464 (N_2464,In_2200,In_2087);
nand U2465 (N_2465,In_328,In_1168);
xnor U2466 (N_2466,In_2393,In_233);
or U2467 (N_2467,In_18,In_830);
and U2468 (N_2468,In_1167,In_2293);
nand U2469 (N_2469,In_2040,In_536);
xor U2470 (N_2470,In_1471,In_1235);
nor U2471 (N_2471,In_1535,In_1299);
nor U2472 (N_2472,In_1164,In_684);
nor U2473 (N_2473,In_1331,In_101);
nand U2474 (N_2474,In_379,In_1551);
and U2475 (N_2475,In_876,In_1819);
nor U2476 (N_2476,In_31,In_2484);
xnor U2477 (N_2477,In_1334,In_1010);
xor U2478 (N_2478,In_1671,In_1721);
or U2479 (N_2479,In_1001,In_14);
nor U2480 (N_2480,In_1032,In_1848);
or U2481 (N_2481,In_1971,In_609);
and U2482 (N_2482,In_1421,In_579);
nor U2483 (N_2483,In_349,In_84);
or U2484 (N_2484,In_457,In_193);
or U2485 (N_2485,In_2440,In_598);
nand U2486 (N_2486,In_2226,In_66);
or U2487 (N_2487,In_1681,In_1938);
or U2488 (N_2488,In_909,In_596);
nor U2489 (N_2489,In_1380,In_383);
nand U2490 (N_2490,In_895,In_4);
nand U2491 (N_2491,In_519,In_342);
or U2492 (N_2492,In_744,In_1489);
or U2493 (N_2493,In_67,In_984);
xnor U2494 (N_2494,In_1967,In_1985);
and U2495 (N_2495,In_665,In_924);
nand U2496 (N_2496,In_2058,In_2448);
xnor U2497 (N_2497,In_2226,In_968);
nor U2498 (N_2498,In_2366,In_200);
nor U2499 (N_2499,In_1361,In_2473);
nor U2500 (N_2500,N_860,N_1616);
and U2501 (N_2501,N_1950,N_1964);
nand U2502 (N_2502,N_1325,N_733);
and U2503 (N_2503,N_1215,N_430);
nor U2504 (N_2504,N_1329,N_1338);
nor U2505 (N_2505,N_2332,N_1822);
and U2506 (N_2506,N_1821,N_799);
nand U2507 (N_2507,N_1013,N_605);
nand U2508 (N_2508,N_1566,N_1496);
nor U2509 (N_2509,N_2484,N_2373);
xor U2510 (N_2510,N_1607,N_388);
or U2511 (N_2511,N_1728,N_1836);
nor U2512 (N_2512,N_1135,N_574);
nand U2513 (N_2513,N_1777,N_1384);
and U2514 (N_2514,N_1605,N_2094);
xnor U2515 (N_2515,N_177,N_1889);
or U2516 (N_2516,N_1312,N_2463);
nand U2517 (N_2517,N_612,N_1517);
or U2518 (N_2518,N_532,N_1952);
xor U2519 (N_2519,N_812,N_1596);
or U2520 (N_2520,N_764,N_1352);
nor U2521 (N_2521,N_1511,N_2177);
nand U2522 (N_2522,N_1880,N_1983);
nand U2523 (N_2523,N_1005,N_2004);
nand U2524 (N_2524,N_1411,N_93);
nand U2525 (N_2525,N_1606,N_1675);
xor U2526 (N_2526,N_1038,N_499);
nand U2527 (N_2527,N_1297,N_1724);
nand U2528 (N_2528,N_1590,N_2308);
and U2529 (N_2529,N_8,N_880);
nor U2530 (N_2530,N_2456,N_776);
xnor U2531 (N_2531,N_1594,N_1418);
and U2532 (N_2532,N_1377,N_1049);
nand U2533 (N_2533,N_15,N_2488);
nor U2534 (N_2534,N_398,N_1505);
nand U2535 (N_2535,N_644,N_929);
nor U2536 (N_2536,N_2050,N_707);
xnor U2537 (N_2537,N_990,N_2196);
or U2538 (N_2538,N_88,N_276);
xnor U2539 (N_2539,N_908,N_766);
nand U2540 (N_2540,N_145,N_1421);
xnor U2541 (N_2541,N_1318,N_2096);
nand U2542 (N_2542,N_1404,N_932);
nor U2543 (N_2543,N_789,N_2175);
nand U2544 (N_2544,N_508,N_1916);
nand U2545 (N_2545,N_474,N_2181);
and U2546 (N_2546,N_1472,N_435);
xor U2547 (N_2547,N_2281,N_1962);
xnor U2548 (N_2548,N_39,N_782);
nand U2549 (N_2549,N_993,N_1798);
nor U2550 (N_2550,N_592,N_709);
nand U2551 (N_2551,N_1931,N_510);
and U2552 (N_2552,N_2126,N_655);
nand U2553 (N_2553,N_852,N_610);
xor U2554 (N_2554,N_1165,N_2228);
or U2555 (N_2555,N_1294,N_2295);
xnor U2556 (N_2556,N_118,N_1579);
or U2557 (N_2557,N_280,N_2122);
and U2558 (N_2558,N_2118,N_1541);
nand U2559 (N_2559,N_42,N_1035);
and U2560 (N_2560,N_1126,N_101);
or U2561 (N_2561,N_1848,N_397);
or U2562 (N_2562,N_2345,N_127);
nor U2563 (N_2563,N_1401,N_2365);
or U2564 (N_2564,N_300,N_1920);
or U2565 (N_2565,N_1892,N_2315);
nand U2566 (N_2566,N_1858,N_985);
or U2567 (N_2567,N_30,N_1900);
nand U2568 (N_2568,N_673,N_1857);
and U2569 (N_2569,N_1768,N_2452);
nand U2570 (N_2570,N_2042,N_1520);
or U2571 (N_2571,N_1844,N_1122);
xnor U2572 (N_2572,N_1965,N_1519);
nand U2573 (N_2573,N_2113,N_2271);
nand U2574 (N_2574,N_495,N_914);
nor U2575 (N_2575,N_1899,N_69);
and U2576 (N_2576,N_1568,N_110);
nor U2577 (N_2577,N_164,N_0);
xor U2578 (N_2578,N_1080,N_197);
and U2579 (N_2579,N_1308,N_432);
and U2580 (N_2580,N_311,N_103);
nand U2581 (N_2581,N_1361,N_218);
and U2582 (N_2582,N_232,N_146);
xor U2583 (N_2583,N_1641,N_2013);
and U2584 (N_2584,N_2162,N_729);
nor U2585 (N_2585,N_1694,N_333);
xor U2586 (N_2586,N_1640,N_1451);
or U2587 (N_2587,N_994,N_426);
xnor U2588 (N_2588,N_423,N_1226);
or U2589 (N_2589,N_669,N_948);
xnor U2590 (N_2590,N_1056,N_1570);
and U2591 (N_2591,N_702,N_215);
xnor U2592 (N_2592,N_978,N_711);
and U2593 (N_2593,N_570,N_1033);
nand U2594 (N_2594,N_1551,N_1879);
xor U2595 (N_2595,N_1207,N_445);
and U2596 (N_2596,N_2427,N_1604);
xnor U2597 (N_2597,N_2421,N_964);
nand U2598 (N_2598,N_571,N_1054);
or U2599 (N_2599,N_1015,N_2286);
and U2600 (N_2600,N_105,N_730);
or U2601 (N_2601,N_336,N_1389);
xnor U2602 (N_2602,N_1524,N_1250);
or U2603 (N_2603,N_1462,N_420);
or U2604 (N_2604,N_2375,N_1549);
nand U2605 (N_2605,N_1529,N_1647);
xnor U2606 (N_2606,N_556,N_791);
xnor U2607 (N_2607,N_77,N_181);
or U2608 (N_2608,N_469,N_1940);
or U2609 (N_2609,N_1837,N_1202);
nor U2610 (N_2610,N_1275,N_2193);
nor U2611 (N_2611,N_2076,N_1749);
nand U2612 (N_2612,N_316,N_1907);
and U2613 (N_2613,N_477,N_2259);
and U2614 (N_2614,N_62,N_384);
and U2615 (N_2615,N_1637,N_493);
or U2616 (N_2616,N_2248,N_35);
and U2617 (N_2617,N_987,N_2104);
nand U2618 (N_2618,N_1181,N_1695);
nand U2619 (N_2619,N_868,N_1809);
and U2620 (N_2620,N_2361,N_1435);
nor U2621 (N_2621,N_2357,N_1058);
or U2622 (N_2622,N_1939,N_2448);
nor U2623 (N_2623,N_1806,N_1718);
nand U2624 (N_2624,N_1097,N_1494);
or U2625 (N_2625,N_1351,N_43);
nand U2626 (N_2626,N_1769,N_596);
or U2627 (N_2627,N_599,N_1373);
xnor U2628 (N_2628,N_2416,N_200);
or U2629 (N_2629,N_1774,N_583);
xor U2630 (N_2630,N_684,N_19);
xor U2631 (N_2631,N_1265,N_958);
xnor U2632 (N_2632,N_1930,N_1738);
and U2633 (N_2633,N_433,N_170);
and U2634 (N_2634,N_235,N_554);
xnor U2635 (N_2635,N_98,N_1788);
or U2636 (N_2636,N_2316,N_1781);
nand U2637 (N_2637,N_1201,N_1881);
and U2638 (N_2638,N_1565,N_66);
and U2639 (N_2639,N_1129,N_32);
nand U2640 (N_2640,N_338,N_2163);
and U2641 (N_2641,N_1146,N_1386);
or U2642 (N_2642,N_1757,N_1317);
nand U2643 (N_2643,N_380,N_2433);
xor U2644 (N_2644,N_1395,N_2238);
nand U2645 (N_2645,N_503,N_1855);
or U2646 (N_2646,N_1152,N_535);
and U2647 (N_2647,N_34,N_1089);
and U2648 (N_2648,N_2097,N_1330);
xnor U2649 (N_2649,N_143,N_1556);
nor U2650 (N_2650,N_717,N_1131);
nand U2651 (N_2651,N_1743,N_2307);
nor U2652 (N_2652,N_1052,N_1751);
nand U2653 (N_2653,N_378,N_869);
nor U2654 (N_2654,N_2413,N_2465);
xnor U2655 (N_2655,N_1113,N_642);
or U2656 (N_2656,N_1702,N_838);
or U2657 (N_2657,N_2366,N_1984);
nor U2658 (N_2658,N_74,N_2026);
nand U2659 (N_2659,N_418,N_2233);
or U2660 (N_2660,N_1854,N_255);
and U2661 (N_2661,N_2401,N_1018);
or U2662 (N_2662,N_2222,N_873);
xor U2663 (N_2663,N_2207,N_370);
nand U2664 (N_2664,N_1353,N_1526);
nand U2665 (N_2665,N_2493,N_810);
and U2666 (N_2666,N_1633,N_1614);
xnor U2667 (N_2667,N_1211,N_509);
or U2668 (N_2668,N_2420,N_390);
nor U2669 (N_2669,N_2187,N_1117);
or U2670 (N_2670,N_847,N_462);
and U2671 (N_2671,N_1234,N_1929);
nand U2672 (N_2672,N_213,N_885);
xor U2673 (N_2673,N_1954,N_476);
xnor U2674 (N_2674,N_1229,N_2393);
or U2675 (N_2675,N_1658,N_1994);
and U2676 (N_2676,N_1499,N_2123);
nand U2677 (N_2677,N_394,N_792);
xor U2678 (N_2678,N_1742,N_1471);
xor U2679 (N_2679,N_2344,N_392);
nor U2680 (N_2680,N_2061,N_162);
nor U2681 (N_2681,N_1368,N_154);
nor U2682 (N_2682,N_1167,N_1066);
and U2683 (N_2683,N_1942,N_23);
nand U2684 (N_2684,N_2125,N_2204);
and U2685 (N_2685,N_1729,N_1895);
and U2686 (N_2686,N_2329,N_1163);
or U2687 (N_2687,N_2184,N_220);
xnor U2688 (N_2688,N_1528,N_1592);
and U2689 (N_2689,N_1642,N_1871);
and U2690 (N_2690,N_1951,N_1655);
nor U2691 (N_2691,N_2343,N_168);
nand U2692 (N_2692,N_70,N_153);
or U2693 (N_2693,N_1651,N_1919);
xnor U2694 (N_2694,N_1103,N_1423);
nand U2695 (N_2695,N_1648,N_2230);
or U2696 (N_2696,N_2284,N_102);
or U2697 (N_2697,N_750,N_193);
xnor U2698 (N_2698,N_536,N_1691);
or U2699 (N_2699,N_1241,N_134);
nand U2700 (N_2700,N_2431,N_1230);
nand U2701 (N_2701,N_478,N_1470);
and U2702 (N_2702,N_225,N_119);
nor U2703 (N_2703,N_158,N_1772);
xnor U2704 (N_2704,N_259,N_857);
and U2705 (N_2705,N_1006,N_1620);
nand U2706 (N_2706,N_2009,N_1510);
or U2707 (N_2707,N_892,N_1646);
nor U2708 (N_2708,N_2263,N_1001);
and U2709 (N_2709,N_449,N_2270);
and U2710 (N_2710,N_975,N_1838);
nand U2711 (N_2711,N_2149,N_2132);
nor U2712 (N_2712,N_1552,N_443);
or U2713 (N_2713,N_302,N_683);
xnor U2714 (N_2714,N_2291,N_1007);
or U2715 (N_2715,N_331,N_1224);
nand U2716 (N_2716,N_204,N_2102);
xor U2717 (N_2717,N_1959,N_613);
and U2718 (N_2718,N_356,N_1652);
or U2719 (N_2719,N_521,N_1703);
and U2720 (N_2720,N_1783,N_2156);
nand U2721 (N_2721,N_620,N_1990);
xnor U2722 (N_2722,N_231,N_586);
nand U2723 (N_2723,N_245,N_2227);
nand U2724 (N_2724,N_1561,N_1626);
nor U2725 (N_2725,N_827,N_1328);
and U2726 (N_2726,N_494,N_822);
xor U2727 (N_2727,N_1321,N_2188);
or U2728 (N_2728,N_1461,N_1672);
nand U2729 (N_2729,N_910,N_770);
nor U2730 (N_2730,N_2048,N_1782);
xnor U2731 (N_2731,N_2453,N_2392);
nand U2732 (N_2732,N_1019,N_560);
nor U2733 (N_2733,N_1660,N_242);
or U2734 (N_2734,N_486,N_1078);
or U2735 (N_2735,N_171,N_1824);
nand U2736 (N_2736,N_2014,N_2245);
xnor U2737 (N_2737,N_344,N_2110);
or U2738 (N_2738,N_1589,N_679);
nand U2739 (N_2739,N_45,N_920);
or U2740 (N_2740,N_630,N_1567);
nor U2741 (N_2741,N_1903,N_51);
and U2742 (N_2742,N_90,N_38);
nand U2743 (N_2743,N_2243,N_1831);
and U2744 (N_2744,N_685,N_715);
or U2745 (N_2745,N_1797,N_272);
xor U2746 (N_2746,N_1323,N_2112);
xnor U2747 (N_2747,N_523,N_1346);
xor U2748 (N_2748,N_1828,N_1300);
and U2749 (N_2749,N_1538,N_1755);
nor U2750 (N_2750,N_1185,N_754);
nor U2751 (N_2751,N_135,N_44);
xor U2752 (N_2752,N_624,N_1850);
and U2753 (N_2753,N_253,N_755);
nor U2754 (N_2754,N_1509,N_1114);
nand U2755 (N_2755,N_1843,N_1989);
or U2756 (N_2756,N_2334,N_2246);
nand U2757 (N_2757,N_2103,N_2041);
nand U2758 (N_2758,N_2328,N_1140);
and U2759 (N_2759,N_2157,N_1302);
xor U2760 (N_2760,N_2016,N_1814);
nand U2761 (N_2761,N_954,N_1970);
xnor U2762 (N_2762,N_2449,N_2027);
or U2763 (N_2763,N_1905,N_1009);
nor U2764 (N_2764,N_1064,N_796);
xnor U2765 (N_2765,N_840,N_1921);
nor U2766 (N_2766,N_1192,N_81);
nand U2767 (N_2767,N_788,N_1177);
nor U2768 (N_2768,N_2310,N_1223);
and U2769 (N_2769,N_1186,N_16);
nand U2770 (N_2770,N_55,N_1148);
nand U2771 (N_2771,N_515,N_322);
nand U2772 (N_2772,N_537,N_2020);
nor U2773 (N_2773,N_678,N_1041);
nand U2774 (N_2774,N_1799,N_848);
or U2775 (N_2775,N_1915,N_2317);
xnor U2776 (N_2776,N_1073,N_1305);
and U2777 (N_2777,N_894,N_2485);
or U2778 (N_2778,N_1688,N_2073);
xor U2779 (N_2779,N_1971,N_1834);
nor U2780 (N_2780,N_1170,N_653);
and U2781 (N_2781,N_1206,N_1287);
and U2782 (N_2782,N_1422,N_2134);
and U2783 (N_2783,N_1099,N_2079);
nand U2784 (N_2784,N_377,N_1761);
nor U2785 (N_2785,N_863,N_2491);
nor U2786 (N_2786,N_1725,N_1946);
and U2787 (N_2787,N_1363,N_833);
nor U2788 (N_2788,N_917,N_1277);
nand U2789 (N_2789,N_60,N_1639);
and U2790 (N_2790,N_636,N_1051);
and U2791 (N_2791,N_2487,N_1296);
and U2792 (N_2792,N_297,N_1608);
and U2793 (N_2793,N_1654,N_1877);
or U2794 (N_2794,N_1543,N_444);
nor U2795 (N_2795,N_968,N_909);
or U2796 (N_2796,N_1508,N_1853);
xor U2797 (N_2797,N_2075,N_721);
and U2798 (N_2798,N_309,N_434);
nand U2799 (N_2799,N_593,N_1886);
or U2800 (N_2800,N_104,N_549);
or U2801 (N_2801,N_1130,N_224);
xnor U2802 (N_2802,N_1020,N_1488);
nand U2803 (N_2803,N_313,N_745);
xnor U2804 (N_2804,N_1102,N_2250);
or U2805 (N_2805,N_282,N_1671);
or U2806 (N_2806,N_1412,N_199);
nand U2807 (N_2807,N_2160,N_1469);
xnor U2808 (N_2808,N_2235,N_828);
nand U2809 (N_2809,N_1092,N_436);
or U2810 (N_2810,N_552,N_1248);
nand U2811 (N_2811,N_241,N_2064);
or U2812 (N_2812,N_606,N_117);
or U2813 (N_2813,N_175,N_500);
xnor U2814 (N_2814,N_1280,N_1966);
nor U2815 (N_2815,N_1174,N_981);
or U2816 (N_2816,N_1826,N_790);
and U2817 (N_2817,N_1586,N_1100);
or U2818 (N_2818,N_2147,N_1887);
and U2819 (N_2819,N_2273,N_712);
or U2820 (N_2820,N_2011,N_293);
nand U2821 (N_2821,N_1766,N_191);
xor U2822 (N_2822,N_744,N_1467);
xor U2823 (N_2823,N_617,N_279);
xor U2824 (N_2824,N_957,N_835);
xnor U2825 (N_2825,N_126,N_1399);
xnor U2826 (N_2826,N_1453,N_308);
or U2827 (N_2827,N_841,N_2335);
nand U2828 (N_2828,N_188,N_58);
xor U2829 (N_2829,N_1866,N_2483);
and U2830 (N_2830,N_1869,N_2037);
xnor U2831 (N_2831,N_516,N_2339);
nor U2832 (N_2832,N_1062,N_292);
and U2833 (N_2833,N_1872,N_2494);
nor U2834 (N_2834,N_1303,N_2171);
or U2835 (N_2835,N_1358,N_1618);
and U2836 (N_2836,N_1173,N_727);
or U2837 (N_2837,N_122,N_1835);
and U2838 (N_2838,N_1823,N_1406);
or U2839 (N_2839,N_1283,N_68);
xor U2840 (N_2840,N_1164,N_1115);
or U2841 (N_2841,N_1255,N_1686);
nand U2842 (N_2842,N_741,N_2178);
nand U2843 (N_2843,N_821,N_1744);
or U2844 (N_2844,N_1995,N_460);
and U2845 (N_2845,N_648,N_619);
or U2846 (N_2846,N_2060,N_2199);
nand U2847 (N_2847,N_889,N_473);
or U2848 (N_2848,N_2100,N_2425);
nor U2849 (N_2849,N_797,N_115);
and U2850 (N_2850,N_1290,N_611);
and U2851 (N_2851,N_1091,N_618);
and U2852 (N_2852,N_2022,N_298);
nand U2853 (N_2853,N_1619,N_1452);
or U2854 (N_2854,N_913,N_2210);
or U2855 (N_2855,N_466,N_2442);
nor U2856 (N_2856,N_1546,N_2017);
or U2857 (N_2857,N_1678,N_1390);
or U2858 (N_2858,N_1884,N_1021);
xnor U2859 (N_2859,N_912,N_937);
or U2860 (N_2860,N_299,N_984);
xnor U2861 (N_2861,N_690,N_654);
and U2862 (N_2862,N_260,N_1663);
or U2863 (N_2863,N_1554,N_2349);
and U2864 (N_2864,N_2362,N_1210);
xnor U2865 (N_2865,N_2066,N_1839);
and U2866 (N_2866,N_456,N_1053);
nor U2867 (N_2867,N_1810,N_323);
or U2868 (N_2868,N_374,N_97);
or U2869 (N_2869,N_2430,N_875);
and U2870 (N_2870,N_538,N_584);
and U2871 (N_2871,N_2404,N_99);
nor U2872 (N_2872,N_1521,N_2353);
xor U2873 (N_2873,N_73,N_632);
nand U2874 (N_2874,N_1118,N_2168);
and U2875 (N_2875,N_2261,N_1096);
nand U2876 (N_2876,N_1754,N_772);
nor U2877 (N_2877,N_1301,N_1106);
or U2878 (N_2878,N_1503,N_785);
nor U2879 (N_2879,N_2220,N_1832);
nor U2880 (N_2880,N_1104,N_986);
nor U2881 (N_2881,N_33,N_3);
nand U2882 (N_2882,N_656,N_1924);
nand U2883 (N_2883,N_1630,N_1901);
nand U2884 (N_2884,N_1233,N_971);
and U2885 (N_2885,N_1455,N_1004);
or U2886 (N_2886,N_427,N_930);
nand U2887 (N_2887,N_2234,N_625);
xor U2888 (N_2888,N_132,N_1577);
and U2889 (N_2889,N_2285,N_1912);
and U2890 (N_2890,N_448,N_1536);
or U2891 (N_2891,N_1196,N_351);
nor U2892 (N_2892,N_1161,N_1304);
nor U2893 (N_2893,N_2005,N_482);
and U2894 (N_2894,N_933,N_2381);
nand U2895 (N_2895,N_2313,N_289);
nand U2896 (N_2896,N_1251,N_907);
and U2897 (N_2897,N_2260,N_1890);
xor U2898 (N_2898,N_2081,N_890);
or U2899 (N_2899,N_1217,N_566);
or U2900 (N_2900,N_79,N_185);
or U2901 (N_2901,N_2320,N_1157);
xor U2902 (N_2902,N_1627,N_1231);
xnor U2903 (N_2903,N_726,N_222);
or U2904 (N_2904,N_956,N_998);
and U2905 (N_2905,N_735,N_594);
and U2906 (N_2906,N_2256,N_1711);
xnor U2907 (N_2907,N_1057,N_1269);
xor U2908 (N_2908,N_977,N_762);
nor U2909 (N_2909,N_1977,N_725);
nand U2910 (N_2910,N_2202,N_1896);
xnor U2911 (N_2911,N_603,N_1846);
or U2912 (N_2912,N_1506,N_1910);
xnor U2913 (N_2913,N_555,N_262);
and U2914 (N_2914,N_1200,N_1086);
or U2915 (N_2915,N_595,N_410);
xnor U2916 (N_2916,N_2165,N_1827);
or U2917 (N_2917,N_2387,N_992);
or U2918 (N_2918,N_1840,N_1168);
xnor U2919 (N_2919,N_507,N_2206);
xnor U2920 (N_2920,N_1746,N_2194);
xor U2921 (N_2921,N_2476,N_668);
nand U2922 (N_2922,N_439,N_1136);
nor U2923 (N_2923,N_1059,N_393);
nand U2924 (N_2924,N_425,N_1868);
xor U2925 (N_2925,N_2489,N_91);
and U2926 (N_2926,N_2333,N_2305);
nand U2927 (N_2927,N_809,N_455);
and U2928 (N_2928,N_581,N_1862);
nor U2929 (N_2929,N_2192,N_1539);
nand U2930 (N_2930,N_1578,N_2144);
and U2931 (N_2931,N_2380,N_1343);
or U2932 (N_2932,N_2498,N_1046);
xnor U2933 (N_2933,N_697,N_1450);
nor U2934 (N_2934,N_1732,N_1547);
xor U2935 (N_2935,N_962,N_421);
and U2936 (N_2936,N_2180,N_1125);
and U2937 (N_2937,N_1927,N_609);
nand U2938 (N_2938,N_2237,N_1601);
xnor U2939 (N_2939,N_1645,N_614);
and U2940 (N_2940,N_1527,N_219);
nand U2941 (N_2941,N_1339,N_740);
xor U2942 (N_2942,N_641,N_517);
xor U2943 (N_2943,N_1085,N_252);
nor U2944 (N_2944,N_1805,N_1758);
or U2945 (N_2945,N_2265,N_2330);
and U2946 (N_2946,N_736,N_2240);
and U2947 (N_2947,N_303,N_1531);
and U2948 (N_2948,N_1923,N_2030);
or U2949 (N_2949,N_454,N_1322);
or U2950 (N_2950,N_1143,N_1025);
xnor U2951 (N_2951,N_896,N_72);
nor U2952 (N_2952,N_1629,N_1544);
xor U2953 (N_2953,N_775,N_1699);
nand U2954 (N_2954,N_665,N_1516);
xnor U2955 (N_2955,N_2277,N_2475);
or U2956 (N_2956,N_1176,N_327);
nand U2957 (N_2957,N_17,N_1818);
nor U2958 (N_2958,N_1609,N_543);
and U2959 (N_2959,N_2438,N_2407);
and U2960 (N_2960,N_2267,N_2296);
and U2961 (N_2961,N_2153,N_1825);
or U2962 (N_2962,N_1650,N_2124);
nand U2963 (N_2963,N_86,N_661);
and U2964 (N_2964,N_2053,N_811);
nand U2965 (N_2965,N_317,N_341);
or U2966 (N_2966,N_1750,N_487);
and U2967 (N_2967,N_1888,N_1815);
and U2968 (N_2968,N_780,N_203);
nand U2969 (N_2969,N_2289,N_1679);
and U2970 (N_2970,N_506,N_1705);
nand U2971 (N_2971,N_321,N_1657);
or U2972 (N_2972,N_467,N_720);
or U2973 (N_2973,N_675,N_1740);
and U2974 (N_2974,N_1491,N_2223);
nor U2975 (N_2975,N_352,N_1417);
nor U2976 (N_2976,N_2001,N_179);
xor U2977 (N_2977,N_2455,N_2169);
and U2978 (N_2978,N_214,N_579);
xnor U2979 (N_2979,N_381,N_442);
nand U2980 (N_2980,N_1383,N_1523);
xnor U2981 (N_2981,N_1029,N_501);
or U2982 (N_2982,N_823,N_404);
nor U2983 (N_2983,N_2136,N_2351);
xor U2984 (N_2984,N_1918,N_2067);
and U2985 (N_2985,N_2283,N_1008);
and U2986 (N_2986,N_1374,N_236);
nor U2987 (N_2987,N_1974,N_1685);
nor U2988 (N_2988,N_1714,N_1767);
and U2989 (N_2989,N_284,N_2225);
nor U2990 (N_2990,N_1048,N_825);
nor U2991 (N_2991,N_1350,N_2382);
nand U2992 (N_2992,N_1026,N_1416);
xnor U2993 (N_2993,N_1980,N_346);
xor U2994 (N_2994,N_853,N_814);
nor U2995 (N_2995,N_149,N_261);
and U2996 (N_2996,N_943,N_874);
xnor U2997 (N_2997,N_148,N_1332);
nor U2998 (N_2998,N_5,N_2107);
nor U2999 (N_2999,N_876,N_2065);
nor U3000 (N_3000,N_891,N_2109);
or U3001 (N_3001,N_1497,N_1716);
nor U3002 (N_3002,N_1199,N_2255);
or U3003 (N_3003,N_1958,N_1747);
or U3004 (N_3004,N_2327,N_1137);
and U3005 (N_3005,N_1534,N_813);
and U3006 (N_3006,N_2106,N_11);
nand U3007 (N_3007,N_737,N_882);
nor U3008 (N_3008,N_803,N_767);
nor U3009 (N_3009,N_771,N_1498);
nand U3010 (N_3010,N_407,N_2319);
nand U3011 (N_3011,N_1182,N_2143);
nor U3012 (N_3012,N_2473,N_264);
nand U3013 (N_3013,N_1953,N_999);
nand U3014 (N_3014,N_2028,N_2376);
nor U3015 (N_3015,N_938,N_2195);
nand U3016 (N_3016,N_1439,N_447);
xnor U3017 (N_3017,N_238,N_1717);
xnor U3018 (N_3018,N_598,N_1504);
or U3019 (N_3019,N_2336,N_1357);
nor U3020 (N_3020,N_496,N_1925);
or U3021 (N_3021,N_1220,N_2116);
and U3022 (N_3022,N_1037,N_1047);
and U3023 (N_3023,N_793,N_1267);
and U3024 (N_3024,N_672,N_1518);
xor U3025 (N_3025,N_734,N_257);
and U3026 (N_3026,N_109,N_82);
xnor U3027 (N_3027,N_884,N_942);
nor U3028 (N_3028,N_2088,N_2383);
and U3029 (N_3029,N_575,N_1628);
xnor U3030 (N_3030,N_777,N_1108);
nor U3031 (N_3031,N_2428,N_820);
and U3032 (N_3032,N_1748,N_1370);
and U3033 (N_3033,N_355,N_1935);
xnor U3034 (N_3034,N_1119,N_1445);
xnor U3035 (N_3035,N_2043,N_92);
and U3036 (N_3036,N_2386,N_2480);
nand U3037 (N_3037,N_290,N_1050);
or U3038 (N_3038,N_1263,N_2253);
or U3039 (N_3039,N_634,N_692);
xnor U3040 (N_3040,N_1987,N_1429);
and U3041 (N_3041,N_1535,N_36);
xor U3042 (N_3042,N_904,N_761);
nand U3043 (N_3043,N_1643,N_2141);
xnor U3044 (N_3044,N_2244,N_2364);
nand U3045 (N_3045,N_247,N_1636);
and U3046 (N_3046,N_46,N_1582);
nor U3047 (N_3047,N_226,N_320);
nand U3048 (N_3048,N_1817,N_1409);
and U3049 (N_3049,N_965,N_633);
or U3050 (N_3050,N_1337,N_1438);
nand U3051 (N_3051,N_1473,N_895);
and U3052 (N_3052,N_587,N_361);
nand U3053 (N_3053,N_1222,N_722);
xnor U3054 (N_3054,N_781,N_1434);
nand U3055 (N_3055,N_1816,N_2298);
nand U3056 (N_3056,N_686,N_2040);
nor U3057 (N_3057,N_879,N_1891);
nand U3058 (N_3058,N_1677,N_1842);
xor U3059 (N_3059,N_952,N_815);
nand U3060 (N_3060,N_2085,N_1967);
nor U3061 (N_3061,N_899,N_905);
nand U3062 (N_3062,N_1955,N_2497);
nor U3063 (N_3063,N_2409,N_1885);
nand U3064 (N_3064,N_1457,N_1068);
or U3065 (N_3065,N_1945,N_1286);
and U3066 (N_3066,N_2024,N_419);
nand U3067 (N_3067,N_513,N_939);
or U3068 (N_3068,N_804,N_2051);
xnor U3069 (N_3069,N_2355,N_816);
xor U3070 (N_3070,N_2403,N_2044);
xor U3071 (N_3071,N_738,N_2290);
nor U3072 (N_3072,N_1841,N_768);
xnor U3073 (N_3073,N_1803,N_1993);
nor U3074 (N_3074,N_1800,N_1145);
nor U3075 (N_3075,N_136,N_1036);
nor U3076 (N_3076,N_137,N_40);
or U3077 (N_3077,N_1334,N_1533);
nor U3078 (N_3078,N_1205,N_1882);
and U3079 (N_3079,N_2390,N_2176);
xor U3080 (N_3080,N_1433,N_207);
nor U3081 (N_3081,N_267,N_1288);
xnor U3082 (N_3082,N_2470,N_1860);
nor U3083 (N_3083,N_1466,N_2117);
xor U3084 (N_3084,N_1415,N_2221);
xnor U3085 (N_3085,N_2032,N_1465);
and U3086 (N_3086,N_2127,N_728);
nand U3087 (N_3087,N_1956,N_1479);
nand U3088 (N_3088,N_1014,N_2262);
and U3089 (N_3089,N_237,N_1254);
nand U3090 (N_3090,N_1142,N_1349);
nor U3091 (N_3091,N_1934,N_528);
and U3092 (N_3092,N_1715,N_2350);
nor U3093 (N_3093,N_129,N_491);
or U3094 (N_3094,N_244,N_1690);
or U3095 (N_3095,N_1669,N_1313);
nor U3096 (N_3096,N_1123,N_1653);
and U3097 (N_3097,N_1414,N_2077);
xnor U3098 (N_3098,N_1446,N_1316);
or U3099 (N_3099,N_1124,N_960);
nand U3100 (N_3100,N_2249,N_2010);
and U3101 (N_3101,N_1069,N_1621);
nor U3102 (N_3102,N_723,N_22);
nand U3103 (N_3103,N_2105,N_1730);
or U3104 (N_3104,N_453,N_2395);
nand U3105 (N_3105,N_2495,N_1807);
xnor U3106 (N_3106,N_2346,N_982);
nor U3107 (N_3107,N_2341,N_1030);
nor U3108 (N_3108,N_941,N_1088);
nor U3109 (N_3109,N_877,N_2191);
and U3110 (N_3110,N_1371,N_2137);
nand U3111 (N_3111,N_2008,N_778);
and U3112 (N_3112,N_2279,N_128);
xor U3113 (N_3113,N_693,N_1588);
or U3114 (N_3114,N_2391,N_208);
nor U3115 (N_3115,N_1111,N_924);
nor U3116 (N_3116,N_485,N_307);
nand U3117 (N_3117,N_997,N_1775);
and U3118 (N_3118,N_855,N_1213);
nor U3119 (N_3119,N_967,N_2422);
or U3120 (N_3120,N_1107,N_2046);
nand U3121 (N_3121,N_2326,N_2231);
xnor U3122 (N_3122,N_1514,N_1340);
or U3123 (N_3123,N_1997,N_1179);
xor U3124 (N_3124,N_1474,N_1319);
and U3125 (N_3125,N_1878,N_1698);
or U3126 (N_3126,N_989,N_463);
and U3127 (N_3127,N_502,N_2083);
xnor U3128 (N_3128,N_1109,N_1559);
nand U3129 (N_3129,N_607,N_1365);
nor U3130 (N_3130,N_980,N_1072);
nand U3131 (N_3131,N_2215,N_1726);
and U3132 (N_3132,N_818,N_2303);
or U3133 (N_3133,N_312,N_413);
and U3134 (N_3134,N_386,N_2324);
nand U3135 (N_3135,N_1863,N_1665);
xor U3136 (N_3136,N_2185,N_1948);
nor U3137 (N_3137,N_1991,N_1364);
nand U3138 (N_3138,N_1408,N_836);
or U3139 (N_3139,N_2229,N_724);
nand U3140 (N_3140,N_2139,N_623);
xnor U3141 (N_3141,N_856,N_250);
xnor U3142 (N_3142,N_429,N_2314);
nand U3143 (N_3143,N_1067,N_54);
and U3144 (N_3144,N_139,N_1584);
nand U3145 (N_3145,N_401,N_1259);
or U3146 (N_3146,N_2200,N_2197);
or U3147 (N_3147,N_281,N_1710);
nor U3148 (N_3148,N_837,N_1366);
nor U3149 (N_3149,N_2414,N_1262);
nor U3150 (N_3150,N_1603,N_1396);
or U3151 (N_3151,N_1225,N_1292);
nor U3152 (N_3152,N_363,N_140);
and U3153 (N_3153,N_2457,N_1680);
xnor U3154 (N_3154,N_1973,N_1550);
nor U3155 (N_3155,N_786,N_1933);
or U3156 (N_3156,N_1481,N_2367);
and U3157 (N_3157,N_1074,N_1625);
or U3158 (N_3158,N_152,N_1507);
nand U3159 (N_3159,N_406,N_2415);
nor U3160 (N_3160,N_2216,N_80);
nor U3161 (N_3161,N_2274,N_490);
nand U3162 (N_3162,N_2128,N_657);
and U3163 (N_3163,N_2130,N_878);
xnor U3164 (N_3164,N_849,N_629);
xor U3165 (N_3165,N_540,N_438);
xnor U3166 (N_3166,N_133,N_2115);
and U3167 (N_3167,N_529,N_519);
and U3168 (N_3168,N_1382,N_1661);
and U3169 (N_3169,N_851,N_1281);
or U3170 (N_3170,N_651,N_1375);
nand U3171 (N_3171,N_116,N_1734);
xor U3172 (N_3172,N_1084,N_1553);
xor U3173 (N_3173,N_2172,N_846);
nor U3174 (N_3174,N_437,N_2190);
nor U3175 (N_3175,N_1149,N_1792);
and U3176 (N_3176,N_1941,N_21);
nor U3177 (N_3177,N_966,N_1162);
nor U3178 (N_3178,N_759,N_1023);
nor U3179 (N_3179,N_1475,N_1090);
or U3180 (N_3180,N_2209,N_1083);
nand U3181 (N_3181,N_2241,N_970);
or U3182 (N_3182,N_2189,N_628);
nor U3183 (N_3183,N_1065,N_1355);
or U3184 (N_3184,N_2426,N_2212);
and U3185 (N_3185,N_1564,N_169);
or U3186 (N_3186,N_1420,N_2039);
xnor U3187 (N_3187,N_254,N_1082);
nand U3188 (N_3188,N_1791,N_916);
nor U3189 (N_3189,N_1402,N_769);
and U3190 (N_3190,N_534,N_1770);
and U3191 (N_3191,N_1105,N_1443);
xnor U3192 (N_3192,N_739,N_1602);
nand U3193 (N_3193,N_138,N_1771);
or U3194 (N_3194,N_1278,N_325);
nor U3195 (N_3195,N_520,N_843);
and U3196 (N_3196,N_1513,N_1558);
xor U3197 (N_3197,N_921,N_234);
nor U3198 (N_3198,N_949,N_1883);
or U3199 (N_3199,N_1156,N_831);
nor U3200 (N_3200,N_416,N_2492);
nand U3201 (N_3201,N_31,N_258);
or U3202 (N_3202,N_2150,N_2278);
and U3203 (N_3203,N_2252,N_1356);
or U3204 (N_3204,N_1793,N_524);
and U3205 (N_3205,N_1043,N_2301);
xor U3206 (N_3206,N_2486,N_1314);
xor U3207 (N_3207,N_2434,N_559);
or U3208 (N_3208,N_533,N_2078);
xor U3209 (N_3209,N_794,N_1512);
nand U3210 (N_3210,N_27,N_542);
nor U3211 (N_3211,N_1682,N_2211);
and U3212 (N_3212,N_87,N_2140);
nand U3213 (N_3213,N_1360,N_2429);
nand U3214 (N_3214,N_306,N_2146);
nor U3215 (N_3215,N_2183,N_1147);
xor U3216 (N_3216,N_1284,N_2445);
xnor U3217 (N_3217,N_1960,N_1739);
nand U3218 (N_3218,N_649,N_52);
nor U3219 (N_3219,N_590,N_947);
nand U3220 (N_3220,N_1175,N_2311);
and U3221 (N_3221,N_2084,N_263);
or U3222 (N_3222,N_1345,N_1203);
nor U3223 (N_3223,N_558,N_94);
nor U3224 (N_3224,N_2242,N_37);
nor U3225 (N_3225,N_2131,N_53);
nor U3226 (N_3226,N_2297,N_41);
nor U3227 (N_3227,N_1737,N_2173);
xor U3228 (N_3228,N_512,N_372);
nand U3229 (N_3229,N_578,N_972);
nand U3230 (N_3230,N_1155,N_2054);
or U3231 (N_3231,N_995,N_604);
or U3232 (N_3232,N_1985,N_1937);
nor U3233 (N_3233,N_198,N_1610);
nand U3234 (N_3234,N_1359,N_2031);
nor U3235 (N_3235,N_2477,N_1996);
nand U3236 (N_3236,N_2045,N_996);
xor U3237 (N_3237,N_2254,N_2441);
and U3238 (N_3238,N_2232,N_340);
nor U3239 (N_3239,N_1486,N_461);
nor U3240 (N_3240,N_391,N_1865);
nor U3241 (N_3241,N_2440,N_2481);
xnor U3242 (N_3242,N_582,N_687);
nor U3243 (N_3243,N_760,N_1151);
and U3244 (N_3244,N_2293,N_2379);
and U3245 (N_3245,N_805,N_621);
nand U3246 (N_3246,N_1394,N_159);
nand U3247 (N_3247,N_1477,N_286);
nand U3248 (N_3248,N_2003,N_695);
xor U3249 (N_3249,N_1159,N_1776);
or U3250 (N_3250,N_2213,N_862);
nor U3251 (N_3251,N_328,N_787);
and U3252 (N_3252,N_703,N_806);
and U3253 (N_3253,N_2342,N_522);
xnor U3254 (N_3254,N_2306,N_96);
or U3255 (N_3255,N_1598,N_1969);
or U3256 (N_3256,N_1859,N_897);
nand U3257 (N_3257,N_573,N_2082);
nor U3258 (N_3258,N_1127,N_511);
and U3259 (N_3259,N_626,N_705);
nor U3260 (N_3260,N_2264,N_1012);
and U3261 (N_3261,N_646,N_1820);
nor U3262 (N_3262,N_365,N_2482);
and U3263 (N_3263,N_2074,N_29);
nand U3264 (N_3264,N_1542,N_2062);
or U3265 (N_3265,N_1833,N_492);
nand U3266 (N_3266,N_1502,N_713);
xor U3267 (N_3267,N_704,N_569);
or U3268 (N_3268,N_2347,N_1478);
xor U3269 (N_3269,N_1393,N_2406);
and U3270 (N_3270,N_2059,N_1397);
and U3271 (N_3271,N_864,N_1999);
or U3272 (N_3272,N_1615,N_2411);
nor U3273 (N_3273,N_1169,N_1936);
nor U3274 (N_3274,N_2025,N_652);
and U3275 (N_3275,N_699,N_631);
nand U3276 (N_3276,N_1388,N_1273);
or U3277 (N_3277,N_1988,N_314);
or U3278 (N_3278,N_1595,N_428);
and U3279 (N_3279,N_1908,N_1362);
or U3280 (N_3280,N_1922,N_839);
nor U3281 (N_3281,N_1722,N_1656);
xor U3282 (N_3282,N_209,N_212);
xor U3283 (N_3283,N_576,N_202);
xor U3284 (N_3284,N_1635,N_2142);
nor U3285 (N_3285,N_2236,N_1632);
nand U3286 (N_3286,N_376,N_2217);
xor U3287 (N_3287,N_1271,N_834);
or U3288 (N_3288,N_2282,N_123);
xor U3289 (N_3289,N_2219,N_680);
and U3290 (N_3290,N_2443,N_1709);
nor U3291 (N_3291,N_2338,N_468);
or U3292 (N_3292,N_1236,N_67);
xor U3293 (N_3293,N_278,N_1171);
and U3294 (N_3294,N_1662,N_1902);
nand U3295 (N_3295,N_1765,N_906);
and U3296 (N_3296,N_1279,N_1431);
and U3297 (N_3297,N_2466,N_472);
nor U3298 (N_3298,N_57,N_1696);
nor U3299 (N_3299,N_901,N_2399);
nor U3300 (N_3300,N_1449,N_2340);
nor U3301 (N_3301,N_1522,N_1400);
nor U3302 (N_3302,N_1042,N_1454);
nand U3303 (N_3303,N_1276,N_1495);
nand U3304 (N_3304,N_172,N_229);
or U3305 (N_3305,N_131,N_1460);
and U3306 (N_3306,N_1379,N_451);
or U3307 (N_3307,N_2055,N_1687);
nand U3308 (N_3308,N_1333,N_1407);
nand U3309 (N_3309,N_1039,N_1134);
xor U3310 (N_3310,N_1232,N_1501);
nor U3311 (N_3311,N_1121,N_1311);
nor U3312 (N_3312,N_76,N_903);
nor U3313 (N_3313,N_2154,N_1909);
and U3314 (N_3314,N_922,N_2388);
nand U3315 (N_3315,N_867,N_640);
xnor U3316 (N_3316,N_1190,N_18);
nand U3317 (N_3317,N_1845,N_125);
nand U3318 (N_3318,N_616,N_795);
nor U3319 (N_3319,N_1246,N_694);
or U3320 (N_3320,N_1258,N_845);
nand U3321 (N_3321,N_414,N_547);
nor U3322 (N_3322,N_498,N_1193);
xnor U3323 (N_3323,N_269,N_1);
nor U3324 (N_3324,N_1410,N_2461);
xor U3325 (N_3325,N_1209,N_2356);
or U3326 (N_3326,N_25,N_842);
nand U3327 (N_3327,N_888,N_1309);
xnor U3328 (N_3328,N_963,N_1095);
nand U3329 (N_3329,N_1720,N_2167);
or U3330 (N_3330,N_2089,N_1468);
xnor U3331 (N_3331,N_2450,N_1243);
or U3332 (N_3332,N_157,N_330);
xor U3333 (N_3333,N_504,N_417);
and U3334 (N_3334,N_1847,N_1327);
xnor U3335 (N_3335,N_677,N_1372);
or U3336 (N_3336,N_1098,N_893);
nand U3337 (N_3337,N_525,N_2023);
xor U3338 (N_3338,N_1978,N_411);
or U3339 (N_3339,N_488,N_243);
nand U3340 (N_3340,N_1998,N_622);
or U3341 (N_3341,N_2467,N_2070);
or U3342 (N_3342,N_2437,N_4);
or U3343 (N_3343,N_1295,N_230);
nor U3344 (N_3344,N_251,N_698);
nor U3345 (N_3345,N_65,N_1195);
or U3346 (N_3346,N_682,N_2397);
and U3347 (N_3347,N_1144,N_83);
nor U3348 (N_3348,N_870,N_1555);
xnor U3349 (N_3349,N_1659,N_296);
nand U3350 (N_3350,N_49,N_1055);
nor U3351 (N_3351,N_1444,N_2418);
or U3352 (N_3352,N_807,N_424);
nor U3353 (N_3353,N_1413,N_1458);
xnor U3354 (N_3354,N_953,N_2372);
nor U3355 (N_3355,N_926,N_635);
xor U3356 (N_3356,N_1347,N_2208);
or U3357 (N_3357,N_459,N_1576);
nor U3358 (N_3358,N_2164,N_1893);
or U3359 (N_3359,N_249,N_2432);
xor U3360 (N_3360,N_402,N_1437);
xor U3361 (N_3361,N_1681,N_256);
or U3362 (N_3362,N_1320,N_973);
and U3363 (N_3363,N_1282,N_329);
nor U3364 (N_3364,N_526,N_934);
nor U3365 (N_3365,N_347,N_911);
xor U3366 (N_3366,N_2439,N_2435);
and U3367 (N_3367,N_89,N_1571);
xnor U3368 (N_3368,N_1247,N_190);
or U3369 (N_3369,N_24,N_415);
nor U3370 (N_3370,N_2419,N_1154);
and U3371 (N_3371,N_1683,N_1856);
or U3372 (N_3372,N_1802,N_859);
or U3373 (N_3373,N_1622,N_84);
and U3374 (N_3374,N_240,N_1214);
xnor U3375 (N_3375,N_1867,N_1745);
nor U3376 (N_3376,N_1024,N_923);
xor U3377 (N_3377,N_2239,N_580);
nor U3378 (N_3378,N_663,N_2182);
or U3379 (N_3379,N_178,N_1331);
and U3380 (N_3380,N_400,N_1208);
or U3381 (N_3381,N_2462,N_2405);
nor U3382 (N_3382,N_205,N_1076);
xor U3383 (N_3383,N_991,N_1306);
and U3384 (N_3384,N_861,N_375);
xnor U3385 (N_3385,N_2490,N_464);
xor U3386 (N_3386,N_2038,N_1569);
nor U3387 (N_3387,N_1753,N_446);
or U3388 (N_3388,N_1759,N_751);
and U3389 (N_3389,N_192,N_1385);
and U3390 (N_3390,N_951,N_1666);
or U3391 (N_3391,N_142,N_2321);
xor U3392 (N_3392,N_546,N_288);
nor U3393 (N_3393,N_577,N_1253);
nand U3394 (N_3394,N_1778,N_763);
xor U3395 (N_3395,N_6,N_824);
and U3396 (N_3396,N_2036,N_273);
and U3397 (N_3397,N_1315,N_779);
nand U3398 (N_3398,N_681,N_1992);
nand U3399 (N_3399,N_480,N_1260);
nand U3400 (N_3400,N_2258,N_2374);
nor U3401 (N_3401,N_1932,N_749);
xnor U3402 (N_3402,N_1708,N_718);
or U3403 (N_3403,N_2058,N_561);
xor U3404 (N_3404,N_1963,N_2359);
xor U3405 (N_3405,N_141,N_1638);
xor U3406 (N_3406,N_2063,N_1975);
nand U3407 (N_3407,N_1184,N_1428);
xor U3408 (N_3408,N_1911,N_1442);
or U3409 (N_3409,N_2331,N_1419);
and U3410 (N_3410,N_2479,N_1897);
nand U3411 (N_3411,N_12,N_1490);
nor U3412 (N_3412,N_349,N_1485);
nand U3413 (N_3413,N_1735,N_753);
nand U3414 (N_3414,N_1938,N_1133);
nand U3415 (N_3415,N_189,N_1060);
nor U3416 (N_3416,N_1463,N_550);
and U3417 (N_3417,N_1299,N_1138);
or U3418 (N_3418,N_1684,N_1110);
nand U3419 (N_3419,N_1093,N_396);
and U3420 (N_3420,N_2402,N_1075);
or U3421 (N_3421,N_2166,N_1492);
xnor U3422 (N_3422,N_1873,N_2034);
nand U3423 (N_3423,N_1427,N_514);
nor U3424 (N_3424,N_2111,N_2389);
and U3425 (N_3425,N_2323,N_483);
nand U3426 (N_3426,N_2352,N_176);
or U3427 (N_3427,N_2148,N_1139);
and U3428 (N_3428,N_1011,N_1189);
nor U3429 (N_3429,N_239,N_530);
or U3430 (N_3430,N_2052,N_1017);
or U3431 (N_3431,N_2071,N_883);
nand U3432 (N_3432,N_976,N_2159);
and U3433 (N_3433,N_2087,N_2396);
xor U3434 (N_3434,N_700,N_1116);
nand U3435 (N_3435,N_56,N_567);
nor U3436 (N_3436,N_2446,N_2371);
and U3437 (N_3437,N_928,N_1849);
nand U3438 (N_3438,N_2447,N_2385);
nor U3439 (N_3439,N_1274,N_800);
xnor U3440 (N_3440,N_2226,N_2471);
nand U3441 (N_3441,N_1087,N_206);
xnor U3442 (N_3442,N_1487,N_1574);
or U3443 (N_3443,N_2266,N_568);
nand U3444 (N_3444,N_563,N_194);
xor U3445 (N_3445,N_1212,N_2318);
nor U3446 (N_3446,N_310,N_155);
and U3447 (N_3447,N_1081,N_2247);
and U3448 (N_3448,N_1218,N_100);
nand U3449 (N_3449,N_866,N_1674);
or U3450 (N_3450,N_1010,N_564);
xor U3451 (N_3451,N_676,N_1244);
and U3452 (N_3452,N_399,N_1972);
xnor U3453 (N_3453,N_548,N_1405);
nor U3454 (N_3454,N_531,N_784);
nand U3455 (N_3455,N_1027,N_1986);
xor U3456 (N_3456,N_589,N_2002);
xnor U3457 (N_3457,N_113,N_731);
and U3458 (N_3458,N_2035,N_1898);
nand U3459 (N_3459,N_871,N_1976);
xor U3460 (N_3460,N_527,N_638);
nand U3461 (N_3461,N_1580,N_1668);
nand U3462 (N_3462,N_20,N_475);
nor U3463 (N_3463,N_2312,N_379);
xor U3464 (N_3464,N_1804,N_2068);
or U3465 (N_3465,N_1572,N_1071);
and U3466 (N_3466,N_1644,N_1456);
xnor U3467 (N_3467,N_440,N_2135);
nor U3468 (N_3468,N_301,N_1707);
and U3469 (N_3469,N_403,N_927);
or U3470 (N_3470,N_395,N_1968);
or U3471 (N_3471,N_389,N_1874);
and U3472 (N_3472,N_1756,N_1000);
xor U3473 (N_3473,N_1545,N_688);
nor U3474 (N_3474,N_2186,N_2384);
nand U3475 (N_3475,N_1611,N_597);
xor U3476 (N_3476,N_1961,N_332);
nor U3477 (N_3477,N_343,N_1180);
xor U3478 (N_3478,N_130,N_1132);
and U3479 (N_3479,N_1575,N_1562);
or U3480 (N_3480,N_1354,N_1369);
nor U3481 (N_3481,N_183,N_441);
and U3482 (N_3482,N_408,N_2424);
or U3483 (N_3483,N_1700,N_647);
and U3484 (N_3484,N_1813,N_1563);
xor U3485 (N_3485,N_1692,N_1649);
and U3486 (N_3486,N_1298,N_1166);
and U3487 (N_3487,N_2029,N_1153);
nor U3488 (N_3488,N_1240,N_886);
nor U3489 (N_3489,N_1044,N_184);
and U3490 (N_3490,N_246,N_2474);
xnor U3491 (N_3491,N_1022,N_187);
xor U3492 (N_3492,N_2049,N_1219);
or U3493 (N_3493,N_1829,N_2369);
or U3494 (N_3494,N_1795,N_2170);
nor U3495 (N_3495,N_2300,N_844);
and U3496 (N_3496,N_2280,N_2091);
nor U3497 (N_3497,N_710,N_544);
nor U3498 (N_3498,N_1733,N_2114);
and U3499 (N_3499,N_1876,N_1392);
xor U3500 (N_3500,N_2214,N_1380);
nor U3501 (N_3501,N_1624,N_1198);
xnor U3502 (N_3502,N_1784,N_452);
and U3503 (N_3503,N_479,N_335);
xor U3504 (N_3504,N_505,N_2145);
and U3505 (N_3505,N_925,N_2000);
xor U3506 (N_3506,N_95,N_2138);
nor U3507 (N_3507,N_1237,N_742);
nor U3508 (N_3508,N_1070,N_2288);
xor U3509 (N_3509,N_2423,N_174);
and U3510 (N_3510,N_1257,N_166);
xnor U3511 (N_3511,N_1943,N_353);
and U3512 (N_3512,N_227,N_881);
or U3513 (N_3513,N_539,N_955);
nand U3514 (N_3514,N_1381,N_2033);
nand U3515 (N_3515,N_345,N_50);
nand U3516 (N_3516,N_1861,N_2090);
xor U3517 (N_3517,N_405,N_1028);
and U3518 (N_3518,N_2394,N_371);
nor U3519 (N_3519,N_915,N_1530);
and U3520 (N_3520,N_2358,N_173);
or U3521 (N_3521,N_1926,N_659);
or U3522 (N_3522,N_732,N_484);
or U3523 (N_3523,N_2121,N_944);
and U3524 (N_3524,N_1560,N_1664);
xnor U3525 (N_3525,N_774,N_716);
or U3526 (N_3526,N_144,N_1034);
xnor U3527 (N_3527,N_2072,N_664);
nor U3528 (N_3528,N_2155,N_2436);
nand U3529 (N_3529,N_1476,N_602);
nand U3530 (N_3530,N_2007,N_1913);
nor U3531 (N_3531,N_2496,N_1819);
xor U3532 (N_3532,N_367,N_458);
nor U3533 (N_3533,N_2108,N_1573);
nand U3534 (N_3534,N_518,N_387);
nor U3535 (N_3535,N_1061,N_637);
and U3536 (N_3536,N_2464,N_124);
nor U3537 (N_3537,N_354,N_706);
nand U3538 (N_3538,N_2019,N_111);
or U3539 (N_3539,N_935,N_946);
nand U3540 (N_3540,N_1599,N_645);
and U3541 (N_3541,N_1706,N_2459);
and U3542 (N_3542,N_832,N_1128);
or U3543 (N_3543,N_1425,N_383);
xor U3544 (N_3544,N_1704,N_674);
or U3545 (N_3545,N_988,N_1270);
or U3546 (N_3546,N_270,N_1762);
and U3547 (N_3547,N_2093,N_608);
and U3548 (N_3548,N_1256,N_1183);
nand U3549 (N_3549,N_1440,N_748);
or U3550 (N_3550,N_1851,N_615);
nor U3551 (N_3551,N_872,N_643);
or U3552 (N_3552,N_1727,N_696);
nor U3553 (N_3553,N_1721,N_1613);
and U3554 (N_3554,N_2292,N_1631);
and U3555 (N_3555,N_1982,N_1713);
xor U3556 (N_3556,N_662,N_2224);
nand U3557 (N_3557,N_572,N_1464);
nand U3558 (N_3558,N_112,N_1101);
nand U3559 (N_3559,N_1701,N_1917);
xor U3560 (N_3560,N_940,N_1500);
nand U3561 (N_3561,N_1150,N_1676);
nor U3562 (N_3562,N_660,N_2309);
and U3563 (N_3563,N_1426,N_1307);
and U3564 (N_3564,N_265,N_326);
and U3565 (N_3565,N_1597,N_2412);
nor U3566 (N_3566,N_108,N_1904);
xnor U3567 (N_3567,N_1981,N_271);
and U3568 (N_3568,N_1403,N_182);
xor U3569 (N_3569,N_1268,N_295);
nand U3570 (N_3570,N_1187,N_357);
nor U3571 (N_3571,N_557,N_223);
nand U3572 (N_3572,N_1587,N_2201);
and U3573 (N_3573,N_2047,N_1216);
or U3574 (N_3574,N_2092,N_1077);
nor U3575 (N_3575,N_950,N_1326);
or U3576 (N_3576,N_471,N_2);
and U3577 (N_3577,N_1693,N_1376);
xnor U3578 (N_3578,N_2268,N_348);
or U3579 (N_3579,N_1245,N_1063);
nor U3580 (N_3580,N_1324,N_1581);
xnor U3581 (N_3581,N_2458,N_708);
and U3582 (N_3582,N_431,N_2069);
nand U3583 (N_3583,N_195,N_305);
xnor U3584 (N_3584,N_691,N_64);
nor U3585 (N_3585,N_422,N_359);
and U3586 (N_3586,N_898,N_714);
or U3587 (N_3587,N_1525,N_1432);
or U3588 (N_3588,N_61,N_2101);
nor U3589 (N_3589,N_75,N_2276);
xor U3590 (N_3590,N_1031,N_974);
nand U3591 (N_3591,N_285,N_1448);
nor U3592 (N_3592,N_47,N_1112);
nor U3593 (N_3593,N_1045,N_1348);
or U3594 (N_3594,N_658,N_1249);
xor U3595 (N_3595,N_601,N_773);
and U3596 (N_3596,N_1944,N_801);
nor U3597 (N_3597,N_196,N_1870);
or U3598 (N_3598,N_1341,N_1141);
nand U3599 (N_3599,N_945,N_59);
nor U3600 (N_3600,N_1623,N_1906);
xnor U3601 (N_3601,N_1773,N_210);
nor U3602 (N_3602,N_983,N_2468);
nand U3603 (N_3603,N_9,N_2179);
or U3604 (N_3604,N_854,N_819);
nor U3605 (N_3605,N_2158,N_701);
and U3606 (N_3606,N_2360,N_1191);
and U3607 (N_3607,N_541,N_1367);
and U3608 (N_3608,N_2129,N_221);
xnor U3609 (N_3609,N_1160,N_28);
nand U3610 (N_3610,N_1079,N_1424);
nand U3611 (N_3611,N_1808,N_1787);
nand U3612 (N_3612,N_2218,N_26);
nor U3613 (N_3613,N_979,N_228);
nand U3614 (N_3614,N_2294,N_319);
and U3615 (N_3615,N_588,N_373);
nand U3616 (N_3616,N_71,N_1852);
nor U3617 (N_3617,N_362,N_798);
nor U3618 (N_3618,N_627,N_121);
or U3619 (N_3619,N_757,N_1235);
or U3620 (N_3620,N_2021,N_1515);
or U3621 (N_3621,N_2348,N_1480);
nor U3622 (N_3622,N_382,N_1760);
nand U3623 (N_3623,N_1242,N_551);
or U3624 (N_3624,N_120,N_1875);
xnor U3625 (N_3625,N_1585,N_553);
nand U3626 (N_3626,N_1667,N_2363);
nand U3627 (N_3627,N_1801,N_1723);
or U3628 (N_3628,N_2444,N_2205);
nand U3629 (N_3629,N_165,N_497);
and U3630 (N_3630,N_1779,N_2099);
and U3631 (N_3631,N_2057,N_2454);
nor U3632 (N_3632,N_1459,N_481);
xnor U3633 (N_3633,N_1003,N_756);
and U3634 (N_3634,N_1532,N_1789);
nor U3635 (N_3635,N_287,N_368);
nor U3636 (N_3636,N_2451,N_1600);
or U3637 (N_3637,N_1238,N_1591);
xor U3638 (N_3638,N_1830,N_337);
xor U3639 (N_3639,N_1764,N_817);
and U3640 (N_3640,N_2151,N_902);
or U3641 (N_3641,N_2161,N_2368);
or U3642 (N_3642,N_2119,N_2354);
nand U3643 (N_3643,N_1763,N_918);
nor U3644 (N_3644,N_1285,N_1794);
and U3645 (N_3645,N_1612,N_2203);
nor U3646 (N_3646,N_1228,N_1634);
and U3647 (N_3647,N_743,N_826);
xnor U3648 (N_3648,N_156,N_1864);
or U3649 (N_3649,N_248,N_2120);
or U3650 (N_3650,N_2398,N_358);
and U3651 (N_3651,N_1252,N_1158);
nor U3652 (N_3652,N_752,N_1032);
and U3653 (N_3653,N_1261,N_1583);
xor U3654 (N_3654,N_670,N_1780);
xor U3655 (N_3655,N_369,N_211);
nand U3656 (N_3656,N_1719,N_2257);
or U3657 (N_3657,N_163,N_1344);
nand U3658 (N_3658,N_2337,N_48);
xnor U3659 (N_3659,N_85,N_1040);
nor U3660 (N_3660,N_565,N_585);
and U3661 (N_3661,N_1172,N_865);
nor U3662 (N_3662,N_2080,N_150);
nand U3663 (N_3663,N_2370,N_858);
xor U3664 (N_3664,N_2499,N_1178);
or U3665 (N_3665,N_1548,N_1016);
nand U3666 (N_3666,N_186,N_2478);
nand U3667 (N_3667,N_2287,N_1914);
and U3668 (N_3668,N_1221,N_1790);
or U3669 (N_3669,N_412,N_1689);
and U3670 (N_3670,N_1441,N_78);
nor U3671 (N_3671,N_1002,N_600);
xor U3672 (N_3672,N_1378,N_1188);
xnor U3673 (N_3673,N_1310,N_2469);
xnor U3674 (N_3674,N_360,N_180);
and U3675 (N_3675,N_765,N_931);
and U3676 (N_3676,N_7,N_450);
and U3677 (N_3677,N_1673,N_1928);
nor U3678 (N_3678,N_1617,N_114);
and U3679 (N_3679,N_1387,N_591);
nand U3680 (N_3680,N_1291,N_1447);
nor U3681 (N_3681,N_1811,N_802);
or U3682 (N_3682,N_1812,N_639);
nor U3683 (N_3683,N_2198,N_489);
or U3684 (N_3684,N_1979,N_1785);
and U3685 (N_3685,N_339,N_201);
nand U3686 (N_3686,N_161,N_959);
or U3687 (N_3687,N_2417,N_1537);
or U3688 (N_3688,N_318,N_887);
xor U3689 (N_3689,N_969,N_2400);
xnor U3690 (N_3690,N_2095,N_650);
or U3691 (N_3691,N_1489,N_1670);
nand U3692 (N_3692,N_1557,N_274);
nand U3693 (N_3693,N_2056,N_666);
and U3694 (N_3694,N_268,N_689);
nor U3695 (N_3695,N_275,N_107);
nand U3696 (N_3696,N_1949,N_315);
nor U3697 (N_3697,N_2377,N_2098);
nor U3698 (N_3698,N_1731,N_2015);
nor U3699 (N_3699,N_2304,N_2275);
nand U3700 (N_3700,N_1484,N_850);
nor U3701 (N_3701,N_1786,N_808);
nor U3702 (N_3702,N_1204,N_2472);
xor U3703 (N_3703,N_758,N_2378);
nand U3704 (N_3704,N_63,N_1697);
xnor U3705 (N_3705,N_1593,N_1336);
or U3706 (N_3706,N_1120,N_147);
nor U3707 (N_3707,N_277,N_2325);
xor U3708 (N_3708,N_2408,N_1094);
or U3709 (N_3709,N_919,N_936);
nand U3710 (N_3710,N_14,N_1335);
nand U3711 (N_3711,N_2152,N_562);
xor U3712 (N_3712,N_2018,N_1493);
or U3713 (N_3713,N_1436,N_746);
nor U3714 (N_3714,N_470,N_2006);
xnor U3715 (N_3715,N_10,N_1482);
nor U3716 (N_3716,N_830,N_2302);
nand U3717 (N_3717,N_350,N_1483);
or U3718 (N_3718,N_1197,N_409);
and U3719 (N_3719,N_2269,N_1957);
nor U3720 (N_3720,N_366,N_2086);
nor U3721 (N_3721,N_2251,N_747);
nand U3722 (N_3722,N_291,N_1293);
and U3723 (N_3723,N_151,N_1741);
or U3724 (N_3724,N_961,N_1266);
or U3725 (N_3725,N_266,N_1227);
or U3726 (N_3726,N_217,N_283);
nor U3727 (N_3727,N_106,N_2410);
or U3728 (N_3728,N_1712,N_160);
nand U3729 (N_3729,N_364,N_1391);
nor U3730 (N_3730,N_2322,N_1342);
xnor U3731 (N_3731,N_829,N_1752);
or U3732 (N_3732,N_2012,N_2133);
nand U3733 (N_3733,N_667,N_900);
and U3734 (N_3734,N_2174,N_2460);
nand U3735 (N_3735,N_342,N_1264);
nor U3736 (N_3736,N_457,N_324);
nor U3737 (N_3737,N_1796,N_304);
or U3738 (N_3738,N_294,N_233);
xor U3739 (N_3739,N_783,N_1272);
or U3740 (N_3740,N_1540,N_13);
xor U3741 (N_3741,N_1947,N_465);
and U3742 (N_3742,N_1894,N_167);
and U3743 (N_3743,N_1736,N_1430);
nand U3744 (N_3744,N_1398,N_719);
nand U3745 (N_3745,N_2272,N_1289);
xnor U3746 (N_3746,N_385,N_1239);
nand U3747 (N_3747,N_1194,N_545);
or U3748 (N_3748,N_334,N_216);
or U3749 (N_3749,N_671,N_2299);
and U3750 (N_3750,N_938,N_1828);
nand U3751 (N_3751,N_1464,N_2080);
nand U3752 (N_3752,N_1064,N_1482);
and U3753 (N_3753,N_1184,N_289);
and U3754 (N_3754,N_498,N_1532);
nand U3755 (N_3755,N_1903,N_1465);
nand U3756 (N_3756,N_1646,N_1048);
nor U3757 (N_3757,N_1252,N_1215);
nand U3758 (N_3758,N_2300,N_600);
xor U3759 (N_3759,N_826,N_2154);
nor U3760 (N_3760,N_886,N_67);
nand U3761 (N_3761,N_895,N_2054);
and U3762 (N_3762,N_1225,N_2261);
xor U3763 (N_3763,N_1480,N_1523);
or U3764 (N_3764,N_1742,N_1115);
and U3765 (N_3765,N_1361,N_1074);
nand U3766 (N_3766,N_2066,N_651);
nand U3767 (N_3767,N_3,N_688);
or U3768 (N_3768,N_1069,N_1013);
xor U3769 (N_3769,N_797,N_808);
and U3770 (N_3770,N_689,N_1103);
xnor U3771 (N_3771,N_1985,N_1039);
xnor U3772 (N_3772,N_1361,N_99);
xnor U3773 (N_3773,N_1931,N_1129);
and U3774 (N_3774,N_1934,N_1682);
or U3775 (N_3775,N_1047,N_1413);
and U3776 (N_3776,N_1372,N_169);
xnor U3777 (N_3777,N_110,N_537);
xor U3778 (N_3778,N_1969,N_2057);
xor U3779 (N_3779,N_1590,N_450);
or U3780 (N_3780,N_2333,N_698);
nor U3781 (N_3781,N_2063,N_439);
xor U3782 (N_3782,N_1672,N_2227);
or U3783 (N_3783,N_1131,N_2254);
and U3784 (N_3784,N_1351,N_1510);
nor U3785 (N_3785,N_1417,N_1684);
or U3786 (N_3786,N_236,N_258);
or U3787 (N_3787,N_2317,N_237);
nand U3788 (N_3788,N_1422,N_1401);
nand U3789 (N_3789,N_1654,N_1292);
nor U3790 (N_3790,N_1458,N_730);
nand U3791 (N_3791,N_2254,N_850);
or U3792 (N_3792,N_1470,N_2219);
and U3793 (N_3793,N_2187,N_898);
nand U3794 (N_3794,N_1580,N_1489);
nand U3795 (N_3795,N_438,N_455);
xnor U3796 (N_3796,N_1640,N_523);
xnor U3797 (N_3797,N_1973,N_2300);
nand U3798 (N_3798,N_538,N_1542);
or U3799 (N_3799,N_1395,N_2423);
nor U3800 (N_3800,N_582,N_2259);
nand U3801 (N_3801,N_697,N_713);
xor U3802 (N_3802,N_616,N_1390);
and U3803 (N_3803,N_683,N_777);
xnor U3804 (N_3804,N_111,N_1100);
xnor U3805 (N_3805,N_1778,N_1360);
and U3806 (N_3806,N_622,N_629);
nand U3807 (N_3807,N_1428,N_2143);
and U3808 (N_3808,N_782,N_1770);
and U3809 (N_3809,N_2386,N_2371);
xnor U3810 (N_3810,N_1584,N_1522);
and U3811 (N_3811,N_936,N_2292);
or U3812 (N_3812,N_2440,N_929);
and U3813 (N_3813,N_1551,N_1153);
xor U3814 (N_3814,N_1387,N_2254);
and U3815 (N_3815,N_21,N_1102);
nand U3816 (N_3816,N_216,N_941);
nor U3817 (N_3817,N_574,N_2234);
xnor U3818 (N_3818,N_1377,N_2070);
xor U3819 (N_3819,N_137,N_1398);
nand U3820 (N_3820,N_1359,N_2047);
nand U3821 (N_3821,N_135,N_1336);
nand U3822 (N_3822,N_1455,N_1203);
and U3823 (N_3823,N_2155,N_2120);
or U3824 (N_3824,N_1288,N_792);
and U3825 (N_3825,N_1306,N_523);
xnor U3826 (N_3826,N_135,N_175);
nand U3827 (N_3827,N_2466,N_992);
xor U3828 (N_3828,N_1341,N_2428);
and U3829 (N_3829,N_450,N_1020);
nor U3830 (N_3830,N_2318,N_615);
or U3831 (N_3831,N_2275,N_1616);
or U3832 (N_3832,N_1607,N_2063);
and U3833 (N_3833,N_2459,N_2181);
nor U3834 (N_3834,N_1418,N_910);
nand U3835 (N_3835,N_553,N_113);
or U3836 (N_3836,N_904,N_1336);
nand U3837 (N_3837,N_765,N_1265);
nor U3838 (N_3838,N_2489,N_1657);
and U3839 (N_3839,N_302,N_904);
nor U3840 (N_3840,N_321,N_2155);
nand U3841 (N_3841,N_1984,N_1737);
xor U3842 (N_3842,N_101,N_553);
or U3843 (N_3843,N_676,N_1568);
nand U3844 (N_3844,N_2276,N_2028);
and U3845 (N_3845,N_2143,N_2371);
nand U3846 (N_3846,N_564,N_124);
or U3847 (N_3847,N_1469,N_756);
xnor U3848 (N_3848,N_801,N_1825);
nor U3849 (N_3849,N_206,N_999);
nand U3850 (N_3850,N_1352,N_689);
and U3851 (N_3851,N_1020,N_2285);
or U3852 (N_3852,N_1477,N_1350);
xnor U3853 (N_3853,N_2313,N_896);
and U3854 (N_3854,N_152,N_592);
nand U3855 (N_3855,N_1707,N_2208);
nand U3856 (N_3856,N_586,N_1718);
xnor U3857 (N_3857,N_839,N_476);
nor U3858 (N_3858,N_1429,N_350);
and U3859 (N_3859,N_1238,N_1392);
and U3860 (N_3860,N_1428,N_2180);
and U3861 (N_3861,N_1894,N_144);
xnor U3862 (N_3862,N_1813,N_1015);
xnor U3863 (N_3863,N_1962,N_744);
and U3864 (N_3864,N_1363,N_785);
or U3865 (N_3865,N_2429,N_824);
xnor U3866 (N_3866,N_2212,N_310);
or U3867 (N_3867,N_2098,N_2402);
or U3868 (N_3868,N_1345,N_2493);
or U3869 (N_3869,N_1829,N_541);
or U3870 (N_3870,N_918,N_1235);
nand U3871 (N_3871,N_260,N_1147);
or U3872 (N_3872,N_1880,N_2210);
nor U3873 (N_3873,N_2093,N_1214);
nor U3874 (N_3874,N_2218,N_439);
nand U3875 (N_3875,N_2179,N_560);
or U3876 (N_3876,N_96,N_2280);
and U3877 (N_3877,N_978,N_2311);
or U3878 (N_3878,N_2059,N_2227);
xnor U3879 (N_3879,N_713,N_603);
nor U3880 (N_3880,N_1474,N_2150);
xnor U3881 (N_3881,N_31,N_2427);
nor U3882 (N_3882,N_2498,N_1993);
nor U3883 (N_3883,N_1859,N_1692);
xnor U3884 (N_3884,N_999,N_1275);
or U3885 (N_3885,N_2227,N_1469);
and U3886 (N_3886,N_495,N_1653);
xor U3887 (N_3887,N_2395,N_2378);
nor U3888 (N_3888,N_120,N_1867);
or U3889 (N_3889,N_464,N_954);
nand U3890 (N_3890,N_1370,N_2098);
or U3891 (N_3891,N_2232,N_1040);
nor U3892 (N_3892,N_1025,N_1906);
and U3893 (N_3893,N_198,N_2076);
nor U3894 (N_3894,N_1445,N_1472);
and U3895 (N_3895,N_932,N_1513);
xnor U3896 (N_3896,N_2160,N_181);
nor U3897 (N_3897,N_962,N_56);
nand U3898 (N_3898,N_412,N_1583);
nor U3899 (N_3899,N_1533,N_805);
or U3900 (N_3900,N_257,N_860);
nor U3901 (N_3901,N_248,N_1578);
or U3902 (N_3902,N_1564,N_2047);
and U3903 (N_3903,N_2397,N_1118);
xnor U3904 (N_3904,N_2238,N_2045);
and U3905 (N_3905,N_2374,N_1679);
and U3906 (N_3906,N_2016,N_636);
xnor U3907 (N_3907,N_616,N_1617);
or U3908 (N_3908,N_2129,N_1591);
xor U3909 (N_3909,N_1846,N_283);
and U3910 (N_3910,N_803,N_162);
nand U3911 (N_3911,N_1360,N_775);
xor U3912 (N_3912,N_1162,N_1651);
and U3913 (N_3913,N_1317,N_575);
or U3914 (N_3914,N_581,N_1323);
and U3915 (N_3915,N_1317,N_819);
and U3916 (N_3916,N_579,N_1117);
nand U3917 (N_3917,N_293,N_2194);
and U3918 (N_3918,N_2188,N_2376);
nor U3919 (N_3919,N_2299,N_1708);
nor U3920 (N_3920,N_103,N_1524);
nor U3921 (N_3921,N_1493,N_1710);
or U3922 (N_3922,N_315,N_831);
and U3923 (N_3923,N_2241,N_1484);
nand U3924 (N_3924,N_1742,N_706);
or U3925 (N_3925,N_1375,N_984);
nor U3926 (N_3926,N_815,N_1269);
nor U3927 (N_3927,N_806,N_365);
xnor U3928 (N_3928,N_1214,N_428);
nand U3929 (N_3929,N_1488,N_2119);
or U3930 (N_3930,N_1990,N_983);
xnor U3931 (N_3931,N_1096,N_1760);
and U3932 (N_3932,N_8,N_1411);
nor U3933 (N_3933,N_1850,N_1591);
or U3934 (N_3934,N_1748,N_2436);
nand U3935 (N_3935,N_2430,N_1663);
and U3936 (N_3936,N_488,N_2211);
nor U3937 (N_3937,N_829,N_1502);
nand U3938 (N_3938,N_1795,N_2487);
nor U3939 (N_3939,N_1244,N_2121);
and U3940 (N_3940,N_678,N_249);
and U3941 (N_3941,N_115,N_1782);
nor U3942 (N_3942,N_1262,N_2210);
nand U3943 (N_3943,N_1347,N_234);
and U3944 (N_3944,N_1911,N_2043);
xnor U3945 (N_3945,N_2462,N_821);
and U3946 (N_3946,N_2325,N_1477);
nand U3947 (N_3947,N_1785,N_668);
nor U3948 (N_3948,N_2376,N_99);
xor U3949 (N_3949,N_1180,N_585);
nand U3950 (N_3950,N_1472,N_1070);
or U3951 (N_3951,N_1367,N_777);
or U3952 (N_3952,N_1229,N_1890);
nor U3953 (N_3953,N_1584,N_1341);
or U3954 (N_3954,N_823,N_243);
or U3955 (N_3955,N_133,N_63);
nor U3956 (N_3956,N_376,N_2424);
nand U3957 (N_3957,N_2464,N_86);
and U3958 (N_3958,N_2158,N_661);
xor U3959 (N_3959,N_368,N_1797);
or U3960 (N_3960,N_1996,N_633);
xnor U3961 (N_3961,N_1741,N_589);
and U3962 (N_3962,N_2280,N_801);
nand U3963 (N_3963,N_925,N_598);
and U3964 (N_3964,N_183,N_1293);
nor U3965 (N_3965,N_2485,N_1987);
nand U3966 (N_3966,N_263,N_1847);
nand U3967 (N_3967,N_86,N_834);
nand U3968 (N_3968,N_2340,N_2288);
xnor U3969 (N_3969,N_1261,N_1391);
xor U3970 (N_3970,N_686,N_1044);
or U3971 (N_3971,N_696,N_785);
nor U3972 (N_3972,N_694,N_211);
and U3973 (N_3973,N_2202,N_2362);
xnor U3974 (N_3974,N_1805,N_476);
nand U3975 (N_3975,N_567,N_1222);
or U3976 (N_3976,N_276,N_287);
nor U3977 (N_3977,N_384,N_1182);
nor U3978 (N_3978,N_1356,N_1282);
or U3979 (N_3979,N_1115,N_2187);
and U3980 (N_3980,N_885,N_115);
nand U3981 (N_3981,N_2262,N_1801);
nor U3982 (N_3982,N_733,N_1381);
nand U3983 (N_3983,N_1331,N_1792);
nor U3984 (N_3984,N_989,N_1384);
nor U3985 (N_3985,N_1035,N_207);
nor U3986 (N_3986,N_1633,N_250);
and U3987 (N_3987,N_501,N_448);
nor U3988 (N_3988,N_1023,N_1340);
or U3989 (N_3989,N_1542,N_1001);
and U3990 (N_3990,N_715,N_1511);
nor U3991 (N_3991,N_650,N_839);
nand U3992 (N_3992,N_882,N_2375);
or U3993 (N_3993,N_911,N_1097);
nand U3994 (N_3994,N_1708,N_256);
xor U3995 (N_3995,N_1191,N_624);
nor U3996 (N_3996,N_777,N_1650);
xor U3997 (N_3997,N_1797,N_580);
xor U3998 (N_3998,N_342,N_634);
or U3999 (N_3999,N_747,N_886);
nor U4000 (N_4000,N_1736,N_1268);
nor U4001 (N_4001,N_2387,N_1439);
and U4002 (N_4002,N_1306,N_1929);
and U4003 (N_4003,N_914,N_1429);
nand U4004 (N_4004,N_2179,N_2088);
xor U4005 (N_4005,N_2131,N_721);
or U4006 (N_4006,N_1677,N_2044);
xnor U4007 (N_4007,N_52,N_1438);
nor U4008 (N_4008,N_1200,N_2055);
or U4009 (N_4009,N_1142,N_2467);
or U4010 (N_4010,N_1871,N_1467);
xnor U4011 (N_4011,N_691,N_1804);
and U4012 (N_4012,N_820,N_181);
nand U4013 (N_4013,N_805,N_269);
xnor U4014 (N_4014,N_1534,N_308);
nand U4015 (N_4015,N_1861,N_1412);
or U4016 (N_4016,N_1496,N_1492);
nand U4017 (N_4017,N_205,N_880);
and U4018 (N_4018,N_1658,N_2460);
nand U4019 (N_4019,N_2491,N_1005);
nor U4020 (N_4020,N_1753,N_363);
nor U4021 (N_4021,N_194,N_1276);
or U4022 (N_4022,N_2293,N_1128);
xnor U4023 (N_4023,N_1818,N_221);
nand U4024 (N_4024,N_556,N_1);
or U4025 (N_4025,N_710,N_913);
xor U4026 (N_4026,N_1828,N_1018);
and U4027 (N_4027,N_1645,N_74);
and U4028 (N_4028,N_189,N_137);
and U4029 (N_4029,N_284,N_1717);
xor U4030 (N_4030,N_549,N_305);
xor U4031 (N_4031,N_23,N_1637);
xnor U4032 (N_4032,N_606,N_160);
nand U4033 (N_4033,N_1880,N_784);
or U4034 (N_4034,N_1161,N_2176);
xnor U4035 (N_4035,N_2055,N_323);
nor U4036 (N_4036,N_1176,N_1256);
or U4037 (N_4037,N_1981,N_481);
or U4038 (N_4038,N_1037,N_1154);
and U4039 (N_4039,N_2000,N_2360);
xnor U4040 (N_4040,N_291,N_2179);
or U4041 (N_4041,N_196,N_2319);
and U4042 (N_4042,N_1501,N_1001);
xor U4043 (N_4043,N_1992,N_2201);
nor U4044 (N_4044,N_439,N_2037);
or U4045 (N_4045,N_1518,N_977);
or U4046 (N_4046,N_959,N_1495);
nor U4047 (N_4047,N_1621,N_2282);
or U4048 (N_4048,N_302,N_1135);
nand U4049 (N_4049,N_1488,N_38);
nand U4050 (N_4050,N_1842,N_1756);
or U4051 (N_4051,N_545,N_1940);
or U4052 (N_4052,N_1757,N_1697);
nand U4053 (N_4053,N_1857,N_650);
nor U4054 (N_4054,N_181,N_1023);
or U4055 (N_4055,N_1638,N_1340);
nor U4056 (N_4056,N_1019,N_840);
nor U4057 (N_4057,N_1650,N_1336);
nor U4058 (N_4058,N_254,N_900);
xnor U4059 (N_4059,N_1682,N_779);
xnor U4060 (N_4060,N_1684,N_788);
and U4061 (N_4061,N_1719,N_314);
and U4062 (N_4062,N_1644,N_612);
nor U4063 (N_4063,N_2162,N_412);
or U4064 (N_4064,N_345,N_865);
nand U4065 (N_4065,N_1652,N_1964);
or U4066 (N_4066,N_53,N_595);
or U4067 (N_4067,N_682,N_1489);
and U4068 (N_4068,N_1910,N_1984);
xnor U4069 (N_4069,N_669,N_525);
nor U4070 (N_4070,N_439,N_442);
or U4071 (N_4071,N_1340,N_1708);
or U4072 (N_4072,N_1214,N_1284);
nor U4073 (N_4073,N_880,N_744);
nor U4074 (N_4074,N_2044,N_555);
and U4075 (N_4075,N_372,N_910);
and U4076 (N_4076,N_548,N_1251);
xnor U4077 (N_4077,N_207,N_580);
nand U4078 (N_4078,N_1638,N_2291);
nand U4079 (N_4079,N_2182,N_1172);
and U4080 (N_4080,N_1564,N_745);
or U4081 (N_4081,N_455,N_2301);
or U4082 (N_4082,N_248,N_1538);
xor U4083 (N_4083,N_353,N_2073);
nand U4084 (N_4084,N_905,N_1050);
or U4085 (N_4085,N_238,N_1844);
or U4086 (N_4086,N_310,N_302);
or U4087 (N_4087,N_459,N_671);
xnor U4088 (N_4088,N_1731,N_795);
nand U4089 (N_4089,N_2260,N_247);
and U4090 (N_4090,N_1621,N_2185);
nor U4091 (N_4091,N_1107,N_1348);
or U4092 (N_4092,N_874,N_778);
nor U4093 (N_4093,N_1724,N_1695);
or U4094 (N_4094,N_1658,N_1908);
or U4095 (N_4095,N_46,N_522);
nand U4096 (N_4096,N_2160,N_1549);
or U4097 (N_4097,N_581,N_0);
and U4098 (N_4098,N_1767,N_490);
nand U4099 (N_4099,N_2489,N_328);
xor U4100 (N_4100,N_488,N_1653);
nand U4101 (N_4101,N_2373,N_850);
xor U4102 (N_4102,N_2180,N_2481);
or U4103 (N_4103,N_2312,N_1192);
nand U4104 (N_4104,N_2133,N_867);
nor U4105 (N_4105,N_1721,N_2472);
and U4106 (N_4106,N_1685,N_1589);
xnor U4107 (N_4107,N_1607,N_446);
nor U4108 (N_4108,N_1475,N_1069);
nor U4109 (N_4109,N_1141,N_758);
or U4110 (N_4110,N_2297,N_764);
xor U4111 (N_4111,N_1970,N_569);
nor U4112 (N_4112,N_149,N_378);
or U4113 (N_4113,N_378,N_272);
nand U4114 (N_4114,N_1278,N_2335);
nand U4115 (N_4115,N_518,N_1685);
xnor U4116 (N_4116,N_873,N_2130);
or U4117 (N_4117,N_820,N_183);
and U4118 (N_4118,N_234,N_2398);
and U4119 (N_4119,N_1353,N_2219);
or U4120 (N_4120,N_2174,N_1770);
xnor U4121 (N_4121,N_1336,N_1714);
or U4122 (N_4122,N_1542,N_327);
or U4123 (N_4123,N_223,N_786);
xor U4124 (N_4124,N_550,N_2321);
and U4125 (N_4125,N_2464,N_174);
xor U4126 (N_4126,N_1688,N_1357);
nand U4127 (N_4127,N_322,N_573);
xnor U4128 (N_4128,N_2219,N_568);
and U4129 (N_4129,N_2123,N_61);
nand U4130 (N_4130,N_1829,N_289);
nand U4131 (N_4131,N_703,N_555);
or U4132 (N_4132,N_1898,N_352);
nor U4133 (N_4133,N_1577,N_2294);
nand U4134 (N_4134,N_2443,N_1549);
xnor U4135 (N_4135,N_2310,N_1726);
nor U4136 (N_4136,N_865,N_804);
nand U4137 (N_4137,N_1509,N_1957);
nor U4138 (N_4138,N_2370,N_1636);
and U4139 (N_4139,N_2183,N_339);
and U4140 (N_4140,N_1961,N_1288);
or U4141 (N_4141,N_1417,N_1780);
and U4142 (N_4142,N_651,N_2129);
or U4143 (N_4143,N_2248,N_64);
and U4144 (N_4144,N_1049,N_1347);
nand U4145 (N_4145,N_1075,N_2403);
xnor U4146 (N_4146,N_1598,N_92);
nor U4147 (N_4147,N_2432,N_1898);
nand U4148 (N_4148,N_1976,N_1065);
or U4149 (N_4149,N_1804,N_699);
nor U4150 (N_4150,N_477,N_1422);
nor U4151 (N_4151,N_777,N_1029);
and U4152 (N_4152,N_401,N_2059);
and U4153 (N_4153,N_2172,N_2048);
nand U4154 (N_4154,N_1301,N_1664);
nand U4155 (N_4155,N_1274,N_655);
nand U4156 (N_4156,N_1695,N_1335);
nor U4157 (N_4157,N_1727,N_2289);
xor U4158 (N_4158,N_1095,N_1669);
or U4159 (N_4159,N_203,N_793);
xor U4160 (N_4160,N_219,N_904);
nand U4161 (N_4161,N_1036,N_1291);
nor U4162 (N_4162,N_578,N_1868);
nand U4163 (N_4163,N_1450,N_1933);
nor U4164 (N_4164,N_1272,N_643);
or U4165 (N_4165,N_538,N_2132);
nor U4166 (N_4166,N_1570,N_1849);
or U4167 (N_4167,N_1906,N_838);
nand U4168 (N_4168,N_1943,N_1931);
and U4169 (N_4169,N_743,N_858);
and U4170 (N_4170,N_174,N_1273);
or U4171 (N_4171,N_1001,N_2145);
or U4172 (N_4172,N_401,N_1773);
or U4173 (N_4173,N_2273,N_1197);
nor U4174 (N_4174,N_2291,N_1741);
nand U4175 (N_4175,N_109,N_1349);
nor U4176 (N_4176,N_2229,N_87);
nand U4177 (N_4177,N_178,N_1726);
or U4178 (N_4178,N_906,N_1057);
or U4179 (N_4179,N_2376,N_722);
nor U4180 (N_4180,N_651,N_251);
nand U4181 (N_4181,N_529,N_1545);
xnor U4182 (N_4182,N_1451,N_718);
nand U4183 (N_4183,N_468,N_40);
nand U4184 (N_4184,N_856,N_1561);
or U4185 (N_4185,N_435,N_253);
or U4186 (N_4186,N_423,N_1911);
or U4187 (N_4187,N_308,N_1343);
xnor U4188 (N_4188,N_2370,N_881);
nor U4189 (N_4189,N_1372,N_1120);
nand U4190 (N_4190,N_2264,N_118);
nor U4191 (N_4191,N_1081,N_1859);
nor U4192 (N_4192,N_1729,N_91);
or U4193 (N_4193,N_543,N_1921);
nor U4194 (N_4194,N_1054,N_2423);
nor U4195 (N_4195,N_143,N_1087);
nor U4196 (N_4196,N_235,N_774);
and U4197 (N_4197,N_635,N_2183);
and U4198 (N_4198,N_2254,N_2059);
xnor U4199 (N_4199,N_1882,N_1385);
nor U4200 (N_4200,N_412,N_1167);
nor U4201 (N_4201,N_1814,N_657);
or U4202 (N_4202,N_2012,N_503);
nor U4203 (N_4203,N_2005,N_695);
and U4204 (N_4204,N_569,N_435);
or U4205 (N_4205,N_1309,N_1369);
and U4206 (N_4206,N_1122,N_731);
nand U4207 (N_4207,N_135,N_1896);
and U4208 (N_4208,N_1811,N_853);
and U4209 (N_4209,N_1233,N_362);
nand U4210 (N_4210,N_405,N_2479);
or U4211 (N_4211,N_519,N_2287);
xor U4212 (N_4212,N_1845,N_2354);
xor U4213 (N_4213,N_2200,N_653);
xnor U4214 (N_4214,N_577,N_1071);
nor U4215 (N_4215,N_623,N_1433);
and U4216 (N_4216,N_327,N_364);
xnor U4217 (N_4217,N_61,N_1280);
nand U4218 (N_4218,N_1736,N_611);
and U4219 (N_4219,N_301,N_269);
and U4220 (N_4220,N_197,N_1588);
xor U4221 (N_4221,N_871,N_308);
nor U4222 (N_4222,N_2032,N_737);
nor U4223 (N_4223,N_384,N_1787);
nand U4224 (N_4224,N_848,N_231);
and U4225 (N_4225,N_1275,N_727);
or U4226 (N_4226,N_1068,N_1398);
nor U4227 (N_4227,N_694,N_2385);
or U4228 (N_4228,N_1914,N_355);
xnor U4229 (N_4229,N_2448,N_1933);
or U4230 (N_4230,N_1276,N_2022);
and U4231 (N_4231,N_1508,N_873);
and U4232 (N_4232,N_227,N_134);
nand U4233 (N_4233,N_1218,N_997);
or U4234 (N_4234,N_1686,N_51);
or U4235 (N_4235,N_783,N_2019);
or U4236 (N_4236,N_1828,N_1338);
and U4237 (N_4237,N_2287,N_1423);
xnor U4238 (N_4238,N_1455,N_471);
xnor U4239 (N_4239,N_1831,N_139);
and U4240 (N_4240,N_12,N_872);
xor U4241 (N_4241,N_1802,N_551);
and U4242 (N_4242,N_1388,N_2075);
nor U4243 (N_4243,N_1869,N_1482);
and U4244 (N_4244,N_545,N_1599);
nor U4245 (N_4245,N_704,N_1393);
xor U4246 (N_4246,N_2269,N_1337);
and U4247 (N_4247,N_1861,N_23);
xnor U4248 (N_4248,N_830,N_1274);
and U4249 (N_4249,N_1038,N_288);
nor U4250 (N_4250,N_1363,N_633);
xor U4251 (N_4251,N_2178,N_1731);
or U4252 (N_4252,N_1041,N_1770);
or U4253 (N_4253,N_1982,N_2158);
xor U4254 (N_4254,N_2338,N_1214);
nand U4255 (N_4255,N_1776,N_2065);
xor U4256 (N_4256,N_690,N_1610);
xnor U4257 (N_4257,N_1880,N_862);
or U4258 (N_4258,N_2158,N_321);
xnor U4259 (N_4259,N_2147,N_2066);
or U4260 (N_4260,N_220,N_432);
nand U4261 (N_4261,N_2131,N_1365);
nand U4262 (N_4262,N_944,N_2342);
and U4263 (N_4263,N_2357,N_1000);
nor U4264 (N_4264,N_2462,N_1055);
xnor U4265 (N_4265,N_2398,N_1890);
nand U4266 (N_4266,N_115,N_2281);
xnor U4267 (N_4267,N_1474,N_576);
or U4268 (N_4268,N_1904,N_838);
nand U4269 (N_4269,N_765,N_118);
xnor U4270 (N_4270,N_1969,N_2143);
nor U4271 (N_4271,N_1506,N_2183);
xnor U4272 (N_4272,N_926,N_2449);
and U4273 (N_4273,N_1078,N_1555);
or U4274 (N_4274,N_2193,N_1972);
nand U4275 (N_4275,N_659,N_1865);
or U4276 (N_4276,N_1010,N_1701);
nor U4277 (N_4277,N_1437,N_134);
xnor U4278 (N_4278,N_399,N_2087);
and U4279 (N_4279,N_1464,N_1430);
or U4280 (N_4280,N_2475,N_721);
or U4281 (N_4281,N_913,N_1863);
nor U4282 (N_4282,N_1897,N_2214);
nand U4283 (N_4283,N_1328,N_295);
nand U4284 (N_4284,N_1695,N_1102);
or U4285 (N_4285,N_1422,N_783);
nand U4286 (N_4286,N_610,N_615);
or U4287 (N_4287,N_1319,N_2119);
and U4288 (N_4288,N_250,N_2329);
xnor U4289 (N_4289,N_1256,N_2333);
or U4290 (N_4290,N_2016,N_1555);
and U4291 (N_4291,N_2396,N_2100);
or U4292 (N_4292,N_194,N_912);
nor U4293 (N_4293,N_2280,N_218);
nand U4294 (N_4294,N_379,N_1185);
xnor U4295 (N_4295,N_2132,N_328);
xor U4296 (N_4296,N_1890,N_1991);
nor U4297 (N_4297,N_166,N_1335);
nor U4298 (N_4298,N_1890,N_1269);
and U4299 (N_4299,N_2364,N_1572);
nor U4300 (N_4300,N_1138,N_1179);
xnor U4301 (N_4301,N_2121,N_1657);
or U4302 (N_4302,N_115,N_2334);
nand U4303 (N_4303,N_1815,N_1454);
xnor U4304 (N_4304,N_1294,N_2006);
or U4305 (N_4305,N_1598,N_549);
xor U4306 (N_4306,N_1698,N_238);
and U4307 (N_4307,N_252,N_1031);
xor U4308 (N_4308,N_6,N_1303);
nor U4309 (N_4309,N_460,N_1186);
nand U4310 (N_4310,N_601,N_2285);
or U4311 (N_4311,N_1721,N_718);
or U4312 (N_4312,N_1910,N_1680);
nand U4313 (N_4313,N_1471,N_2235);
and U4314 (N_4314,N_1988,N_2470);
nand U4315 (N_4315,N_49,N_1943);
nand U4316 (N_4316,N_1410,N_1557);
and U4317 (N_4317,N_2088,N_537);
nor U4318 (N_4318,N_2135,N_1883);
nor U4319 (N_4319,N_1174,N_508);
nand U4320 (N_4320,N_1033,N_2193);
nand U4321 (N_4321,N_2439,N_335);
and U4322 (N_4322,N_2326,N_1107);
and U4323 (N_4323,N_185,N_2312);
nor U4324 (N_4324,N_206,N_1146);
nor U4325 (N_4325,N_2499,N_1319);
nand U4326 (N_4326,N_2385,N_1286);
xnor U4327 (N_4327,N_271,N_1043);
nor U4328 (N_4328,N_1512,N_1398);
and U4329 (N_4329,N_2347,N_1391);
and U4330 (N_4330,N_1113,N_51);
nand U4331 (N_4331,N_1043,N_1799);
or U4332 (N_4332,N_782,N_2234);
xnor U4333 (N_4333,N_1669,N_922);
and U4334 (N_4334,N_1879,N_1022);
xnor U4335 (N_4335,N_1381,N_1129);
nand U4336 (N_4336,N_1854,N_1601);
nand U4337 (N_4337,N_93,N_1660);
and U4338 (N_4338,N_187,N_404);
and U4339 (N_4339,N_1221,N_2484);
nor U4340 (N_4340,N_677,N_87);
nand U4341 (N_4341,N_1162,N_1393);
or U4342 (N_4342,N_1632,N_1857);
and U4343 (N_4343,N_2446,N_1359);
and U4344 (N_4344,N_2159,N_2301);
and U4345 (N_4345,N_2083,N_1024);
nor U4346 (N_4346,N_798,N_2144);
nand U4347 (N_4347,N_57,N_1483);
nand U4348 (N_4348,N_214,N_1436);
nand U4349 (N_4349,N_459,N_2217);
nor U4350 (N_4350,N_1225,N_1821);
or U4351 (N_4351,N_1799,N_2398);
nand U4352 (N_4352,N_1060,N_2003);
or U4353 (N_4353,N_1079,N_1815);
or U4354 (N_4354,N_584,N_433);
and U4355 (N_4355,N_1993,N_2197);
or U4356 (N_4356,N_78,N_1859);
and U4357 (N_4357,N_984,N_1870);
nor U4358 (N_4358,N_287,N_1265);
and U4359 (N_4359,N_2184,N_2469);
and U4360 (N_4360,N_3,N_883);
and U4361 (N_4361,N_1956,N_108);
nor U4362 (N_4362,N_1063,N_1124);
xor U4363 (N_4363,N_2352,N_340);
or U4364 (N_4364,N_672,N_25);
nor U4365 (N_4365,N_568,N_2142);
nand U4366 (N_4366,N_1281,N_1848);
and U4367 (N_4367,N_2011,N_486);
and U4368 (N_4368,N_448,N_1781);
and U4369 (N_4369,N_1511,N_1134);
xor U4370 (N_4370,N_112,N_1181);
nor U4371 (N_4371,N_2189,N_1721);
xor U4372 (N_4372,N_177,N_1268);
xnor U4373 (N_4373,N_1333,N_688);
xor U4374 (N_4374,N_1914,N_1490);
nor U4375 (N_4375,N_391,N_2344);
xnor U4376 (N_4376,N_2260,N_689);
xnor U4377 (N_4377,N_1631,N_758);
and U4378 (N_4378,N_1710,N_917);
and U4379 (N_4379,N_1687,N_1432);
and U4380 (N_4380,N_1833,N_845);
xor U4381 (N_4381,N_1916,N_826);
xor U4382 (N_4382,N_2003,N_2143);
or U4383 (N_4383,N_787,N_486);
or U4384 (N_4384,N_2225,N_1220);
nand U4385 (N_4385,N_680,N_1287);
or U4386 (N_4386,N_1756,N_1489);
xor U4387 (N_4387,N_2466,N_891);
or U4388 (N_4388,N_419,N_1822);
or U4389 (N_4389,N_2393,N_1413);
nor U4390 (N_4390,N_1762,N_1082);
or U4391 (N_4391,N_376,N_35);
nand U4392 (N_4392,N_405,N_1968);
or U4393 (N_4393,N_1800,N_842);
xor U4394 (N_4394,N_940,N_1303);
nand U4395 (N_4395,N_84,N_1737);
nor U4396 (N_4396,N_2278,N_2162);
and U4397 (N_4397,N_1743,N_552);
or U4398 (N_4398,N_1264,N_1656);
nand U4399 (N_4399,N_723,N_1341);
xnor U4400 (N_4400,N_691,N_1184);
nor U4401 (N_4401,N_2040,N_2131);
nand U4402 (N_4402,N_2269,N_1133);
xor U4403 (N_4403,N_313,N_1838);
and U4404 (N_4404,N_2480,N_1202);
or U4405 (N_4405,N_1597,N_1252);
nor U4406 (N_4406,N_1528,N_817);
nand U4407 (N_4407,N_47,N_818);
and U4408 (N_4408,N_1560,N_1271);
nand U4409 (N_4409,N_1100,N_957);
nor U4410 (N_4410,N_681,N_2351);
or U4411 (N_4411,N_113,N_567);
nor U4412 (N_4412,N_537,N_2464);
and U4413 (N_4413,N_120,N_1607);
or U4414 (N_4414,N_1647,N_796);
xnor U4415 (N_4415,N_2198,N_760);
and U4416 (N_4416,N_222,N_1921);
nor U4417 (N_4417,N_1219,N_70);
nand U4418 (N_4418,N_1658,N_1221);
nor U4419 (N_4419,N_50,N_1821);
or U4420 (N_4420,N_1668,N_2187);
and U4421 (N_4421,N_1021,N_1893);
nand U4422 (N_4422,N_2224,N_668);
nor U4423 (N_4423,N_236,N_1822);
or U4424 (N_4424,N_905,N_2458);
nand U4425 (N_4425,N_1790,N_2136);
xnor U4426 (N_4426,N_1043,N_2185);
xnor U4427 (N_4427,N_1038,N_1975);
xnor U4428 (N_4428,N_1855,N_963);
nand U4429 (N_4429,N_1934,N_2116);
nor U4430 (N_4430,N_405,N_2052);
or U4431 (N_4431,N_2010,N_1346);
nand U4432 (N_4432,N_1684,N_1295);
or U4433 (N_4433,N_1606,N_2403);
nand U4434 (N_4434,N_1192,N_821);
nor U4435 (N_4435,N_300,N_964);
or U4436 (N_4436,N_1974,N_758);
or U4437 (N_4437,N_2070,N_217);
or U4438 (N_4438,N_2232,N_1846);
nor U4439 (N_4439,N_418,N_532);
nor U4440 (N_4440,N_1328,N_247);
and U4441 (N_4441,N_2,N_368);
nand U4442 (N_4442,N_1365,N_1746);
and U4443 (N_4443,N_469,N_696);
xnor U4444 (N_4444,N_1986,N_1203);
and U4445 (N_4445,N_2259,N_1216);
xnor U4446 (N_4446,N_197,N_671);
xnor U4447 (N_4447,N_1042,N_1596);
and U4448 (N_4448,N_2083,N_1020);
nand U4449 (N_4449,N_1243,N_1813);
xnor U4450 (N_4450,N_2352,N_618);
and U4451 (N_4451,N_1247,N_1357);
xnor U4452 (N_4452,N_349,N_1505);
nor U4453 (N_4453,N_2331,N_996);
and U4454 (N_4454,N_1455,N_1156);
nor U4455 (N_4455,N_1019,N_1720);
and U4456 (N_4456,N_586,N_297);
nor U4457 (N_4457,N_1404,N_1952);
and U4458 (N_4458,N_1252,N_172);
and U4459 (N_4459,N_2431,N_2240);
and U4460 (N_4460,N_317,N_2042);
or U4461 (N_4461,N_678,N_664);
or U4462 (N_4462,N_2208,N_1087);
or U4463 (N_4463,N_23,N_2080);
and U4464 (N_4464,N_1880,N_2402);
nor U4465 (N_4465,N_430,N_1283);
xnor U4466 (N_4466,N_2489,N_364);
and U4467 (N_4467,N_1788,N_1252);
nand U4468 (N_4468,N_1370,N_1951);
and U4469 (N_4469,N_1810,N_370);
or U4470 (N_4470,N_2456,N_2150);
nand U4471 (N_4471,N_1786,N_1925);
or U4472 (N_4472,N_2078,N_1654);
or U4473 (N_4473,N_2263,N_805);
xor U4474 (N_4474,N_185,N_1522);
nand U4475 (N_4475,N_587,N_1465);
or U4476 (N_4476,N_1465,N_1374);
and U4477 (N_4477,N_91,N_953);
nor U4478 (N_4478,N_2042,N_1839);
nor U4479 (N_4479,N_1975,N_1665);
nand U4480 (N_4480,N_214,N_637);
nor U4481 (N_4481,N_1814,N_1649);
xor U4482 (N_4482,N_1611,N_1089);
and U4483 (N_4483,N_429,N_916);
and U4484 (N_4484,N_1856,N_333);
nor U4485 (N_4485,N_1193,N_746);
or U4486 (N_4486,N_611,N_2478);
nand U4487 (N_4487,N_2305,N_445);
nor U4488 (N_4488,N_1156,N_2395);
nand U4489 (N_4489,N_1686,N_1699);
xnor U4490 (N_4490,N_2070,N_726);
and U4491 (N_4491,N_337,N_2204);
xor U4492 (N_4492,N_364,N_605);
and U4493 (N_4493,N_992,N_1008);
nand U4494 (N_4494,N_1888,N_312);
and U4495 (N_4495,N_1123,N_1787);
and U4496 (N_4496,N_1447,N_1721);
xnor U4497 (N_4497,N_2227,N_1869);
and U4498 (N_4498,N_1361,N_300);
and U4499 (N_4499,N_1709,N_2410);
nand U4500 (N_4500,N_1737,N_868);
nand U4501 (N_4501,N_162,N_1045);
and U4502 (N_4502,N_1348,N_1577);
nand U4503 (N_4503,N_691,N_525);
and U4504 (N_4504,N_714,N_173);
or U4505 (N_4505,N_343,N_1055);
and U4506 (N_4506,N_2131,N_1817);
nor U4507 (N_4507,N_2076,N_2015);
and U4508 (N_4508,N_2467,N_1625);
xnor U4509 (N_4509,N_1182,N_845);
nor U4510 (N_4510,N_417,N_1003);
nor U4511 (N_4511,N_2112,N_410);
nand U4512 (N_4512,N_2458,N_2464);
nand U4513 (N_4513,N_885,N_834);
nand U4514 (N_4514,N_1725,N_99);
and U4515 (N_4515,N_2388,N_1213);
nand U4516 (N_4516,N_2008,N_178);
nor U4517 (N_4517,N_786,N_1186);
xor U4518 (N_4518,N_1132,N_2354);
or U4519 (N_4519,N_277,N_1511);
xnor U4520 (N_4520,N_191,N_2428);
and U4521 (N_4521,N_317,N_1833);
and U4522 (N_4522,N_1621,N_37);
nor U4523 (N_4523,N_1186,N_868);
or U4524 (N_4524,N_145,N_1758);
nand U4525 (N_4525,N_1009,N_148);
nand U4526 (N_4526,N_657,N_1296);
nor U4527 (N_4527,N_795,N_2109);
and U4528 (N_4528,N_121,N_2242);
nor U4529 (N_4529,N_3,N_1218);
nand U4530 (N_4530,N_2054,N_1597);
nand U4531 (N_4531,N_1816,N_852);
xnor U4532 (N_4532,N_1008,N_2012);
nor U4533 (N_4533,N_2275,N_888);
nor U4534 (N_4534,N_2354,N_2280);
xnor U4535 (N_4535,N_172,N_1920);
and U4536 (N_4536,N_2109,N_1121);
nand U4537 (N_4537,N_2275,N_436);
nor U4538 (N_4538,N_2038,N_287);
xor U4539 (N_4539,N_1730,N_1428);
and U4540 (N_4540,N_423,N_776);
nand U4541 (N_4541,N_1225,N_858);
nor U4542 (N_4542,N_30,N_2468);
or U4543 (N_4543,N_226,N_512);
and U4544 (N_4544,N_647,N_1178);
and U4545 (N_4545,N_2374,N_28);
nor U4546 (N_4546,N_2414,N_2149);
xnor U4547 (N_4547,N_1215,N_1643);
or U4548 (N_4548,N_589,N_1129);
nand U4549 (N_4549,N_1123,N_264);
nor U4550 (N_4550,N_176,N_1892);
nand U4551 (N_4551,N_2043,N_2206);
nand U4552 (N_4552,N_1124,N_2281);
nand U4553 (N_4553,N_720,N_624);
nor U4554 (N_4554,N_1408,N_1127);
xor U4555 (N_4555,N_1267,N_2263);
nand U4556 (N_4556,N_1068,N_538);
nor U4557 (N_4557,N_74,N_2051);
xor U4558 (N_4558,N_375,N_2350);
nor U4559 (N_4559,N_1483,N_2127);
and U4560 (N_4560,N_793,N_1382);
xor U4561 (N_4561,N_1811,N_1010);
or U4562 (N_4562,N_284,N_1778);
nand U4563 (N_4563,N_1975,N_1318);
and U4564 (N_4564,N_1900,N_1168);
xnor U4565 (N_4565,N_1096,N_2429);
or U4566 (N_4566,N_2188,N_1764);
and U4567 (N_4567,N_1456,N_1756);
and U4568 (N_4568,N_856,N_337);
or U4569 (N_4569,N_1498,N_1752);
nor U4570 (N_4570,N_2174,N_288);
nor U4571 (N_4571,N_716,N_2071);
xnor U4572 (N_4572,N_755,N_943);
nor U4573 (N_4573,N_2376,N_1247);
nand U4574 (N_4574,N_1610,N_591);
xnor U4575 (N_4575,N_1509,N_119);
and U4576 (N_4576,N_263,N_22);
and U4577 (N_4577,N_1069,N_2031);
nand U4578 (N_4578,N_1040,N_1797);
or U4579 (N_4579,N_195,N_1479);
and U4580 (N_4580,N_1786,N_1791);
nor U4581 (N_4581,N_1518,N_635);
and U4582 (N_4582,N_1312,N_2218);
or U4583 (N_4583,N_2088,N_1668);
nor U4584 (N_4584,N_1403,N_965);
or U4585 (N_4585,N_1065,N_1300);
nand U4586 (N_4586,N_1459,N_2106);
nand U4587 (N_4587,N_876,N_1049);
and U4588 (N_4588,N_1162,N_2009);
nand U4589 (N_4589,N_1951,N_1427);
or U4590 (N_4590,N_1854,N_1948);
and U4591 (N_4591,N_1738,N_932);
nand U4592 (N_4592,N_1159,N_172);
nand U4593 (N_4593,N_114,N_2442);
and U4594 (N_4594,N_311,N_2272);
nand U4595 (N_4595,N_2186,N_2397);
xor U4596 (N_4596,N_1142,N_227);
nand U4597 (N_4597,N_2208,N_974);
nand U4598 (N_4598,N_463,N_1059);
nand U4599 (N_4599,N_2111,N_162);
or U4600 (N_4600,N_1816,N_21);
xor U4601 (N_4601,N_994,N_1354);
nor U4602 (N_4602,N_992,N_743);
xnor U4603 (N_4603,N_2202,N_765);
nor U4604 (N_4604,N_713,N_1945);
nand U4605 (N_4605,N_2274,N_1266);
and U4606 (N_4606,N_1395,N_592);
nand U4607 (N_4607,N_1430,N_1701);
nand U4608 (N_4608,N_2315,N_2181);
or U4609 (N_4609,N_619,N_1015);
and U4610 (N_4610,N_2369,N_1903);
nand U4611 (N_4611,N_257,N_2461);
nor U4612 (N_4612,N_959,N_756);
and U4613 (N_4613,N_981,N_2314);
nor U4614 (N_4614,N_135,N_1513);
and U4615 (N_4615,N_651,N_122);
xnor U4616 (N_4616,N_2301,N_1451);
nor U4617 (N_4617,N_2159,N_1348);
nor U4618 (N_4618,N_1632,N_1859);
or U4619 (N_4619,N_2402,N_1983);
xor U4620 (N_4620,N_2373,N_126);
and U4621 (N_4621,N_185,N_1896);
xnor U4622 (N_4622,N_1314,N_137);
and U4623 (N_4623,N_1151,N_37);
nor U4624 (N_4624,N_1482,N_1481);
xor U4625 (N_4625,N_2036,N_2384);
nor U4626 (N_4626,N_2272,N_2391);
or U4627 (N_4627,N_0,N_695);
and U4628 (N_4628,N_1860,N_762);
and U4629 (N_4629,N_1451,N_1051);
or U4630 (N_4630,N_2223,N_2018);
nor U4631 (N_4631,N_2486,N_1983);
nor U4632 (N_4632,N_2110,N_1174);
xnor U4633 (N_4633,N_2134,N_944);
xnor U4634 (N_4634,N_2080,N_106);
xnor U4635 (N_4635,N_711,N_1710);
xor U4636 (N_4636,N_2488,N_818);
and U4637 (N_4637,N_2274,N_1895);
nand U4638 (N_4638,N_123,N_1057);
nor U4639 (N_4639,N_898,N_336);
nand U4640 (N_4640,N_2192,N_475);
or U4641 (N_4641,N_1639,N_711);
nor U4642 (N_4642,N_1739,N_1254);
or U4643 (N_4643,N_2470,N_2474);
or U4644 (N_4644,N_2093,N_1089);
or U4645 (N_4645,N_1813,N_1096);
nand U4646 (N_4646,N_25,N_988);
and U4647 (N_4647,N_988,N_2135);
and U4648 (N_4648,N_694,N_1915);
nand U4649 (N_4649,N_1826,N_978);
xnor U4650 (N_4650,N_904,N_1026);
and U4651 (N_4651,N_1951,N_1311);
nand U4652 (N_4652,N_2093,N_1469);
xnor U4653 (N_4653,N_2320,N_2286);
nor U4654 (N_4654,N_2049,N_1057);
nand U4655 (N_4655,N_460,N_74);
xnor U4656 (N_4656,N_1781,N_2010);
xor U4657 (N_4657,N_1318,N_1159);
or U4658 (N_4658,N_2184,N_609);
and U4659 (N_4659,N_1019,N_1648);
or U4660 (N_4660,N_2062,N_2437);
nand U4661 (N_4661,N_674,N_1017);
nand U4662 (N_4662,N_258,N_629);
nor U4663 (N_4663,N_2091,N_2061);
xnor U4664 (N_4664,N_1665,N_25);
nand U4665 (N_4665,N_1835,N_796);
nor U4666 (N_4666,N_2493,N_512);
nor U4667 (N_4667,N_809,N_775);
or U4668 (N_4668,N_1412,N_479);
xor U4669 (N_4669,N_381,N_1246);
or U4670 (N_4670,N_625,N_240);
or U4671 (N_4671,N_1243,N_2026);
or U4672 (N_4672,N_2146,N_367);
nand U4673 (N_4673,N_2076,N_447);
xnor U4674 (N_4674,N_1344,N_840);
and U4675 (N_4675,N_1001,N_316);
or U4676 (N_4676,N_635,N_107);
nand U4677 (N_4677,N_2349,N_1081);
and U4678 (N_4678,N_1049,N_812);
or U4679 (N_4679,N_1516,N_1019);
nand U4680 (N_4680,N_1992,N_372);
nor U4681 (N_4681,N_362,N_2030);
or U4682 (N_4682,N_2216,N_2021);
xor U4683 (N_4683,N_1056,N_823);
and U4684 (N_4684,N_841,N_579);
nor U4685 (N_4685,N_1760,N_2311);
xnor U4686 (N_4686,N_1358,N_377);
xnor U4687 (N_4687,N_2279,N_99);
or U4688 (N_4688,N_2034,N_967);
and U4689 (N_4689,N_1607,N_619);
or U4690 (N_4690,N_229,N_1487);
and U4691 (N_4691,N_198,N_891);
nand U4692 (N_4692,N_824,N_1396);
nor U4693 (N_4693,N_1520,N_59);
nor U4694 (N_4694,N_2080,N_2045);
or U4695 (N_4695,N_771,N_1260);
nand U4696 (N_4696,N_1378,N_1480);
xnor U4697 (N_4697,N_45,N_1855);
nor U4698 (N_4698,N_964,N_842);
xnor U4699 (N_4699,N_673,N_1674);
or U4700 (N_4700,N_621,N_1152);
nor U4701 (N_4701,N_1771,N_2244);
nor U4702 (N_4702,N_360,N_2475);
nand U4703 (N_4703,N_377,N_1233);
and U4704 (N_4704,N_946,N_239);
xnor U4705 (N_4705,N_277,N_1027);
and U4706 (N_4706,N_571,N_582);
nand U4707 (N_4707,N_2382,N_1215);
nand U4708 (N_4708,N_103,N_353);
nor U4709 (N_4709,N_2368,N_206);
nand U4710 (N_4710,N_911,N_1299);
and U4711 (N_4711,N_1282,N_1243);
nor U4712 (N_4712,N_817,N_1540);
or U4713 (N_4713,N_640,N_940);
xor U4714 (N_4714,N_1942,N_2046);
xnor U4715 (N_4715,N_1038,N_2037);
xor U4716 (N_4716,N_2032,N_2076);
nor U4717 (N_4717,N_1097,N_2285);
xnor U4718 (N_4718,N_357,N_1140);
nor U4719 (N_4719,N_1773,N_697);
nand U4720 (N_4720,N_1396,N_748);
xor U4721 (N_4721,N_2305,N_2070);
or U4722 (N_4722,N_2237,N_2343);
and U4723 (N_4723,N_1833,N_1326);
and U4724 (N_4724,N_1191,N_206);
or U4725 (N_4725,N_2278,N_483);
nor U4726 (N_4726,N_1741,N_1844);
nor U4727 (N_4727,N_217,N_878);
nand U4728 (N_4728,N_14,N_382);
nand U4729 (N_4729,N_672,N_1887);
nand U4730 (N_4730,N_333,N_1093);
xor U4731 (N_4731,N_256,N_2335);
and U4732 (N_4732,N_823,N_1272);
nor U4733 (N_4733,N_1246,N_1225);
and U4734 (N_4734,N_2190,N_1753);
or U4735 (N_4735,N_570,N_491);
nor U4736 (N_4736,N_320,N_1226);
nor U4737 (N_4737,N_1911,N_298);
nand U4738 (N_4738,N_1693,N_2178);
or U4739 (N_4739,N_1139,N_2365);
nor U4740 (N_4740,N_12,N_420);
nor U4741 (N_4741,N_1958,N_2352);
xnor U4742 (N_4742,N_805,N_272);
xor U4743 (N_4743,N_1067,N_320);
xor U4744 (N_4744,N_961,N_1410);
or U4745 (N_4745,N_1908,N_1681);
nand U4746 (N_4746,N_1057,N_1557);
or U4747 (N_4747,N_958,N_236);
nor U4748 (N_4748,N_504,N_1807);
nor U4749 (N_4749,N_817,N_1329);
xor U4750 (N_4750,N_136,N_86);
nand U4751 (N_4751,N_713,N_172);
nor U4752 (N_4752,N_2160,N_1359);
or U4753 (N_4753,N_1166,N_1820);
xor U4754 (N_4754,N_712,N_1153);
nand U4755 (N_4755,N_956,N_187);
nor U4756 (N_4756,N_1307,N_2453);
and U4757 (N_4757,N_853,N_620);
or U4758 (N_4758,N_613,N_2239);
and U4759 (N_4759,N_1024,N_2278);
nor U4760 (N_4760,N_1273,N_450);
xnor U4761 (N_4761,N_1520,N_378);
xnor U4762 (N_4762,N_556,N_725);
or U4763 (N_4763,N_1235,N_2452);
nand U4764 (N_4764,N_2031,N_1992);
or U4765 (N_4765,N_1336,N_2337);
and U4766 (N_4766,N_2350,N_1553);
nor U4767 (N_4767,N_816,N_2391);
or U4768 (N_4768,N_714,N_196);
and U4769 (N_4769,N_161,N_1063);
nor U4770 (N_4770,N_247,N_1046);
or U4771 (N_4771,N_319,N_1250);
nand U4772 (N_4772,N_1673,N_2362);
xor U4773 (N_4773,N_223,N_2446);
nand U4774 (N_4774,N_1254,N_147);
nor U4775 (N_4775,N_778,N_81);
nand U4776 (N_4776,N_2370,N_104);
nor U4777 (N_4777,N_1312,N_425);
and U4778 (N_4778,N_2041,N_2127);
nor U4779 (N_4779,N_1017,N_477);
and U4780 (N_4780,N_218,N_2121);
nand U4781 (N_4781,N_2145,N_1016);
nand U4782 (N_4782,N_1688,N_1912);
or U4783 (N_4783,N_1334,N_1655);
or U4784 (N_4784,N_1682,N_1145);
and U4785 (N_4785,N_1286,N_80);
xnor U4786 (N_4786,N_934,N_1149);
nor U4787 (N_4787,N_1567,N_864);
nor U4788 (N_4788,N_772,N_2293);
and U4789 (N_4789,N_460,N_497);
and U4790 (N_4790,N_479,N_1195);
or U4791 (N_4791,N_2153,N_432);
nor U4792 (N_4792,N_854,N_954);
nor U4793 (N_4793,N_1842,N_1811);
xor U4794 (N_4794,N_894,N_652);
nand U4795 (N_4795,N_1328,N_417);
xor U4796 (N_4796,N_1055,N_2108);
and U4797 (N_4797,N_1576,N_474);
and U4798 (N_4798,N_1570,N_1388);
xnor U4799 (N_4799,N_42,N_1392);
and U4800 (N_4800,N_1179,N_1431);
and U4801 (N_4801,N_1031,N_862);
nor U4802 (N_4802,N_979,N_704);
nor U4803 (N_4803,N_91,N_1631);
and U4804 (N_4804,N_677,N_1885);
xnor U4805 (N_4805,N_1621,N_1213);
or U4806 (N_4806,N_1366,N_273);
and U4807 (N_4807,N_1094,N_1342);
or U4808 (N_4808,N_510,N_1032);
xor U4809 (N_4809,N_1441,N_917);
and U4810 (N_4810,N_1677,N_1222);
nor U4811 (N_4811,N_1119,N_58);
nor U4812 (N_4812,N_677,N_1262);
xor U4813 (N_4813,N_1364,N_1774);
and U4814 (N_4814,N_285,N_1833);
nand U4815 (N_4815,N_2047,N_427);
or U4816 (N_4816,N_459,N_759);
or U4817 (N_4817,N_687,N_596);
nand U4818 (N_4818,N_2068,N_214);
and U4819 (N_4819,N_1164,N_1017);
nor U4820 (N_4820,N_829,N_229);
xor U4821 (N_4821,N_639,N_2);
xnor U4822 (N_4822,N_2120,N_745);
xor U4823 (N_4823,N_1245,N_636);
xnor U4824 (N_4824,N_610,N_1259);
and U4825 (N_4825,N_354,N_538);
xnor U4826 (N_4826,N_38,N_2229);
nor U4827 (N_4827,N_1239,N_2409);
xnor U4828 (N_4828,N_333,N_215);
nand U4829 (N_4829,N_436,N_159);
nor U4830 (N_4830,N_24,N_710);
xor U4831 (N_4831,N_449,N_895);
nand U4832 (N_4832,N_991,N_1331);
or U4833 (N_4833,N_397,N_2227);
and U4834 (N_4834,N_535,N_1294);
nor U4835 (N_4835,N_1501,N_185);
or U4836 (N_4836,N_1422,N_2033);
or U4837 (N_4837,N_308,N_1657);
nand U4838 (N_4838,N_588,N_1523);
xnor U4839 (N_4839,N_761,N_388);
nand U4840 (N_4840,N_107,N_412);
and U4841 (N_4841,N_1824,N_352);
or U4842 (N_4842,N_170,N_2462);
xor U4843 (N_4843,N_2345,N_755);
xor U4844 (N_4844,N_1872,N_694);
nor U4845 (N_4845,N_692,N_568);
nand U4846 (N_4846,N_1834,N_2009);
or U4847 (N_4847,N_645,N_1235);
nand U4848 (N_4848,N_2184,N_1840);
xor U4849 (N_4849,N_2303,N_2122);
xnor U4850 (N_4850,N_2487,N_1967);
nor U4851 (N_4851,N_1670,N_2194);
nor U4852 (N_4852,N_1490,N_44);
or U4853 (N_4853,N_1152,N_1913);
nor U4854 (N_4854,N_1749,N_1124);
nand U4855 (N_4855,N_2340,N_1227);
or U4856 (N_4856,N_2032,N_1213);
nor U4857 (N_4857,N_1877,N_863);
and U4858 (N_4858,N_788,N_1440);
xnor U4859 (N_4859,N_1660,N_446);
xor U4860 (N_4860,N_2322,N_536);
or U4861 (N_4861,N_355,N_1294);
and U4862 (N_4862,N_113,N_2424);
or U4863 (N_4863,N_2330,N_718);
and U4864 (N_4864,N_1991,N_670);
or U4865 (N_4865,N_568,N_1081);
nor U4866 (N_4866,N_81,N_1902);
and U4867 (N_4867,N_1313,N_1391);
nand U4868 (N_4868,N_2084,N_361);
xor U4869 (N_4869,N_2342,N_1980);
or U4870 (N_4870,N_1287,N_1167);
and U4871 (N_4871,N_1441,N_1427);
or U4872 (N_4872,N_1368,N_1514);
nor U4873 (N_4873,N_1989,N_1422);
nand U4874 (N_4874,N_2045,N_2443);
and U4875 (N_4875,N_1172,N_1647);
nor U4876 (N_4876,N_1956,N_1172);
xnor U4877 (N_4877,N_320,N_1135);
xnor U4878 (N_4878,N_103,N_1766);
nand U4879 (N_4879,N_1874,N_1611);
and U4880 (N_4880,N_1993,N_1154);
or U4881 (N_4881,N_1271,N_159);
or U4882 (N_4882,N_653,N_2055);
xnor U4883 (N_4883,N_489,N_524);
or U4884 (N_4884,N_1198,N_286);
or U4885 (N_4885,N_241,N_2431);
or U4886 (N_4886,N_1472,N_506);
nand U4887 (N_4887,N_1802,N_282);
and U4888 (N_4888,N_833,N_355);
nor U4889 (N_4889,N_928,N_2372);
nor U4890 (N_4890,N_1800,N_1212);
or U4891 (N_4891,N_284,N_599);
and U4892 (N_4892,N_550,N_652);
or U4893 (N_4893,N_261,N_140);
nor U4894 (N_4894,N_343,N_192);
xnor U4895 (N_4895,N_2221,N_2300);
nand U4896 (N_4896,N_2050,N_1806);
nand U4897 (N_4897,N_1182,N_1978);
and U4898 (N_4898,N_1813,N_1026);
xnor U4899 (N_4899,N_658,N_2059);
nor U4900 (N_4900,N_2412,N_2064);
xor U4901 (N_4901,N_1916,N_712);
xnor U4902 (N_4902,N_1828,N_1693);
or U4903 (N_4903,N_1471,N_250);
and U4904 (N_4904,N_1342,N_128);
xnor U4905 (N_4905,N_2,N_2192);
xor U4906 (N_4906,N_515,N_2075);
and U4907 (N_4907,N_463,N_2377);
nor U4908 (N_4908,N_1226,N_634);
or U4909 (N_4909,N_1892,N_1431);
nor U4910 (N_4910,N_395,N_235);
xor U4911 (N_4911,N_2422,N_1761);
nor U4912 (N_4912,N_2242,N_13);
and U4913 (N_4913,N_1565,N_2463);
and U4914 (N_4914,N_65,N_2496);
nor U4915 (N_4915,N_1009,N_23);
and U4916 (N_4916,N_2430,N_328);
nor U4917 (N_4917,N_1380,N_2103);
nor U4918 (N_4918,N_1224,N_1488);
nand U4919 (N_4919,N_2473,N_194);
nand U4920 (N_4920,N_1664,N_508);
nand U4921 (N_4921,N_1580,N_646);
xor U4922 (N_4922,N_534,N_1413);
and U4923 (N_4923,N_1289,N_2461);
and U4924 (N_4924,N_1256,N_1676);
xnor U4925 (N_4925,N_1238,N_2027);
nand U4926 (N_4926,N_234,N_898);
or U4927 (N_4927,N_1327,N_1099);
or U4928 (N_4928,N_1377,N_63);
and U4929 (N_4929,N_2268,N_1282);
or U4930 (N_4930,N_1824,N_1546);
and U4931 (N_4931,N_1645,N_1827);
xnor U4932 (N_4932,N_271,N_1059);
xor U4933 (N_4933,N_229,N_2495);
and U4934 (N_4934,N_1562,N_490);
nand U4935 (N_4935,N_2195,N_960);
nor U4936 (N_4936,N_161,N_2442);
nand U4937 (N_4937,N_1156,N_807);
nor U4938 (N_4938,N_2256,N_466);
nor U4939 (N_4939,N_491,N_720);
or U4940 (N_4940,N_1578,N_2260);
nor U4941 (N_4941,N_1797,N_455);
and U4942 (N_4942,N_590,N_887);
nor U4943 (N_4943,N_2203,N_267);
xnor U4944 (N_4944,N_1564,N_2208);
nor U4945 (N_4945,N_18,N_2403);
nand U4946 (N_4946,N_1211,N_2070);
nor U4947 (N_4947,N_1624,N_1628);
or U4948 (N_4948,N_979,N_1142);
nand U4949 (N_4949,N_409,N_538);
xor U4950 (N_4950,N_1062,N_1532);
xor U4951 (N_4951,N_1540,N_651);
nor U4952 (N_4952,N_2383,N_1332);
nor U4953 (N_4953,N_587,N_1568);
nor U4954 (N_4954,N_2049,N_841);
and U4955 (N_4955,N_2463,N_2284);
nor U4956 (N_4956,N_37,N_122);
and U4957 (N_4957,N_583,N_993);
or U4958 (N_4958,N_890,N_1285);
xnor U4959 (N_4959,N_1749,N_1108);
nor U4960 (N_4960,N_566,N_2047);
and U4961 (N_4961,N_421,N_2494);
and U4962 (N_4962,N_69,N_539);
and U4963 (N_4963,N_2045,N_2137);
nand U4964 (N_4964,N_2094,N_1648);
xor U4965 (N_4965,N_921,N_1193);
nor U4966 (N_4966,N_145,N_1130);
and U4967 (N_4967,N_761,N_1526);
xnor U4968 (N_4968,N_1006,N_852);
nor U4969 (N_4969,N_1354,N_2335);
or U4970 (N_4970,N_1761,N_392);
xor U4971 (N_4971,N_1570,N_263);
nand U4972 (N_4972,N_648,N_171);
nor U4973 (N_4973,N_113,N_839);
or U4974 (N_4974,N_812,N_805);
or U4975 (N_4975,N_221,N_1810);
nand U4976 (N_4976,N_804,N_2389);
nand U4977 (N_4977,N_2061,N_1140);
nor U4978 (N_4978,N_820,N_1408);
xor U4979 (N_4979,N_548,N_545);
or U4980 (N_4980,N_51,N_1044);
nand U4981 (N_4981,N_1062,N_1695);
nor U4982 (N_4982,N_1600,N_296);
nor U4983 (N_4983,N_688,N_2139);
nand U4984 (N_4984,N_1507,N_1725);
nor U4985 (N_4985,N_1674,N_1407);
nor U4986 (N_4986,N_666,N_1199);
nor U4987 (N_4987,N_2120,N_1997);
or U4988 (N_4988,N_568,N_52);
and U4989 (N_4989,N_2297,N_104);
or U4990 (N_4990,N_1733,N_212);
or U4991 (N_4991,N_665,N_1486);
or U4992 (N_4992,N_1849,N_2386);
xor U4993 (N_4993,N_947,N_1250);
xnor U4994 (N_4994,N_1949,N_102);
xnor U4995 (N_4995,N_697,N_1177);
and U4996 (N_4996,N_1894,N_2110);
and U4997 (N_4997,N_633,N_101);
nand U4998 (N_4998,N_1748,N_846);
nand U4999 (N_4999,N_1766,N_736);
xor U5000 (N_5000,N_3805,N_4149);
nand U5001 (N_5001,N_2563,N_3787);
or U5002 (N_5002,N_3737,N_2709);
xor U5003 (N_5003,N_4825,N_2706);
and U5004 (N_5004,N_3840,N_2605);
xnor U5005 (N_5005,N_3899,N_2717);
or U5006 (N_5006,N_2946,N_3161);
or U5007 (N_5007,N_4027,N_3584);
nand U5008 (N_5008,N_3814,N_3617);
nand U5009 (N_5009,N_4864,N_3363);
nand U5010 (N_5010,N_4764,N_3104);
or U5011 (N_5011,N_3693,N_2512);
nor U5012 (N_5012,N_3644,N_4925);
or U5013 (N_5013,N_3373,N_4097);
and U5014 (N_5014,N_2708,N_4932);
and U5015 (N_5015,N_4496,N_4677);
nor U5016 (N_5016,N_3258,N_4719);
nor U5017 (N_5017,N_2726,N_4237);
xor U5018 (N_5018,N_2772,N_4566);
and U5019 (N_5019,N_2812,N_3388);
nor U5020 (N_5020,N_3222,N_4740);
and U5021 (N_5021,N_4125,N_3521);
or U5022 (N_5022,N_2634,N_3543);
xnor U5023 (N_5023,N_2588,N_2650);
or U5024 (N_5024,N_4300,N_4054);
xor U5025 (N_5025,N_4669,N_3582);
and U5026 (N_5026,N_4734,N_3763);
nand U5027 (N_5027,N_3485,N_3205);
nand U5028 (N_5028,N_4281,N_4470);
xor U5029 (N_5029,N_3869,N_4327);
xnor U5030 (N_5030,N_4851,N_4235);
or U5031 (N_5031,N_3507,N_2527);
and U5032 (N_5032,N_3371,N_2889);
xor U5033 (N_5033,N_3483,N_3106);
and U5034 (N_5034,N_4041,N_2851);
nand U5035 (N_5035,N_2682,N_3756);
nand U5036 (N_5036,N_3623,N_4941);
or U5037 (N_5037,N_3727,N_4874);
or U5038 (N_5038,N_2674,N_3921);
and U5039 (N_5039,N_3083,N_2891);
or U5040 (N_5040,N_4642,N_4778);
or U5041 (N_5041,N_3826,N_4152);
nor U5042 (N_5042,N_4631,N_3908);
and U5043 (N_5043,N_3895,N_3233);
nor U5044 (N_5044,N_3070,N_3073);
or U5045 (N_5045,N_3094,N_3467);
nor U5046 (N_5046,N_3568,N_3360);
and U5047 (N_5047,N_3802,N_3912);
and U5048 (N_5048,N_4559,N_3384);
or U5049 (N_5049,N_4294,N_2737);
nor U5050 (N_5050,N_3559,N_3565);
and U5051 (N_5051,N_3036,N_2947);
xnor U5052 (N_5052,N_4929,N_3675);
nand U5053 (N_5053,N_4543,N_4093);
and U5054 (N_5054,N_3628,N_4164);
and U5055 (N_5055,N_4179,N_3063);
or U5056 (N_5056,N_4022,N_3116);
nor U5057 (N_5057,N_3374,N_4107);
and U5058 (N_5058,N_4563,N_3410);
nor U5059 (N_5059,N_3976,N_3223);
or U5060 (N_5060,N_4920,N_3798);
nor U5061 (N_5061,N_3468,N_4945);
xor U5062 (N_5062,N_3757,N_3361);
nor U5063 (N_5063,N_3231,N_4910);
or U5064 (N_5064,N_2585,N_2752);
xnor U5065 (N_5065,N_3602,N_4103);
nand U5066 (N_5066,N_4005,N_2562);
xnor U5067 (N_5067,N_4341,N_3867);
nor U5068 (N_5068,N_4254,N_3438);
or U5069 (N_5069,N_4167,N_3042);
and U5070 (N_5070,N_4940,N_4224);
nor U5071 (N_5071,N_2932,N_2804);
xnor U5072 (N_5072,N_3989,N_3389);
or U5073 (N_5073,N_3387,N_2616);
and U5074 (N_5074,N_3301,N_4445);
or U5075 (N_5075,N_4405,N_3055);
nand U5076 (N_5076,N_3093,N_3303);
xor U5077 (N_5077,N_2557,N_4819);
nor U5078 (N_5078,N_4935,N_4183);
nand U5079 (N_5079,N_3133,N_2956);
or U5080 (N_5080,N_4219,N_3206);
nor U5081 (N_5081,N_4367,N_2978);
nand U5082 (N_5082,N_3679,N_4700);
xor U5083 (N_5083,N_2698,N_4619);
nor U5084 (N_5084,N_3536,N_4936);
xor U5085 (N_5085,N_3624,N_4604);
xor U5086 (N_5086,N_3350,N_4142);
or U5087 (N_5087,N_2710,N_3605);
nor U5088 (N_5088,N_2846,N_3382);
nand U5089 (N_5089,N_4443,N_3829);
and U5090 (N_5090,N_4964,N_4261);
nand U5091 (N_5091,N_4453,N_3843);
nand U5092 (N_5092,N_4966,N_4109);
xor U5093 (N_5093,N_3777,N_4476);
or U5094 (N_5094,N_3851,N_2509);
nor U5095 (N_5095,N_2874,N_4564);
xor U5096 (N_5096,N_3909,N_3316);
nor U5097 (N_5097,N_4113,N_4086);
nand U5098 (N_5098,N_4413,N_4870);
nor U5099 (N_5099,N_3721,N_2644);
or U5100 (N_5100,N_4462,N_3689);
nand U5101 (N_5101,N_3978,N_2856);
and U5102 (N_5102,N_4833,N_3393);
and U5103 (N_5103,N_2511,N_4065);
nand U5104 (N_5104,N_4270,N_3033);
xor U5105 (N_5105,N_4577,N_2763);
and U5106 (N_5106,N_2522,N_4494);
and U5107 (N_5107,N_4360,N_3118);
nor U5108 (N_5108,N_4205,N_3060);
or U5109 (N_5109,N_3232,N_3749);
xor U5110 (N_5110,N_4781,N_2739);
xnor U5111 (N_5111,N_3918,N_4776);
xnor U5112 (N_5112,N_3834,N_3186);
nand U5113 (N_5113,N_3383,N_3764);
or U5114 (N_5114,N_3669,N_4807);
nor U5115 (N_5115,N_3923,N_4621);
xnor U5116 (N_5116,N_3882,N_2906);
or U5117 (N_5117,N_3012,N_3920);
xor U5118 (N_5118,N_4542,N_4601);
xnor U5119 (N_5119,N_2681,N_2952);
nand U5120 (N_5120,N_2530,N_2529);
xnor U5121 (N_5121,N_3422,N_3919);
or U5122 (N_5122,N_3202,N_4288);
nand U5123 (N_5123,N_3611,N_3001);
or U5124 (N_5124,N_3889,N_3088);
xnor U5125 (N_5125,N_3026,N_4722);
nor U5126 (N_5126,N_4575,N_2531);
or U5127 (N_5127,N_2842,N_4772);
xor U5128 (N_5128,N_2535,N_4828);
nor U5129 (N_5129,N_3121,N_4909);
nor U5130 (N_5130,N_3459,N_3961);
or U5131 (N_5131,N_4188,N_4197);
or U5132 (N_5132,N_2673,N_4387);
nor U5133 (N_5133,N_3520,N_3509);
nand U5134 (N_5134,N_2643,N_3250);
nand U5135 (N_5135,N_4049,N_2518);
nor U5136 (N_5136,N_4531,N_4757);
nor U5137 (N_5137,N_4510,N_3988);
nand U5138 (N_5138,N_3898,N_3537);
xor U5139 (N_5139,N_3246,N_4505);
nor U5140 (N_5140,N_3181,N_3442);
nand U5141 (N_5141,N_3977,N_4970);
or U5142 (N_5142,N_4344,N_3254);
and U5143 (N_5143,N_3030,N_4804);
or U5144 (N_5144,N_3200,N_4641);
xnor U5145 (N_5145,N_4115,N_2596);
xor U5146 (N_5146,N_2555,N_4884);
and U5147 (N_5147,N_4056,N_3691);
and U5148 (N_5148,N_3610,N_3220);
and U5149 (N_5149,N_4253,N_2676);
nand U5150 (N_5150,N_2750,N_3453);
nor U5151 (N_5151,N_4245,N_3684);
xnor U5152 (N_5152,N_2994,N_2897);
xor U5153 (N_5153,N_4878,N_4763);
xnor U5154 (N_5154,N_3658,N_2927);
and U5155 (N_5155,N_2707,N_4528);
or U5156 (N_5156,N_4195,N_3115);
or U5157 (N_5157,N_3355,N_4385);
nand U5158 (N_5158,N_2930,N_3883);
xnor U5159 (N_5159,N_4745,N_3569);
nand U5160 (N_5160,N_3928,N_3759);
or U5161 (N_5161,N_3991,N_3709);
xor U5162 (N_5162,N_3852,N_4368);
xor U5163 (N_5163,N_2951,N_2558);
nand U5164 (N_5164,N_4530,N_4014);
or U5165 (N_5165,N_2547,N_4068);
or U5166 (N_5166,N_2798,N_4892);
or U5167 (N_5167,N_2918,N_3000);
nand U5168 (N_5168,N_4267,N_2971);
xnor U5169 (N_5169,N_4287,N_3212);
and U5170 (N_5170,N_2655,N_3279);
and U5171 (N_5171,N_4608,N_4006);
and U5172 (N_5172,N_4317,N_4981);
and U5173 (N_5173,N_4104,N_4003);
xor U5174 (N_5174,N_4436,N_4334);
or U5175 (N_5175,N_4928,N_2975);
xnor U5176 (N_5176,N_3681,N_3514);
nor U5177 (N_5177,N_3622,N_3994);
xnor U5178 (N_5178,N_2913,N_3966);
nor U5179 (N_5179,N_2546,N_3170);
nand U5180 (N_5180,N_4428,N_3642);
nor U5181 (N_5181,N_4343,N_3803);
nor U5182 (N_5182,N_4364,N_4536);
and U5183 (N_5183,N_2669,N_4656);
and U5184 (N_5184,N_3261,N_4043);
nor U5185 (N_5185,N_3445,N_4371);
or U5186 (N_5186,N_4643,N_4708);
xnor U5187 (N_5187,N_4401,N_3513);
nand U5188 (N_5188,N_4816,N_3005);
nor U5189 (N_5189,N_2955,N_4144);
and U5190 (N_5190,N_4626,N_3390);
or U5191 (N_5191,N_3735,N_4122);
nor U5192 (N_5192,N_4544,N_4280);
and U5193 (N_5193,N_3169,N_2735);
xnor U5194 (N_5194,N_4948,N_4310);
xnor U5195 (N_5195,N_4241,N_4567);
nand U5196 (N_5196,N_2705,N_3431);
nand U5197 (N_5197,N_3424,N_4551);
nand U5198 (N_5198,N_4859,N_3992);
and U5199 (N_5199,N_4001,N_3105);
nand U5200 (N_5200,N_3493,N_2774);
and U5201 (N_5201,N_2582,N_3217);
and U5202 (N_5202,N_3810,N_4308);
and U5203 (N_5203,N_2861,N_3340);
or U5204 (N_5204,N_3574,N_3465);
xnor U5205 (N_5205,N_4046,N_3187);
nand U5206 (N_5206,N_4244,N_3392);
xnor U5207 (N_5207,N_3017,N_3213);
nor U5208 (N_5208,N_2755,N_4926);
and U5209 (N_5209,N_4934,N_3227);
xor U5210 (N_5210,N_3315,N_4016);
and U5211 (N_5211,N_4432,N_3462);
and U5212 (N_5212,N_2506,N_4206);
and U5213 (N_5213,N_3915,N_3469);
xnor U5214 (N_5214,N_3307,N_2614);
or U5215 (N_5215,N_2924,N_3694);
nor U5216 (N_5216,N_3114,N_2981);
nand U5217 (N_5217,N_4134,N_3690);
xnor U5218 (N_5218,N_4584,N_2607);
nor U5219 (N_5219,N_3306,N_3646);
nor U5220 (N_5220,N_2618,N_3761);
nor U5221 (N_5221,N_4562,N_3818);
nand U5222 (N_5222,N_4974,N_3224);
or U5223 (N_5223,N_4227,N_2890);
nand U5224 (N_5224,N_3823,N_3583);
xor U5225 (N_5225,N_3504,N_2896);
nand U5226 (N_5226,N_2830,N_4318);
or U5227 (N_5227,N_4306,N_4486);
or U5228 (N_5228,N_4750,N_4073);
and U5229 (N_5229,N_4408,N_4667);
nor U5230 (N_5230,N_4618,N_3201);
nand U5231 (N_5231,N_4571,N_3348);
nor U5232 (N_5232,N_2699,N_4855);
or U5233 (N_5233,N_3796,N_3386);
nor U5234 (N_5234,N_3308,N_3241);
or U5235 (N_5235,N_4037,N_4760);
or U5236 (N_5236,N_3952,N_4507);
xnor U5237 (N_5237,N_3771,N_4611);
nand U5238 (N_5238,N_2559,N_2844);
xor U5239 (N_5239,N_4574,N_4877);
and U5240 (N_5240,N_4256,N_3656);
xnor U5241 (N_5241,N_3828,N_4379);
nor U5242 (N_5242,N_4495,N_3865);
nor U5243 (N_5243,N_4943,N_3497);
and U5244 (N_5244,N_4013,N_4250);
or U5245 (N_5245,N_2756,N_4370);
nor U5246 (N_5246,N_4490,N_4117);
and U5247 (N_5247,N_2568,N_2664);
nand U5248 (N_5248,N_3337,N_3282);
nand U5249 (N_5249,N_4994,N_2769);
nor U5250 (N_5250,N_4305,N_4140);
nor U5251 (N_5251,N_3550,N_3578);
or U5252 (N_5252,N_2933,N_3564);
nor U5253 (N_5253,N_2868,N_4890);
nor U5254 (N_5254,N_2865,N_4808);
or U5255 (N_5255,N_4578,N_4896);
or U5256 (N_5256,N_4595,N_2575);
nand U5257 (N_5257,N_4707,N_3357);
xnor U5258 (N_5258,N_2524,N_4148);
nand U5259 (N_5259,N_3238,N_3334);
nor U5260 (N_5260,N_3318,N_4463);
nand U5261 (N_5261,N_4191,N_4102);
and U5262 (N_5262,N_2803,N_2824);
xnor U5263 (N_5263,N_4441,N_4228);
and U5264 (N_5264,N_2572,N_3451);
nor U5265 (N_5265,N_3524,N_4678);
or U5266 (N_5266,N_3893,N_4025);
xor U5267 (N_5267,N_3714,N_4587);
xnor U5268 (N_5268,N_3144,N_3738);
and U5269 (N_5269,N_2734,N_4609);
or U5270 (N_5270,N_4127,N_3519);
and U5271 (N_5271,N_4946,N_2802);
or U5272 (N_5272,N_3715,N_4735);
and U5273 (N_5273,N_4849,N_3833);
and U5274 (N_5274,N_4889,N_4454);
or U5275 (N_5275,N_2791,N_4957);
nor U5276 (N_5276,N_4547,N_2731);
xor U5277 (N_5277,N_3148,N_4481);
or U5278 (N_5278,N_2711,N_2600);
xnor U5279 (N_5279,N_3653,N_3180);
or U5280 (N_5280,N_4581,N_4111);
or U5281 (N_5281,N_3417,N_2520);
or U5282 (N_5282,N_4984,N_3874);
nand U5283 (N_5283,N_3147,N_4171);
and U5284 (N_5284,N_3322,N_3960);
xnor U5285 (N_5285,N_3845,N_2730);
nand U5286 (N_5286,N_3054,N_3203);
nor U5287 (N_5287,N_3102,N_4472);
nor U5288 (N_5288,N_4246,N_4777);
nand U5289 (N_5289,N_3758,N_3103);
and U5290 (N_5290,N_3290,N_3585);
and U5291 (N_5291,N_3275,N_3077);
nand U5292 (N_5292,N_2881,N_3100);
or U5293 (N_5293,N_3508,N_3765);
xor U5294 (N_5294,N_4147,N_4683);
and U5295 (N_5295,N_4434,N_2980);
and U5296 (N_5296,N_2725,N_2622);
nand U5297 (N_5297,N_3941,N_2903);
xnor U5298 (N_5298,N_4602,N_4491);
xnor U5299 (N_5299,N_3214,N_3950);
or U5300 (N_5300,N_3153,N_2795);
nand U5301 (N_5301,N_3437,N_3518);
nor U5302 (N_5302,N_4450,N_3996);
nand U5303 (N_5303,N_4837,N_3376);
nand U5304 (N_5304,N_4610,N_3041);
nor U5305 (N_5305,N_2539,N_3910);
or U5306 (N_5306,N_4185,N_4458);
xor U5307 (N_5307,N_2991,N_4215);
and U5308 (N_5308,N_3902,N_4817);
nand U5309 (N_5309,N_4336,N_4688);
nor U5310 (N_5310,N_4502,N_3625);
or U5311 (N_5311,N_3481,N_4868);
nand U5312 (N_5312,N_4794,N_3473);
nor U5313 (N_5313,N_4924,N_3792);
xnor U5314 (N_5314,N_3860,N_4954);
or U5315 (N_5315,N_3414,N_3712);
nor U5316 (N_5316,N_3745,N_3654);
or U5317 (N_5317,N_3659,N_2768);
and U5318 (N_5318,N_4949,N_2758);
xor U5319 (N_5319,N_2678,N_3171);
nand U5320 (N_5320,N_3827,N_4863);
or U5321 (N_5321,N_2992,N_3630);
or U5322 (N_5322,N_3907,N_3420);
nor U5323 (N_5323,N_3166,N_2797);
xnor U5324 (N_5324,N_3040,N_4951);
and U5325 (N_5325,N_4200,N_4325);
or U5326 (N_5326,N_3130,N_2592);
xor U5327 (N_5327,N_3606,N_3844);
or U5328 (N_5328,N_2999,N_3380);
xnor U5329 (N_5329,N_4121,N_2727);
nand U5330 (N_5330,N_3052,N_4266);
or U5331 (N_5331,N_4057,N_3651);
nand U5332 (N_5332,N_3149,N_2863);
nand U5333 (N_5333,N_4239,N_3773);
nor U5334 (N_5334,N_3973,N_4154);
and U5335 (N_5335,N_4881,N_3464);
xnor U5336 (N_5336,N_4233,N_4739);
or U5337 (N_5337,N_4499,N_4651);
xnor U5338 (N_5338,N_2806,N_2516);
and U5339 (N_5339,N_3885,N_3762);
xnor U5340 (N_5340,N_4591,N_4321);
or U5341 (N_5341,N_4682,N_4208);
xnor U5342 (N_5342,N_3239,N_3356);
nand U5343 (N_5343,N_3312,N_2603);
and U5344 (N_5344,N_3434,N_3047);
nand U5345 (N_5345,N_4229,N_3378);
or U5346 (N_5346,N_2579,N_4758);
nand U5347 (N_5347,N_2670,N_4299);
nor U5348 (N_5348,N_3426,N_3639);
xor U5349 (N_5349,N_3779,N_2508);
and U5350 (N_5350,N_3726,N_4552);
or U5351 (N_5351,N_3947,N_4997);
or U5352 (N_5352,N_4440,N_4252);
xnor U5353 (N_5353,N_3471,N_3008);
xor U5354 (N_5354,N_4406,N_2675);
nand U5355 (N_5355,N_3351,N_3364);
or U5356 (N_5356,N_3511,N_3285);
nor U5357 (N_5357,N_3234,N_3441);
nor U5358 (N_5358,N_2996,N_2817);
xnor U5359 (N_5359,N_3456,N_3491);
nand U5360 (N_5360,N_3488,N_2612);
or U5361 (N_5361,N_4882,N_3046);
nand U5362 (N_5362,N_4617,N_2642);
or U5363 (N_5363,N_3397,N_3365);
or U5364 (N_5364,N_3278,N_3789);
nor U5365 (N_5365,N_4520,N_3271);
xnor U5366 (N_5366,N_3806,N_4383);
nor U5367 (N_5367,N_2777,N_2716);
and U5368 (N_5368,N_2982,N_3815);
nor U5369 (N_5369,N_4840,N_3986);
and U5370 (N_5370,N_3255,N_4720);
and U5371 (N_5371,N_4062,N_3967);
or U5372 (N_5372,N_3589,N_2858);
or U5373 (N_5373,N_2884,N_4589);
nor U5374 (N_5374,N_4193,N_3281);
and U5375 (N_5375,N_3782,N_3440);
and U5376 (N_5376,N_2764,N_4907);
xor U5377 (N_5377,N_4083,N_3160);
and U5378 (N_5378,N_4324,N_3412);
nand U5379 (N_5379,N_4059,N_3649);
or U5380 (N_5380,N_4084,N_3859);
xnor U5381 (N_5381,N_4876,N_3185);
nand U5382 (N_5382,N_4684,N_2507);
nor U5383 (N_5383,N_3097,N_2500);
or U5384 (N_5384,N_3951,N_3731);
nand U5385 (N_5385,N_3825,N_4931);
nor U5386 (N_5386,N_2745,N_4349);
xor U5387 (N_5387,N_4426,N_4715);
or U5388 (N_5388,N_4355,N_3221);
and U5389 (N_5389,N_4255,N_2569);
and U5390 (N_5390,N_3489,N_3189);
nor U5391 (N_5391,N_2986,N_3573);
and U5392 (N_5392,N_4369,N_2781);
and U5393 (N_5393,N_3723,N_4826);
or U5394 (N_5394,N_2829,N_2660);
xnor U5395 (N_5395,N_3525,N_4232);
or U5396 (N_5396,N_4960,N_3652);
nor U5397 (N_5397,N_3124,N_4754);
and U5398 (N_5398,N_3167,N_4363);
nand U5399 (N_5399,N_3522,N_3870);
nand U5400 (N_5400,N_2624,N_4917);
nand U5401 (N_5401,N_3512,N_4854);
or U5402 (N_5402,N_3595,N_2598);
nor U5403 (N_5403,N_4357,N_4635);
and U5404 (N_5404,N_3016,N_4460);
or U5405 (N_5405,N_3942,N_2519);
nor U5406 (N_5406,N_4021,N_4397);
nor U5407 (N_5407,N_4328,N_4846);
nor U5408 (N_5408,N_2788,N_2898);
nor U5409 (N_5409,N_3470,N_2746);
nand U5410 (N_5410,N_3269,N_4466);
nor U5411 (N_5411,N_2887,N_4222);
nor U5412 (N_5412,N_2873,N_3999);
or U5413 (N_5413,N_3940,N_4633);
nand U5414 (N_5414,N_3517,N_3927);
or U5415 (N_5415,N_4112,N_2875);
or U5416 (N_5416,N_3381,N_2894);
or U5417 (N_5417,N_3120,N_4705);
nor U5418 (N_5418,N_3753,N_4961);
and U5419 (N_5419,N_2591,N_3498);
nand U5420 (N_5420,N_3868,N_4091);
nand U5421 (N_5421,N_4801,N_4430);
nor U5422 (N_5422,N_2733,N_4785);
or U5423 (N_5423,N_3816,N_4756);
or U5424 (N_5424,N_3747,N_4967);
xnor U5425 (N_5425,N_4751,N_4717);
nor U5426 (N_5426,N_3890,N_2862);
xor U5427 (N_5427,N_3929,N_2835);
and U5428 (N_5428,N_3528,N_4749);
nand U5429 (N_5429,N_3643,N_2538);
xor U5430 (N_5430,N_2827,N_4314);
or U5431 (N_5431,N_2895,N_4032);
nand U5432 (N_5432,N_3028,N_3607);
or U5433 (N_5433,N_4672,N_2893);
and U5434 (N_5434,N_3964,N_2528);
and U5435 (N_5435,N_4431,N_4908);
and U5436 (N_5436,N_4987,N_3391);
and U5437 (N_5437,N_4276,N_4911);
nor U5438 (N_5438,N_3957,N_2521);
or U5439 (N_5439,N_4307,N_3081);
nor U5440 (N_5440,N_4290,N_4784);
nand U5441 (N_5441,N_4251,N_3039);
xor U5442 (N_5442,N_4962,N_4774);
xnor U5443 (N_5443,N_3195,N_3229);
nor U5444 (N_5444,N_2821,N_3068);
and U5445 (N_5445,N_3219,N_3276);
xnor U5446 (N_5446,N_3107,N_3225);
or U5447 (N_5447,N_3329,N_4654);
or U5448 (N_5448,N_3847,N_4337);
or U5449 (N_5449,N_4625,N_3136);
and U5450 (N_5450,N_4927,N_4204);
or U5451 (N_5451,N_4417,N_4741);
nand U5452 (N_5452,N_4410,N_3178);
nand U5453 (N_5453,N_4339,N_4085);
and U5454 (N_5454,N_4067,N_2566);
or U5455 (N_5455,N_3310,N_3627);
and U5456 (N_5456,N_3159,N_3419);
or U5457 (N_5457,N_4242,N_4956);
nor U5458 (N_5458,N_4407,N_4131);
nand U5459 (N_5459,N_2985,N_4323);
and U5460 (N_5460,N_4898,N_3480);
xor U5461 (N_5461,N_4079,N_3396);
or U5462 (N_5462,N_4897,N_4302);
xnor U5463 (N_5463,N_3953,N_3023);
xor U5464 (N_5464,N_2594,N_2611);
xor U5465 (N_5465,N_2595,N_2641);
and U5466 (N_5466,N_3861,N_4451);
nand U5467 (N_5467,N_2537,N_3257);
xnor U5468 (N_5468,N_4503,N_3085);
xor U5469 (N_5469,N_3836,N_2646);
and U5470 (N_5470,N_4175,N_3067);
nand U5471 (N_5471,N_3176,N_2586);
nor U5472 (N_5472,N_3140,N_4585);
or U5473 (N_5473,N_3193,N_3479);
and U5474 (N_5474,N_4033,N_4783);
xor U5475 (N_5475,N_2964,N_4165);
and U5476 (N_5476,N_3475,N_3172);
or U5477 (N_5477,N_4146,N_3249);
or U5478 (N_5478,N_3795,N_2601);
xor U5479 (N_5479,N_2721,N_2661);
nor U5480 (N_5480,N_3900,N_3638);
xor U5481 (N_5481,N_4090,N_2937);
xnor U5482 (N_5482,N_2948,N_4380);
nand U5483 (N_5483,N_2584,N_4468);
nand U5484 (N_5484,N_4540,N_3010);
xnor U5485 (N_5485,N_4768,N_4706);
and U5486 (N_5486,N_4933,N_2550);
or U5487 (N_5487,N_3551,N_2608);
and U5488 (N_5488,N_3812,N_3680);
nor U5489 (N_5489,N_4518,N_4671);
nor U5490 (N_5490,N_3824,N_3596);
and U5491 (N_5491,N_4657,N_3808);
or U5492 (N_5492,N_3003,N_3065);
nand U5493 (N_5493,N_3494,N_2686);
or U5494 (N_5494,N_4640,N_4545);
xor U5495 (N_5495,N_4108,N_3640);
or U5496 (N_5496,N_3822,N_4202);
nor U5497 (N_5497,N_4028,N_2939);
xor U5498 (N_5498,N_4143,N_3015);
or U5499 (N_5499,N_3132,N_3954);
nor U5500 (N_5500,N_4105,N_3987);
and U5501 (N_5501,N_3615,N_2688);
nand U5502 (N_5502,N_4767,N_2943);
and U5503 (N_5503,N_4081,N_4480);
and U5504 (N_5504,N_4478,N_2787);
xor U5505 (N_5505,N_4612,N_2816);
nand U5506 (N_5506,N_2515,N_4990);
nor U5507 (N_5507,N_4919,N_2685);
and U5508 (N_5508,N_3095,N_4020);
nor U5509 (N_5509,N_2548,N_4880);
or U5510 (N_5510,N_4723,N_3216);
and U5511 (N_5511,N_4861,N_2929);
nor U5512 (N_5512,N_3708,N_2847);
xnor U5513 (N_5513,N_3794,N_2749);
nor U5514 (N_5514,N_3620,N_4074);
nand U5515 (N_5515,N_4178,N_3699);
xnor U5516 (N_5516,N_3862,N_2694);
nand U5517 (N_5517,N_3982,N_2867);
xor U5518 (N_5518,N_2854,N_4560);
and U5519 (N_5519,N_2915,N_3352);
or U5520 (N_5520,N_2910,N_3495);
or U5521 (N_5521,N_4332,N_4404);
or U5522 (N_5522,N_2715,N_3260);
nand U5523 (N_5523,N_3074,N_3330);
nor U5524 (N_5524,N_3425,N_3204);
xor U5525 (N_5525,N_4393,N_2617);
and U5526 (N_5526,N_4007,N_4627);
xnor U5527 (N_5527,N_4572,N_3506);
nor U5528 (N_5528,N_3766,N_4524);
nor U5529 (N_5529,N_4123,N_3020);
xnor U5530 (N_5530,N_4249,N_4141);
or U5531 (N_5531,N_3235,N_4196);
xor U5532 (N_5532,N_3552,N_3891);
xor U5533 (N_5533,N_4479,N_3700);
nand U5534 (N_5534,N_4549,N_4331);
or U5535 (N_5535,N_2567,N_4993);
nor U5536 (N_5536,N_4265,N_3969);
or U5537 (N_5537,N_2619,N_3354);
nand U5538 (N_5538,N_4110,N_2517);
nand U5539 (N_5539,N_3838,N_2696);
and U5540 (N_5540,N_4992,N_4972);
or U5541 (N_5541,N_3139,N_3956);
and U5542 (N_5542,N_4319,N_3786);
nand U5543 (N_5543,N_4713,N_3251);
nor U5544 (N_5544,N_2784,N_3811);
xor U5545 (N_5545,N_4095,N_4883);
nor U5546 (N_5546,N_3087,N_3797);
or U5547 (N_5547,N_2917,N_4303);
and U5548 (N_5548,N_2973,N_2583);
or U5549 (N_5549,N_3482,N_3353);
xnor U5550 (N_5550,N_3038,N_2852);
xnor U5551 (N_5551,N_3314,N_4569);
nor U5552 (N_5552,N_2811,N_2657);
nand U5553 (N_5553,N_3993,N_4351);
nand U5554 (N_5554,N_4703,N_4834);
nand U5555 (N_5555,N_4588,N_2815);
nor U5556 (N_5556,N_3682,N_4823);
nor U5557 (N_5557,N_2738,N_4210);
or U5558 (N_5558,N_4348,N_4978);
xnor U5559 (N_5559,N_4616,N_3686);
or U5560 (N_5560,N_2790,N_4311);
nand U5561 (N_5561,N_3084,N_4283);
nand U5562 (N_5562,N_4207,N_4743);
nor U5563 (N_5563,N_4099,N_2905);
nor U5564 (N_5564,N_4561,N_2689);
or U5565 (N_5565,N_3979,N_3190);
nor U5566 (N_5566,N_4670,N_4975);
xor U5567 (N_5567,N_2526,N_2628);
nand U5568 (N_5568,N_4999,N_2860);
xor U5569 (N_5569,N_3327,N_3922);
nand U5570 (N_5570,N_4010,N_4162);
xor U5571 (N_5571,N_3864,N_2704);
xnor U5572 (N_5572,N_4398,N_4008);
xor U5573 (N_5573,N_4976,N_4273);
xnor U5574 (N_5574,N_3558,N_4691);
xor U5575 (N_5575,N_4879,N_2921);
xnor U5576 (N_5576,N_4375,N_4170);
nand U5577 (N_5577,N_2623,N_2773);
nand U5578 (N_5578,N_4391,N_4965);
nor U5579 (N_5579,N_2969,N_4579);
or U5580 (N_5580,N_4145,N_2869);
and U5581 (N_5581,N_3059,N_4513);
and U5582 (N_5582,N_3970,N_3857);
nor U5583 (N_5583,N_2502,N_3541);
xor U5584 (N_5584,N_3886,N_2722);
xnor U5585 (N_5585,N_4977,N_3678);
or U5586 (N_5586,N_2525,N_3660);
or U5587 (N_5587,N_4345,N_4501);
and U5588 (N_5588,N_2695,N_4847);
nor U5589 (N_5589,N_4464,N_2631);
xnor U5590 (N_5590,N_4923,N_2638);
or U5591 (N_5591,N_2532,N_4268);
nand U5592 (N_5592,N_3372,N_3608);
xor U5593 (N_5593,N_3066,N_3586);
nand U5594 (N_5594,N_4469,N_2785);
nand U5595 (N_5595,N_3398,N_4755);
or U5596 (N_5596,N_3533,N_2635);
nand U5597 (N_5597,N_3198,N_3336);
nor U5598 (N_5598,N_2807,N_3741);
nor U5599 (N_5599,N_2720,N_4746);
or U5600 (N_5600,N_2718,N_3409);
nor U5601 (N_5601,N_3633,N_4077);
or U5602 (N_5602,N_2945,N_4554);
and U5603 (N_5603,N_4514,N_4172);
or U5604 (N_5604,N_3487,N_3856);
or U5605 (N_5605,N_3648,N_3706);
nand U5606 (N_5606,N_3974,N_3711);
or U5607 (N_5607,N_4092,N_4615);
nand U5608 (N_5608,N_3134,N_4029);
nor U5609 (N_5609,N_4026,N_2958);
nor U5610 (N_5610,N_4403,N_4394);
and U5611 (N_5611,N_4690,N_4361);
or U5612 (N_5612,N_3734,N_4069);
or U5613 (N_5613,N_3963,N_2581);
xnor U5614 (N_5614,N_3618,N_3553);
or U5615 (N_5615,N_3240,N_3184);
xor U5616 (N_5616,N_4996,N_4326);
and U5617 (N_5617,N_4181,N_3549);
nor U5618 (N_5618,N_2859,N_4624);
xnor U5619 (N_5619,N_4129,N_4203);
or U5620 (N_5620,N_4382,N_3879);
nor U5621 (N_5621,N_3671,N_3021);
xnor U5622 (N_5622,N_3035,N_3692);
xnor U5623 (N_5623,N_3127,N_3368);
nor U5624 (N_5624,N_4291,N_2935);
xor U5625 (N_5625,N_3903,N_4634);
nor U5626 (N_5626,N_2665,N_3740);
and U5627 (N_5627,N_3292,N_3914);
nand U5628 (N_5628,N_4770,N_4971);
or U5629 (N_5629,N_4820,N_3767);
xnor U5630 (N_5630,N_3177,N_4875);
or U5631 (N_5631,N_4214,N_4666);
and U5632 (N_5632,N_3086,N_4487);
xor U5633 (N_5633,N_4446,N_2931);
nand U5634 (N_5634,N_4852,N_4821);
xnor U5635 (N_5635,N_4721,N_4680);
and U5636 (N_5636,N_3701,N_2902);
or U5637 (N_5637,N_3892,N_4004);
xnor U5638 (N_5638,N_2831,N_4712);
nand U5639 (N_5639,N_3415,N_3273);
and U5640 (N_5640,N_4630,N_2900);
or U5641 (N_5641,N_4947,N_3113);
xnor U5642 (N_5642,N_2602,N_3472);
or U5643 (N_5643,N_3218,N_3359);
or U5644 (N_5644,N_4733,N_3129);
or U5645 (N_5645,N_4457,N_4805);
xor U5646 (N_5646,N_4632,N_3770);
or U5647 (N_5647,N_3496,N_3295);
or U5648 (N_5648,N_4922,N_3256);
nand U5649 (N_5649,N_4150,N_4221);
or U5650 (N_5650,N_3975,N_3500);
nand U5651 (N_5651,N_3875,N_2963);
nand U5652 (N_5652,N_4132,N_3577);
xor U5653 (N_5653,N_3138,N_4135);
or U5654 (N_5654,N_4824,N_2697);
and U5655 (N_5655,N_2988,N_3252);
or U5656 (N_5656,N_2809,N_2967);
nand U5657 (N_5657,N_3887,N_3405);
and U5658 (N_5658,N_2926,N_3729);
nor U5659 (N_5659,N_2663,N_2848);
or U5660 (N_5660,N_4568,N_3849);
nor U5661 (N_5661,N_3450,N_3501);
nor U5662 (N_5662,N_4659,N_2892);
and U5663 (N_5663,N_3502,N_2613);
or U5664 (N_5664,N_4187,N_3333);
nor U5665 (N_5665,N_3801,N_2983);
or U5666 (N_5666,N_4894,N_4765);
xor U5667 (N_5667,N_2552,N_4198);
nand U5668 (N_5668,N_4726,N_4988);
or U5669 (N_5669,N_4614,N_2671);
or U5670 (N_5670,N_4769,N_4153);
and U5671 (N_5671,N_4211,N_3277);
nor U5672 (N_5672,N_3191,N_4374);
and U5673 (N_5673,N_4736,N_3695);
nand U5674 (N_5674,N_4356,N_4298);
or U5675 (N_5675,N_2593,N_4704);
and U5676 (N_5676,N_3666,N_2748);
nor U5677 (N_5677,N_3780,N_3636);
xnor U5678 (N_5678,N_4329,N_4728);
xor U5679 (N_5679,N_3613,N_2580);
nor U5680 (N_5680,N_4613,N_2683);
nand U5681 (N_5681,N_2972,N_2677);
or U5682 (N_5682,N_2736,N_3056);
or U5683 (N_5683,N_4015,N_3367);
nand U5684 (N_5684,N_3645,N_4841);
and U5685 (N_5685,N_3288,N_3122);
nand U5686 (N_5686,N_4168,N_4448);
nand U5687 (N_5687,N_4293,N_4040);
and U5688 (N_5688,N_3265,N_4573);
and U5689 (N_5689,N_2565,N_2504);
and U5690 (N_5690,N_3298,N_3990);
xor U5691 (N_5691,N_3598,N_4045);
and U5692 (N_5692,N_3800,N_3539);
xnor U5693 (N_5693,N_3813,N_3032);
or U5694 (N_5694,N_4648,N_4159);
xor U5695 (N_5695,N_3732,N_3566);
nor U5696 (N_5696,N_4189,N_4260);
nand U5697 (N_5697,N_3486,N_4201);
nor U5698 (N_5698,N_3446,N_4096);
or U5699 (N_5699,N_3784,N_4906);
and U5700 (N_5700,N_3548,N_3211);
nor U5701 (N_5701,N_3253,N_3452);
and U5702 (N_5702,N_2668,N_4485);
or U5703 (N_5703,N_3427,N_3670);
xor U5704 (N_5704,N_2658,N_3604);
xor U5705 (N_5705,N_4070,N_4019);
xor U5706 (N_5706,N_3580,N_3461);
and U5707 (N_5707,N_3283,N_4660);
xor U5708 (N_5708,N_4047,N_3984);
nor U5709 (N_5709,N_4258,N_3478);
and U5710 (N_5710,N_3280,N_4508);
or U5711 (N_5711,N_4504,N_4710);
nor U5712 (N_5712,N_4217,N_3128);
xor U5713 (N_5713,N_4586,N_4791);
and U5714 (N_5714,N_3946,N_3965);
nor U5715 (N_5715,N_3082,N_3099);
and U5716 (N_5716,N_2757,N_3936);
or U5717 (N_5717,N_4304,N_4687);
or U5718 (N_5718,N_2684,N_3968);
or U5719 (N_5719,N_4813,N_2997);
or U5720 (N_5720,N_3981,N_3848);
and U5721 (N_5721,N_3338,N_4762);
or U5722 (N_5722,N_3750,N_4685);
xnor U5723 (N_5723,N_3730,N_4199);
nand U5724 (N_5724,N_2590,N_2632);
xnor U5725 (N_5725,N_2672,N_2882);
and U5726 (N_5726,N_4275,N_3510);
nor U5727 (N_5727,N_3901,N_3443);
nor U5728 (N_5728,N_3719,N_3157);
or U5729 (N_5729,N_2556,N_3145);
and U5730 (N_5730,N_3647,N_4322);
xnor U5731 (N_5731,N_3702,N_3109);
nor U5732 (N_5732,N_3268,N_4930);
or U5733 (N_5733,N_3532,N_3004);
nand U5734 (N_5734,N_3600,N_2870);
xnor U5735 (N_5735,N_2928,N_4161);
or U5736 (N_5736,N_3629,N_3665);
or U5737 (N_5737,N_3799,N_4555);
and U5738 (N_5738,N_4895,N_2653);
nand U5739 (N_5739,N_3309,N_4166);
xor U5740 (N_5740,N_4623,N_3436);
and U5741 (N_5741,N_2759,N_4439);
xnor U5742 (N_5742,N_3683,N_2942);
nand U5743 (N_5743,N_4163,N_3400);
or U5744 (N_5744,N_4018,N_4689);
and U5745 (N_5745,N_3022,N_2693);
xor U5746 (N_5746,N_4435,N_4419);
xnor U5747 (N_5747,N_3394,N_2834);
and U5748 (N_5748,N_3404,N_2626);
nand U5749 (N_5749,N_3943,N_3293);
xor U5750 (N_5750,N_4796,N_4456);
or U5751 (N_5751,N_3326,N_4118);
or U5752 (N_5752,N_3855,N_2761);
xor U5753 (N_5753,N_3311,N_3401);
nor U5754 (N_5754,N_2776,N_3897);
nand U5755 (N_5755,N_2837,N_4012);
nor U5756 (N_5756,N_4985,N_4952);
or U5757 (N_5757,N_3194,N_2850);
nor U5758 (N_5758,N_4184,N_2762);
nand U5759 (N_5759,N_4887,N_3119);
nor U5760 (N_5760,N_2789,N_2753);
nor U5761 (N_5761,N_4653,N_2651);
xnor U5762 (N_5762,N_4583,N_4904);
and U5763 (N_5763,N_4449,N_2960);
xor U5764 (N_5764,N_4388,N_3018);
and U5765 (N_5765,N_2794,N_4031);
or U5766 (N_5766,N_4871,N_3096);
nand U5767 (N_5767,N_4958,N_2801);
and U5768 (N_5768,N_3916,N_3294);
or U5769 (N_5769,N_4078,N_3614);
and U5770 (N_5770,N_3877,N_2553);
and U5771 (N_5771,N_4644,N_4400);
nor U5772 (N_5772,N_3460,N_4793);
nand U5773 (N_5773,N_4050,N_4271);
xor U5774 (N_5774,N_4461,N_3561);
xnor U5775 (N_5775,N_2843,N_2878);
and U5776 (N_5776,N_3089,N_3876);
nand U5777 (N_5777,N_3112,N_3014);
nand U5778 (N_5778,N_3781,N_4521);
nand U5779 (N_5779,N_4647,N_4309);
or U5780 (N_5780,N_4212,N_3407);
and U5781 (N_5781,N_3045,N_4452);
nor U5782 (N_5782,N_2615,N_2640);
xnor U5783 (N_5783,N_3674,N_3108);
xnor U5784 (N_5784,N_3335,N_4411);
nor U5785 (N_5785,N_4853,N_2656);
nand U5786 (N_5786,N_4790,N_4437);
nor U5787 (N_5787,N_4590,N_4106);
and U5788 (N_5788,N_4565,N_4664);
nand U5789 (N_5789,N_3143,N_4433);
and U5790 (N_5790,N_4515,N_3641);
or U5791 (N_5791,N_4582,N_2880);
xnor U5792 (N_5792,N_3291,N_4247);
nor U5793 (N_5793,N_3101,N_3944);
nor U5794 (N_5794,N_4998,N_3044);
and U5795 (N_5795,N_3332,N_4788);
xor U5796 (N_5796,N_3704,N_2793);
nor U5797 (N_5797,N_4139,N_2953);
nor U5798 (N_5798,N_2523,N_4916);
nand U5799 (N_5799,N_4292,N_4983);
nand U5800 (N_5800,N_3748,N_3677);
nor U5801 (N_5801,N_4353,N_3632);
and U5802 (N_5802,N_3053,N_2534);
xor U5803 (N_5803,N_4156,N_4969);
nand U5804 (N_5804,N_2907,N_3621);
nor U5805 (N_5805,N_4396,N_4297);
nand U5806 (N_5806,N_3881,N_4731);
xnor U5807 (N_5807,N_4596,N_3262);
nor U5808 (N_5808,N_4986,N_4637);
nor U5809 (N_5809,N_4606,N_3599);
nor U5810 (N_5810,N_3878,N_3057);
and U5811 (N_5811,N_4009,N_3616);
nand U5812 (N_5812,N_4489,N_4060);
and U5813 (N_5813,N_3718,N_3554);
and U5814 (N_5814,N_4753,N_3775);
and U5815 (N_5815,N_2934,N_2587);
nor U5816 (N_5816,N_3264,N_4537);
nor U5817 (N_5817,N_4340,N_2904);
and U5818 (N_5818,N_4392,N_2574);
and U5819 (N_5819,N_4607,N_2877);
and U5820 (N_5820,N_4937,N_3503);
and U5821 (N_5821,N_4263,N_4315);
and U5822 (N_5822,N_4527,N_4000);
xor U5823 (N_5823,N_3006,N_4711);
xnor U5824 (N_5824,N_3299,N_2633);
and U5825 (N_5825,N_3634,N_3575);
or U5826 (N_5826,N_4044,N_4629);
xnor U5827 (N_5827,N_4905,N_3938);
nor U5828 (N_5828,N_3948,N_4511);
or U5829 (N_5829,N_4277,N_4693);
xor U5830 (N_5830,N_4550,N_4752);
xor U5831 (N_5831,N_3328,N_2786);
xnor U5832 (N_5832,N_2578,N_4120);
xnor U5833 (N_5833,N_2810,N_3962);
or U5834 (N_5834,N_4580,N_4991);
nor U5835 (N_5835,N_4498,N_4802);
nand U5836 (N_5836,N_4335,N_4529);
xnor U5837 (N_5837,N_4158,N_3817);
nand U5838 (N_5838,N_2589,N_3048);
xor U5839 (N_5839,N_3540,N_3321);
nand U5840 (N_5840,N_3601,N_4603);
xnor U5841 (N_5841,N_3408,N_4338);
nor U5842 (N_5842,N_2922,N_4893);
nand U5843 (N_5843,N_3662,N_3609);
and U5844 (N_5844,N_2554,N_3924);
and U5845 (N_5845,N_2919,N_4301);
nand U5846 (N_5846,N_3791,N_4484);
or U5847 (N_5847,N_2560,N_3839);
and U5848 (N_5848,N_4248,N_2923);
and U5849 (N_5849,N_4850,N_3011);
nor U5850 (N_5850,N_4835,N_3466);
nor U5851 (N_5851,N_3164,N_4030);
nand U5852 (N_5852,N_4223,N_4858);
nor U5853 (N_5853,N_3421,N_3156);
nand U5854 (N_5854,N_3567,N_3590);
nand U5855 (N_5855,N_4128,N_2855);
nand U5856 (N_5856,N_2636,N_4218);
nor U5857 (N_5857,N_2542,N_3743);
and U5858 (N_5858,N_3423,N_4101);
nand U5859 (N_5859,N_4488,N_4867);
and U5860 (N_5860,N_3809,N_3663);
xor U5861 (N_5861,N_3774,N_4725);
nor U5862 (N_5862,N_2514,N_2961);
xnor U5863 (N_5863,N_3165,N_4558);
or U5864 (N_5864,N_4412,N_3141);
or U5865 (N_5865,N_2766,N_3432);
and U5866 (N_5866,N_3685,N_3587);
or U5867 (N_5867,N_4320,N_3939);
nand U5868 (N_5868,N_4240,N_3331);
nand U5869 (N_5869,N_3534,N_4886);
or U5870 (N_5870,N_3888,N_3937);
xnor U5871 (N_5871,N_2729,N_4422);
xnor U5872 (N_5872,N_4541,N_3790);
or U5873 (N_5873,N_3661,N_3069);
nand U5874 (N_5874,N_3284,N_2621);
xnor U5875 (N_5875,N_3631,N_3842);
xor U5876 (N_5876,N_4786,N_3894);
xor U5877 (N_5877,N_3050,N_4151);
or U5878 (N_5878,N_2645,N_4652);
or U5879 (N_5879,N_2629,N_2549);
and U5880 (N_5880,N_4226,N_3183);
or U5881 (N_5881,N_3123,N_4465);
xnor U5882 (N_5882,N_2783,N_3182);
nand U5883 (N_5883,N_3687,N_3413);
or U5884 (N_5884,N_4597,N_3772);
nor U5885 (N_5885,N_3672,N_2866);
nand U5886 (N_5886,N_2654,N_2828);
and U5887 (N_5887,N_3934,N_3418);
nor U5888 (N_5888,N_4679,N_4857);
xor U5889 (N_5889,N_3072,N_4546);
xor U5890 (N_5890,N_2944,N_2680);
and U5891 (N_5891,N_2778,N_3430);
nand U5892 (N_5892,N_3137,N_4702);
and U5893 (N_5893,N_3049,N_2702);
or U5894 (N_5894,N_2836,N_3545);
nor U5895 (N_5895,N_3896,N_4346);
nand U5896 (N_5896,N_3515,N_2818);
nor U5897 (N_5897,N_3698,N_4532);
xnor U5898 (N_5898,N_4668,N_3345);
or U5899 (N_5899,N_4605,N_4269);
nor U5900 (N_5900,N_3751,N_4686);
and U5901 (N_5901,N_3243,N_3320);
nand U5902 (N_5902,N_3819,N_3433);
nor U5903 (N_5903,N_3173,N_3926);
xor U5904 (N_5904,N_2938,N_4856);
and U5905 (N_5905,N_4525,N_4636);
nor U5906 (N_5906,N_4860,N_3572);
xor U5907 (N_5907,N_3591,N_3820);
nor U5908 (N_5908,N_4114,N_3377);
and U5909 (N_5909,N_4534,N_2839);
xor U5910 (N_5910,N_3476,N_3542);
or U5911 (N_5911,N_3742,N_3406);
nor U5912 (N_5912,N_3027,N_3831);
and U5913 (N_5913,N_4839,N_3319);
and U5914 (N_5914,N_3092,N_4938);
nand U5915 (N_5915,N_3230,N_3455);
nand U5916 (N_5916,N_2501,N_4535);
and U5917 (N_5917,N_3958,N_4011);
and U5918 (N_5918,N_2743,N_3588);
or U5919 (N_5919,N_2719,N_3248);
nand U5920 (N_5920,N_3579,N_3626);
nand U5921 (N_5921,N_4284,N_3444);
nor U5922 (N_5922,N_4716,N_4133);
nand U5923 (N_5923,N_2840,N_2979);
xnor U5924 (N_5924,N_4420,N_4136);
nand U5925 (N_5925,N_2544,N_2540);
and U5926 (N_5926,N_3267,N_4780);
nor U5927 (N_5927,N_4395,N_3526);
nand U5928 (N_5928,N_3785,N_2648);
or U5929 (N_5929,N_3752,N_4557);
nor U5930 (N_5930,N_4126,N_2822);
nor U5931 (N_5931,N_4973,N_3339);
or U5932 (N_5932,N_2888,N_2545);
nand U5933 (N_5933,N_2576,N_3527);
nor U5934 (N_5934,N_4216,N_3720);
or U5935 (N_5935,N_3594,N_3576);
xnor U5936 (N_5936,N_2883,N_3673);
nand U5937 (N_5937,N_4342,N_3846);
nor U5938 (N_5938,N_4243,N_4425);
xnor U5939 (N_5939,N_3571,N_4089);
or U5940 (N_5940,N_4264,N_3142);
or U5941 (N_5941,N_4843,N_3037);
nand U5942 (N_5942,N_4814,N_4130);
or U5943 (N_5943,N_2968,N_4830);
xnor U5944 (N_5944,N_3581,N_4942);
nand U5945 (N_5945,N_3272,N_4803);
nor U5946 (N_5946,N_4742,N_2976);
xor U5947 (N_5947,N_2864,N_3226);
nor U5948 (N_5948,N_3245,N_4526);
and U5949 (N_5949,N_4076,N_4186);
or U5950 (N_5950,N_4209,N_4098);
and U5951 (N_5951,N_3302,N_4598);
and U5952 (N_5952,N_4968,N_3324);
xnor U5953 (N_5953,N_4225,N_3841);
and U5954 (N_5954,N_4160,N_3557);
nand U5955 (N_5955,N_4718,N_3612);
xor U5956 (N_5956,N_4873,N_4475);
nand U5957 (N_5957,N_2775,N_4442);
nor U5958 (N_5958,N_3375,N_4730);
and U5959 (N_5959,N_3725,N_3402);
or U5960 (N_5960,N_4600,N_4628);
or U5961 (N_5961,N_4709,N_2751);
nor U5962 (N_5962,N_2610,N_4312);
and U5963 (N_5963,N_4795,N_2690);
or U5964 (N_5964,N_3349,N_3215);
nor U5965 (N_5965,N_3385,N_4455);
nand U5966 (N_5966,N_3009,N_4424);
and U5967 (N_5967,N_4500,N_3025);
nor U5968 (N_5968,N_4497,N_4194);
nor U5969 (N_5969,N_4865,N_3544);
xor U5970 (N_5970,N_4982,N_4799);
nor U5971 (N_5971,N_3448,N_3793);
and U5972 (N_5972,N_2987,N_2742);
nand U5973 (N_5973,N_4034,N_4918);
or U5974 (N_5974,N_4378,N_4646);
xor U5975 (N_5975,N_3736,N_3174);
xor U5976 (N_5976,N_3031,N_3703);
and U5977 (N_5977,N_4729,N_3237);
xor U5978 (N_5978,N_3858,N_3696);
and U5979 (N_5979,N_4539,N_4921);
and U5980 (N_5980,N_4415,N_2872);
nand U5981 (N_5981,N_3930,N_3029);
nor U5982 (N_5982,N_4950,N_3716);
nor U5983 (N_5983,N_4944,N_2536);
or U5984 (N_5984,N_4272,N_3911);
or U5985 (N_5985,N_2936,N_2609);
nand U5986 (N_5986,N_3832,N_3778);
xor U5987 (N_5987,N_3210,N_4051);
or U5988 (N_5988,N_3739,N_2974);
nor U5989 (N_5989,N_2970,N_3188);
xnor U5990 (N_5990,N_2724,N_3296);
and U5991 (N_5991,N_3071,N_4100);
nor U5992 (N_5992,N_3286,N_2914);
or U5993 (N_5993,N_4023,N_3175);
nand U5994 (N_5994,N_4673,N_4622);
xnor U5995 (N_5995,N_3091,N_3872);
xor U5996 (N_5996,N_3325,N_2962);
xor U5997 (N_5997,N_4477,N_4017);
nor U5998 (N_5998,N_3935,N_3854);
or U5999 (N_5999,N_4474,N_4279);
nor U6000 (N_6000,N_4330,N_4655);
xor U6001 (N_6001,N_3523,N_4822);
nor U6002 (N_6002,N_3297,N_4888);
nor U6003 (N_6003,N_4553,N_4533);
xnor U6004 (N_6004,N_3051,N_4492);
nand U6005 (N_6005,N_4509,N_3477);
and U6006 (N_6006,N_4955,N_3925);
xor U6007 (N_6007,N_4831,N_3850);
nand U6008 (N_6008,N_4116,N_4989);
and U6009 (N_6009,N_4959,N_4800);
nor U6010 (N_6010,N_4570,N_3274);
and U6011 (N_6011,N_4862,N_2679);
nor U6012 (N_6012,N_4696,N_2760);
nor U6013 (N_6013,N_4381,N_4359);
and U6014 (N_6014,N_4438,N_3555);
and U6015 (N_6015,N_4891,N_2659);
nand U6016 (N_6016,N_3664,N_4176);
and U6017 (N_6017,N_4414,N_2899);
and U6018 (N_6018,N_2792,N_4316);
or U6019 (N_6019,N_4838,N_4389);
or U6020 (N_6020,N_4467,N_4812);
and U6021 (N_6021,N_4697,N_4333);
xor U6022 (N_6022,N_4714,N_3236);
xnor U6023 (N_6023,N_3931,N_4053);
nand U6024 (N_6024,N_4842,N_4675);
nand U6025 (N_6025,N_4516,N_2627);
xnor U6026 (N_6026,N_4362,N_4901);
nand U6027 (N_6027,N_4913,N_3863);
nand U6028 (N_6028,N_3932,N_3744);
and U6029 (N_6029,N_3945,N_4354);
nor U6030 (N_6030,N_3997,N_4517);
and U6031 (N_6031,N_4390,N_4278);
or U6032 (N_6032,N_4177,N_3263);
and U6033 (N_6033,N_3313,N_3196);
nor U6034 (N_6034,N_3492,N_3906);
or U6035 (N_6035,N_2959,N_2703);
or U6036 (N_6036,N_4295,N_2780);
and U6037 (N_6037,N_2849,N_2541);
nor U6038 (N_6038,N_4869,N_3505);
and U6039 (N_6039,N_4832,N_3995);
xnor U6040 (N_6040,N_3168,N_3955);
or U6041 (N_6041,N_4296,N_2754);
or U6042 (N_6042,N_4282,N_3454);
xor U6043 (N_6043,N_4061,N_2723);
nor U6044 (N_6044,N_4416,N_2796);
nand U6045 (N_6045,N_3917,N_3776);
nand U6046 (N_6046,N_4072,N_4182);
or U6047 (N_6047,N_4836,N_3002);
nor U6048 (N_6048,N_4493,N_4638);
nand U6049 (N_6049,N_3668,N_4230);
nor U6050 (N_6050,N_3546,N_3346);
and U6051 (N_6051,N_4192,N_3197);
nand U6052 (N_6052,N_2701,N_3980);
or U6053 (N_6053,N_3676,N_3317);
and U6054 (N_6054,N_3746,N_4157);
nor U6055 (N_6055,N_2741,N_2879);
nand U6056 (N_6056,N_3529,N_4737);
and U6057 (N_6057,N_4732,N_3971);
or U6058 (N_6058,N_4699,N_2647);
nand U6059 (N_6059,N_4747,N_4447);
nor U6060 (N_6060,N_3358,N_3788);
xor U6061 (N_6061,N_4939,N_4903);
or U6062 (N_6062,N_3342,N_3705);
and U6063 (N_6063,N_4429,N_3428);
nor U6064 (N_6064,N_4779,N_3323);
or U6065 (N_6065,N_4512,N_2916);
and U6066 (N_6066,N_4376,N_2782);
nand U6067 (N_6067,N_2637,N_3760);
xor U6068 (N_6068,N_2620,N_4071);
xor U6069 (N_6069,N_4052,N_3835);
nand U6070 (N_6070,N_2920,N_2564);
nand U6071 (N_6071,N_4002,N_4386);
nand U6072 (N_6072,N_4180,N_3728);
and U6073 (N_6073,N_3603,N_2832);
xnor U6074 (N_6074,N_3754,N_3474);
or U6075 (N_6075,N_2950,N_3804);
and U6076 (N_6076,N_3597,N_2820);
and U6077 (N_6077,N_3013,N_4039);
and U6078 (N_6078,N_3192,N_3369);
nand U6079 (N_6079,N_3019,N_3152);
or U6080 (N_6080,N_2533,N_3007);
or U6081 (N_6081,N_4771,N_3090);
xor U6082 (N_6082,N_2940,N_4262);
nand U6083 (N_6083,N_3768,N_3366);
nor U6084 (N_6084,N_4519,N_3913);
nand U6085 (N_6085,N_4082,N_3807);
nand U6086 (N_6086,N_3061,N_3208);
xnor U6087 (N_6087,N_4872,N_3287);
nand U6088 (N_6088,N_2912,N_4358);
nor U6089 (N_6089,N_4231,N_3362);
and U6090 (N_6090,N_4274,N_3080);
nand U6091 (N_6091,N_2667,N_4038);
and U6092 (N_6092,N_2925,N_2728);
or U6093 (N_6093,N_4902,N_3076);
xnor U6094 (N_6094,N_3688,N_2957);
xnor U6095 (N_6095,N_2770,N_2639);
nand U6096 (N_6096,N_4169,N_2995);
nor U6097 (N_6097,N_2771,N_4665);
xnor U6098 (N_6098,N_3650,N_3266);
xnor U6099 (N_6099,N_4042,N_4459);
and U6100 (N_6100,N_2800,N_3075);
and U6101 (N_6101,N_3150,N_4556);
xnor U6102 (N_6102,N_2993,N_3416);
and U6103 (N_6103,N_2712,N_2808);
xnor U6104 (N_6104,N_2505,N_2977);
nor U6105 (N_6105,N_2966,N_2732);
nand U6106 (N_6106,N_4692,N_4066);
nand U6107 (N_6107,N_2597,N_3619);
or U6108 (N_6108,N_4676,N_4782);
xnor U6109 (N_6109,N_2857,N_3985);
nor U6110 (N_6110,N_3871,N_3490);
nor U6111 (N_6111,N_4829,N_3830);
nand U6112 (N_6112,N_3707,N_2713);
and U6113 (N_6113,N_4064,N_4576);
xor U6114 (N_6114,N_3530,N_2799);
nand U6115 (N_6115,N_3463,N_2813);
nor U6116 (N_6116,N_3499,N_4124);
xor U6117 (N_6117,N_3484,N_2876);
xor U6118 (N_6118,N_4662,N_4900);
and U6119 (N_6119,N_4811,N_3535);
or U6120 (N_6120,N_3657,N_4286);
or U6121 (N_6121,N_3560,N_3769);
or U6122 (N_6122,N_3163,N_2649);
nand U6123 (N_6123,N_2691,N_2989);
or U6124 (N_6124,N_3429,N_2666);
xor U6125 (N_6125,N_4775,N_4236);
or U6126 (N_6126,N_2853,N_3722);
nand U6127 (N_6127,N_2885,N_3724);
xor U6128 (N_6128,N_3837,N_4522);
nor U6129 (N_6129,N_2886,N_4365);
or U6130 (N_6130,N_4080,N_2845);
xor U6131 (N_6131,N_3458,N_2599);
or U6132 (N_6132,N_2871,N_4427);
nand U6133 (N_6133,N_3158,N_3131);
nand U6134 (N_6134,N_4055,N_2954);
xor U6135 (N_6135,N_2833,N_3300);
and U6136 (N_6136,N_3344,N_3983);
xnor U6137 (N_6137,N_3516,N_3710);
and U6138 (N_6138,N_4035,N_3242);
and U6139 (N_6139,N_2740,N_2901);
xnor U6140 (N_6140,N_2814,N_3717);
nand U6141 (N_6141,N_3078,N_3209);
nor U6142 (N_6142,N_2747,N_4058);
nand U6143 (N_6143,N_2826,N_4523);
nor U6144 (N_6144,N_4538,N_3270);
nor U6145 (N_6145,N_4384,N_4173);
nand U6146 (N_6146,N_4373,N_3399);
and U6147 (N_6147,N_4797,N_4366);
nand U6148 (N_6148,N_4844,N_3998);
nor U6149 (N_6149,N_4810,N_3959);
and U6150 (N_6150,N_3783,N_4792);
nand U6151 (N_6151,N_4809,N_4352);
xnor U6152 (N_6152,N_3635,N_2692);
xor U6153 (N_6153,N_4806,N_3697);
nor U6154 (N_6154,N_2573,N_3058);
nand U6155 (N_6155,N_3866,N_2965);
nor U6156 (N_6156,N_4761,N_3570);
nand U6157 (N_6157,N_2543,N_2662);
xnor U6158 (N_6158,N_3259,N_4137);
nor U6159 (N_6159,N_3151,N_3449);
nor U6160 (N_6160,N_4347,N_3370);
and U6161 (N_6161,N_4190,N_3154);
nand U6162 (N_6162,N_2949,N_4698);
or U6163 (N_6163,N_4259,N_4372);
nand U6164 (N_6164,N_2823,N_4963);
xnor U6165 (N_6165,N_4639,N_3155);
or U6166 (N_6166,N_3135,N_2984);
nor U6167 (N_6167,N_3755,N_4418);
or U6168 (N_6168,N_4506,N_4421);
nand U6169 (N_6169,N_2625,N_3873);
or U6170 (N_6170,N_4238,N_4409);
nand U6171 (N_6171,N_4620,N_3949);
nand U6172 (N_6172,N_4094,N_4866);
and U6173 (N_6173,N_2570,N_4914);
or U6174 (N_6174,N_3228,N_3447);
xnor U6175 (N_6175,N_4885,N_4727);
nand U6176 (N_6176,N_3439,N_3531);
nor U6177 (N_6177,N_4289,N_3904);
nor U6178 (N_6178,N_4701,N_4661);
nand U6179 (N_6179,N_4473,N_3162);
and U6180 (N_6180,N_3395,N_3179);
xor U6181 (N_6181,N_4599,N_2652);
and U6182 (N_6182,N_4350,N_4313);
and U6183 (N_6183,N_4995,N_3199);
or U6184 (N_6184,N_2767,N_4787);
and U6185 (N_6185,N_2990,N_3079);
xor U6186 (N_6186,N_4402,N_4285);
or U6187 (N_6187,N_3667,N_4980);
xnor U6188 (N_6188,N_3592,N_3111);
nor U6189 (N_6189,N_4444,N_4694);
nand U6190 (N_6190,N_4724,N_3435);
xnor U6191 (N_6191,N_3655,N_4377);
nand U6192 (N_6192,N_4815,N_3905);
and U6193 (N_6193,N_3305,N_3411);
nor U6194 (N_6194,N_3024,N_4789);
nor U6195 (N_6195,N_4399,N_3379);
nand U6196 (N_6196,N_2503,N_3126);
nor U6197 (N_6197,N_2841,N_2630);
nor U6198 (N_6198,N_3563,N_4663);
nor U6199 (N_6199,N_4483,N_3733);
nand U6200 (N_6200,N_3125,N_3247);
nand U6201 (N_6201,N_2561,N_4593);
and U6202 (N_6202,N_3933,N_4912);
or U6203 (N_6203,N_2779,N_4024);
or U6204 (N_6204,N_3853,N_4471);
xnor U6205 (N_6205,N_3304,N_2908);
and U6206 (N_6206,N_4063,N_2687);
nand U6207 (N_6207,N_4798,N_3117);
nand U6208 (N_6208,N_3341,N_4818);
xor U6209 (N_6209,N_3034,N_4087);
xnor U6210 (N_6210,N_3110,N_2513);
and U6211 (N_6211,N_4744,N_2714);
xnor U6212 (N_6212,N_4482,N_4848);
xor U6213 (N_6213,N_4645,N_3098);
or U6214 (N_6214,N_4827,N_4695);
xnor U6215 (N_6215,N_3880,N_2941);
xnor U6216 (N_6216,N_4075,N_4594);
nand U6217 (N_6217,N_4766,N_3593);
xor U6218 (N_6218,N_3064,N_4915);
and U6219 (N_6219,N_2998,N_4681);
nand U6220 (N_6220,N_4650,N_3821);
nand U6221 (N_6221,N_4845,N_2805);
and U6222 (N_6222,N_3343,N_4423);
and U6223 (N_6223,N_2604,N_3347);
xor U6224 (N_6224,N_4048,N_2700);
and U6225 (N_6225,N_2909,N_2577);
or U6226 (N_6226,N_3884,N_3547);
or U6227 (N_6227,N_3062,N_3637);
nand U6228 (N_6228,N_4088,N_3403);
or U6229 (N_6229,N_3289,N_4592);
and U6230 (N_6230,N_4899,N_4979);
nor U6231 (N_6231,N_4174,N_4953);
or U6232 (N_6232,N_4738,N_2551);
nor U6233 (N_6233,N_3713,N_3043);
nor U6234 (N_6234,N_4036,N_2571);
and U6235 (N_6235,N_4658,N_3207);
nand U6236 (N_6236,N_2510,N_4138);
nand U6237 (N_6237,N_4773,N_2838);
or U6238 (N_6238,N_4649,N_4674);
or U6239 (N_6239,N_4155,N_4759);
or U6240 (N_6240,N_4257,N_2765);
or U6241 (N_6241,N_3457,N_4548);
and U6242 (N_6242,N_4220,N_4234);
nor U6243 (N_6243,N_2606,N_2744);
nand U6244 (N_6244,N_3538,N_3562);
nor U6245 (N_6245,N_2819,N_4119);
or U6246 (N_6246,N_3244,N_3972);
nand U6247 (N_6247,N_3556,N_2911);
xnor U6248 (N_6248,N_4748,N_2825);
xnor U6249 (N_6249,N_4213,N_3146);
nor U6250 (N_6250,N_4321,N_3081);
xnor U6251 (N_6251,N_4438,N_3043);
nand U6252 (N_6252,N_3131,N_3682);
xnor U6253 (N_6253,N_4346,N_3649);
nand U6254 (N_6254,N_3275,N_4868);
nand U6255 (N_6255,N_4282,N_2516);
xnor U6256 (N_6256,N_4905,N_4398);
nand U6257 (N_6257,N_2916,N_3747);
nand U6258 (N_6258,N_4996,N_3668);
and U6259 (N_6259,N_3857,N_4426);
nor U6260 (N_6260,N_3018,N_4395);
nor U6261 (N_6261,N_4902,N_4817);
and U6262 (N_6262,N_3567,N_4048);
nand U6263 (N_6263,N_2897,N_4515);
nand U6264 (N_6264,N_3862,N_2708);
or U6265 (N_6265,N_4794,N_2852);
nor U6266 (N_6266,N_2826,N_4046);
xor U6267 (N_6267,N_2517,N_4644);
nand U6268 (N_6268,N_4916,N_4364);
nand U6269 (N_6269,N_3705,N_2898);
nand U6270 (N_6270,N_3398,N_2511);
xnor U6271 (N_6271,N_4685,N_2544);
xnor U6272 (N_6272,N_4283,N_4528);
nor U6273 (N_6273,N_4649,N_4501);
and U6274 (N_6274,N_3887,N_4031);
or U6275 (N_6275,N_4817,N_2936);
nor U6276 (N_6276,N_2748,N_4391);
and U6277 (N_6277,N_3702,N_2553);
xnor U6278 (N_6278,N_3252,N_3374);
nand U6279 (N_6279,N_2678,N_4585);
nor U6280 (N_6280,N_3866,N_2940);
nor U6281 (N_6281,N_4747,N_3537);
nand U6282 (N_6282,N_3490,N_3986);
xnor U6283 (N_6283,N_3319,N_3484);
nand U6284 (N_6284,N_4808,N_4545);
nand U6285 (N_6285,N_4219,N_3023);
xor U6286 (N_6286,N_4347,N_2568);
nand U6287 (N_6287,N_3346,N_3311);
or U6288 (N_6288,N_3731,N_4742);
nor U6289 (N_6289,N_2806,N_3658);
nor U6290 (N_6290,N_2746,N_4079);
nand U6291 (N_6291,N_4817,N_2804);
xnor U6292 (N_6292,N_2856,N_4526);
nand U6293 (N_6293,N_4208,N_4235);
xor U6294 (N_6294,N_4843,N_3752);
nor U6295 (N_6295,N_3550,N_3941);
nor U6296 (N_6296,N_4093,N_4917);
and U6297 (N_6297,N_3120,N_3937);
xnor U6298 (N_6298,N_3909,N_3472);
nand U6299 (N_6299,N_4347,N_4044);
xor U6300 (N_6300,N_4504,N_2526);
or U6301 (N_6301,N_4177,N_2546);
nor U6302 (N_6302,N_4707,N_4128);
and U6303 (N_6303,N_3194,N_2993);
or U6304 (N_6304,N_4509,N_3930);
or U6305 (N_6305,N_4693,N_4304);
nand U6306 (N_6306,N_4144,N_3481);
and U6307 (N_6307,N_4783,N_4037);
nor U6308 (N_6308,N_4057,N_4278);
xnor U6309 (N_6309,N_3629,N_4787);
xor U6310 (N_6310,N_2980,N_3855);
or U6311 (N_6311,N_4633,N_4632);
nor U6312 (N_6312,N_3397,N_4933);
nand U6313 (N_6313,N_3214,N_3510);
or U6314 (N_6314,N_4777,N_3561);
nand U6315 (N_6315,N_3538,N_2799);
and U6316 (N_6316,N_3441,N_3077);
or U6317 (N_6317,N_4728,N_4812);
and U6318 (N_6318,N_3131,N_3403);
nor U6319 (N_6319,N_4232,N_2597);
nor U6320 (N_6320,N_4325,N_2580);
nor U6321 (N_6321,N_4145,N_2873);
or U6322 (N_6322,N_4768,N_3361);
nor U6323 (N_6323,N_4639,N_3256);
xnor U6324 (N_6324,N_4208,N_2995);
and U6325 (N_6325,N_2733,N_2711);
and U6326 (N_6326,N_4786,N_3918);
and U6327 (N_6327,N_2614,N_4603);
or U6328 (N_6328,N_3664,N_2999);
xor U6329 (N_6329,N_3434,N_4150);
and U6330 (N_6330,N_3213,N_4885);
xnor U6331 (N_6331,N_4446,N_3349);
and U6332 (N_6332,N_4971,N_4218);
or U6333 (N_6333,N_3125,N_2868);
or U6334 (N_6334,N_3446,N_4150);
nor U6335 (N_6335,N_2793,N_3968);
nor U6336 (N_6336,N_3155,N_2687);
nand U6337 (N_6337,N_4741,N_4738);
or U6338 (N_6338,N_3598,N_3316);
nor U6339 (N_6339,N_4967,N_3317);
nor U6340 (N_6340,N_4693,N_3364);
nand U6341 (N_6341,N_4240,N_4150);
or U6342 (N_6342,N_3853,N_3190);
nor U6343 (N_6343,N_3928,N_3805);
nor U6344 (N_6344,N_4762,N_3220);
nand U6345 (N_6345,N_3860,N_3141);
xor U6346 (N_6346,N_2768,N_2838);
nor U6347 (N_6347,N_4814,N_4041);
and U6348 (N_6348,N_4789,N_4233);
nand U6349 (N_6349,N_3059,N_4054);
nand U6350 (N_6350,N_4016,N_4317);
nand U6351 (N_6351,N_2710,N_4215);
or U6352 (N_6352,N_3191,N_3335);
nor U6353 (N_6353,N_2670,N_4754);
nand U6354 (N_6354,N_4505,N_4064);
or U6355 (N_6355,N_3754,N_2913);
xnor U6356 (N_6356,N_3847,N_3317);
nor U6357 (N_6357,N_4517,N_3606);
or U6358 (N_6358,N_3710,N_4245);
and U6359 (N_6359,N_3780,N_3242);
nor U6360 (N_6360,N_3025,N_2975);
xnor U6361 (N_6361,N_3419,N_4624);
xnor U6362 (N_6362,N_4720,N_4861);
and U6363 (N_6363,N_2678,N_4482);
xor U6364 (N_6364,N_4733,N_4874);
or U6365 (N_6365,N_3603,N_4390);
nor U6366 (N_6366,N_3768,N_3607);
xnor U6367 (N_6367,N_4445,N_4230);
or U6368 (N_6368,N_3628,N_4598);
or U6369 (N_6369,N_3509,N_4695);
and U6370 (N_6370,N_4022,N_4313);
nor U6371 (N_6371,N_4347,N_4918);
or U6372 (N_6372,N_3822,N_2521);
or U6373 (N_6373,N_3610,N_3269);
nor U6374 (N_6374,N_4057,N_3422);
or U6375 (N_6375,N_2516,N_2572);
nor U6376 (N_6376,N_3785,N_4905);
nor U6377 (N_6377,N_3862,N_4930);
xor U6378 (N_6378,N_2904,N_3164);
xnor U6379 (N_6379,N_4953,N_4220);
xnor U6380 (N_6380,N_4531,N_4048);
and U6381 (N_6381,N_3210,N_3069);
xnor U6382 (N_6382,N_2958,N_3730);
nand U6383 (N_6383,N_4537,N_3141);
or U6384 (N_6384,N_3254,N_2737);
and U6385 (N_6385,N_3141,N_3662);
xor U6386 (N_6386,N_4802,N_2686);
xor U6387 (N_6387,N_2990,N_2561);
and U6388 (N_6388,N_4065,N_4094);
xnor U6389 (N_6389,N_4126,N_4629);
xnor U6390 (N_6390,N_3289,N_4869);
or U6391 (N_6391,N_4562,N_4717);
and U6392 (N_6392,N_3116,N_3851);
xor U6393 (N_6393,N_2981,N_4694);
or U6394 (N_6394,N_4325,N_2830);
nor U6395 (N_6395,N_3612,N_4106);
nor U6396 (N_6396,N_3088,N_2625);
nor U6397 (N_6397,N_4750,N_3402);
xnor U6398 (N_6398,N_4504,N_3934);
nor U6399 (N_6399,N_4403,N_4708);
or U6400 (N_6400,N_3166,N_4236);
nand U6401 (N_6401,N_3797,N_4151);
nor U6402 (N_6402,N_2759,N_4705);
xor U6403 (N_6403,N_3659,N_3407);
nand U6404 (N_6404,N_4440,N_4303);
or U6405 (N_6405,N_4912,N_2821);
or U6406 (N_6406,N_4553,N_4388);
or U6407 (N_6407,N_2711,N_3635);
nor U6408 (N_6408,N_4825,N_4165);
nor U6409 (N_6409,N_3209,N_2964);
nand U6410 (N_6410,N_4938,N_4870);
or U6411 (N_6411,N_4966,N_2726);
nor U6412 (N_6412,N_3951,N_4416);
nor U6413 (N_6413,N_2691,N_3672);
nor U6414 (N_6414,N_2946,N_4399);
and U6415 (N_6415,N_2614,N_2695);
xor U6416 (N_6416,N_4801,N_4606);
xnor U6417 (N_6417,N_4119,N_3717);
xor U6418 (N_6418,N_4275,N_4835);
nand U6419 (N_6419,N_3042,N_4473);
xnor U6420 (N_6420,N_4219,N_3310);
or U6421 (N_6421,N_4407,N_3581);
or U6422 (N_6422,N_4928,N_3905);
or U6423 (N_6423,N_3395,N_3358);
and U6424 (N_6424,N_3631,N_3122);
or U6425 (N_6425,N_4904,N_3247);
or U6426 (N_6426,N_4563,N_4069);
or U6427 (N_6427,N_4145,N_4815);
nor U6428 (N_6428,N_4030,N_2791);
and U6429 (N_6429,N_3344,N_3871);
nor U6430 (N_6430,N_3272,N_2586);
xor U6431 (N_6431,N_4681,N_4811);
xor U6432 (N_6432,N_4977,N_4430);
xnor U6433 (N_6433,N_2846,N_4036);
nor U6434 (N_6434,N_4337,N_3241);
xor U6435 (N_6435,N_2691,N_4409);
xor U6436 (N_6436,N_3570,N_3003);
nand U6437 (N_6437,N_4053,N_3225);
nor U6438 (N_6438,N_4750,N_2754);
or U6439 (N_6439,N_4502,N_4070);
and U6440 (N_6440,N_4089,N_3748);
nor U6441 (N_6441,N_3883,N_3783);
nand U6442 (N_6442,N_3305,N_3920);
nand U6443 (N_6443,N_3799,N_3303);
nor U6444 (N_6444,N_3089,N_4467);
or U6445 (N_6445,N_4036,N_2776);
nand U6446 (N_6446,N_4057,N_4428);
or U6447 (N_6447,N_3032,N_4081);
xor U6448 (N_6448,N_3640,N_3816);
and U6449 (N_6449,N_2545,N_4842);
and U6450 (N_6450,N_3276,N_4968);
nand U6451 (N_6451,N_3720,N_4094);
nand U6452 (N_6452,N_3585,N_4111);
or U6453 (N_6453,N_3447,N_4531);
and U6454 (N_6454,N_4505,N_2724);
and U6455 (N_6455,N_2584,N_3021);
nor U6456 (N_6456,N_3784,N_3063);
and U6457 (N_6457,N_4094,N_3893);
or U6458 (N_6458,N_4301,N_2869);
or U6459 (N_6459,N_3798,N_4313);
or U6460 (N_6460,N_2901,N_3366);
nand U6461 (N_6461,N_2706,N_2958);
and U6462 (N_6462,N_4951,N_3309);
and U6463 (N_6463,N_2798,N_4554);
nand U6464 (N_6464,N_4638,N_4321);
xor U6465 (N_6465,N_3363,N_3626);
nand U6466 (N_6466,N_4607,N_4169);
nand U6467 (N_6467,N_3290,N_2779);
nand U6468 (N_6468,N_4635,N_3713);
nor U6469 (N_6469,N_4445,N_2741);
nor U6470 (N_6470,N_3074,N_3413);
xor U6471 (N_6471,N_3401,N_4598);
nor U6472 (N_6472,N_4896,N_3695);
nand U6473 (N_6473,N_4178,N_4673);
or U6474 (N_6474,N_2793,N_4493);
xor U6475 (N_6475,N_3726,N_4594);
xor U6476 (N_6476,N_3419,N_3494);
xor U6477 (N_6477,N_2538,N_4952);
nand U6478 (N_6478,N_4907,N_4658);
and U6479 (N_6479,N_4167,N_2586);
and U6480 (N_6480,N_2610,N_3419);
and U6481 (N_6481,N_2939,N_3866);
or U6482 (N_6482,N_4008,N_4967);
xor U6483 (N_6483,N_3478,N_4340);
nor U6484 (N_6484,N_4139,N_3770);
nor U6485 (N_6485,N_2698,N_3527);
xor U6486 (N_6486,N_4915,N_3602);
or U6487 (N_6487,N_3560,N_4974);
or U6488 (N_6488,N_2571,N_3004);
nor U6489 (N_6489,N_3422,N_4422);
nor U6490 (N_6490,N_3175,N_4056);
xor U6491 (N_6491,N_3234,N_2999);
xor U6492 (N_6492,N_2516,N_3099);
or U6493 (N_6493,N_3538,N_3079);
xor U6494 (N_6494,N_3653,N_4678);
nand U6495 (N_6495,N_2663,N_3203);
and U6496 (N_6496,N_4662,N_3387);
and U6497 (N_6497,N_4718,N_4562);
xnor U6498 (N_6498,N_4793,N_4442);
or U6499 (N_6499,N_3275,N_4123);
xor U6500 (N_6500,N_2667,N_3369);
xnor U6501 (N_6501,N_4864,N_4094);
nor U6502 (N_6502,N_3912,N_4874);
nor U6503 (N_6503,N_4043,N_4210);
nor U6504 (N_6504,N_3291,N_2538);
nand U6505 (N_6505,N_2631,N_3321);
and U6506 (N_6506,N_3417,N_3038);
and U6507 (N_6507,N_4719,N_2507);
xnor U6508 (N_6508,N_4956,N_3827);
xor U6509 (N_6509,N_2933,N_3599);
and U6510 (N_6510,N_2900,N_3108);
nor U6511 (N_6511,N_4326,N_3735);
nor U6512 (N_6512,N_3270,N_2711);
nand U6513 (N_6513,N_3418,N_2500);
and U6514 (N_6514,N_4353,N_3648);
xnor U6515 (N_6515,N_2891,N_4450);
and U6516 (N_6516,N_3303,N_4758);
nand U6517 (N_6517,N_3110,N_2936);
nor U6518 (N_6518,N_4255,N_4843);
or U6519 (N_6519,N_3078,N_4230);
or U6520 (N_6520,N_3633,N_2846);
or U6521 (N_6521,N_4569,N_4045);
nand U6522 (N_6522,N_2762,N_3408);
or U6523 (N_6523,N_3020,N_4148);
or U6524 (N_6524,N_4614,N_4320);
nor U6525 (N_6525,N_4334,N_3862);
and U6526 (N_6526,N_3430,N_2751);
nand U6527 (N_6527,N_4360,N_3852);
nand U6528 (N_6528,N_2863,N_3487);
nand U6529 (N_6529,N_4137,N_4390);
and U6530 (N_6530,N_2794,N_3201);
nor U6531 (N_6531,N_3314,N_3080);
nand U6532 (N_6532,N_3154,N_3869);
xnor U6533 (N_6533,N_4181,N_4937);
or U6534 (N_6534,N_3321,N_4697);
xnor U6535 (N_6535,N_4964,N_2500);
or U6536 (N_6536,N_4706,N_4602);
and U6537 (N_6537,N_4823,N_3028);
nor U6538 (N_6538,N_3249,N_2880);
xor U6539 (N_6539,N_3470,N_3594);
nor U6540 (N_6540,N_4863,N_4473);
or U6541 (N_6541,N_3688,N_2574);
xor U6542 (N_6542,N_3424,N_3558);
nor U6543 (N_6543,N_3614,N_3736);
nor U6544 (N_6544,N_3872,N_4159);
nand U6545 (N_6545,N_4985,N_2863);
xor U6546 (N_6546,N_3319,N_3331);
and U6547 (N_6547,N_4698,N_4813);
xor U6548 (N_6548,N_2851,N_2569);
and U6549 (N_6549,N_4104,N_2632);
nor U6550 (N_6550,N_3609,N_3222);
xor U6551 (N_6551,N_4483,N_3258);
xnor U6552 (N_6552,N_3403,N_3453);
or U6553 (N_6553,N_3667,N_4995);
nor U6554 (N_6554,N_4614,N_3156);
nand U6555 (N_6555,N_4480,N_2924);
nor U6556 (N_6556,N_3294,N_3686);
nor U6557 (N_6557,N_4787,N_3443);
nor U6558 (N_6558,N_3622,N_3730);
nor U6559 (N_6559,N_3666,N_3802);
nor U6560 (N_6560,N_3498,N_3302);
nor U6561 (N_6561,N_3712,N_3011);
nor U6562 (N_6562,N_4695,N_4564);
xnor U6563 (N_6563,N_4730,N_4801);
nor U6564 (N_6564,N_3914,N_3142);
nor U6565 (N_6565,N_3211,N_3521);
nand U6566 (N_6566,N_4944,N_3355);
or U6567 (N_6567,N_2537,N_4722);
or U6568 (N_6568,N_3213,N_4808);
xor U6569 (N_6569,N_4027,N_4284);
or U6570 (N_6570,N_2533,N_3818);
nor U6571 (N_6571,N_2569,N_4365);
and U6572 (N_6572,N_4580,N_3022);
or U6573 (N_6573,N_4473,N_4325);
and U6574 (N_6574,N_2626,N_4675);
or U6575 (N_6575,N_4322,N_3506);
xor U6576 (N_6576,N_2727,N_3413);
and U6577 (N_6577,N_3062,N_2575);
or U6578 (N_6578,N_3742,N_3290);
or U6579 (N_6579,N_3122,N_4606);
or U6580 (N_6580,N_3104,N_3357);
xor U6581 (N_6581,N_4795,N_4699);
and U6582 (N_6582,N_3149,N_3506);
nor U6583 (N_6583,N_4821,N_4302);
and U6584 (N_6584,N_4276,N_3561);
nor U6585 (N_6585,N_4579,N_3721);
xnor U6586 (N_6586,N_3353,N_3086);
nand U6587 (N_6587,N_2945,N_4102);
and U6588 (N_6588,N_3612,N_4031);
and U6589 (N_6589,N_3607,N_4812);
xnor U6590 (N_6590,N_2909,N_4544);
and U6591 (N_6591,N_2672,N_3037);
and U6592 (N_6592,N_3448,N_3527);
nand U6593 (N_6593,N_4519,N_3904);
nor U6594 (N_6594,N_4484,N_3380);
nand U6595 (N_6595,N_3607,N_3256);
nor U6596 (N_6596,N_4887,N_3753);
and U6597 (N_6597,N_3874,N_4256);
or U6598 (N_6598,N_4835,N_4505);
and U6599 (N_6599,N_4499,N_3815);
xnor U6600 (N_6600,N_4579,N_2617);
nand U6601 (N_6601,N_4857,N_4582);
nor U6602 (N_6602,N_3059,N_4868);
or U6603 (N_6603,N_3465,N_4489);
xnor U6604 (N_6604,N_2840,N_4304);
nand U6605 (N_6605,N_3503,N_3598);
nor U6606 (N_6606,N_4742,N_3568);
and U6607 (N_6607,N_3273,N_4002);
or U6608 (N_6608,N_2984,N_3726);
or U6609 (N_6609,N_4129,N_4164);
nor U6610 (N_6610,N_4549,N_4121);
or U6611 (N_6611,N_4773,N_3099);
and U6612 (N_6612,N_4194,N_4277);
nand U6613 (N_6613,N_4071,N_3897);
or U6614 (N_6614,N_3702,N_4933);
or U6615 (N_6615,N_3625,N_3007);
nor U6616 (N_6616,N_4127,N_4666);
nor U6617 (N_6617,N_4888,N_3126);
and U6618 (N_6618,N_4388,N_4211);
nand U6619 (N_6619,N_2972,N_4451);
nand U6620 (N_6620,N_4617,N_3461);
and U6621 (N_6621,N_3538,N_2571);
and U6622 (N_6622,N_3184,N_3428);
nor U6623 (N_6623,N_2842,N_4939);
xor U6624 (N_6624,N_2673,N_4551);
nand U6625 (N_6625,N_3809,N_2988);
xnor U6626 (N_6626,N_2600,N_3851);
or U6627 (N_6627,N_4298,N_4672);
nor U6628 (N_6628,N_3629,N_4454);
nand U6629 (N_6629,N_3204,N_4452);
or U6630 (N_6630,N_4964,N_4522);
nor U6631 (N_6631,N_3496,N_2589);
xnor U6632 (N_6632,N_4824,N_4291);
nand U6633 (N_6633,N_4935,N_3136);
nand U6634 (N_6634,N_4237,N_2560);
or U6635 (N_6635,N_3192,N_2637);
nand U6636 (N_6636,N_4101,N_4502);
xor U6637 (N_6637,N_4190,N_3391);
xnor U6638 (N_6638,N_3680,N_2942);
nand U6639 (N_6639,N_3880,N_3162);
or U6640 (N_6640,N_4858,N_3194);
nor U6641 (N_6641,N_2517,N_3068);
nand U6642 (N_6642,N_3067,N_3824);
nor U6643 (N_6643,N_4244,N_3922);
nand U6644 (N_6644,N_4967,N_2993);
and U6645 (N_6645,N_3523,N_2908);
nand U6646 (N_6646,N_3525,N_3673);
and U6647 (N_6647,N_4987,N_3096);
xor U6648 (N_6648,N_4175,N_4049);
nand U6649 (N_6649,N_3013,N_3208);
xnor U6650 (N_6650,N_4670,N_4442);
nand U6651 (N_6651,N_2500,N_2899);
nor U6652 (N_6652,N_3385,N_2665);
nor U6653 (N_6653,N_2576,N_4872);
nand U6654 (N_6654,N_3291,N_3033);
nand U6655 (N_6655,N_3979,N_4024);
or U6656 (N_6656,N_3767,N_2673);
nand U6657 (N_6657,N_4408,N_4983);
nand U6658 (N_6658,N_4893,N_3007);
or U6659 (N_6659,N_4669,N_3900);
and U6660 (N_6660,N_4167,N_3568);
nand U6661 (N_6661,N_3347,N_4155);
or U6662 (N_6662,N_3229,N_2656);
xor U6663 (N_6663,N_2618,N_4473);
xnor U6664 (N_6664,N_3263,N_4319);
xnor U6665 (N_6665,N_3883,N_3777);
nor U6666 (N_6666,N_2795,N_4987);
nand U6667 (N_6667,N_4396,N_4475);
and U6668 (N_6668,N_4209,N_3231);
or U6669 (N_6669,N_4319,N_3497);
and U6670 (N_6670,N_3219,N_3394);
nor U6671 (N_6671,N_4387,N_4339);
and U6672 (N_6672,N_2830,N_3764);
nand U6673 (N_6673,N_4243,N_4475);
nor U6674 (N_6674,N_3509,N_3120);
xor U6675 (N_6675,N_2674,N_3784);
nor U6676 (N_6676,N_2963,N_4801);
xnor U6677 (N_6677,N_3129,N_4461);
xor U6678 (N_6678,N_4701,N_3873);
nor U6679 (N_6679,N_4528,N_3985);
and U6680 (N_6680,N_2853,N_3699);
or U6681 (N_6681,N_3262,N_4860);
or U6682 (N_6682,N_4361,N_4549);
nor U6683 (N_6683,N_3657,N_2735);
and U6684 (N_6684,N_3701,N_4701);
xnor U6685 (N_6685,N_3322,N_3767);
or U6686 (N_6686,N_4386,N_2919);
nand U6687 (N_6687,N_3868,N_3428);
xor U6688 (N_6688,N_2797,N_2627);
and U6689 (N_6689,N_4778,N_2874);
xor U6690 (N_6690,N_3397,N_3324);
nand U6691 (N_6691,N_4224,N_3512);
xor U6692 (N_6692,N_2598,N_4849);
nand U6693 (N_6693,N_3492,N_3768);
or U6694 (N_6694,N_2570,N_3333);
and U6695 (N_6695,N_4845,N_3239);
or U6696 (N_6696,N_3143,N_3071);
nor U6697 (N_6697,N_4318,N_4756);
or U6698 (N_6698,N_4417,N_3869);
nand U6699 (N_6699,N_2675,N_4009);
xor U6700 (N_6700,N_3985,N_4985);
nor U6701 (N_6701,N_4872,N_4453);
nand U6702 (N_6702,N_4210,N_3386);
and U6703 (N_6703,N_4879,N_3906);
and U6704 (N_6704,N_2632,N_4902);
nand U6705 (N_6705,N_4954,N_3743);
or U6706 (N_6706,N_2588,N_4829);
xnor U6707 (N_6707,N_3273,N_4320);
and U6708 (N_6708,N_2532,N_4984);
and U6709 (N_6709,N_4018,N_2870);
nor U6710 (N_6710,N_2823,N_3917);
or U6711 (N_6711,N_4039,N_4121);
or U6712 (N_6712,N_4034,N_3409);
xor U6713 (N_6713,N_3439,N_3174);
xor U6714 (N_6714,N_3525,N_3191);
or U6715 (N_6715,N_3570,N_3099);
and U6716 (N_6716,N_2655,N_4280);
nand U6717 (N_6717,N_3853,N_2814);
or U6718 (N_6718,N_4265,N_4811);
xnor U6719 (N_6719,N_3639,N_3276);
and U6720 (N_6720,N_4277,N_4581);
nor U6721 (N_6721,N_2624,N_2874);
nor U6722 (N_6722,N_3290,N_4205);
or U6723 (N_6723,N_4065,N_4025);
xor U6724 (N_6724,N_4373,N_3119);
xor U6725 (N_6725,N_4182,N_2774);
nand U6726 (N_6726,N_2851,N_4314);
nand U6727 (N_6727,N_2957,N_4971);
xnor U6728 (N_6728,N_3714,N_4487);
and U6729 (N_6729,N_3731,N_2877);
xnor U6730 (N_6730,N_3454,N_4241);
and U6731 (N_6731,N_4275,N_4178);
or U6732 (N_6732,N_3376,N_3928);
nand U6733 (N_6733,N_4787,N_2558);
and U6734 (N_6734,N_2836,N_4760);
and U6735 (N_6735,N_4551,N_3095);
xnor U6736 (N_6736,N_3669,N_2897);
nor U6737 (N_6737,N_4206,N_2906);
or U6738 (N_6738,N_4121,N_4489);
or U6739 (N_6739,N_2747,N_3412);
and U6740 (N_6740,N_2843,N_3241);
and U6741 (N_6741,N_2589,N_3818);
nand U6742 (N_6742,N_2925,N_2662);
xnor U6743 (N_6743,N_4674,N_3503);
nor U6744 (N_6744,N_3056,N_3137);
or U6745 (N_6745,N_2584,N_4243);
or U6746 (N_6746,N_3448,N_4389);
xor U6747 (N_6747,N_3914,N_3170);
or U6748 (N_6748,N_4408,N_4801);
nor U6749 (N_6749,N_3596,N_4314);
and U6750 (N_6750,N_3330,N_3419);
and U6751 (N_6751,N_2949,N_3843);
nand U6752 (N_6752,N_2938,N_3843);
nor U6753 (N_6753,N_4967,N_3753);
nand U6754 (N_6754,N_2575,N_2929);
xnor U6755 (N_6755,N_2658,N_3981);
xnor U6756 (N_6756,N_4289,N_2772);
nand U6757 (N_6757,N_4734,N_2694);
and U6758 (N_6758,N_4573,N_3007);
xor U6759 (N_6759,N_3504,N_3589);
nand U6760 (N_6760,N_2692,N_2567);
or U6761 (N_6761,N_3959,N_3081);
and U6762 (N_6762,N_2527,N_4087);
and U6763 (N_6763,N_3237,N_3216);
nor U6764 (N_6764,N_3369,N_2634);
and U6765 (N_6765,N_4284,N_4195);
xor U6766 (N_6766,N_3638,N_2736);
xor U6767 (N_6767,N_2524,N_2750);
and U6768 (N_6768,N_2546,N_4734);
nand U6769 (N_6769,N_4135,N_4783);
nand U6770 (N_6770,N_4126,N_4868);
and U6771 (N_6771,N_3888,N_4645);
or U6772 (N_6772,N_4640,N_3648);
and U6773 (N_6773,N_4486,N_2966);
nand U6774 (N_6774,N_2840,N_4476);
nand U6775 (N_6775,N_3017,N_4131);
nand U6776 (N_6776,N_3250,N_3388);
nor U6777 (N_6777,N_4523,N_4481);
nand U6778 (N_6778,N_3581,N_2568);
nor U6779 (N_6779,N_2627,N_4371);
nand U6780 (N_6780,N_3730,N_3721);
nor U6781 (N_6781,N_2911,N_4507);
nor U6782 (N_6782,N_3868,N_3092);
nor U6783 (N_6783,N_2607,N_4286);
xor U6784 (N_6784,N_4795,N_2939);
xor U6785 (N_6785,N_2601,N_4736);
xnor U6786 (N_6786,N_3334,N_4910);
or U6787 (N_6787,N_3501,N_3363);
or U6788 (N_6788,N_4672,N_2574);
nor U6789 (N_6789,N_3898,N_2509);
nor U6790 (N_6790,N_4453,N_3802);
and U6791 (N_6791,N_4883,N_2867);
nand U6792 (N_6792,N_4275,N_3575);
and U6793 (N_6793,N_3454,N_3583);
nor U6794 (N_6794,N_4974,N_4705);
and U6795 (N_6795,N_4836,N_3643);
nand U6796 (N_6796,N_4147,N_2912);
or U6797 (N_6797,N_4267,N_3697);
xor U6798 (N_6798,N_2641,N_4813);
nor U6799 (N_6799,N_2644,N_4909);
nor U6800 (N_6800,N_4524,N_4879);
and U6801 (N_6801,N_4580,N_3949);
nand U6802 (N_6802,N_2997,N_3162);
nor U6803 (N_6803,N_2735,N_4224);
or U6804 (N_6804,N_4158,N_2567);
and U6805 (N_6805,N_3907,N_2522);
nand U6806 (N_6806,N_4952,N_3027);
or U6807 (N_6807,N_3044,N_2667);
nor U6808 (N_6808,N_2824,N_3671);
and U6809 (N_6809,N_4626,N_3188);
xor U6810 (N_6810,N_3928,N_4882);
nand U6811 (N_6811,N_3626,N_3865);
nand U6812 (N_6812,N_4164,N_3516);
and U6813 (N_6813,N_2553,N_2834);
xor U6814 (N_6814,N_3901,N_3479);
nor U6815 (N_6815,N_3802,N_4593);
or U6816 (N_6816,N_4725,N_3047);
xnor U6817 (N_6817,N_4513,N_3396);
xnor U6818 (N_6818,N_2980,N_4466);
and U6819 (N_6819,N_3317,N_4570);
nand U6820 (N_6820,N_4244,N_4869);
nand U6821 (N_6821,N_4108,N_3730);
nor U6822 (N_6822,N_2592,N_3665);
and U6823 (N_6823,N_3354,N_4253);
xnor U6824 (N_6824,N_3361,N_2931);
xnor U6825 (N_6825,N_3224,N_4480);
xnor U6826 (N_6826,N_3584,N_3639);
and U6827 (N_6827,N_3984,N_3028);
nand U6828 (N_6828,N_2624,N_3987);
xnor U6829 (N_6829,N_3223,N_3761);
nor U6830 (N_6830,N_4921,N_4894);
or U6831 (N_6831,N_3607,N_4414);
and U6832 (N_6832,N_3288,N_4937);
nand U6833 (N_6833,N_4348,N_3776);
or U6834 (N_6834,N_2579,N_4355);
and U6835 (N_6835,N_2658,N_2989);
xnor U6836 (N_6836,N_4704,N_2803);
nor U6837 (N_6837,N_4226,N_3193);
and U6838 (N_6838,N_3445,N_2637);
xnor U6839 (N_6839,N_4128,N_3332);
or U6840 (N_6840,N_4913,N_2720);
nand U6841 (N_6841,N_2626,N_2593);
or U6842 (N_6842,N_3563,N_4910);
xnor U6843 (N_6843,N_4367,N_3208);
and U6844 (N_6844,N_4948,N_4629);
and U6845 (N_6845,N_3041,N_3754);
or U6846 (N_6846,N_4876,N_3533);
and U6847 (N_6847,N_4163,N_3397);
xor U6848 (N_6848,N_2558,N_4993);
and U6849 (N_6849,N_3456,N_3441);
and U6850 (N_6850,N_2856,N_4594);
and U6851 (N_6851,N_4663,N_3853);
and U6852 (N_6852,N_4477,N_3766);
xnor U6853 (N_6853,N_2782,N_3503);
or U6854 (N_6854,N_4864,N_4302);
and U6855 (N_6855,N_3805,N_3578);
xor U6856 (N_6856,N_4937,N_3582);
nand U6857 (N_6857,N_3678,N_4983);
and U6858 (N_6858,N_3022,N_3725);
nor U6859 (N_6859,N_4309,N_4272);
nand U6860 (N_6860,N_4515,N_3760);
nor U6861 (N_6861,N_4298,N_3239);
nor U6862 (N_6862,N_4332,N_4451);
and U6863 (N_6863,N_3867,N_3943);
and U6864 (N_6864,N_3692,N_2869);
nand U6865 (N_6865,N_4296,N_4395);
nand U6866 (N_6866,N_4545,N_2673);
nand U6867 (N_6867,N_3694,N_3568);
or U6868 (N_6868,N_4024,N_2748);
nand U6869 (N_6869,N_3623,N_4037);
nand U6870 (N_6870,N_4242,N_2878);
nor U6871 (N_6871,N_3607,N_4593);
xnor U6872 (N_6872,N_2966,N_3797);
nor U6873 (N_6873,N_4454,N_3298);
nand U6874 (N_6874,N_4707,N_3735);
xnor U6875 (N_6875,N_4159,N_4409);
nand U6876 (N_6876,N_3830,N_4860);
nand U6877 (N_6877,N_3051,N_4198);
xnor U6878 (N_6878,N_4575,N_3687);
xnor U6879 (N_6879,N_3900,N_4144);
nand U6880 (N_6880,N_2568,N_2634);
nor U6881 (N_6881,N_4921,N_2880);
and U6882 (N_6882,N_2718,N_4970);
or U6883 (N_6883,N_3976,N_4202);
nor U6884 (N_6884,N_3124,N_4091);
nand U6885 (N_6885,N_3532,N_4201);
and U6886 (N_6886,N_4288,N_4393);
or U6887 (N_6887,N_4281,N_4882);
nor U6888 (N_6888,N_4270,N_4998);
nor U6889 (N_6889,N_3972,N_4879);
or U6890 (N_6890,N_2506,N_4687);
nor U6891 (N_6891,N_3861,N_4895);
or U6892 (N_6892,N_3947,N_3348);
or U6893 (N_6893,N_4631,N_2515);
or U6894 (N_6894,N_2576,N_3533);
or U6895 (N_6895,N_3349,N_3441);
nand U6896 (N_6896,N_2611,N_4934);
nor U6897 (N_6897,N_3615,N_4167);
xnor U6898 (N_6898,N_3444,N_4361);
nor U6899 (N_6899,N_4331,N_3413);
or U6900 (N_6900,N_3233,N_2762);
nand U6901 (N_6901,N_2656,N_4360);
xor U6902 (N_6902,N_4388,N_2692);
xor U6903 (N_6903,N_3747,N_3133);
and U6904 (N_6904,N_3436,N_2649);
nand U6905 (N_6905,N_3997,N_3975);
nor U6906 (N_6906,N_4554,N_2899);
nor U6907 (N_6907,N_3297,N_3864);
or U6908 (N_6908,N_3538,N_3583);
nand U6909 (N_6909,N_3645,N_3051);
nand U6910 (N_6910,N_2606,N_4347);
nand U6911 (N_6911,N_3375,N_3362);
and U6912 (N_6912,N_4898,N_4189);
nor U6913 (N_6913,N_2567,N_2701);
xor U6914 (N_6914,N_2656,N_3837);
nand U6915 (N_6915,N_4032,N_3343);
or U6916 (N_6916,N_4592,N_4509);
and U6917 (N_6917,N_2507,N_4299);
xnor U6918 (N_6918,N_3656,N_3321);
xnor U6919 (N_6919,N_4036,N_3156);
and U6920 (N_6920,N_2806,N_2696);
and U6921 (N_6921,N_4710,N_3080);
nand U6922 (N_6922,N_4124,N_3935);
xnor U6923 (N_6923,N_2772,N_4679);
and U6924 (N_6924,N_4659,N_3197);
and U6925 (N_6925,N_2767,N_4101);
and U6926 (N_6926,N_4670,N_3129);
and U6927 (N_6927,N_3687,N_3992);
nor U6928 (N_6928,N_4542,N_3435);
xor U6929 (N_6929,N_2848,N_4214);
nor U6930 (N_6930,N_2965,N_4579);
nand U6931 (N_6931,N_2805,N_3914);
nor U6932 (N_6932,N_3057,N_2641);
or U6933 (N_6933,N_3789,N_4874);
and U6934 (N_6934,N_4763,N_4794);
nand U6935 (N_6935,N_3065,N_2696);
or U6936 (N_6936,N_3330,N_4480);
nor U6937 (N_6937,N_4742,N_4263);
and U6938 (N_6938,N_2920,N_3224);
or U6939 (N_6939,N_3821,N_4328);
nor U6940 (N_6940,N_4017,N_2853);
xnor U6941 (N_6941,N_4569,N_3190);
or U6942 (N_6942,N_3549,N_3085);
xor U6943 (N_6943,N_2756,N_4445);
and U6944 (N_6944,N_4898,N_2550);
or U6945 (N_6945,N_4202,N_3384);
and U6946 (N_6946,N_4896,N_3421);
nand U6947 (N_6947,N_4764,N_3010);
nor U6948 (N_6948,N_4486,N_2700);
nor U6949 (N_6949,N_4814,N_4233);
or U6950 (N_6950,N_2545,N_3270);
nand U6951 (N_6951,N_4167,N_3381);
xnor U6952 (N_6952,N_4896,N_2747);
and U6953 (N_6953,N_3374,N_2960);
nor U6954 (N_6954,N_2979,N_3320);
or U6955 (N_6955,N_2644,N_4135);
or U6956 (N_6956,N_3775,N_3686);
or U6957 (N_6957,N_4968,N_4772);
nand U6958 (N_6958,N_3522,N_3279);
nand U6959 (N_6959,N_3329,N_3257);
nor U6960 (N_6960,N_2524,N_2624);
or U6961 (N_6961,N_2574,N_3837);
nor U6962 (N_6962,N_4403,N_3747);
xor U6963 (N_6963,N_4424,N_3897);
nand U6964 (N_6964,N_4246,N_3741);
and U6965 (N_6965,N_4392,N_4533);
and U6966 (N_6966,N_4787,N_3540);
nand U6967 (N_6967,N_4759,N_4114);
nand U6968 (N_6968,N_2538,N_4297);
nand U6969 (N_6969,N_3680,N_3978);
and U6970 (N_6970,N_3862,N_3122);
nor U6971 (N_6971,N_2999,N_2510);
or U6972 (N_6972,N_3298,N_3311);
nand U6973 (N_6973,N_4896,N_3345);
xor U6974 (N_6974,N_2661,N_2838);
or U6975 (N_6975,N_4663,N_3940);
nor U6976 (N_6976,N_4984,N_4269);
nand U6977 (N_6977,N_3169,N_4132);
nor U6978 (N_6978,N_2608,N_3976);
or U6979 (N_6979,N_2927,N_4854);
xnor U6980 (N_6980,N_3710,N_2517);
or U6981 (N_6981,N_3199,N_4998);
xor U6982 (N_6982,N_2595,N_4847);
or U6983 (N_6983,N_2926,N_3268);
and U6984 (N_6984,N_3044,N_3973);
nor U6985 (N_6985,N_3602,N_4346);
xor U6986 (N_6986,N_3436,N_3977);
nand U6987 (N_6987,N_3597,N_4441);
xor U6988 (N_6988,N_4776,N_4399);
xnor U6989 (N_6989,N_3285,N_3236);
nor U6990 (N_6990,N_2857,N_2624);
or U6991 (N_6991,N_2814,N_4402);
or U6992 (N_6992,N_4698,N_4447);
or U6993 (N_6993,N_4929,N_4825);
and U6994 (N_6994,N_4079,N_3148);
nand U6995 (N_6995,N_3109,N_4923);
xnor U6996 (N_6996,N_4883,N_4508);
nand U6997 (N_6997,N_3417,N_4638);
or U6998 (N_6998,N_4838,N_3587);
xor U6999 (N_6999,N_4891,N_3039);
and U7000 (N_7000,N_4640,N_3112);
and U7001 (N_7001,N_3551,N_3198);
xnor U7002 (N_7002,N_2535,N_3394);
nor U7003 (N_7003,N_2687,N_3581);
and U7004 (N_7004,N_2886,N_2782);
and U7005 (N_7005,N_3684,N_4062);
xnor U7006 (N_7006,N_3260,N_4197);
xor U7007 (N_7007,N_2726,N_2644);
nand U7008 (N_7008,N_3240,N_2679);
nand U7009 (N_7009,N_4914,N_4372);
nor U7010 (N_7010,N_3715,N_2508);
xnor U7011 (N_7011,N_4595,N_4541);
or U7012 (N_7012,N_4062,N_3424);
nor U7013 (N_7013,N_4886,N_4577);
or U7014 (N_7014,N_3112,N_3024);
or U7015 (N_7015,N_3402,N_3124);
and U7016 (N_7016,N_4091,N_3622);
and U7017 (N_7017,N_4703,N_2511);
nor U7018 (N_7018,N_3847,N_3249);
nand U7019 (N_7019,N_4517,N_3825);
and U7020 (N_7020,N_4294,N_3488);
or U7021 (N_7021,N_2799,N_3239);
xnor U7022 (N_7022,N_3090,N_4241);
nor U7023 (N_7023,N_3953,N_3153);
and U7024 (N_7024,N_3866,N_3968);
nor U7025 (N_7025,N_2927,N_4705);
xor U7026 (N_7026,N_4408,N_4327);
and U7027 (N_7027,N_2676,N_4319);
nor U7028 (N_7028,N_4447,N_3654);
nor U7029 (N_7029,N_2608,N_2512);
nand U7030 (N_7030,N_3396,N_2975);
or U7031 (N_7031,N_3934,N_3730);
and U7032 (N_7032,N_3045,N_3933);
xor U7033 (N_7033,N_4073,N_4996);
nand U7034 (N_7034,N_4722,N_2501);
nand U7035 (N_7035,N_4783,N_4812);
nand U7036 (N_7036,N_4048,N_4974);
xor U7037 (N_7037,N_4185,N_4031);
xor U7038 (N_7038,N_3731,N_3952);
nor U7039 (N_7039,N_3143,N_4977);
and U7040 (N_7040,N_4410,N_2511);
nor U7041 (N_7041,N_2745,N_4503);
and U7042 (N_7042,N_2863,N_4646);
xnor U7043 (N_7043,N_2834,N_2843);
nand U7044 (N_7044,N_4884,N_2535);
xor U7045 (N_7045,N_4244,N_3840);
or U7046 (N_7046,N_4263,N_2944);
and U7047 (N_7047,N_4724,N_3775);
nor U7048 (N_7048,N_3878,N_2850);
nor U7049 (N_7049,N_3571,N_3941);
or U7050 (N_7050,N_2607,N_4112);
nor U7051 (N_7051,N_3094,N_3959);
xnor U7052 (N_7052,N_3838,N_3678);
or U7053 (N_7053,N_3771,N_3303);
nor U7054 (N_7054,N_4029,N_4581);
nand U7055 (N_7055,N_3125,N_4340);
and U7056 (N_7056,N_4441,N_4146);
and U7057 (N_7057,N_2886,N_2518);
or U7058 (N_7058,N_4702,N_4765);
xor U7059 (N_7059,N_3011,N_4904);
xor U7060 (N_7060,N_4360,N_4899);
or U7061 (N_7061,N_3634,N_4357);
or U7062 (N_7062,N_4327,N_4639);
or U7063 (N_7063,N_3760,N_4719);
nor U7064 (N_7064,N_4369,N_3046);
and U7065 (N_7065,N_4776,N_3308);
or U7066 (N_7066,N_4486,N_4271);
nor U7067 (N_7067,N_4382,N_2710);
xor U7068 (N_7068,N_4132,N_3906);
nor U7069 (N_7069,N_2632,N_3665);
and U7070 (N_7070,N_4707,N_3098);
nand U7071 (N_7071,N_2578,N_3446);
and U7072 (N_7072,N_4986,N_3749);
and U7073 (N_7073,N_4275,N_3725);
or U7074 (N_7074,N_3227,N_4314);
nand U7075 (N_7075,N_4200,N_4420);
or U7076 (N_7076,N_4045,N_3126);
or U7077 (N_7077,N_4283,N_3484);
nor U7078 (N_7078,N_2899,N_3896);
or U7079 (N_7079,N_4652,N_4721);
nor U7080 (N_7080,N_3326,N_4582);
xor U7081 (N_7081,N_2745,N_4812);
or U7082 (N_7082,N_3439,N_3820);
and U7083 (N_7083,N_3219,N_4603);
and U7084 (N_7084,N_2568,N_4127);
xor U7085 (N_7085,N_4991,N_3090);
or U7086 (N_7086,N_3021,N_4927);
nand U7087 (N_7087,N_4688,N_3090);
or U7088 (N_7088,N_2811,N_3933);
or U7089 (N_7089,N_4962,N_3866);
nor U7090 (N_7090,N_2722,N_4082);
and U7091 (N_7091,N_3232,N_4503);
nor U7092 (N_7092,N_2898,N_2593);
nor U7093 (N_7093,N_2990,N_4270);
xor U7094 (N_7094,N_2905,N_4240);
and U7095 (N_7095,N_4781,N_3555);
nand U7096 (N_7096,N_3705,N_4368);
or U7097 (N_7097,N_3168,N_4655);
nor U7098 (N_7098,N_2977,N_3370);
nand U7099 (N_7099,N_4438,N_2565);
nand U7100 (N_7100,N_2677,N_4589);
and U7101 (N_7101,N_3492,N_4806);
or U7102 (N_7102,N_3312,N_3144);
xor U7103 (N_7103,N_4084,N_2996);
xnor U7104 (N_7104,N_3384,N_4530);
xnor U7105 (N_7105,N_4185,N_2527);
or U7106 (N_7106,N_4397,N_3448);
xnor U7107 (N_7107,N_3990,N_3714);
xnor U7108 (N_7108,N_4737,N_3281);
or U7109 (N_7109,N_2972,N_3101);
or U7110 (N_7110,N_2770,N_3427);
nor U7111 (N_7111,N_4961,N_3405);
or U7112 (N_7112,N_3298,N_3655);
xor U7113 (N_7113,N_3622,N_4939);
nand U7114 (N_7114,N_4601,N_3361);
and U7115 (N_7115,N_3225,N_4115);
or U7116 (N_7116,N_4405,N_4416);
nand U7117 (N_7117,N_3836,N_2762);
or U7118 (N_7118,N_3126,N_4870);
xor U7119 (N_7119,N_3512,N_4744);
and U7120 (N_7120,N_3929,N_2719);
and U7121 (N_7121,N_3412,N_3436);
xor U7122 (N_7122,N_4405,N_4489);
and U7123 (N_7123,N_4071,N_4061);
or U7124 (N_7124,N_2571,N_4668);
nand U7125 (N_7125,N_4976,N_4606);
nor U7126 (N_7126,N_3518,N_4482);
nand U7127 (N_7127,N_2506,N_2511);
nor U7128 (N_7128,N_3348,N_4904);
or U7129 (N_7129,N_4737,N_2744);
nor U7130 (N_7130,N_3586,N_3238);
xnor U7131 (N_7131,N_4712,N_3540);
xnor U7132 (N_7132,N_4914,N_4847);
and U7133 (N_7133,N_3322,N_2958);
nor U7134 (N_7134,N_3096,N_4291);
nor U7135 (N_7135,N_2660,N_3876);
nand U7136 (N_7136,N_2794,N_3312);
nor U7137 (N_7137,N_4444,N_3490);
or U7138 (N_7138,N_4733,N_2729);
nand U7139 (N_7139,N_4420,N_3824);
nor U7140 (N_7140,N_4912,N_4329);
nor U7141 (N_7141,N_3155,N_4118);
or U7142 (N_7142,N_3354,N_4150);
or U7143 (N_7143,N_2596,N_3234);
and U7144 (N_7144,N_4704,N_3706);
nand U7145 (N_7145,N_3586,N_4700);
or U7146 (N_7146,N_4867,N_4261);
xnor U7147 (N_7147,N_4797,N_4871);
nand U7148 (N_7148,N_4882,N_2535);
or U7149 (N_7149,N_2630,N_4101);
xor U7150 (N_7150,N_2777,N_4868);
and U7151 (N_7151,N_3097,N_4614);
nor U7152 (N_7152,N_3729,N_4164);
and U7153 (N_7153,N_2958,N_3480);
or U7154 (N_7154,N_4649,N_3552);
nor U7155 (N_7155,N_3786,N_3037);
nor U7156 (N_7156,N_3190,N_3604);
nor U7157 (N_7157,N_3415,N_3360);
nand U7158 (N_7158,N_4945,N_3191);
nand U7159 (N_7159,N_4302,N_3291);
and U7160 (N_7160,N_2543,N_2521);
and U7161 (N_7161,N_2941,N_3387);
and U7162 (N_7162,N_3023,N_4009);
nor U7163 (N_7163,N_3337,N_3481);
nor U7164 (N_7164,N_2513,N_4085);
nand U7165 (N_7165,N_3752,N_3316);
nand U7166 (N_7166,N_3556,N_3861);
and U7167 (N_7167,N_2817,N_2522);
and U7168 (N_7168,N_4314,N_2864);
nor U7169 (N_7169,N_4570,N_4617);
nor U7170 (N_7170,N_4286,N_2679);
or U7171 (N_7171,N_3652,N_3595);
nand U7172 (N_7172,N_4122,N_4430);
xor U7173 (N_7173,N_2621,N_2706);
or U7174 (N_7174,N_2563,N_3922);
or U7175 (N_7175,N_4638,N_4301);
nand U7176 (N_7176,N_4739,N_3156);
and U7177 (N_7177,N_2648,N_3587);
nand U7178 (N_7178,N_4887,N_2952);
nor U7179 (N_7179,N_3808,N_3274);
xor U7180 (N_7180,N_4655,N_3198);
and U7181 (N_7181,N_2708,N_4160);
and U7182 (N_7182,N_3904,N_4632);
xor U7183 (N_7183,N_4720,N_3952);
or U7184 (N_7184,N_3713,N_3935);
and U7185 (N_7185,N_4724,N_3345);
nor U7186 (N_7186,N_3474,N_3960);
and U7187 (N_7187,N_2933,N_3842);
xor U7188 (N_7188,N_2974,N_4129);
xor U7189 (N_7189,N_3707,N_3204);
or U7190 (N_7190,N_4809,N_4122);
or U7191 (N_7191,N_3174,N_4922);
or U7192 (N_7192,N_3355,N_3015);
xor U7193 (N_7193,N_3338,N_3219);
nand U7194 (N_7194,N_4591,N_4271);
nand U7195 (N_7195,N_4183,N_2828);
xor U7196 (N_7196,N_4108,N_4901);
or U7197 (N_7197,N_2875,N_3751);
xnor U7198 (N_7198,N_4642,N_3218);
xnor U7199 (N_7199,N_4274,N_3860);
nand U7200 (N_7200,N_2525,N_4394);
or U7201 (N_7201,N_4198,N_4870);
xor U7202 (N_7202,N_3527,N_3557);
or U7203 (N_7203,N_4239,N_3401);
nand U7204 (N_7204,N_3814,N_3192);
nand U7205 (N_7205,N_2749,N_3697);
or U7206 (N_7206,N_2628,N_3789);
or U7207 (N_7207,N_2676,N_2524);
nand U7208 (N_7208,N_2526,N_3138);
and U7209 (N_7209,N_4029,N_3469);
and U7210 (N_7210,N_3939,N_2665);
nor U7211 (N_7211,N_4948,N_2692);
and U7212 (N_7212,N_4443,N_3845);
xnor U7213 (N_7213,N_4655,N_3781);
xnor U7214 (N_7214,N_4553,N_2961);
nand U7215 (N_7215,N_2852,N_4595);
xnor U7216 (N_7216,N_4583,N_3229);
nor U7217 (N_7217,N_4416,N_3067);
or U7218 (N_7218,N_3357,N_4082);
nor U7219 (N_7219,N_2791,N_4306);
nand U7220 (N_7220,N_3235,N_2752);
and U7221 (N_7221,N_2661,N_4654);
nand U7222 (N_7222,N_2538,N_4913);
and U7223 (N_7223,N_4707,N_3712);
and U7224 (N_7224,N_4056,N_4433);
or U7225 (N_7225,N_4962,N_2724);
or U7226 (N_7226,N_2906,N_4540);
xnor U7227 (N_7227,N_2646,N_2681);
nor U7228 (N_7228,N_4544,N_2780);
or U7229 (N_7229,N_3608,N_4397);
nand U7230 (N_7230,N_3504,N_3867);
and U7231 (N_7231,N_3932,N_4301);
or U7232 (N_7232,N_4492,N_4183);
nand U7233 (N_7233,N_4009,N_4795);
nand U7234 (N_7234,N_2611,N_4315);
xnor U7235 (N_7235,N_3797,N_2723);
and U7236 (N_7236,N_2773,N_3598);
xnor U7237 (N_7237,N_3831,N_3307);
and U7238 (N_7238,N_4244,N_4722);
nor U7239 (N_7239,N_4793,N_3785);
and U7240 (N_7240,N_3229,N_2611);
nand U7241 (N_7241,N_3275,N_3570);
and U7242 (N_7242,N_3734,N_3633);
nand U7243 (N_7243,N_3251,N_4879);
nor U7244 (N_7244,N_4134,N_4498);
nand U7245 (N_7245,N_3923,N_4418);
xor U7246 (N_7246,N_4248,N_3996);
and U7247 (N_7247,N_3494,N_2602);
xor U7248 (N_7248,N_2791,N_4274);
nor U7249 (N_7249,N_2854,N_4684);
and U7250 (N_7250,N_4377,N_2553);
xnor U7251 (N_7251,N_4837,N_4623);
or U7252 (N_7252,N_2508,N_2978);
or U7253 (N_7253,N_2925,N_4847);
and U7254 (N_7254,N_4650,N_3503);
xnor U7255 (N_7255,N_4682,N_3819);
nor U7256 (N_7256,N_4484,N_4748);
nand U7257 (N_7257,N_3636,N_3834);
nand U7258 (N_7258,N_4196,N_4324);
nor U7259 (N_7259,N_3337,N_2601);
xor U7260 (N_7260,N_3461,N_4829);
or U7261 (N_7261,N_3084,N_4599);
nor U7262 (N_7262,N_4328,N_3228);
or U7263 (N_7263,N_4978,N_4465);
or U7264 (N_7264,N_2942,N_2939);
or U7265 (N_7265,N_3974,N_4109);
or U7266 (N_7266,N_4857,N_4474);
nor U7267 (N_7267,N_3706,N_3507);
nor U7268 (N_7268,N_3529,N_2523);
nor U7269 (N_7269,N_4856,N_4775);
xor U7270 (N_7270,N_3545,N_4851);
or U7271 (N_7271,N_3540,N_4233);
or U7272 (N_7272,N_3624,N_3153);
and U7273 (N_7273,N_4919,N_3933);
nand U7274 (N_7274,N_4168,N_3841);
nor U7275 (N_7275,N_4218,N_4381);
xnor U7276 (N_7276,N_3142,N_3800);
and U7277 (N_7277,N_3880,N_4575);
and U7278 (N_7278,N_3240,N_3210);
xnor U7279 (N_7279,N_3264,N_4698);
and U7280 (N_7280,N_4643,N_4946);
and U7281 (N_7281,N_3210,N_3047);
xor U7282 (N_7282,N_3616,N_3436);
nor U7283 (N_7283,N_3117,N_4974);
or U7284 (N_7284,N_4552,N_3858);
nor U7285 (N_7285,N_3114,N_3385);
nor U7286 (N_7286,N_4291,N_4670);
or U7287 (N_7287,N_4195,N_2709);
and U7288 (N_7288,N_2676,N_4972);
nand U7289 (N_7289,N_3314,N_4801);
nor U7290 (N_7290,N_4269,N_4635);
xnor U7291 (N_7291,N_2934,N_2878);
xnor U7292 (N_7292,N_3963,N_4765);
xor U7293 (N_7293,N_3684,N_4384);
and U7294 (N_7294,N_4993,N_3616);
nor U7295 (N_7295,N_4707,N_2526);
or U7296 (N_7296,N_3277,N_2880);
nand U7297 (N_7297,N_3172,N_4393);
nand U7298 (N_7298,N_2580,N_4910);
or U7299 (N_7299,N_4625,N_4636);
or U7300 (N_7300,N_3789,N_4193);
and U7301 (N_7301,N_3464,N_3833);
nor U7302 (N_7302,N_3544,N_4537);
nand U7303 (N_7303,N_3515,N_2778);
nand U7304 (N_7304,N_3625,N_4967);
nor U7305 (N_7305,N_4217,N_4804);
xor U7306 (N_7306,N_4241,N_3186);
or U7307 (N_7307,N_4130,N_3510);
nor U7308 (N_7308,N_3268,N_3726);
xor U7309 (N_7309,N_4454,N_4590);
or U7310 (N_7310,N_3104,N_4502);
nor U7311 (N_7311,N_3569,N_3965);
nor U7312 (N_7312,N_3937,N_4578);
xor U7313 (N_7313,N_3939,N_4889);
and U7314 (N_7314,N_4606,N_2567);
or U7315 (N_7315,N_3604,N_3723);
and U7316 (N_7316,N_4469,N_2844);
nor U7317 (N_7317,N_3705,N_3966);
nor U7318 (N_7318,N_3405,N_3522);
or U7319 (N_7319,N_3440,N_4924);
xor U7320 (N_7320,N_3277,N_3858);
nand U7321 (N_7321,N_2593,N_4944);
nor U7322 (N_7322,N_4806,N_2545);
nor U7323 (N_7323,N_3288,N_2601);
and U7324 (N_7324,N_3821,N_4669);
and U7325 (N_7325,N_4395,N_4165);
nor U7326 (N_7326,N_4866,N_4941);
nor U7327 (N_7327,N_3194,N_4965);
nor U7328 (N_7328,N_4126,N_3174);
and U7329 (N_7329,N_4788,N_4351);
and U7330 (N_7330,N_4844,N_3238);
nor U7331 (N_7331,N_4908,N_4577);
nor U7332 (N_7332,N_2821,N_3630);
and U7333 (N_7333,N_2710,N_4834);
and U7334 (N_7334,N_4522,N_2534);
xnor U7335 (N_7335,N_3107,N_4761);
xor U7336 (N_7336,N_4690,N_2689);
xor U7337 (N_7337,N_3099,N_4070);
or U7338 (N_7338,N_4467,N_3856);
nor U7339 (N_7339,N_3737,N_3250);
nor U7340 (N_7340,N_4999,N_4545);
nor U7341 (N_7341,N_4308,N_4595);
or U7342 (N_7342,N_2598,N_2781);
nor U7343 (N_7343,N_2891,N_3745);
nor U7344 (N_7344,N_3169,N_4818);
or U7345 (N_7345,N_4729,N_4153);
nand U7346 (N_7346,N_4882,N_3633);
and U7347 (N_7347,N_2610,N_4924);
xnor U7348 (N_7348,N_4052,N_2650);
or U7349 (N_7349,N_3495,N_4972);
or U7350 (N_7350,N_2698,N_3945);
nand U7351 (N_7351,N_3350,N_4899);
xor U7352 (N_7352,N_3091,N_2751);
or U7353 (N_7353,N_3567,N_3200);
nor U7354 (N_7354,N_3344,N_4248);
nor U7355 (N_7355,N_4472,N_2781);
or U7356 (N_7356,N_3296,N_3500);
xnor U7357 (N_7357,N_3313,N_3871);
nand U7358 (N_7358,N_4827,N_3598);
xnor U7359 (N_7359,N_2901,N_4962);
xor U7360 (N_7360,N_3469,N_2823);
or U7361 (N_7361,N_4971,N_4997);
or U7362 (N_7362,N_3352,N_3929);
xor U7363 (N_7363,N_4666,N_2638);
nor U7364 (N_7364,N_3036,N_3943);
nand U7365 (N_7365,N_3569,N_3239);
nand U7366 (N_7366,N_4737,N_3816);
or U7367 (N_7367,N_4373,N_3063);
or U7368 (N_7368,N_3735,N_3835);
nor U7369 (N_7369,N_3037,N_3700);
or U7370 (N_7370,N_3757,N_3880);
or U7371 (N_7371,N_4649,N_4229);
or U7372 (N_7372,N_3256,N_3349);
nand U7373 (N_7373,N_2746,N_4758);
nor U7374 (N_7374,N_3522,N_3321);
and U7375 (N_7375,N_4170,N_3256);
nand U7376 (N_7376,N_4880,N_4417);
nor U7377 (N_7377,N_4997,N_3819);
xor U7378 (N_7378,N_2754,N_3791);
nand U7379 (N_7379,N_4670,N_4779);
and U7380 (N_7380,N_3072,N_3537);
or U7381 (N_7381,N_3542,N_3366);
nor U7382 (N_7382,N_2766,N_2613);
nand U7383 (N_7383,N_3539,N_4094);
nor U7384 (N_7384,N_4254,N_4374);
xor U7385 (N_7385,N_3541,N_2891);
or U7386 (N_7386,N_4780,N_3464);
nor U7387 (N_7387,N_2905,N_3599);
and U7388 (N_7388,N_3460,N_4429);
xor U7389 (N_7389,N_2791,N_4061);
xnor U7390 (N_7390,N_4898,N_4717);
or U7391 (N_7391,N_2583,N_2546);
nor U7392 (N_7392,N_4345,N_3235);
nand U7393 (N_7393,N_4709,N_3431);
or U7394 (N_7394,N_4981,N_2656);
or U7395 (N_7395,N_4894,N_2964);
and U7396 (N_7396,N_3658,N_2633);
nand U7397 (N_7397,N_4347,N_3632);
and U7398 (N_7398,N_3736,N_4392);
nor U7399 (N_7399,N_3331,N_3887);
and U7400 (N_7400,N_4679,N_4953);
nor U7401 (N_7401,N_3700,N_3746);
or U7402 (N_7402,N_3206,N_2890);
or U7403 (N_7403,N_3096,N_4111);
nor U7404 (N_7404,N_2889,N_4808);
nand U7405 (N_7405,N_3627,N_2509);
xnor U7406 (N_7406,N_4965,N_4450);
or U7407 (N_7407,N_3339,N_3251);
nand U7408 (N_7408,N_4483,N_3963);
nor U7409 (N_7409,N_3570,N_2569);
nor U7410 (N_7410,N_3399,N_4265);
xnor U7411 (N_7411,N_4314,N_4138);
nand U7412 (N_7412,N_4502,N_4053);
or U7413 (N_7413,N_3818,N_3785);
xor U7414 (N_7414,N_3854,N_4490);
and U7415 (N_7415,N_3631,N_3965);
or U7416 (N_7416,N_2982,N_2551);
nand U7417 (N_7417,N_4960,N_4036);
nor U7418 (N_7418,N_2765,N_4564);
nand U7419 (N_7419,N_4670,N_4980);
or U7420 (N_7420,N_2966,N_4577);
or U7421 (N_7421,N_3032,N_2999);
or U7422 (N_7422,N_4107,N_4695);
or U7423 (N_7423,N_2838,N_4118);
xnor U7424 (N_7424,N_3082,N_4849);
nand U7425 (N_7425,N_3227,N_2986);
nand U7426 (N_7426,N_3302,N_3846);
nand U7427 (N_7427,N_4762,N_2816);
xor U7428 (N_7428,N_4145,N_4376);
nor U7429 (N_7429,N_3679,N_3373);
xnor U7430 (N_7430,N_4936,N_4119);
nand U7431 (N_7431,N_3320,N_2667);
or U7432 (N_7432,N_4936,N_4758);
or U7433 (N_7433,N_4642,N_4670);
and U7434 (N_7434,N_3085,N_3772);
xor U7435 (N_7435,N_3207,N_2701);
or U7436 (N_7436,N_3040,N_4075);
or U7437 (N_7437,N_2523,N_3655);
nand U7438 (N_7438,N_2547,N_4161);
xor U7439 (N_7439,N_4709,N_4878);
nand U7440 (N_7440,N_3918,N_3161);
or U7441 (N_7441,N_4144,N_3993);
xnor U7442 (N_7442,N_3837,N_4966);
nand U7443 (N_7443,N_4685,N_3373);
xnor U7444 (N_7444,N_4961,N_3273);
nor U7445 (N_7445,N_2594,N_4775);
or U7446 (N_7446,N_4457,N_4263);
xor U7447 (N_7447,N_2517,N_3800);
and U7448 (N_7448,N_4637,N_4877);
xnor U7449 (N_7449,N_4174,N_2909);
nor U7450 (N_7450,N_4842,N_2795);
and U7451 (N_7451,N_3001,N_4251);
nor U7452 (N_7452,N_4677,N_2801);
nand U7453 (N_7453,N_3376,N_4602);
nand U7454 (N_7454,N_3643,N_4685);
xnor U7455 (N_7455,N_3443,N_3526);
or U7456 (N_7456,N_4316,N_4186);
nor U7457 (N_7457,N_4132,N_3491);
xnor U7458 (N_7458,N_4037,N_4807);
or U7459 (N_7459,N_3849,N_4646);
or U7460 (N_7460,N_4932,N_3897);
or U7461 (N_7461,N_3626,N_2769);
xnor U7462 (N_7462,N_4636,N_4164);
or U7463 (N_7463,N_4220,N_3010);
xor U7464 (N_7464,N_4146,N_4137);
nor U7465 (N_7465,N_4754,N_2525);
and U7466 (N_7466,N_4839,N_2692);
nor U7467 (N_7467,N_4652,N_4747);
and U7468 (N_7468,N_4807,N_3050);
xor U7469 (N_7469,N_3284,N_4864);
nand U7470 (N_7470,N_3977,N_4389);
or U7471 (N_7471,N_3063,N_4511);
nand U7472 (N_7472,N_4722,N_2802);
xnor U7473 (N_7473,N_2784,N_2990);
xnor U7474 (N_7474,N_3705,N_4631);
nor U7475 (N_7475,N_3263,N_4006);
nand U7476 (N_7476,N_4757,N_4231);
xor U7477 (N_7477,N_3825,N_3458);
xnor U7478 (N_7478,N_2538,N_2566);
xnor U7479 (N_7479,N_2549,N_4031);
nor U7480 (N_7480,N_3341,N_4973);
or U7481 (N_7481,N_2512,N_2874);
nand U7482 (N_7482,N_4987,N_3902);
or U7483 (N_7483,N_3902,N_3436);
or U7484 (N_7484,N_4707,N_4225);
nor U7485 (N_7485,N_3498,N_4134);
and U7486 (N_7486,N_4240,N_4253);
nor U7487 (N_7487,N_4766,N_3324);
xor U7488 (N_7488,N_4411,N_4568);
nand U7489 (N_7489,N_3284,N_2684);
nand U7490 (N_7490,N_3572,N_4743);
nand U7491 (N_7491,N_4825,N_3158);
nand U7492 (N_7492,N_4144,N_4036);
nand U7493 (N_7493,N_4582,N_3592);
nor U7494 (N_7494,N_3796,N_4673);
or U7495 (N_7495,N_3713,N_2860);
or U7496 (N_7496,N_2853,N_4297);
or U7497 (N_7497,N_4636,N_2974);
xnor U7498 (N_7498,N_4282,N_4240);
nand U7499 (N_7499,N_2619,N_4585);
xnor U7500 (N_7500,N_7050,N_6869);
nor U7501 (N_7501,N_7246,N_5662);
and U7502 (N_7502,N_7368,N_6488);
nand U7503 (N_7503,N_6893,N_6382);
nand U7504 (N_7504,N_6247,N_5052);
nand U7505 (N_7505,N_6292,N_5113);
or U7506 (N_7506,N_6962,N_6688);
and U7507 (N_7507,N_5191,N_5478);
nor U7508 (N_7508,N_6053,N_6924);
xnor U7509 (N_7509,N_5375,N_5590);
xnor U7510 (N_7510,N_6141,N_5869);
nor U7511 (N_7511,N_5948,N_7414);
xnor U7512 (N_7512,N_7394,N_6862);
xor U7513 (N_7513,N_6128,N_7416);
xnor U7514 (N_7514,N_7242,N_5855);
and U7515 (N_7515,N_7395,N_5990);
and U7516 (N_7516,N_6113,N_6275);
xnor U7517 (N_7517,N_7270,N_5906);
nor U7518 (N_7518,N_5309,N_7439);
nor U7519 (N_7519,N_5148,N_6960);
nor U7520 (N_7520,N_5848,N_5017);
or U7521 (N_7521,N_5237,N_6337);
nand U7522 (N_7522,N_5429,N_7095);
and U7523 (N_7523,N_5835,N_5525);
nand U7524 (N_7524,N_6036,N_5680);
nor U7525 (N_7525,N_6780,N_5588);
and U7526 (N_7526,N_6546,N_5610);
nor U7527 (N_7527,N_6416,N_5838);
and U7528 (N_7528,N_7273,N_6354);
and U7529 (N_7529,N_5614,N_6592);
xnor U7530 (N_7530,N_6238,N_5932);
xnor U7531 (N_7531,N_5401,N_7052);
nand U7532 (N_7532,N_7228,N_5741);
xor U7533 (N_7533,N_6081,N_6925);
and U7534 (N_7534,N_5102,N_5160);
nor U7535 (N_7535,N_6218,N_7472);
and U7536 (N_7536,N_6381,N_5540);
or U7537 (N_7537,N_7140,N_7456);
xor U7538 (N_7538,N_7441,N_5611);
nand U7539 (N_7539,N_6191,N_6796);
and U7540 (N_7540,N_6087,N_5892);
nand U7541 (N_7541,N_7371,N_5004);
or U7542 (N_7542,N_5810,N_5999);
and U7543 (N_7543,N_6037,N_6512);
or U7544 (N_7544,N_6433,N_5231);
or U7545 (N_7545,N_7046,N_6226);
xor U7546 (N_7546,N_5597,N_5171);
and U7547 (N_7547,N_6310,N_6413);
nor U7548 (N_7548,N_7361,N_7265);
or U7549 (N_7549,N_5569,N_6786);
nor U7550 (N_7550,N_6114,N_7451);
nand U7551 (N_7551,N_6207,N_5034);
xor U7552 (N_7552,N_6300,N_7398);
nor U7553 (N_7553,N_6369,N_5937);
xor U7554 (N_7554,N_6561,N_5495);
or U7555 (N_7555,N_7388,N_5824);
and U7556 (N_7556,N_6626,N_7283);
xnor U7557 (N_7557,N_5969,N_5268);
or U7558 (N_7558,N_5441,N_5749);
nor U7559 (N_7559,N_5199,N_6673);
nor U7560 (N_7560,N_5554,N_5747);
nand U7561 (N_7561,N_5370,N_6966);
xor U7562 (N_7562,N_5660,N_6815);
and U7563 (N_7563,N_6825,N_5512);
xor U7564 (N_7564,N_5310,N_5153);
nor U7565 (N_7565,N_5389,N_7300);
xor U7566 (N_7566,N_5816,N_5468);
nand U7567 (N_7567,N_5390,N_6847);
nand U7568 (N_7568,N_6690,N_5057);
nor U7569 (N_7569,N_6415,N_5998);
or U7570 (N_7570,N_7411,N_6432);
or U7571 (N_7571,N_6918,N_5567);
and U7572 (N_7572,N_6770,N_5652);
xnor U7573 (N_7573,N_5950,N_6253);
and U7574 (N_7574,N_5851,N_6172);
and U7575 (N_7575,N_5471,N_6131);
nand U7576 (N_7576,N_7479,N_7212);
nand U7577 (N_7577,N_6027,N_7111);
and U7578 (N_7578,N_5219,N_5323);
nand U7579 (N_7579,N_5155,N_7393);
nor U7580 (N_7580,N_6933,N_5211);
and U7581 (N_7581,N_6232,N_7001);
and U7582 (N_7582,N_6608,N_6981);
nand U7583 (N_7583,N_5924,N_5149);
or U7584 (N_7584,N_6928,N_5533);
and U7585 (N_7585,N_7003,N_6622);
xnor U7586 (N_7586,N_5474,N_5053);
xnor U7587 (N_7587,N_7326,N_7367);
nand U7588 (N_7588,N_5260,N_5142);
nor U7589 (N_7589,N_7267,N_6948);
and U7590 (N_7590,N_5773,N_7178);
xor U7591 (N_7591,N_7440,N_5167);
nor U7592 (N_7592,N_7063,N_5581);
nor U7593 (N_7593,N_7202,N_7028);
nor U7594 (N_7594,N_6464,N_6889);
nand U7595 (N_7595,N_6777,N_6288);
nor U7596 (N_7596,N_5989,N_6767);
and U7597 (N_7597,N_6741,N_6917);
nand U7598 (N_7598,N_6322,N_6628);
or U7599 (N_7599,N_7229,N_6088);
and U7600 (N_7600,N_7215,N_5696);
nor U7601 (N_7601,N_7338,N_6619);
or U7602 (N_7602,N_5762,N_5890);
nor U7603 (N_7603,N_6216,N_7328);
xor U7604 (N_7604,N_7362,N_5695);
nand U7605 (N_7605,N_6186,N_6012);
or U7606 (N_7606,N_7276,N_5328);
nand U7607 (N_7607,N_7094,N_5656);
xnor U7608 (N_7608,N_7185,N_5623);
nand U7609 (N_7609,N_7272,N_5041);
and U7610 (N_7610,N_6240,N_7153);
and U7611 (N_7611,N_5184,N_5538);
xor U7612 (N_7612,N_6892,N_6340);
and U7613 (N_7613,N_5121,N_5952);
nor U7614 (N_7614,N_5802,N_5130);
xnor U7615 (N_7615,N_7399,N_5542);
xnor U7616 (N_7616,N_5265,N_7124);
nand U7617 (N_7617,N_6484,N_6792);
xnor U7618 (N_7618,N_7350,N_5087);
and U7619 (N_7619,N_6522,N_5748);
nor U7620 (N_7620,N_7029,N_5688);
and U7621 (N_7621,N_7415,N_6838);
xnor U7622 (N_7622,N_6364,N_5307);
xnor U7623 (N_7623,N_5535,N_5712);
nand U7624 (N_7624,N_6701,N_6902);
xor U7625 (N_7625,N_6376,N_7288);
nand U7626 (N_7626,N_6738,N_6610);
and U7627 (N_7627,N_6436,N_6570);
or U7628 (N_7628,N_5018,N_5889);
xnor U7629 (N_7629,N_7135,N_7258);
xor U7630 (N_7630,N_5766,N_6691);
or U7631 (N_7631,N_6748,N_7304);
nand U7632 (N_7632,N_6830,N_6900);
nor U7633 (N_7633,N_5676,N_7353);
nand U7634 (N_7634,N_5955,N_6321);
nor U7635 (N_7635,N_6472,N_6239);
nand U7636 (N_7636,N_5863,N_6277);
xnor U7637 (N_7637,N_5876,N_6394);
nor U7638 (N_7638,N_5528,N_7285);
or U7639 (N_7639,N_7167,N_5210);
nand U7640 (N_7640,N_5205,N_5062);
xnor U7641 (N_7641,N_6579,N_6162);
nor U7642 (N_7642,N_7250,N_5875);
and U7643 (N_7643,N_7425,N_5281);
nor U7644 (N_7644,N_7256,N_6035);
or U7645 (N_7645,N_6007,N_6696);
or U7646 (N_7646,N_6564,N_6751);
nor U7647 (N_7647,N_6351,N_5508);
nor U7648 (N_7648,N_5068,N_7133);
xnor U7649 (N_7649,N_6851,N_7237);
xnor U7650 (N_7650,N_6366,N_7157);
xor U7651 (N_7651,N_6174,N_5253);
xnor U7652 (N_7652,N_7310,N_6875);
nand U7653 (N_7653,N_5592,N_5621);
and U7654 (N_7654,N_5391,N_5746);
or U7655 (N_7655,N_5521,N_6912);
nand U7656 (N_7656,N_5685,N_6237);
nor U7657 (N_7657,N_7069,N_5398);
nand U7658 (N_7658,N_7308,N_5591);
nand U7659 (N_7659,N_7171,N_6897);
xor U7660 (N_7660,N_7173,N_5315);
or U7661 (N_7661,N_5853,N_5903);
nand U7662 (N_7662,N_6490,N_6434);
nor U7663 (N_7663,N_6998,N_7142);
and U7664 (N_7664,N_6248,N_5648);
nor U7665 (N_7665,N_6383,N_7421);
xor U7666 (N_7666,N_6812,N_5550);
xnor U7667 (N_7667,N_5861,N_7390);
xor U7668 (N_7668,N_5314,N_5404);
or U7669 (N_7669,N_5966,N_5169);
or U7670 (N_7670,N_6123,N_5934);
xor U7671 (N_7671,N_5161,N_5981);
nor U7672 (N_7672,N_7091,N_6665);
nor U7673 (N_7673,N_5985,N_6894);
nor U7674 (N_7674,N_6806,N_5867);
xor U7675 (N_7675,N_6271,N_6316);
nor U7676 (N_7676,N_5479,N_6934);
nor U7677 (N_7677,N_5120,N_5095);
nand U7678 (N_7678,N_6375,N_6721);
or U7679 (N_7679,N_6221,N_5285);
nor U7680 (N_7680,N_5831,N_6227);
and U7681 (N_7681,N_7305,N_6882);
or U7682 (N_7682,N_7130,N_5176);
and U7683 (N_7683,N_5634,N_5625);
nor U7684 (N_7684,N_5679,N_5322);
and U7685 (N_7685,N_5415,N_5523);
and U7686 (N_7686,N_5514,N_6646);
nand U7687 (N_7687,N_5797,N_7044);
or U7688 (N_7688,N_7365,N_6607);
nor U7689 (N_7689,N_6471,N_5821);
nand U7690 (N_7690,N_6813,N_6683);
nor U7691 (N_7691,N_5560,N_6704);
or U7692 (N_7692,N_5896,N_6142);
nor U7693 (N_7693,N_6408,N_7468);
nand U7694 (N_7694,N_6881,N_7358);
or U7695 (N_7695,N_5984,N_6492);
nor U7696 (N_7696,N_7465,N_5911);
and U7697 (N_7697,N_5438,N_7120);
and U7698 (N_7698,N_6947,N_6595);
and U7699 (N_7699,N_6040,N_5456);
and U7700 (N_7700,N_5243,N_6151);
nand U7701 (N_7701,N_6009,N_5044);
and U7702 (N_7702,N_5227,N_5879);
nor U7703 (N_7703,N_5939,N_6030);
and U7704 (N_7704,N_6693,N_7181);
nor U7705 (N_7705,N_5975,N_6720);
xor U7706 (N_7706,N_5868,N_7322);
xnor U7707 (N_7707,N_6206,N_5392);
or U7708 (N_7708,N_6975,N_6794);
or U7709 (N_7709,N_5991,N_7040);
and U7710 (N_7710,N_6352,N_5419);
or U7711 (N_7711,N_6153,N_5814);
or U7712 (N_7712,N_5453,N_5806);
or U7713 (N_7713,N_6290,N_6306);
and U7714 (N_7714,N_6219,N_5872);
or U7715 (N_7715,N_5234,N_7075);
nand U7716 (N_7716,N_5711,N_5175);
and U7717 (N_7717,N_6637,N_5139);
or U7718 (N_7718,N_6784,N_7147);
or U7719 (N_7719,N_7344,N_6896);
and U7720 (N_7720,N_5048,N_7081);
nor U7721 (N_7721,N_5337,N_6510);
nand U7722 (N_7722,N_5692,N_5393);
nor U7723 (N_7723,N_5181,N_6409);
nand U7724 (N_7724,N_6572,N_5620);
nor U7725 (N_7725,N_6257,N_7168);
or U7726 (N_7726,N_6846,N_5069);
and U7727 (N_7727,N_5757,N_7231);
nand U7728 (N_7728,N_6709,N_5953);
nand U7729 (N_7729,N_7461,N_5137);
nor U7730 (N_7730,N_6022,N_5426);
nor U7731 (N_7731,N_5925,N_6656);
nor U7732 (N_7732,N_5815,N_7331);
or U7733 (N_7733,N_5229,N_7027);
nor U7734 (N_7734,N_6001,N_5763);
nor U7735 (N_7735,N_7192,N_6612);
and U7736 (N_7736,N_5024,N_6119);
nor U7737 (N_7737,N_5582,N_6495);
nand U7738 (N_7738,N_6308,N_7352);
nor U7739 (N_7739,N_7249,N_6583);
nand U7740 (N_7740,N_6029,N_6718);
nand U7741 (N_7741,N_5603,N_6980);
xnor U7742 (N_7742,N_6988,N_6230);
xnor U7743 (N_7743,N_5724,N_5269);
nand U7744 (N_7744,N_5992,N_7418);
nand U7745 (N_7745,N_5589,N_5854);
nand U7746 (N_7746,N_6742,N_6251);
and U7747 (N_7747,N_7221,N_5271);
nor U7748 (N_7748,N_5015,N_5382);
or U7749 (N_7749,N_5795,N_6568);
nor U7750 (N_7750,N_6549,N_5794);
nand U7751 (N_7751,N_7125,N_5670);
and U7752 (N_7752,N_7491,N_5104);
nand U7753 (N_7753,N_5127,N_5788);
nor U7754 (N_7754,N_7422,N_5403);
xnor U7755 (N_7755,N_6362,N_6563);
nor U7756 (N_7756,N_5201,N_6294);
nor U7757 (N_7757,N_6299,N_7420);
or U7758 (N_7758,N_7301,N_5021);
or U7759 (N_7759,N_6342,N_5699);
or U7760 (N_7760,N_6942,N_7093);
xnor U7761 (N_7761,N_5064,N_6580);
and U7762 (N_7762,N_5073,N_6148);
xnor U7763 (N_7763,N_6098,N_6745);
nand U7764 (N_7764,N_6614,N_6267);
or U7765 (N_7765,N_6843,N_5248);
nand U7766 (N_7766,N_5881,N_6063);
nor U7767 (N_7767,N_6883,N_7233);
and U7768 (N_7768,N_5172,N_6328);
and U7769 (N_7769,N_5974,N_6903);
xnor U7770 (N_7770,N_7189,N_6145);
nand U7771 (N_7771,N_6067,N_5728);
nand U7772 (N_7772,N_6929,N_5481);
or U7773 (N_7773,N_6655,N_6454);
xor U7774 (N_7774,N_6169,N_5530);
and U7775 (N_7775,N_7449,N_6807);
and U7776 (N_7776,N_6167,N_6258);
nand U7777 (N_7777,N_5672,N_7132);
nand U7778 (N_7778,N_6422,N_6789);
nor U7779 (N_7779,N_5830,N_6938);
nand U7780 (N_7780,N_5000,N_5440);
or U7781 (N_7781,N_5808,N_5183);
and U7782 (N_7782,N_7049,N_5963);
nor U7783 (N_7783,N_5078,N_6031);
or U7784 (N_7784,N_6986,N_6190);
and U7785 (N_7785,N_6641,N_6809);
or U7786 (N_7786,N_5743,N_6915);
xor U7787 (N_7787,N_7030,N_5319);
and U7788 (N_7788,N_6404,N_6594);
or U7789 (N_7789,N_5507,N_7260);
nor U7790 (N_7790,N_5895,N_7110);
xor U7791 (N_7791,N_6010,N_7086);
and U7792 (N_7792,N_5045,N_6241);
nand U7793 (N_7793,N_6757,N_6927);
nand U7794 (N_7794,N_7478,N_6831);
and U7795 (N_7795,N_6201,N_6481);
nand U7796 (N_7796,N_5764,N_5131);
nor U7797 (N_7797,N_5026,N_6707);
xnor U7798 (N_7798,N_7281,N_5196);
xor U7799 (N_7799,N_5972,N_7196);
or U7800 (N_7800,N_6250,N_6097);
and U7801 (N_7801,N_6129,N_5050);
nand U7802 (N_7802,N_6558,N_5408);
or U7803 (N_7803,N_5433,N_7201);
nand U7804 (N_7804,N_7376,N_5860);
nand U7805 (N_7805,N_5626,N_7407);
or U7806 (N_7806,N_5631,N_6817);
nand U7807 (N_7807,N_6544,N_5332);
and U7808 (N_7808,N_5255,N_6543);
nand U7809 (N_7809,N_5263,N_6841);
xnor U7810 (N_7810,N_6615,N_7060);
nor U7811 (N_7811,N_5076,N_7222);
and U7812 (N_7812,N_5931,N_5358);
nand U7813 (N_7813,N_5090,N_7127);
or U7814 (N_7814,N_5510,N_5945);
nand U7815 (N_7815,N_5612,N_6995);
nor U7816 (N_7816,N_6104,N_6747);
or U7817 (N_7817,N_5163,N_6913);
and U7818 (N_7818,N_5106,N_6100);
xor U7819 (N_7819,N_6618,N_6970);
nor U7820 (N_7820,N_7155,N_6005);
and U7821 (N_7821,N_5553,N_5386);
xor U7822 (N_7822,N_5038,N_7444);
or U7823 (N_7823,N_6771,N_7483);
xor U7824 (N_7824,N_5771,N_6943);
nand U7825 (N_7825,N_5883,N_5075);
nor U7826 (N_7826,N_7442,N_7072);
xor U7827 (N_7827,N_6735,N_5336);
xnor U7828 (N_7828,N_5497,N_6477);
nor U7829 (N_7829,N_6587,N_5689);
nor U7830 (N_7830,N_7453,N_6959);
and U7831 (N_7831,N_5424,N_5649);
nand U7832 (N_7832,N_7492,N_6393);
xor U7833 (N_7833,N_5970,N_6750);
or U7834 (N_7834,N_6565,N_6043);
or U7835 (N_7835,N_5862,N_6672);
and U7836 (N_7836,N_5786,N_6138);
and U7837 (N_7837,N_5641,N_6950);
or U7838 (N_7838,N_5813,N_5980);
and U7839 (N_7839,N_6449,N_6629);
nor U7840 (N_7840,N_6776,N_5225);
xnor U7841 (N_7841,N_6289,N_6055);
xor U7842 (N_7842,N_6179,N_6837);
nand U7843 (N_7843,N_6633,N_6888);
or U7844 (N_7844,N_5477,N_7097);
and U7845 (N_7845,N_6386,N_5228);
xor U7846 (N_7846,N_7204,N_5295);
nor U7847 (N_7847,N_6157,N_6575);
and U7848 (N_7848,N_6154,N_7199);
or U7849 (N_7849,N_5736,N_5112);
nor U7850 (N_7850,N_6121,N_6092);
and U7851 (N_7851,N_6410,N_6474);
and U7852 (N_7852,N_7187,N_5347);
or U7853 (N_7853,N_6723,N_6758);
or U7854 (N_7854,N_5028,N_6684);
nor U7855 (N_7855,N_7443,N_6215);
nand U7856 (N_7856,N_5212,N_5572);
or U7857 (N_7857,N_5461,N_6527);
xor U7858 (N_7858,N_5576,N_5914);
or U7859 (N_7859,N_5718,N_5381);
and U7860 (N_7860,N_6229,N_5236);
xor U7861 (N_7861,N_6374,N_6165);
and U7862 (N_7862,N_5146,N_5504);
and U7863 (N_7863,N_5061,N_5674);
nor U7864 (N_7864,N_5402,N_6754);
or U7865 (N_7865,N_5907,N_7137);
and U7866 (N_7866,N_5579,N_5564);
nand U7867 (N_7867,N_5344,N_6095);
or U7868 (N_7868,N_5060,N_5362);
and U7869 (N_7869,N_6181,N_7005);
and U7870 (N_7870,N_6150,N_5252);
or U7871 (N_7871,N_6214,N_5030);
nand U7872 (N_7872,N_5361,N_6367);
nand U7873 (N_7873,N_5006,N_5288);
xor U7874 (N_7874,N_5058,N_6973);
and U7875 (N_7875,N_7116,N_6463);
nor U7876 (N_7876,N_5178,N_6057);
nor U7877 (N_7877,N_6996,N_5709);
or U7878 (N_7878,N_5013,N_5618);
and U7879 (N_7879,N_6122,N_7471);
xor U7880 (N_7880,N_6158,N_6799);
nand U7881 (N_7881,N_6795,N_6597);
nand U7882 (N_7882,N_6402,N_5317);
nand U7883 (N_7883,N_6706,N_5291);
nand U7884 (N_7884,N_5812,N_6945);
nor U7885 (N_7885,N_5458,N_6657);
or U7886 (N_7886,N_5449,N_5070);
and U7887 (N_7887,N_6156,N_7314);
xor U7888 (N_7888,N_5040,N_7016);
or U7889 (N_7889,N_6120,N_7218);
xnor U7890 (N_7890,N_6804,N_6109);
xor U7891 (N_7891,N_6076,N_6245);
nor U7892 (N_7892,N_5943,N_6428);
nand U7893 (N_7893,N_6103,N_5632);
or U7894 (N_7894,N_5186,N_5502);
nor U7895 (N_7895,N_6282,N_6640);
nor U7896 (N_7896,N_5051,N_6976);
nor U7897 (N_7897,N_6370,N_5059);
or U7898 (N_7898,N_7405,N_7000);
nor U7899 (N_7899,N_6476,N_6648);
and U7900 (N_7900,N_5527,N_6593);
or U7901 (N_7901,N_5593,N_5713);
nand U7902 (N_7902,N_7271,N_6183);
xor U7903 (N_7903,N_7397,N_6631);
nand U7904 (N_7904,N_6724,N_6203);
nor U7905 (N_7905,N_5671,N_5270);
nor U7906 (N_7906,N_6635,N_7056);
xor U7907 (N_7907,N_7136,N_7291);
xnor U7908 (N_7908,N_6021,N_6430);
or U7909 (N_7909,N_5077,N_5432);
nor U7910 (N_7910,N_6163,N_5298);
and U7911 (N_7911,N_5958,N_5485);
nor U7912 (N_7912,N_6365,N_5166);
or U7913 (N_7913,N_5664,N_5509);
nand U7914 (N_7914,N_6687,N_5123);
and U7915 (N_7915,N_5330,N_6028);
and U7916 (N_7916,N_6397,N_5141);
or U7917 (N_7917,N_6772,N_5194);
nor U7918 (N_7918,N_6774,N_6677);
nor U7919 (N_7919,N_5817,N_7074);
nor U7920 (N_7920,N_5729,N_7105);
or U7921 (N_7921,N_7051,N_5129);
or U7922 (N_7922,N_6264,N_5339);
or U7923 (N_7923,N_5177,N_6054);
nand U7924 (N_7924,N_6538,N_5321);
xor U7925 (N_7925,N_7239,N_5546);
nor U7926 (N_7926,N_6307,N_6731);
nor U7927 (N_7927,N_5744,N_7404);
or U7928 (N_7928,N_6161,N_5733);
and U7929 (N_7929,N_7311,N_5107);
xnor U7930 (N_7930,N_7345,N_6884);
nor U7931 (N_7931,N_5500,N_6852);
or U7932 (N_7932,N_7011,N_5425);
or U7933 (N_7933,N_6301,N_6254);
nand U7934 (N_7934,N_6205,N_5598);
xor U7935 (N_7935,N_6620,N_7334);
nor U7936 (N_7936,N_6359,N_6042);
xor U7937 (N_7937,N_6761,N_6318);
or U7938 (N_7938,N_6797,N_5434);
xor U7939 (N_7939,N_7190,N_6050);
and U7940 (N_7940,N_5673,N_5266);
nand U7941 (N_7941,N_7089,N_6578);
and U7942 (N_7942,N_6930,N_7152);
xnor U7943 (N_7943,N_6828,N_5930);
xor U7944 (N_7944,N_7145,N_6854);
and U7945 (N_7945,N_6038,N_6286);
nand U7946 (N_7946,N_5946,N_6378);
and U7947 (N_7947,N_6480,N_6255);
or U7948 (N_7948,N_6333,N_6905);
nor U7949 (N_7949,N_6468,N_5047);
xor U7950 (N_7950,N_6462,N_5927);
nor U7951 (N_7951,N_5608,N_5511);
nand U7952 (N_7952,N_6524,N_5442);
nor U7953 (N_7953,N_5377,N_5306);
or U7954 (N_7954,N_6170,N_7156);
xnor U7955 (N_7955,N_5214,N_5857);
or U7956 (N_7956,N_5333,N_6379);
or U7957 (N_7957,N_6589,N_5202);
nor U7958 (N_7958,N_5010,N_5367);
and U7959 (N_7959,N_6764,N_6315);
nand U7960 (N_7960,N_5494,N_6083);
and U7961 (N_7961,N_6319,N_6802);
xor U7962 (N_7962,N_5846,N_6552);
and U7963 (N_7963,N_7485,N_5331);
nor U7964 (N_7964,N_5505,N_6392);
nor U7965 (N_7965,N_7419,N_7054);
nand U7966 (N_7966,N_7437,N_5462);
or U7967 (N_7967,N_5739,N_5165);
nand U7968 (N_7968,N_6242,N_6719);
xnor U7969 (N_7969,N_5880,N_6391);
nor U7970 (N_7970,N_6094,N_6753);
or U7971 (N_7971,N_5758,N_6448);
or U7972 (N_7972,N_5463,N_5368);
nor U7973 (N_7973,N_7266,N_5893);
nand U7974 (N_7974,N_6399,N_5168);
nand U7975 (N_7975,N_6773,N_5208);
or U7976 (N_7976,N_6458,N_5725);
or U7977 (N_7977,N_7269,N_6668);
nor U7978 (N_7978,N_7232,N_5837);
nand U7979 (N_7979,N_7217,N_6496);
nor U7980 (N_7980,N_5562,N_5369);
or U7981 (N_7981,N_6361,N_5785);
xnor U7982 (N_7982,N_5353,N_6539);
nor U7983 (N_7983,N_7428,N_7457);
and U7984 (N_7984,N_6909,N_6541);
and U7985 (N_7985,N_6760,N_6818);
and U7986 (N_7986,N_6291,N_6456);
xor U7987 (N_7987,N_5455,N_7245);
and U7988 (N_7988,N_6395,N_6406);
nand U7989 (N_7989,N_5717,N_6500);
nand U7990 (N_7990,N_5483,N_7332);
and U7991 (N_7991,N_6279,N_6664);
nand U7992 (N_7992,N_6473,N_5427);
and U7993 (N_7993,N_6647,N_5378);
or U7994 (N_7994,N_5035,N_5967);
nor U7995 (N_7995,N_6863,N_6680);
or U7996 (N_7996,N_6136,N_7131);
xnor U7997 (N_7997,N_6630,N_7340);
nand U7998 (N_7998,N_6396,N_5420);
nor U7999 (N_7999,N_7452,N_5083);
nand U8000 (N_8000,N_6555,N_5702);
or U8001 (N_8001,N_7293,N_5944);
xnor U8002 (N_8002,N_5094,N_5138);
nand U8003 (N_8003,N_6173,N_7435);
xnor U8004 (N_8004,N_6372,N_6714);
and U8005 (N_8005,N_6708,N_6293);
xor U8006 (N_8006,N_6494,N_6732);
nand U8007 (N_8007,N_6209,N_5994);
xnor U8008 (N_8008,N_5900,N_5103);
or U8009 (N_8009,N_6344,N_5681);
nand U8010 (N_8010,N_7210,N_5811);
nor U8011 (N_8011,N_5556,N_7348);
and U8012 (N_8012,N_6600,N_5223);
and U8013 (N_8013,N_6590,N_5902);
or U8014 (N_8014,N_6526,N_6702);
and U8015 (N_8015,N_5318,N_7170);
or U8016 (N_8016,N_5850,N_6478);
nand U8017 (N_8017,N_7033,N_5126);
nand U8018 (N_8018,N_7409,N_7417);
and U8019 (N_8019,N_7255,N_5311);
and U8020 (N_8020,N_5936,N_5529);
nor U8021 (N_8021,N_6411,N_7101);
nor U8022 (N_8022,N_6327,N_6911);
nor U8023 (N_8023,N_5293,N_6553);
nand U8024 (N_8024,N_6112,N_6919);
nor U8025 (N_8025,N_7317,N_6762);
xor U8026 (N_8026,N_5345,N_5842);
xor U8027 (N_8027,N_6280,N_7268);
or U8028 (N_8028,N_6509,N_7071);
nand U8029 (N_8029,N_7315,N_5677);
xnor U8030 (N_8030,N_7445,N_5767);
nor U8031 (N_8031,N_7039,N_5586);
xnor U8032 (N_8032,N_5118,N_6144);
and U8033 (N_8033,N_6969,N_5559);
nand U8034 (N_8034,N_6908,N_6537);
xor U8035 (N_8035,N_7227,N_5878);
and U8036 (N_8036,N_7299,N_5905);
xor U8037 (N_8037,N_6877,N_6827);
nor U8038 (N_8038,N_5715,N_5239);
xnor U8039 (N_8039,N_6444,N_7289);
nor U8040 (N_8040,N_7088,N_6065);
nor U8041 (N_8041,N_6783,N_6438);
xnor U8042 (N_8042,N_5374,N_7129);
xnor U8043 (N_8043,N_7477,N_6699);
nand U8044 (N_8044,N_5092,N_7224);
and U8045 (N_8045,N_5250,N_6075);
and U8046 (N_8046,N_6921,N_6263);
and U8047 (N_8047,N_7223,N_6069);
or U8048 (N_8048,N_7287,N_5222);
and U8049 (N_8049,N_7454,N_7172);
nand U8050 (N_8050,N_5645,N_7104);
nor U8051 (N_8051,N_5154,N_6111);
and U8052 (N_8052,N_5385,N_6634);
xnor U8053 (N_8053,N_5159,N_7355);
nand U8054 (N_8054,N_5187,N_6535);
xor U8055 (N_8055,N_6147,N_7475);
and U8056 (N_8056,N_7403,N_7082);
or U8057 (N_8057,N_5661,N_6503);
nand U8058 (N_8058,N_6864,N_5431);
nand U8059 (N_8059,N_7290,N_5957);
xor U8060 (N_8060,N_6274,N_5418);
xnor U8061 (N_8061,N_6584,N_6159);
or U8062 (N_8062,N_6814,N_6086);
xnor U8063 (N_8063,N_6024,N_5350);
and U8064 (N_8064,N_7100,N_6499);
or U8065 (N_8065,N_7042,N_5723);
nor U8066 (N_8066,N_6937,N_6332);
nand U8067 (N_8067,N_7480,N_7474);
and U8068 (N_8068,N_6052,N_6426);
xnor U8069 (N_8069,N_6632,N_7154);
or U8070 (N_8070,N_7076,N_7008);
and U8071 (N_8071,N_5690,N_6452);
xor U8072 (N_8072,N_5951,N_5647);
xnor U8073 (N_8073,N_5247,N_6417);
nand U8074 (N_8074,N_5708,N_7354);
nand U8075 (N_8075,N_6971,N_5466);
nand U8076 (N_8076,N_5745,N_5982);
and U8077 (N_8077,N_5093,N_7103);
nand U8078 (N_8078,N_5439,N_5085);
nor U8079 (N_8079,N_7389,N_6574);
nor U8080 (N_8080,N_6681,N_6560);
nor U8081 (N_8081,N_5988,N_7020);
or U8082 (N_8082,N_6349,N_6978);
nor U8083 (N_8083,N_7427,N_5871);
xnor U8084 (N_8084,N_5299,N_6623);
or U8085 (N_8085,N_5949,N_6779);
nand U8086 (N_8086,N_5490,N_5959);
nor U8087 (N_8087,N_5825,N_6994);
nor U8088 (N_8088,N_5864,N_7024);
xor U8089 (N_8089,N_6189,N_5666);
xor U8090 (N_8090,N_7436,N_7061);
nor U8091 (N_8091,N_5793,N_5629);
or U8092 (N_8092,N_5259,N_5873);
xor U8093 (N_8093,N_5359,N_6682);
and U8094 (N_8094,N_5908,N_5570);
and U8095 (N_8095,N_6273,N_6920);
nand U8096 (N_8096,N_7434,N_6130);
or U8097 (N_8097,N_5340,N_6914);
xor U8098 (N_8098,N_6388,N_5348);
nand U8099 (N_8099,N_5324,N_5173);
xnor U8100 (N_8100,N_7372,N_7077);
or U8101 (N_8101,N_5548,N_6046);
nand U8102 (N_8102,N_6441,N_6599);
nand U8103 (N_8103,N_6652,N_5043);
nand U8104 (N_8104,N_6060,N_7146);
or U8105 (N_8105,N_5224,N_5066);
nand U8106 (N_8106,N_6901,N_5238);
xnor U8107 (N_8107,N_5840,N_7375);
nand U8108 (N_8108,N_7236,N_6431);
or U8109 (N_8109,N_5755,N_6931);
or U8110 (N_8110,N_6347,N_7490);
nand U8111 (N_8111,N_7343,N_5859);
nor U8112 (N_8112,N_6801,N_6991);
and U8113 (N_8113,N_6793,N_7113);
nand U8114 (N_8114,N_7379,N_7333);
nor U8115 (N_8115,N_6856,N_5644);
nand U8116 (N_8116,N_5979,N_7112);
nor U8117 (N_8117,N_5448,N_5198);
nor U8118 (N_8118,N_7066,N_6768);
and U8119 (N_8119,N_6910,N_6530);
nand U8120 (N_8120,N_5935,N_7183);
nand U8121 (N_8121,N_6963,N_6106);
xor U8122 (N_8122,N_5101,N_7484);
nand U8123 (N_8123,N_5396,N_6550);
nor U8124 (N_8124,N_7080,N_7296);
and U8125 (N_8125,N_7235,N_5843);
nor U8126 (N_8126,N_6698,N_6497);
and U8127 (N_8127,N_5254,N_6833);
and U8128 (N_8128,N_6338,N_6210);
nor U8129 (N_8129,N_6602,N_6217);
nand U8130 (N_8130,N_5360,N_5193);
nor U8131 (N_8131,N_7230,N_5557);
and U8132 (N_8132,N_5190,N_7092);
and U8133 (N_8133,N_5942,N_6115);
or U8134 (N_8134,N_6671,N_5732);
or U8135 (N_8135,N_6124,N_6137);
or U8136 (N_8136,N_5473,N_5105);
or U8137 (N_8137,N_5675,N_7481);
and U8138 (N_8138,N_5517,N_6222);
and U8139 (N_8139,N_7488,N_6077);
or U8140 (N_8140,N_6317,N_5776);
and U8141 (N_8141,N_5819,N_7209);
nand U8142 (N_8142,N_5537,N_5657);
nand U8143 (N_8143,N_5841,N_5067);
nand U8144 (N_8144,N_6491,N_6126);
or U8145 (N_8145,N_6697,N_5206);
or U8146 (N_8146,N_5642,N_5726);
or U8147 (N_8147,N_7378,N_7423);
and U8148 (N_8148,N_6166,N_6644);
nor U8149 (N_8149,N_5262,N_5290);
or U8150 (N_8150,N_6178,N_5737);
or U8151 (N_8151,N_5575,N_7166);
nor U8152 (N_8152,N_7370,N_6617);
nor U8153 (N_8153,N_5313,N_6339);
xnor U8154 (N_8154,N_5678,N_6765);
nor U8155 (N_8155,N_6135,N_5475);
nand U8156 (N_8156,N_5325,N_6335);
nand U8157 (N_8157,N_7119,N_6132);
or U8158 (N_8158,N_5973,N_6756);
nor U8159 (N_8159,N_6769,N_6459);
nor U8160 (N_8160,N_6689,N_5659);
nor U8161 (N_8161,N_7225,N_6958);
nor U8162 (N_8162,N_5110,N_5513);
nand U8163 (N_8163,N_5791,N_5301);
and U8164 (N_8164,N_7458,N_5849);
nand U8165 (N_8165,N_5738,N_6514);
xnor U8166 (N_8166,N_6755,N_7083);
nand U8167 (N_8167,N_5405,N_7324);
xnor U8168 (N_8168,N_6999,N_6049);
xnor U8169 (N_8169,N_5524,N_6325);
xor U8170 (N_8170,N_7312,N_5596);
nand U8171 (N_8171,N_5624,N_7366);
or U8172 (N_8172,N_6204,N_5910);
and U8173 (N_8173,N_5820,N_7022);
xnor U8174 (N_8174,N_7035,N_7176);
xnor U8175 (N_8175,N_7194,N_5719);
nand U8176 (N_8176,N_7047,N_7360);
nor U8177 (N_8177,N_6044,N_5651);
nor U8178 (N_8178,N_5491,N_7134);
nor U8179 (N_8179,N_6133,N_6728);
nand U8180 (N_8180,N_5140,N_5029);
or U8181 (N_8181,N_7438,N_6498);
nand U8182 (N_8182,N_6220,N_5541);
nand U8183 (N_8183,N_7169,N_6387);
or U8184 (N_8184,N_5583,N_5472);
xnor U8185 (N_8185,N_6276,N_6961);
nor U8186 (N_8186,N_5874,N_6525);
and U8187 (N_8187,N_6256,N_6302);
nor U8188 (N_8188,N_6749,N_6974);
or U8189 (N_8189,N_6733,N_7377);
xor U8190 (N_8190,N_5799,N_5486);
and U8191 (N_8191,N_6466,N_5001);
nor U8192 (N_8192,N_6152,N_6836);
and U8193 (N_8193,N_7219,N_6661);
xnor U8194 (N_8194,N_6865,N_5135);
and U8195 (N_8195,N_7161,N_6643);
or U8196 (N_8196,N_7470,N_6692);
xor U8197 (N_8197,N_5303,N_5601);
nand U8198 (N_8198,N_5283,N_6650);
nor U8199 (N_8199,N_7381,N_6611);
xnor U8200 (N_8200,N_6283,N_7195);
and U8201 (N_8201,N_7380,N_6548);
xnor U8202 (N_8202,N_7151,N_6246);
nor U8203 (N_8203,N_6816,N_5384);
nand U8204 (N_8204,N_6829,N_6573);
nand U8205 (N_8205,N_7018,N_5055);
nand U8206 (N_8206,N_6225,N_6529);
xnor U8207 (N_8207,N_6177,N_6923);
xnor U8208 (N_8208,N_7031,N_6763);
xor U8209 (N_8209,N_5488,N_5111);
or U8210 (N_8210,N_7374,N_6737);
xor U8211 (N_8211,N_5919,N_6211);
nand U8212 (N_8212,N_7295,N_6601);
and U8213 (N_8213,N_6858,N_5351);
xnor U8214 (N_8214,N_5638,N_6139);
xnor U8215 (N_8215,N_7117,N_7010);
and U8216 (N_8216,N_6084,N_7126);
nor U8217 (N_8217,N_5503,N_7459);
nor U8218 (N_8218,N_6070,N_6000);
and U8219 (N_8219,N_6542,N_5904);
and U8220 (N_8220,N_7424,N_6118);
and U8221 (N_8221,N_5230,N_6822);
nand U8222 (N_8222,N_5915,N_5011);
nor U8223 (N_8223,N_6285,N_7158);
and U8224 (N_8224,N_5007,N_5577);
xnor U8225 (N_8225,N_7213,N_6685);
nor U8226 (N_8226,N_5452,N_6531);
nand U8227 (N_8227,N_5151,N_5428);
and U8228 (N_8228,N_7118,N_5365);
or U8229 (N_8229,N_5888,N_5185);
nand U8230 (N_8230,N_7433,N_6678);
nand U8231 (N_8231,N_7247,N_6676);
nand U8232 (N_8232,N_6185,N_6532);
nand U8233 (N_8233,N_6891,N_5499);
and U8234 (N_8234,N_7025,N_6649);
or U8235 (N_8235,N_5207,N_6278);
xor U8236 (N_8236,N_6906,N_5636);
nand U8237 (N_8237,N_5197,N_7017);
nor U8238 (N_8238,N_5706,N_6455);
or U8239 (N_8239,N_7387,N_6990);
nor U8240 (N_8240,N_6326,N_5444);
or U8241 (N_8241,N_5639,N_6419);
nor U8242 (N_8242,N_5658,N_6604);
xnor U8243 (N_8243,N_5578,N_5833);
nand U8244 (N_8244,N_5257,N_5584);
nand U8245 (N_8245,N_5327,N_5595);
nor U8246 (N_8246,N_6373,N_5705);
and U8247 (N_8247,N_6824,N_5552);
nor U8248 (N_8248,N_7406,N_5751);
xor U8249 (N_8249,N_7396,N_7002);
nor U8250 (N_8250,N_6890,N_6939);
and U8251 (N_8251,N_6625,N_6427);
xor U8252 (N_8252,N_6356,N_5887);
nand U8253 (N_8253,N_6746,N_6465);
xnor U8254 (N_8254,N_6596,N_5704);
nand U8255 (N_8255,N_6439,N_5019);
or U8256 (N_8256,N_6523,N_5489);
and U8257 (N_8257,N_5251,N_5009);
xnor U8258 (N_8258,N_5754,N_5005);
or U8259 (N_8259,N_5536,N_5834);
nand U8260 (N_8260,N_6904,N_5798);
or U8261 (N_8261,N_5772,N_5865);
nor U8262 (N_8262,N_7303,N_5563);
nand U8263 (N_8263,N_6567,N_6298);
xnor U8264 (N_8264,N_7294,N_6199);
or U8265 (N_8265,N_6932,N_6341);
nand U8266 (N_8266,N_7109,N_5818);
xnor U8267 (N_8267,N_5800,N_7298);
nand U8268 (N_8268,N_7043,N_7400);
and U8269 (N_8269,N_6380,N_6168);
nand U8270 (N_8270,N_5960,N_6785);
nand U8271 (N_8271,N_5920,N_7341);
and U8272 (N_8272,N_5602,N_6946);
nand U8273 (N_8273,N_7408,N_6062);
and U8274 (N_8274,N_5686,N_5296);
xor U8275 (N_8275,N_6686,N_6213);
xnor U8276 (N_8276,N_5707,N_5962);
nor U8277 (N_8277,N_7432,N_5742);
xor U8278 (N_8278,N_5371,N_5244);
nor U8279 (N_8279,N_7412,N_5447);
and U8280 (N_8280,N_7108,N_5354);
and U8281 (N_8281,N_6146,N_6639);
xnor U8282 (N_8282,N_5787,N_6717);
and U8283 (N_8283,N_5684,N_5774);
nand U8284 (N_8284,N_6808,N_7252);
nor U8285 (N_8285,N_6423,N_6134);
nand U8286 (N_8286,N_6669,N_6457);
or U8287 (N_8287,N_6636,N_6790);
nand U8288 (N_8288,N_6725,N_6821);
or U8289 (N_8289,N_6143,N_5761);
and U8290 (N_8290,N_5769,N_6823);
xnor U8291 (N_8291,N_6528,N_7139);
nor U8292 (N_8292,N_5300,N_6066);
nor U8293 (N_8293,N_5464,N_7259);
or U8294 (N_8294,N_6323,N_6485);
and U8295 (N_8295,N_5221,N_6244);
and U8296 (N_8296,N_5355,N_6048);
nand U8297 (N_8297,N_7357,N_6743);
or U8298 (N_8298,N_6521,N_5088);
nand U8299 (N_8299,N_6019,N_5822);
or U8300 (N_8300,N_5274,N_6330);
and U8301 (N_8301,N_5752,N_5555);
nor U8302 (N_8302,N_5947,N_6926);
and U8303 (N_8303,N_5518,N_7251);
and U8304 (N_8304,N_6502,N_6074);
and U8305 (N_8305,N_6101,N_7068);
nor U8306 (N_8306,N_5826,N_5150);
xnor U8307 (N_8307,N_5363,N_5394);
and U8308 (N_8308,N_6171,N_6401);
nor U8309 (N_8309,N_6102,N_7102);
and U8310 (N_8310,N_5731,N_7455);
and U8311 (N_8311,N_5667,N_6231);
nand U8312 (N_8312,N_7013,N_5926);
nand U8313 (N_8313,N_6047,N_6016);
nor U8314 (N_8314,N_5996,N_6068);
or U8315 (N_8315,N_7263,N_7336);
nor U8316 (N_8316,N_6297,N_6734);
nor U8317 (N_8317,N_5768,N_5276);
xnor U8318 (N_8318,N_6710,N_6006);
nand U8319 (N_8319,N_5722,N_5501);
xnor U8320 (N_8320,N_7021,N_6002);
nor U8321 (N_8321,N_5421,N_5571);
or U8322 (N_8322,N_5122,N_6188);
nor U8323 (N_8323,N_5233,N_6609);
nor U8324 (N_8324,N_5923,N_5839);
and U8325 (N_8325,N_5532,N_6554);
nand U8326 (N_8326,N_6073,N_5036);
nand U8327 (N_8327,N_6249,N_6703);
and U8328 (N_8328,N_5832,N_5779);
and U8329 (N_8329,N_5279,N_6429);
nor U8330 (N_8330,N_6968,N_7282);
nand U8331 (N_8331,N_5897,N_7410);
and U8332 (N_8332,N_6582,N_5566);
and U8333 (N_8333,N_6348,N_6446);
nor U8334 (N_8334,N_6309,N_6819);
xnor U8335 (N_8335,N_5770,N_6533);
or U8336 (N_8336,N_5170,N_6874);
nand U8337 (N_8337,N_7128,N_6513);
or U8338 (N_8338,N_5278,N_5484);
and U8339 (N_8339,N_7059,N_5682);
or U8340 (N_8340,N_5014,N_7323);
or U8341 (N_8341,N_6726,N_5894);
xnor U8342 (N_8342,N_7413,N_5515);
xor U8343 (N_8343,N_6967,N_6475);
xor U8344 (N_8344,N_5023,N_6559);
and U8345 (N_8345,N_6879,N_7198);
nor U8346 (N_8346,N_7476,N_6694);
or U8347 (N_8347,N_5858,N_5188);
nand U8348 (N_8348,N_6679,N_5387);
or U8349 (N_8349,N_6358,N_5008);
nor U8350 (N_8350,N_6089,N_6516);
nor U8351 (N_8351,N_6407,N_7253);
or U8352 (N_8352,N_6117,N_5242);
xnor U8353 (N_8353,N_7335,N_7106);
and U8354 (N_8354,N_5082,N_7023);
nand U8355 (N_8355,N_7160,N_7275);
or U8356 (N_8356,N_6844,N_7292);
nand U8357 (N_8357,N_5072,N_5071);
nand U8358 (N_8358,N_5961,N_6944);
xnor U8359 (N_8359,N_5522,N_5132);
xnor U8360 (N_8360,N_6412,N_6461);
and U8361 (N_8361,N_5108,N_6591);
nor U8362 (N_8362,N_6885,N_6371);
nor U8363 (N_8363,N_7359,N_5622);
or U8364 (N_8364,N_6435,N_6965);
or U8365 (N_8365,N_5117,N_6957);
xnor U8366 (N_8366,N_5870,N_6935);
and U8367 (N_8367,N_6483,N_7026);
xor U8368 (N_8368,N_5232,N_7121);
nand U8369 (N_8369,N_5258,N_6895);
or U8370 (N_8370,N_5916,N_6020);
nand U8371 (N_8371,N_6848,N_7261);
nand U8372 (N_8372,N_5086,N_5099);
nor U8373 (N_8373,N_7346,N_5789);
nand U8374 (N_8374,N_6982,N_6547);
and U8375 (N_8375,N_6058,N_5909);
nor U8376 (N_8376,N_6357,N_6778);
or U8377 (N_8377,N_5273,N_5277);
xnor U8378 (N_8378,N_5506,N_5097);
nand U8379 (N_8379,N_6993,N_6992);
xnor U8380 (N_8380,N_6184,N_6588);
or U8381 (N_8381,N_6985,N_5089);
xor U8382 (N_8382,N_5335,N_5613);
xor U8383 (N_8383,N_5346,N_7257);
nand U8384 (N_8384,N_5587,N_6091);
or U8385 (N_8385,N_7200,N_6566);
xor U8386 (N_8386,N_6198,N_5380);
and U8387 (N_8387,N_7099,N_6451);
or U8388 (N_8388,N_6295,N_5446);
or U8389 (N_8389,N_6008,N_5109);
nor U8390 (N_8390,N_6303,N_6739);
xor U8391 (N_8391,N_7062,N_7205);
or U8392 (N_8392,N_6236,N_5423);
nand U8393 (N_8393,N_5801,N_5760);
or U8394 (N_8394,N_6713,N_7085);
xor U8395 (N_8395,N_5780,N_6941);
xor U8396 (N_8396,N_7497,N_6662);
nand U8397 (N_8397,N_5192,N_6078);
nor U8398 (N_8398,N_6674,N_5759);
nand U8399 (N_8399,N_6059,N_5480);
nand U8400 (N_8400,N_5968,N_6855);
nor U8401 (N_8401,N_6390,N_7243);
nand U8402 (N_8402,N_5383,N_7115);
nand U8403 (N_8403,N_7320,N_6056);
xnor U8404 (N_8404,N_5735,N_6011);
xor U8405 (N_8405,N_5286,N_5565);
xnor U8406 (N_8406,N_5287,N_6125);
or U8407 (N_8407,N_6336,N_7431);
or U8408 (N_8408,N_5828,N_6695);
xnor U8409 (N_8409,N_6977,N_5899);
nor U8410 (N_8410,N_6964,N_7055);
or U8411 (N_8411,N_5539,N_5877);
and U8412 (N_8412,N_5136,N_5580);
or U8413 (N_8413,N_5100,N_5379);
xnor U8414 (N_8414,N_6268,N_6868);
nor U8415 (N_8415,N_6034,N_5416);
nand U8416 (N_8416,N_5545,N_5349);
or U8417 (N_8417,N_5436,N_6320);
nand U8418 (N_8418,N_6045,N_7469);
or U8419 (N_8419,N_6265,N_6149);
or U8420 (N_8420,N_7012,N_5986);
nor U8421 (N_8421,N_7184,N_6840);
xnor U8422 (N_8422,N_7384,N_5267);
xnor U8423 (N_8423,N_5235,N_6916);
and U8424 (N_8424,N_5366,N_7342);
or U8425 (N_8425,N_7450,N_5407);
nor U8426 (N_8426,N_6954,N_5457);
and U8427 (N_8427,N_5997,N_5049);
nand U8428 (N_8428,N_5633,N_5465);
nor U8429 (N_8429,N_7065,N_7122);
or U8430 (N_8430,N_5180,N_6788);
nor U8431 (N_8431,N_5054,N_6820);
nor U8432 (N_8432,N_7337,N_7487);
or U8433 (N_8433,N_5482,N_5305);
xnor U8434 (N_8434,N_5470,N_7448);
and U8435 (N_8435,N_5012,N_5437);
and U8436 (N_8436,N_5397,N_5326);
nor U8437 (N_8437,N_7067,N_5987);
nand U8438 (N_8438,N_7150,N_5856);
and U8439 (N_8439,N_5604,N_6857);
nand U8440 (N_8440,N_5329,N_6108);
xor U8441 (N_8441,N_6107,N_6032);
nor U8442 (N_8442,N_5520,N_6660);
nand U8443 (N_8443,N_6899,N_6140);
xnor U8444 (N_8444,N_7392,N_5124);
xor U8445 (N_8445,N_5498,N_5357);
xnor U8446 (N_8446,N_5901,N_5640);
nor U8447 (N_8447,N_6180,N_6715);
xnor U8448 (N_8448,N_6099,N_5414);
nand U8449 (N_8449,N_7319,N_5605);
xnor U8450 (N_8450,N_5852,N_7203);
and U8451 (N_8451,N_7207,N_7141);
nor U8452 (N_8452,N_5805,N_5217);
nand U8453 (N_8453,N_7241,N_7038);
and U8454 (N_8454,N_7226,N_5493);
and U8455 (N_8455,N_7238,N_6576);
nor U8456 (N_8456,N_6653,N_7248);
or U8457 (N_8457,N_5775,N_5430);
nor U8458 (N_8458,N_7464,N_5056);
xnor U8459 (N_8459,N_6740,N_6425);
and U8460 (N_8460,N_6638,N_6598);
and U8461 (N_8461,N_7234,N_5469);
nor U8462 (N_8462,N_7159,N_5687);
and U8463 (N_8463,N_7220,N_6400);
nand U8464 (N_8464,N_5796,N_7216);
nand U8465 (N_8465,N_5492,N_6014);
or U8466 (N_8466,N_5628,N_6440);
nor U8467 (N_8467,N_6192,N_6705);
and U8468 (N_8468,N_6845,N_6093);
nand U8469 (N_8469,N_6504,N_6116);
xor U8470 (N_8470,N_5585,N_7070);
nor U8471 (N_8471,N_5410,N_5143);
or U8472 (N_8472,N_7149,N_6467);
nor U8473 (N_8473,N_5032,N_5922);
nand U8474 (N_8474,N_5158,N_7186);
xor U8475 (N_8475,N_6880,N_7182);
nor U8476 (N_8476,N_6015,N_7084);
or U8477 (N_8477,N_6898,N_6922);
and U8478 (N_8478,N_6262,N_5025);
xor U8479 (N_8479,N_7349,N_5065);
xnor U8480 (N_8480,N_6489,N_5216);
xor U8481 (N_8481,N_6187,N_6775);
nor U8482 (N_8482,N_7240,N_5256);
nor U8483 (N_8483,N_6072,N_5929);
nor U8484 (N_8484,N_7177,N_6606);
nand U8485 (N_8485,N_6711,N_6536);
nor U8486 (N_8486,N_5882,N_7079);
and U8487 (N_8487,N_7264,N_5179);
nand U8488 (N_8488,N_6013,N_5928);
xor U8489 (N_8489,N_5561,N_5003);
and U8490 (N_8490,N_5756,N_7382);
nand U8491 (N_8491,N_5534,N_6577);
nor U8492 (N_8492,N_6842,N_6469);
and U8493 (N_8493,N_5116,N_6878);
nand U8494 (N_8494,N_7064,N_5020);
and U8495 (N_8495,N_6569,N_6953);
xor U8496 (N_8496,N_5844,N_5218);
or U8497 (N_8497,N_6266,N_7114);
and U8498 (N_8498,N_5079,N_7386);
xor U8499 (N_8499,N_6987,N_6080);
nor U8500 (N_8500,N_6940,N_6805);
nor U8501 (N_8501,N_6506,N_6716);
nand U8502 (N_8502,N_5526,N_5549);
or U8503 (N_8503,N_6270,N_5803);
or U8504 (N_8504,N_6861,N_5002);
nor U8505 (N_8505,N_6501,N_6018);
and U8506 (N_8506,N_5544,N_6624);
nor U8507 (N_8507,N_5289,N_5668);
and U8508 (N_8508,N_5693,N_6195);
xnor U8509 (N_8509,N_6729,N_6853);
nor U8510 (N_8510,N_5884,N_7446);
nor U8511 (N_8511,N_7053,N_5215);
or U8512 (N_8512,N_5836,N_6667);
nand U8513 (N_8513,N_7430,N_6871);
and U8514 (N_8514,N_6508,N_6571);
nor U8515 (N_8515,N_7351,N_6442);
xnor U8516 (N_8516,N_6453,N_6176);
or U8517 (N_8517,N_6224,N_6421);
xnor U8518 (N_8518,N_6389,N_6787);
xnor U8519 (N_8519,N_5125,N_7032);
xor U8520 (N_8520,N_5547,N_6800);
xnor U8521 (N_8521,N_6493,N_7498);
xor U8522 (N_8522,N_6197,N_5643);
xnor U8523 (N_8523,N_5460,N_6363);
or U8524 (N_8524,N_5182,N_5261);
nand U8525 (N_8525,N_6272,N_5302);
nand U8526 (N_8526,N_6782,N_7496);
nor U8527 (N_8527,N_6736,N_5145);
and U8528 (N_8528,N_7191,N_6355);
nor U8529 (N_8529,N_5128,N_6345);
xor U8530 (N_8530,N_6437,N_5241);
nand U8531 (N_8531,N_5189,N_5454);
and U8532 (N_8532,N_6781,N_6556);
or U8533 (N_8533,N_5134,N_5607);
nand U8534 (N_8534,N_6025,N_6811);
xnor U8535 (N_8535,N_5730,N_5941);
and U8536 (N_8536,N_5784,N_6033);
nor U8537 (N_8537,N_7467,N_5203);
nand U8538 (N_8538,N_6164,N_5096);
xor U8539 (N_8539,N_5782,N_5294);
nor U8540 (N_8540,N_5388,N_7144);
or U8541 (N_8541,N_7073,N_6951);
nor U8542 (N_8542,N_7254,N_5635);
nand U8543 (N_8543,N_6832,N_5209);
and U8544 (N_8544,N_6105,N_6269);
nand U8545 (N_8545,N_5027,N_6260);
xnor U8546 (N_8546,N_5917,N_5395);
nor U8547 (N_8547,N_5804,N_7363);
and U8548 (N_8548,N_5694,N_6160);
nand U8549 (N_8549,N_6223,N_5665);
and U8550 (N_8550,N_6955,N_6004);
and U8551 (N_8551,N_7347,N_5195);
and U8552 (N_8552,N_5098,N_5133);
xnor U8553 (N_8553,N_6051,N_5721);
and U8554 (N_8554,N_6585,N_7107);
nor U8555 (N_8555,N_7048,N_5320);
and U8556 (N_8556,N_6350,N_7401);
nor U8557 (N_8557,N_7447,N_7004);
and U8558 (N_8558,N_6447,N_6175);
and U8559 (N_8559,N_6540,N_6443);
nor U8560 (N_8560,N_6551,N_6949);
nand U8561 (N_8561,N_5866,N_5617);
nor U8562 (N_8562,N_5272,N_6243);
xnor U8563 (N_8563,N_5921,N_5954);
nor U8564 (N_8564,N_7313,N_5084);
or U8565 (N_8565,N_6562,N_7466);
nor U8566 (N_8566,N_6581,N_5316);
nor U8567 (N_8567,N_5918,N_7325);
xnor U8568 (N_8568,N_7364,N_5352);
xor U8569 (N_8569,N_6507,N_6860);
xor U8570 (N_8570,N_6722,N_5573);
xor U8571 (N_8571,N_7486,N_6252);
or U8572 (N_8572,N_5308,N_7494);
nor U8573 (N_8573,N_5413,N_7429);
and U8574 (N_8574,N_6096,N_7045);
and U8575 (N_8575,N_6450,N_7179);
or U8576 (N_8576,N_5411,N_6196);
nor U8577 (N_8577,N_6182,N_6403);
or U8578 (N_8578,N_5983,N_7123);
nand U8579 (N_8579,N_6586,N_7402);
and U8580 (N_8580,N_5654,N_6334);
nor U8581 (N_8581,N_6039,N_7058);
nor U8582 (N_8582,N_7302,N_7057);
nor U8583 (N_8583,N_5409,N_5081);
nor U8584 (N_8584,N_7214,N_5697);
and U8585 (N_8585,N_7460,N_7078);
nand U8586 (N_8586,N_5938,N_5343);
nand U8587 (N_8587,N_5372,N_6849);
xnor U8588 (N_8588,N_5627,N_6082);
nand U8589 (N_8589,N_6759,N_7307);
xor U8590 (N_8590,N_5450,N_5280);
xnor U8591 (N_8591,N_5373,N_6194);
or U8592 (N_8592,N_6329,N_7036);
nand U8593 (N_8593,N_5847,N_6368);
nand U8594 (N_8594,N_6470,N_5249);
nor U8595 (N_8595,N_7163,N_5792);
and U8596 (N_8596,N_6377,N_5574);
xnor U8597 (N_8597,N_6826,N_5558);
nand U8598 (N_8598,N_7321,N_5297);
or U8599 (N_8599,N_6870,N_6233);
xor U8600 (N_8600,N_5342,N_5727);
or U8601 (N_8601,N_5115,N_7306);
and U8602 (N_8602,N_5304,N_7006);
nand U8603 (N_8603,N_5074,N_5213);
and U8604 (N_8604,N_5615,N_5568);
or U8605 (N_8605,N_5016,N_5691);
nor U8606 (N_8606,N_5445,N_6155);
and U8607 (N_8607,N_5282,N_5091);
xor U8608 (N_8608,N_6085,N_5940);
nand U8609 (N_8609,N_7297,N_6642);
nand U8610 (N_8610,N_5204,N_5650);
xnor U8611 (N_8611,N_6867,N_5827);
nor U8612 (N_8612,N_7087,N_5157);
xor U8613 (N_8613,N_6859,N_7193);
or U8614 (N_8614,N_6519,N_5594);
nand U8615 (N_8615,N_6983,N_5264);
and U8616 (N_8616,N_5964,N_7373);
nand U8617 (N_8617,N_6003,N_6659);
nand U8618 (N_8618,N_5700,N_6259);
xnor U8619 (N_8619,N_6627,N_6311);
xnor U8620 (N_8620,N_7277,N_5341);
or U8621 (N_8621,N_6866,N_6420);
or U8622 (N_8622,N_5487,N_5734);
nand U8623 (N_8623,N_7330,N_7383);
nor U8624 (N_8624,N_6534,N_5164);
xnor U8625 (N_8625,N_7356,N_6304);
nand U8626 (N_8626,N_5459,N_7309);
nor U8627 (N_8627,N_7482,N_5338);
xor U8628 (N_8628,N_6398,N_6479);
xnor U8629 (N_8629,N_6907,N_5245);
nor U8630 (N_8630,N_7462,N_6312);
nand U8631 (N_8631,N_7211,N_5039);
nor U8632 (N_8632,N_6505,N_7090);
and U8633 (N_8633,N_6700,N_7197);
nor U8634 (N_8634,N_5275,N_5156);
nor U8635 (N_8635,N_7244,N_5422);
or U8636 (N_8636,N_5406,N_7262);
xor U8637 (N_8637,N_6979,N_6228);
or U8638 (N_8638,N_7009,N_6887);
nor U8639 (N_8639,N_5616,N_5031);
nor U8640 (N_8640,N_6384,N_6803);
nand U8641 (N_8641,N_6343,N_6234);
xnor U8642 (N_8642,N_6064,N_5720);
nand U8643 (N_8643,N_6515,N_7426);
nor U8644 (N_8644,N_5144,N_7329);
nand U8645 (N_8645,N_5476,N_5226);
or U8646 (N_8646,N_7162,N_6518);
or U8647 (N_8647,N_5653,N_7041);
xnor U8648 (N_8648,N_5630,N_7493);
and U8649 (N_8649,N_6324,N_6936);
or U8650 (N_8650,N_6666,N_5995);
xnor U8651 (N_8651,N_7473,N_5334);
nand U8652 (N_8652,N_5063,N_5698);
or U8653 (N_8653,N_5663,N_6281);
nand U8654 (N_8654,N_6675,N_5400);
and U8655 (N_8655,N_6385,N_6834);
nor U8656 (N_8656,N_7318,N_6766);
and U8657 (N_8657,N_6956,N_5978);
nand U8658 (N_8658,N_5891,N_6331);
xor U8659 (N_8659,N_5312,N_6090);
or U8660 (N_8660,N_5965,N_6850);
nor U8661 (N_8661,N_7165,N_6663);
or U8662 (N_8662,N_6487,N_6873);
xnor U8663 (N_8663,N_6314,N_5710);
nand U8664 (N_8664,N_7138,N_5701);
nor U8665 (N_8665,N_5716,N_6110);
and U8666 (N_8666,N_7014,N_5609);
and U8667 (N_8667,N_5042,N_5655);
and U8668 (N_8668,N_6482,N_6658);
nor U8669 (N_8669,N_5220,N_6305);
or U8670 (N_8670,N_5912,N_6200);
and U8671 (N_8671,N_7391,N_7034);
xor U8672 (N_8672,N_6261,N_5467);
nor U8673 (N_8673,N_5292,N_6972);
or U8674 (N_8674,N_5750,N_7463);
xor U8675 (N_8675,N_5740,N_7280);
and U8676 (N_8676,N_7188,N_7019);
nor U8677 (N_8677,N_5809,N_7339);
or U8678 (N_8678,N_7148,N_6645);
or U8679 (N_8679,N_6791,N_6212);
xor U8680 (N_8680,N_5046,N_7369);
or U8681 (N_8681,N_5037,N_6605);
nor U8682 (N_8682,N_6798,N_7327);
or U8683 (N_8683,N_6835,N_5033);
or U8684 (N_8684,N_6651,N_5162);
or U8685 (N_8685,N_6886,N_6613);
nor U8686 (N_8686,N_5246,N_5152);
xnor U8687 (N_8687,N_6445,N_7284);
and U8688 (N_8688,N_5993,N_5417);
or U8689 (N_8689,N_5600,N_5933);
and U8690 (N_8690,N_5443,N_6193);
or U8691 (N_8691,N_7499,N_5356);
and U8692 (N_8692,N_5783,N_6360);
nor U8693 (N_8693,N_6545,N_5147);
nor U8694 (N_8694,N_6346,N_7175);
and U8695 (N_8695,N_7180,N_5913);
or U8696 (N_8696,N_5683,N_5519);
or U8697 (N_8697,N_5778,N_6810);
xnor U8698 (N_8698,N_6460,N_5240);
xnor U8699 (N_8699,N_6520,N_5119);
xnor U8700 (N_8700,N_6670,N_5765);
and U8701 (N_8701,N_5114,N_5777);
nor U8702 (N_8702,N_6511,N_5886);
nor U8703 (N_8703,N_7037,N_5200);
or U8704 (N_8704,N_6284,N_5451);
nor U8705 (N_8705,N_5516,N_7278);
xor U8706 (N_8706,N_5807,N_7489);
or U8707 (N_8707,N_5823,N_5885);
or U8708 (N_8708,N_6296,N_5845);
or U8709 (N_8709,N_6872,N_6989);
nand U8710 (N_8710,N_5399,N_6061);
and U8711 (N_8711,N_5829,N_5496);
or U8712 (N_8712,N_6418,N_6727);
xor U8713 (N_8713,N_6202,N_5956);
or U8714 (N_8714,N_6353,N_6752);
or U8715 (N_8715,N_7174,N_7164);
and U8716 (N_8716,N_7274,N_5637);
nand U8717 (N_8717,N_5606,N_6071);
nor U8718 (N_8718,N_6414,N_7495);
xor U8719 (N_8719,N_6997,N_6017);
nor U8720 (N_8720,N_7098,N_6424);
or U8721 (N_8721,N_6621,N_6603);
xor U8722 (N_8722,N_6839,N_6235);
nand U8723 (N_8723,N_5022,N_6876);
and U8724 (N_8724,N_5412,N_5714);
and U8725 (N_8725,N_7143,N_6730);
xnor U8726 (N_8726,N_7015,N_6079);
xnor U8727 (N_8727,N_7279,N_5531);
or U8728 (N_8728,N_5551,N_5284);
or U8729 (N_8729,N_6026,N_6127);
xnor U8730 (N_8730,N_5703,N_5976);
and U8731 (N_8731,N_5435,N_6744);
xor U8732 (N_8732,N_7007,N_6023);
xor U8733 (N_8733,N_6517,N_7316);
nand U8734 (N_8734,N_5619,N_6712);
xnor U8735 (N_8735,N_7385,N_7206);
nor U8736 (N_8736,N_5599,N_5669);
nand U8737 (N_8737,N_6557,N_7286);
or U8738 (N_8738,N_6405,N_5753);
or U8739 (N_8739,N_7208,N_5646);
nor U8740 (N_8740,N_6486,N_6654);
and U8741 (N_8741,N_6952,N_5898);
and U8742 (N_8742,N_5977,N_6313);
and U8743 (N_8743,N_5376,N_5174);
or U8744 (N_8744,N_6287,N_6041);
xor U8745 (N_8745,N_5543,N_5971);
nor U8746 (N_8746,N_6616,N_5080);
and U8747 (N_8747,N_5781,N_6984);
nor U8748 (N_8748,N_5364,N_5790);
xor U8749 (N_8749,N_7096,N_6208);
or U8750 (N_8750,N_5285,N_6522);
xnor U8751 (N_8751,N_7173,N_6033);
xor U8752 (N_8752,N_5038,N_7254);
nand U8753 (N_8753,N_5724,N_5435);
or U8754 (N_8754,N_5839,N_5630);
or U8755 (N_8755,N_5672,N_6867);
nor U8756 (N_8756,N_7271,N_6335);
nand U8757 (N_8757,N_6081,N_7045);
xor U8758 (N_8758,N_7280,N_7400);
and U8759 (N_8759,N_5932,N_7342);
nand U8760 (N_8760,N_5034,N_7437);
nor U8761 (N_8761,N_5851,N_7145);
nor U8762 (N_8762,N_6656,N_6406);
nand U8763 (N_8763,N_6109,N_6334);
xor U8764 (N_8764,N_5783,N_7458);
nor U8765 (N_8765,N_6491,N_7370);
xor U8766 (N_8766,N_6407,N_6202);
nor U8767 (N_8767,N_5562,N_6945);
nand U8768 (N_8768,N_6181,N_6049);
nand U8769 (N_8769,N_5890,N_6476);
and U8770 (N_8770,N_6194,N_5563);
xor U8771 (N_8771,N_5603,N_5431);
and U8772 (N_8772,N_5854,N_6564);
or U8773 (N_8773,N_7054,N_5169);
xnor U8774 (N_8774,N_5399,N_6367);
nand U8775 (N_8775,N_5973,N_5500);
and U8776 (N_8776,N_7458,N_5989);
nand U8777 (N_8777,N_5973,N_7034);
nor U8778 (N_8778,N_7044,N_5653);
nand U8779 (N_8779,N_7104,N_7036);
xor U8780 (N_8780,N_6472,N_5017);
or U8781 (N_8781,N_6838,N_5208);
or U8782 (N_8782,N_7000,N_5471);
or U8783 (N_8783,N_7408,N_6757);
or U8784 (N_8784,N_6759,N_5445);
xor U8785 (N_8785,N_5595,N_5800);
and U8786 (N_8786,N_5520,N_7468);
and U8787 (N_8787,N_5209,N_6372);
or U8788 (N_8788,N_7050,N_6672);
nand U8789 (N_8789,N_5326,N_6989);
or U8790 (N_8790,N_6701,N_5155);
nand U8791 (N_8791,N_7128,N_5746);
or U8792 (N_8792,N_6706,N_5411);
nor U8793 (N_8793,N_5881,N_5716);
and U8794 (N_8794,N_6580,N_6081);
and U8795 (N_8795,N_7293,N_7207);
nand U8796 (N_8796,N_5558,N_6558);
nor U8797 (N_8797,N_6903,N_5200);
nand U8798 (N_8798,N_5436,N_6580);
nor U8799 (N_8799,N_5664,N_6204);
or U8800 (N_8800,N_6614,N_6551);
nand U8801 (N_8801,N_6744,N_6962);
or U8802 (N_8802,N_7329,N_6628);
or U8803 (N_8803,N_6155,N_6083);
nor U8804 (N_8804,N_7482,N_5581);
or U8805 (N_8805,N_6404,N_6893);
and U8806 (N_8806,N_6333,N_5676);
nand U8807 (N_8807,N_5041,N_6334);
xor U8808 (N_8808,N_5996,N_5194);
and U8809 (N_8809,N_5496,N_5521);
xor U8810 (N_8810,N_7322,N_6460);
nand U8811 (N_8811,N_5729,N_6687);
and U8812 (N_8812,N_5259,N_6904);
or U8813 (N_8813,N_5791,N_5089);
nor U8814 (N_8814,N_5615,N_5625);
xor U8815 (N_8815,N_6462,N_5439);
nor U8816 (N_8816,N_6766,N_7445);
and U8817 (N_8817,N_6749,N_5988);
xnor U8818 (N_8818,N_6114,N_6680);
nand U8819 (N_8819,N_7089,N_7298);
nor U8820 (N_8820,N_6522,N_7204);
and U8821 (N_8821,N_5035,N_5847);
nor U8822 (N_8822,N_5208,N_7374);
xor U8823 (N_8823,N_6999,N_5557);
nor U8824 (N_8824,N_7328,N_5579);
nor U8825 (N_8825,N_5876,N_6216);
or U8826 (N_8826,N_7107,N_5369);
xor U8827 (N_8827,N_6674,N_5084);
xnor U8828 (N_8828,N_5053,N_5747);
nand U8829 (N_8829,N_5501,N_5824);
or U8830 (N_8830,N_6944,N_5605);
xnor U8831 (N_8831,N_6835,N_6154);
xnor U8832 (N_8832,N_5205,N_7239);
nand U8833 (N_8833,N_5353,N_6024);
or U8834 (N_8834,N_5679,N_6568);
nor U8835 (N_8835,N_5238,N_6139);
nor U8836 (N_8836,N_6848,N_7040);
xor U8837 (N_8837,N_6650,N_6903);
nor U8838 (N_8838,N_6518,N_5382);
xor U8839 (N_8839,N_6417,N_6574);
nand U8840 (N_8840,N_6759,N_6666);
or U8841 (N_8841,N_6736,N_6517);
nor U8842 (N_8842,N_7316,N_6518);
and U8843 (N_8843,N_5214,N_5312);
nand U8844 (N_8844,N_6367,N_5319);
and U8845 (N_8845,N_5496,N_5107);
or U8846 (N_8846,N_5182,N_6166);
nor U8847 (N_8847,N_7383,N_5379);
xor U8848 (N_8848,N_6195,N_5192);
nand U8849 (N_8849,N_6868,N_6860);
nor U8850 (N_8850,N_5668,N_5150);
and U8851 (N_8851,N_5336,N_7237);
or U8852 (N_8852,N_6664,N_6464);
and U8853 (N_8853,N_5530,N_6127);
and U8854 (N_8854,N_6885,N_6928);
nor U8855 (N_8855,N_7471,N_5253);
nor U8856 (N_8856,N_5069,N_6995);
xor U8857 (N_8857,N_5907,N_6177);
and U8858 (N_8858,N_7280,N_5286);
nor U8859 (N_8859,N_5628,N_6477);
nor U8860 (N_8860,N_5291,N_6137);
xnor U8861 (N_8861,N_6626,N_5369);
nand U8862 (N_8862,N_7154,N_6818);
nor U8863 (N_8863,N_6765,N_5134);
or U8864 (N_8864,N_6340,N_6262);
or U8865 (N_8865,N_5436,N_7040);
and U8866 (N_8866,N_6524,N_5541);
xnor U8867 (N_8867,N_6124,N_5914);
and U8868 (N_8868,N_5673,N_7100);
nor U8869 (N_8869,N_6560,N_5476);
and U8870 (N_8870,N_5628,N_7227);
and U8871 (N_8871,N_6477,N_6333);
and U8872 (N_8872,N_6986,N_7197);
and U8873 (N_8873,N_5087,N_5919);
and U8874 (N_8874,N_7241,N_6417);
or U8875 (N_8875,N_6497,N_7093);
or U8876 (N_8876,N_6767,N_5872);
nand U8877 (N_8877,N_5175,N_5613);
nor U8878 (N_8878,N_5448,N_6715);
nor U8879 (N_8879,N_6466,N_6186);
xor U8880 (N_8880,N_5864,N_5142);
xor U8881 (N_8881,N_7451,N_5828);
nor U8882 (N_8882,N_6983,N_7111);
xor U8883 (N_8883,N_5245,N_5994);
and U8884 (N_8884,N_5012,N_6760);
and U8885 (N_8885,N_6163,N_5256);
nand U8886 (N_8886,N_7336,N_6533);
or U8887 (N_8887,N_7451,N_5638);
nand U8888 (N_8888,N_7089,N_5199);
nand U8889 (N_8889,N_6217,N_6259);
nor U8890 (N_8890,N_6627,N_5467);
xor U8891 (N_8891,N_6879,N_6187);
nand U8892 (N_8892,N_5328,N_6153);
nand U8893 (N_8893,N_5032,N_5318);
nor U8894 (N_8894,N_5475,N_6795);
and U8895 (N_8895,N_6111,N_6450);
xnor U8896 (N_8896,N_6989,N_6643);
nand U8897 (N_8897,N_6594,N_6984);
xnor U8898 (N_8898,N_7187,N_6005);
xnor U8899 (N_8899,N_6215,N_6068);
nand U8900 (N_8900,N_6248,N_6499);
nor U8901 (N_8901,N_7471,N_5983);
nand U8902 (N_8902,N_6375,N_5444);
nor U8903 (N_8903,N_6481,N_5108);
and U8904 (N_8904,N_7131,N_5689);
nand U8905 (N_8905,N_7217,N_5155);
xnor U8906 (N_8906,N_5398,N_5275);
nor U8907 (N_8907,N_5342,N_6686);
or U8908 (N_8908,N_6097,N_6253);
or U8909 (N_8909,N_6081,N_6334);
or U8910 (N_8910,N_7138,N_6759);
nor U8911 (N_8911,N_7040,N_6334);
or U8912 (N_8912,N_5372,N_7430);
and U8913 (N_8913,N_6866,N_7104);
and U8914 (N_8914,N_6144,N_6173);
nor U8915 (N_8915,N_6707,N_5538);
xnor U8916 (N_8916,N_6596,N_5351);
and U8917 (N_8917,N_7229,N_5803);
or U8918 (N_8918,N_7282,N_5649);
and U8919 (N_8919,N_5129,N_5810);
xor U8920 (N_8920,N_6417,N_5585);
or U8921 (N_8921,N_5970,N_5476);
and U8922 (N_8922,N_6491,N_6750);
or U8923 (N_8923,N_6778,N_6558);
nor U8924 (N_8924,N_5914,N_7337);
xor U8925 (N_8925,N_6540,N_5216);
and U8926 (N_8926,N_5238,N_5166);
xor U8927 (N_8927,N_5872,N_7409);
or U8928 (N_8928,N_6222,N_6777);
or U8929 (N_8929,N_6254,N_5278);
nand U8930 (N_8930,N_6907,N_5366);
and U8931 (N_8931,N_6868,N_5208);
and U8932 (N_8932,N_6555,N_6263);
or U8933 (N_8933,N_6405,N_5344);
nand U8934 (N_8934,N_7225,N_6963);
nor U8935 (N_8935,N_5476,N_6909);
and U8936 (N_8936,N_5025,N_6647);
and U8937 (N_8937,N_6105,N_6968);
and U8938 (N_8938,N_6023,N_5151);
nand U8939 (N_8939,N_5555,N_7065);
nor U8940 (N_8940,N_5558,N_6411);
xnor U8941 (N_8941,N_6697,N_7379);
xor U8942 (N_8942,N_6747,N_7387);
nor U8943 (N_8943,N_6335,N_7287);
xor U8944 (N_8944,N_7031,N_5382);
nor U8945 (N_8945,N_6499,N_7394);
or U8946 (N_8946,N_6603,N_7499);
xor U8947 (N_8947,N_6163,N_5904);
or U8948 (N_8948,N_5152,N_7053);
xnor U8949 (N_8949,N_6653,N_6451);
xnor U8950 (N_8950,N_6696,N_5738);
or U8951 (N_8951,N_6152,N_6911);
nor U8952 (N_8952,N_6843,N_7055);
and U8953 (N_8953,N_7047,N_6088);
xor U8954 (N_8954,N_6691,N_6968);
or U8955 (N_8955,N_6425,N_6033);
nand U8956 (N_8956,N_5012,N_6235);
and U8957 (N_8957,N_7254,N_5839);
nand U8958 (N_8958,N_7284,N_5687);
nand U8959 (N_8959,N_6640,N_6142);
nand U8960 (N_8960,N_7344,N_5415);
or U8961 (N_8961,N_5935,N_5550);
xnor U8962 (N_8962,N_7350,N_5486);
or U8963 (N_8963,N_7252,N_5790);
and U8964 (N_8964,N_5410,N_6368);
xor U8965 (N_8965,N_5067,N_6674);
nand U8966 (N_8966,N_7401,N_5528);
xor U8967 (N_8967,N_6569,N_6327);
nand U8968 (N_8968,N_6109,N_5208);
nor U8969 (N_8969,N_6470,N_5947);
and U8970 (N_8970,N_6035,N_5926);
xnor U8971 (N_8971,N_5366,N_6679);
nand U8972 (N_8972,N_7302,N_7300);
or U8973 (N_8973,N_6972,N_6367);
and U8974 (N_8974,N_5991,N_6139);
nand U8975 (N_8975,N_6990,N_5142);
and U8976 (N_8976,N_7443,N_7212);
and U8977 (N_8977,N_7236,N_5144);
nand U8978 (N_8978,N_7406,N_6283);
and U8979 (N_8979,N_7397,N_5280);
nand U8980 (N_8980,N_6300,N_6533);
nand U8981 (N_8981,N_5740,N_6881);
nand U8982 (N_8982,N_6392,N_5660);
and U8983 (N_8983,N_6955,N_6334);
and U8984 (N_8984,N_5096,N_5335);
xor U8985 (N_8985,N_6323,N_5738);
and U8986 (N_8986,N_7425,N_6947);
and U8987 (N_8987,N_5680,N_5620);
and U8988 (N_8988,N_5084,N_5679);
nor U8989 (N_8989,N_5985,N_6616);
and U8990 (N_8990,N_6539,N_7430);
xor U8991 (N_8991,N_6687,N_5798);
nand U8992 (N_8992,N_5389,N_5532);
and U8993 (N_8993,N_6714,N_6425);
xnor U8994 (N_8994,N_5158,N_5073);
and U8995 (N_8995,N_5791,N_6126);
xnor U8996 (N_8996,N_5649,N_6713);
or U8997 (N_8997,N_7304,N_6690);
nand U8998 (N_8998,N_5046,N_6188);
or U8999 (N_8999,N_6319,N_6609);
nand U9000 (N_9000,N_6998,N_5357);
nand U9001 (N_9001,N_5342,N_6482);
xnor U9002 (N_9002,N_7498,N_6243);
nand U9003 (N_9003,N_6315,N_7372);
or U9004 (N_9004,N_6115,N_5931);
or U9005 (N_9005,N_5683,N_5487);
nor U9006 (N_9006,N_7336,N_7348);
or U9007 (N_9007,N_5590,N_6127);
or U9008 (N_9008,N_6322,N_7021);
or U9009 (N_9009,N_6667,N_5842);
or U9010 (N_9010,N_5235,N_6111);
nand U9011 (N_9011,N_5043,N_5449);
and U9012 (N_9012,N_6254,N_6053);
xnor U9013 (N_9013,N_6928,N_7122);
and U9014 (N_9014,N_5466,N_6717);
nor U9015 (N_9015,N_5487,N_6457);
and U9016 (N_9016,N_6817,N_5130);
or U9017 (N_9017,N_6529,N_6082);
or U9018 (N_9018,N_7253,N_6604);
xor U9019 (N_9019,N_7206,N_6124);
nor U9020 (N_9020,N_5588,N_6017);
or U9021 (N_9021,N_6612,N_6825);
xor U9022 (N_9022,N_5741,N_7292);
and U9023 (N_9023,N_5801,N_5557);
and U9024 (N_9024,N_6986,N_5690);
and U9025 (N_9025,N_7010,N_7463);
nand U9026 (N_9026,N_6783,N_5147);
nor U9027 (N_9027,N_6808,N_6181);
nor U9028 (N_9028,N_6569,N_7363);
nor U9029 (N_9029,N_7194,N_5329);
and U9030 (N_9030,N_5187,N_7146);
xor U9031 (N_9031,N_7313,N_5919);
xnor U9032 (N_9032,N_5174,N_7258);
nor U9033 (N_9033,N_7124,N_7011);
nand U9034 (N_9034,N_6450,N_6181);
nor U9035 (N_9035,N_5483,N_5321);
nand U9036 (N_9036,N_7049,N_6452);
xor U9037 (N_9037,N_6366,N_6381);
nor U9038 (N_9038,N_6370,N_5508);
nand U9039 (N_9039,N_5968,N_6213);
nand U9040 (N_9040,N_7467,N_5139);
xor U9041 (N_9041,N_6481,N_6617);
nand U9042 (N_9042,N_5871,N_5397);
or U9043 (N_9043,N_7175,N_6424);
or U9044 (N_9044,N_5776,N_5983);
xor U9045 (N_9045,N_6245,N_5693);
nor U9046 (N_9046,N_6406,N_7005);
xnor U9047 (N_9047,N_5594,N_7112);
xor U9048 (N_9048,N_5743,N_7457);
or U9049 (N_9049,N_6100,N_6544);
nor U9050 (N_9050,N_5780,N_6176);
xnor U9051 (N_9051,N_6942,N_6119);
nor U9052 (N_9052,N_6681,N_5497);
nor U9053 (N_9053,N_6334,N_5367);
nor U9054 (N_9054,N_5053,N_7043);
nor U9055 (N_9055,N_6648,N_6487);
nor U9056 (N_9056,N_7035,N_5140);
xnor U9057 (N_9057,N_7062,N_5289);
xnor U9058 (N_9058,N_7432,N_5983);
or U9059 (N_9059,N_5815,N_7260);
nand U9060 (N_9060,N_6786,N_6705);
nand U9061 (N_9061,N_5709,N_6423);
or U9062 (N_9062,N_6109,N_7218);
xor U9063 (N_9063,N_6705,N_6817);
nor U9064 (N_9064,N_5670,N_7242);
xor U9065 (N_9065,N_6427,N_6495);
nor U9066 (N_9066,N_5660,N_5178);
nand U9067 (N_9067,N_5532,N_5265);
and U9068 (N_9068,N_5807,N_7126);
and U9069 (N_9069,N_6318,N_5074);
nand U9070 (N_9070,N_5170,N_6966);
and U9071 (N_9071,N_5829,N_5832);
nor U9072 (N_9072,N_5770,N_6073);
xnor U9073 (N_9073,N_5648,N_7311);
or U9074 (N_9074,N_7468,N_6858);
nor U9075 (N_9075,N_5159,N_5447);
nand U9076 (N_9076,N_5489,N_5950);
nor U9077 (N_9077,N_5172,N_6304);
nand U9078 (N_9078,N_5444,N_7154);
and U9079 (N_9079,N_5288,N_6124);
nand U9080 (N_9080,N_6458,N_7185);
nor U9081 (N_9081,N_5863,N_5697);
nand U9082 (N_9082,N_6370,N_6042);
and U9083 (N_9083,N_5212,N_5692);
nor U9084 (N_9084,N_7449,N_7489);
or U9085 (N_9085,N_5305,N_5347);
nand U9086 (N_9086,N_5356,N_6518);
and U9087 (N_9087,N_5282,N_6283);
nand U9088 (N_9088,N_6480,N_5026);
xor U9089 (N_9089,N_6698,N_5153);
nand U9090 (N_9090,N_5792,N_6917);
nor U9091 (N_9091,N_7468,N_5437);
and U9092 (N_9092,N_5944,N_5387);
or U9093 (N_9093,N_5662,N_5298);
or U9094 (N_9094,N_5650,N_5113);
nand U9095 (N_9095,N_7423,N_6871);
nand U9096 (N_9096,N_7190,N_6574);
nor U9097 (N_9097,N_5553,N_5090);
xor U9098 (N_9098,N_5542,N_5665);
or U9099 (N_9099,N_5834,N_6266);
nor U9100 (N_9100,N_6408,N_7048);
xnor U9101 (N_9101,N_7474,N_6133);
nand U9102 (N_9102,N_6505,N_5757);
nor U9103 (N_9103,N_7139,N_5667);
nand U9104 (N_9104,N_5546,N_6912);
and U9105 (N_9105,N_7032,N_6246);
and U9106 (N_9106,N_5402,N_5980);
xnor U9107 (N_9107,N_7250,N_6581);
nor U9108 (N_9108,N_5510,N_5283);
nor U9109 (N_9109,N_6998,N_6800);
nand U9110 (N_9110,N_6567,N_5987);
and U9111 (N_9111,N_7202,N_7323);
and U9112 (N_9112,N_7215,N_6754);
or U9113 (N_9113,N_6202,N_5801);
nand U9114 (N_9114,N_5548,N_5765);
xor U9115 (N_9115,N_5406,N_7446);
or U9116 (N_9116,N_5552,N_5975);
or U9117 (N_9117,N_7018,N_6819);
nand U9118 (N_9118,N_7316,N_5501);
or U9119 (N_9119,N_7297,N_6059);
xor U9120 (N_9120,N_5964,N_6427);
or U9121 (N_9121,N_5725,N_5095);
and U9122 (N_9122,N_5051,N_6019);
nor U9123 (N_9123,N_7268,N_6738);
or U9124 (N_9124,N_6414,N_5558);
nand U9125 (N_9125,N_5658,N_6997);
and U9126 (N_9126,N_5499,N_5774);
or U9127 (N_9127,N_6395,N_7427);
xor U9128 (N_9128,N_7380,N_5380);
nor U9129 (N_9129,N_6224,N_7492);
nor U9130 (N_9130,N_5637,N_5542);
xor U9131 (N_9131,N_5131,N_7147);
xor U9132 (N_9132,N_7081,N_5898);
xnor U9133 (N_9133,N_6454,N_7339);
nand U9134 (N_9134,N_7061,N_6681);
and U9135 (N_9135,N_7204,N_6841);
and U9136 (N_9136,N_7154,N_7332);
and U9137 (N_9137,N_6536,N_5266);
or U9138 (N_9138,N_6204,N_5266);
nand U9139 (N_9139,N_6661,N_5538);
or U9140 (N_9140,N_6993,N_5776);
nand U9141 (N_9141,N_6202,N_7233);
xor U9142 (N_9142,N_6686,N_6680);
nand U9143 (N_9143,N_5449,N_7162);
xnor U9144 (N_9144,N_5882,N_7304);
and U9145 (N_9145,N_7301,N_6729);
or U9146 (N_9146,N_6699,N_5194);
xor U9147 (N_9147,N_7445,N_6197);
nand U9148 (N_9148,N_5626,N_5788);
and U9149 (N_9149,N_5833,N_5107);
or U9150 (N_9150,N_6627,N_5047);
or U9151 (N_9151,N_6598,N_5370);
nand U9152 (N_9152,N_5900,N_5700);
or U9153 (N_9153,N_7178,N_7057);
xnor U9154 (N_9154,N_6222,N_5624);
or U9155 (N_9155,N_7441,N_6495);
or U9156 (N_9156,N_7230,N_5160);
and U9157 (N_9157,N_7245,N_5853);
xnor U9158 (N_9158,N_5036,N_5466);
nor U9159 (N_9159,N_6040,N_5232);
and U9160 (N_9160,N_5756,N_5362);
or U9161 (N_9161,N_5854,N_5321);
and U9162 (N_9162,N_7269,N_7452);
and U9163 (N_9163,N_6197,N_5258);
or U9164 (N_9164,N_5864,N_5873);
nand U9165 (N_9165,N_6841,N_6285);
and U9166 (N_9166,N_6205,N_5128);
nor U9167 (N_9167,N_6344,N_6738);
and U9168 (N_9168,N_5488,N_5000);
xor U9169 (N_9169,N_5590,N_5609);
nor U9170 (N_9170,N_5858,N_7388);
nor U9171 (N_9171,N_5711,N_6629);
and U9172 (N_9172,N_6589,N_5989);
nand U9173 (N_9173,N_6796,N_5996);
xnor U9174 (N_9174,N_6193,N_6450);
and U9175 (N_9175,N_5069,N_7010);
xor U9176 (N_9176,N_5708,N_5984);
nand U9177 (N_9177,N_7123,N_5263);
or U9178 (N_9178,N_5676,N_6651);
and U9179 (N_9179,N_7118,N_6859);
nand U9180 (N_9180,N_6273,N_5672);
or U9181 (N_9181,N_6511,N_6714);
or U9182 (N_9182,N_5544,N_7289);
nor U9183 (N_9183,N_5764,N_6172);
nand U9184 (N_9184,N_6007,N_5317);
nor U9185 (N_9185,N_7070,N_6635);
and U9186 (N_9186,N_6907,N_6756);
nand U9187 (N_9187,N_5550,N_6627);
nor U9188 (N_9188,N_5651,N_5150);
xnor U9189 (N_9189,N_6091,N_6674);
nand U9190 (N_9190,N_5921,N_6953);
nor U9191 (N_9191,N_6226,N_5610);
and U9192 (N_9192,N_5165,N_7430);
nor U9193 (N_9193,N_6957,N_6259);
xor U9194 (N_9194,N_7441,N_5078);
nand U9195 (N_9195,N_5648,N_7276);
and U9196 (N_9196,N_6020,N_6041);
xor U9197 (N_9197,N_5018,N_5834);
xor U9198 (N_9198,N_6322,N_7035);
and U9199 (N_9199,N_5867,N_5635);
nor U9200 (N_9200,N_6904,N_5213);
nand U9201 (N_9201,N_5600,N_5509);
nor U9202 (N_9202,N_5117,N_5399);
nand U9203 (N_9203,N_7412,N_7154);
or U9204 (N_9204,N_6654,N_7314);
and U9205 (N_9205,N_5621,N_5129);
xnor U9206 (N_9206,N_5975,N_6552);
nand U9207 (N_9207,N_6535,N_6628);
nor U9208 (N_9208,N_6862,N_5012);
nor U9209 (N_9209,N_6495,N_5765);
and U9210 (N_9210,N_5528,N_6361);
and U9211 (N_9211,N_7191,N_5107);
nand U9212 (N_9212,N_5341,N_6338);
nor U9213 (N_9213,N_6216,N_5361);
nor U9214 (N_9214,N_6543,N_5186);
or U9215 (N_9215,N_5331,N_5065);
nand U9216 (N_9216,N_5652,N_6563);
nand U9217 (N_9217,N_6977,N_6009);
xnor U9218 (N_9218,N_6933,N_7319);
nor U9219 (N_9219,N_6461,N_5423);
xor U9220 (N_9220,N_6683,N_5909);
and U9221 (N_9221,N_5602,N_6250);
and U9222 (N_9222,N_7131,N_6371);
nand U9223 (N_9223,N_6942,N_5915);
nand U9224 (N_9224,N_6450,N_5647);
nor U9225 (N_9225,N_7367,N_5080);
nor U9226 (N_9226,N_6540,N_6390);
xnor U9227 (N_9227,N_7140,N_5466);
xor U9228 (N_9228,N_5640,N_6650);
xnor U9229 (N_9229,N_5346,N_7321);
and U9230 (N_9230,N_6252,N_6360);
or U9231 (N_9231,N_6229,N_6600);
and U9232 (N_9232,N_7230,N_5353);
nand U9233 (N_9233,N_5171,N_6094);
or U9234 (N_9234,N_6717,N_5744);
and U9235 (N_9235,N_6873,N_5232);
and U9236 (N_9236,N_6484,N_5000);
nand U9237 (N_9237,N_7022,N_5814);
xnor U9238 (N_9238,N_6714,N_6936);
nand U9239 (N_9239,N_6314,N_6841);
nor U9240 (N_9240,N_5113,N_6036);
xor U9241 (N_9241,N_6120,N_7248);
or U9242 (N_9242,N_6489,N_6353);
xnor U9243 (N_9243,N_6812,N_7271);
xor U9244 (N_9244,N_6101,N_7398);
nand U9245 (N_9245,N_6270,N_5685);
nand U9246 (N_9246,N_5701,N_5020);
or U9247 (N_9247,N_6607,N_6067);
nand U9248 (N_9248,N_5150,N_7280);
nor U9249 (N_9249,N_6816,N_6974);
and U9250 (N_9250,N_6397,N_6386);
or U9251 (N_9251,N_7298,N_6065);
or U9252 (N_9252,N_6211,N_5072);
nor U9253 (N_9253,N_6416,N_5375);
and U9254 (N_9254,N_5304,N_6981);
xnor U9255 (N_9255,N_6701,N_7005);
nand U9256 (N_9256,N_5123,N_5587);
and U9257 (N_9257,N_7199,N_5633);
nand U9258 (N_9258,N_6627,N_6984);
nand U9259 (N_9259,N_5785,N_6244);
and U9260 (N_9260,N_5148,N_7180);
nor U9261 (N_9261,N_5049,N_6378);
xnor U9262 (N_9262,N_7121,N_5939);
xor U9263 (N_9263,N_7493,N_5426);
xnor U9264 (N_9264,N_6033,N_6168);
nor U9265 (N_9265,N_6649,N_5900);
xnor U9266 (N_9266,N_7188,N_5818);
xnor U9267 (N_9267,N_6363,N_5188);
or U9268 (N_9268,N_6403,N_7225);
nand U9269 (N_9269,N_5742,N_5745);
xnor U9270 (N_9270,N_7167,N_5648);
xor U9271 (N_9271,N_5360,N_7108);
and U9272 (N_9272,N_5693,N_6959);
or U9273 (N_9273,N_5093,N_6902);
and U9274 (N_9274,N_5209,N_5932);
or U9275 (N_9275,N_6916,N_7011);
or U9276 (N_9276,N_6958,N_5054);
nor U9277 (N_9277,N_7408,N_5697);
xnor U9278 (N_9278,N_5450,N_6482);
xnor U9279 (N_9279,N_6394,N_5763);
nor U9280 (N_9280,N_6560,N_6235);
nor U9281 (N_9281,N_5927,N_5233);
nand U9282 (N_9282,N_6230,N_7433);
and U9283 (N_9283,N_5674,N_5214);
xor U9284 (N_9284,N_5614,N_7396);
xor U9285 (N_9285,N_5842,N_7421);
nand U9286 (N_9286,N_5950,N_5297);
nor U9287 (N_9287,N_5352,N_6461);
or U9288 (N_9288,N_7255,N_5066);
or U9289 (N_9289,N_5980,N_5736);
xnor U9290 (N_9290,N_6785,N_6322);
or U9291 (N_9291,N_5560,N_7232);
nor U9292 (N_9292,N_5853,N_6029);
nand U9293 (N_9293,N_6111,N_6093);
xor U9294 (N_9294,N_6206,N_5219);
xor U9295 (N_9295,N_7170,N_5724);
and U9296 (N_9296,N_7037,N_6492);
nor U9297 (N_9297,N_6553,N_5420);
or U9298 (N_9298,N_5545,N_6171);
nand U9299 (N_9299,N_6435,N_5357);
nand U9300 (N_9300,N_5033,N_7025);
or U9301 (N_9301,N_6554,N_5005);
xor U9302 (N_9302,N_5171,N_6029);
nor U9303 (N_9303,N_5247,N_6329);
nor U9304 (N_9304,N_6312,N_6320);
or U9305 (N_9305,N_6864,N_6593);
and U9306 (N_9306,N_6248,N_6582);
xor U9307 (N_9307,N_5919,N_6239);
nand U9308 (N_9308,N_7469,N_7014);
xor U9309 (N_9309,N_5911,N_5750);
nor U9310 (N_9310,N_6206,N_6577);
nor U9311 (N_9311,N_7292,N_5327);
nand U9312 (N_9312,N_7100,N_5265);
and U9313 (N_9313,N_5523,N_6434);
and U9314 (N_9314,N_7135,N_5363);
nor U9315 (N_9315,N_6551,N_6715);
or U9316 (N_9316,N_6882,N_5431);
xnor U9317 (N_9317,N_6163,N_7292);
nand U9318 (N_9318,N_5645,N_7043);
nand U9319 (N_9319,N_7447,N_5235);
or U9320 (N_9320,N_7345,N_7355);
or U9321 (N_9321,N_6300,N_7451);
and U9322 (N_9322,N_7240,N_6592);
nand U9323 (N_9323,N_6143,N_6393);
and U9324 (N_9324,N_6279,N_6694);
nor U9325 (N_9325,N_5647,N_7191);
and U9326 (N_9326,N_5988,N_5530);
and U9327 (N_9327,N_6770,N_5837);
and U9328 (N_9328,N_7321,N_7189);
nand U9329 (N_9329,N_5675,N_5993);
or U9330 (N_9330,N_5200,N_5632);
nand U9331 (N_9331,N_5405,N_5790);
and U9332 (N_9332,N_6907,N_6604);
xor U9333 (N_9333,N_5331,N_7448);
nor U9334 (N_9334,N_7373,N_7408);
and U9335 (N_9335,N_5545,N_6635);
and U9336 (N_9336,N_7197,N_7339);
and U9337 (N_9337,N_6683,N_6884);
and U9338 (N_9338,N_7318,N_5104);
and U9339 (N_9339,N_6373,N_6671);
nor U9340 (N_9340,N_5430,N_7219);
nor U9341 (N_9341,N_6897,N_7087);
nand U9342 (N_9342,N_7160,N_7091);
nand U9343 (N_9343,N_7303,N_5777);
nand U9344 (N_9344,N_7284,N_5495);
nand U9345 (N_9345,N_5508,N_6722);
nand U9346 (N_9346,N_5510,N_6438);
nand U9347 (N_9347,N_5692,N_5366);
and U9348 (N_9348,N_5282,N_7385);
xor U9349 (N_9349,N_7062,N_6784);
xnor U9350 (N_9350,N_7174,N_7236);
and U9351 (N_9351,N_5821,N_6199);
xor U9352 (N_9352,N_6291,N_6715);
nand U9353 (N_9353,N_5493,N_7183);
or U9354 (N_9354,N_6004,N_7364);
and U9355 (N_9355,N_6875,N_5059);
nor U9356 (N_9356,N_7050,N_7085);
and U9357 (N_9357,N_6056,N_5580);
and U9358 (N_9358,N_6140,N_6698);
or U9359 (N_9359,N_6122,N_7350);
nor U9360 (N_9360,N_7100,N_5983);
nand U9361 (N_9361,N_6509,N_6549);
and U9362 (N_9362,N_5604,N_6820);
and U9363 (N_9363,N_7120,N_5564);
xnor U9364 (N_9364,N_6987,N_7209);
xnor U9365 (N_9365,N_7097,N_6862);
nand U9366 (N_9366,N_5220,N_5552);
or U9367 (N_9367,N_6975,N_6388);
and U9368 (N_9368,N_7307,N_6096);
or U9369 (N_9369,N_5133,N_5082);
nand U9370 (N_9370,N_5482,N_6903);
and U9371 (N_9371,N_6063,N_7264);
nand U9372 (N_9372,N_6810,N_5040);
xnor U9373 (N_9373,N_6049,N_7356);
xnor U9374 (N_9374,N_6799,N_5836);
nor U9375 (N_9375,N_6889,N_6401);
nand U9376 (N_9376,N_7104,N_6024);
and U9377 (N_9377,N_6409,N_5122);
nor U9378 (N_9378,N_5324,N_6922);
or U9379 (N_9379,N_7036,N_6246);
and U9380 (N_9380,N_6823,N_5819);
and U9381 (N_9381,N_5262,N_7324);
xor U9382 (N_9382,N_5068,N_6739);
xor U9383 (N_9383,N_7145,N_5899);
xnor U9384 (N_9384,N_5502,N_6244);
nor U9385 (N_9385,N_6951,N_6553);
nand U9386 (N_9386,N_5538,N_6752);
xor U9387 (N_9387,N_7396,N_6080);
xor U9388 (N_9388,N_6829,N_6926);
xor U9389 (N_9389,N_7284,N_6793);
or U9390 (N_9390,N_6038,N_5763);
nor U9391 (N_9391,N_7496,N_6283);
nand U9392 (N_9392,N_5480,N_5311);
and U9393 (N_9393,N_5151,N_6878);
xor U9394 (N_9394,N_6055,N_6606);
and U9395 (N_9395,N_6384,N_5755);
or U9396 (N_9396,N_5314,N_5201);
and U9397 (N_9397,N_6928,N_6320);
xor U9398 (N_9398,N_6039,N_5781);
nor U9399 (N_9399,N_7251,N_5944);
xnor U9400 (N_9400,N_5325,N_7090);
nand U9401 (N_9401,N_6707,N_5698);
or U9402 (N_9402,N_5373,N_7291);
nor U9403 (N_9403,N_6598,N_7204);
nor U9404 (N_9404,N_5813,N_6105);
nand U9405 (N_9405,N_6515,N_5745);
nand U9406 (N_9406,N_6545,N_7229);
nand U9407 (N_9407,N_6500,N_5861);
nand U9408 (N_9408,N_7166,N_7149);
and U9409 (N_9409,N_6415,N_7266);
or U9410 (N_9410,N_6931,N_6311);
nand U9411 (N_9411,N_5701,N_7119);
nand U9412 (N_9412,N_6082,N_6352);
nand U9413 (N_9413,N_6268,N_6661);
or U9414 (N_9414,N_5564,N_6409);
nor U9415 (N_9415,N_6577,N_5520);
and U9416 (N_9416,N_5514,N_6738);
nand U9417 (N_9417,N_7075,N_6611);
xnor U9418 (N_9418,N_5272,N_6974);
nor U9419 (N_9419,N_5008,N_5018);
nand U9420 (N_9420,N_6807,N_7238);
xor U9421 (N_9421,N_6190,N_6311);
and U9422 (N_9422,N_7183,N_6077);
nand U9423 (N_9423,N_5534,N_5115);
or U9424 (N_9424,N_7308,N_6258);
or U9425 (N_9425,N_6576,N_7319);
or U9426 (N_9426,N_6174,N_5548);
or U9427 (N_9427,N_6759,N_6830);
and U9428 (N_9428,N_6786,N_7164);
nand U9429 (N_9429,N_7096,N_6196);
and U9430 (N_9430,N_6823,N_5012);
xnor U9431 (N_9431,N_6314,N_7288);
or U9432 (N_9432,N_5837,N_5533);
and U9433 (N_9433,N_5086,N_6207);
nor U9434 (N_9434,N_6917,N_6635);
nand U9435 (N_9435,N_5044,N_6484);
or U9436 (N_9436,N_6823,N_5109);
and U9437 (N_9437,N_5212,N_6034);
nand U9438 (N_9438,N_6242,N_5859);
and U9439 (N_9439,N_5578,N_5381);
nor U9440 (N_9440,N_6111,N_6119);
xnor U9441 (N_9441,N_6672,N_5596);
nand U9442 (N_9442,N_6260,N_5115);
xor U9443 (N_9443,N_6371,N_6613);
nand U9444 (N_9444,N_6822,N_6185);
nor U9445 (N_9445,N_6787,N_6478);
or U9446 (N_9446,N_5297,N_7106);
xnor U9447 (N_9447,N_7059,N_6320);
and U9448 (N_9448,N_6388,N_5955);
and U9449 (N_9449,N_6419,N_5742);
nand U9450 (N_9450,N_5399,N_6197);
nor U9451 (N_9451,N_6743,N_5762);
nor U9452 (N_9452,N_5362,N_5993);
xor U9453 (N_9453,N_6547,N_5054);
nand U9454 (N_9454,N_5424,N_5934);
or U9455 (N_9455,N_7051,N_5555);
nand U9456 (N_9456,N_5288,N_6543);
nor U9457 (N_9457,N_6654,N_6397);
xnor U9458 (N_9458,N_7261,N_6890);
nor U9459 (N_9459,N_5891,N_6943);
xor U9460 (N_9460,N_6455,N_7077);
xor U9461 (N_9461,N_5608,N_6002);
xor U9462 (N_9462,N_5253,N_6776);
nor U9463 (N_9463,N_6292,N_5124);
xnor U9464 (N_9464,N_7429,N_6459);
nor U9465 (N_9465,N_5331,N_6635);
xor U9466 (N_9466,N_5702,N_6089);
or U9467 (N_9467,N_5082,N_6487);
or U9468 (N_9468,N_5771,N_7137);
nand U9469 (N_9469,N_5204,N_6322);
or U9470 (N_9470,N_5383,N_6144);
or U9471 (N_9471,N_5709,N_5049);
nand U9472 (N_9472,N_5287,N_5259);
nand U9473 (N_9473,N_5985,N_5593);
nand U9474 (N_9474,N_5480,N_5501);
xnor U9475 (N_9475,N_5888,N_5800);
nand U9476 (N_9476,N_7061,N_6834);
and U9477 (N_9477,N_6980,N_7078);
or U9478 (N_9478,N_7221,N_5966);
nor U9479 (N_9479,N_5145,N_6125);
or U9480 (N_9480,N_6141,N_6391);
or U9481 (N_9481,N_5194,N_6072);
and U9482 (N_9482,N_5774,N_6915);
or U9483 (N_9483,N_5773,N_7164);
or U9484 (N_9484,N_7244,N_6786);
xnor U9485 (N_9485,N_7469,N_5980);
or U9486 (N_9486,N_6310,N_5501);
nand U9487 (N_9487,N_5756,N_5759);
nand U9488 (N_9488,N_5693,N_7322);
and U9489 (N_9489,N_5042,N_7112);
nand U9490 (N_9490,N_5643,N_5333);
or U9491 (N_9491,N_7329,N_7441);
xor U9492 (N_9492,N_6036,N_6541);
nand U9493 (N_9493,N_6177,N_6460);
xnor U9494 (N_9494,N_6117,N_5495);
nor U9495 (N_9495,N_5121,N_6273);
xnor U9496 (N_9496,N_7476,N_6534);
xnor U9497 (N_9497,N_6657,N_6114);
or U9498 (N_9498,N_6049,N_6827);
xnor U9499 (N_9499,N_7242,N_5882);
nor U9500 (N_9500,N_5281,N_6084);
and U9501 (N_9501,N_7161,N_6284);
xor U9502 (N_9502,N_6688,N_5985);
or U9503 (N_9503,N_7187,N_5607);
xor U9504 (N_9504,N_7035,N_6362);
and U9505 (N_9505,N_6328,N_6628);
nor U9506 (N_9506,N_6064,N_7024);
or U9507 (N_9507,N_6231,N_6324);
xor U9508 (N_9508,N_5770,N_5346);
xnor U9509 (N_9509,N_6784,N_5057);
and U9510 (N_9510,N_5233,N_5417);
xnor U9511 (N_9511,N_5134,N_5776);
or U9512 (N_9512,N_5247,N_5555);
nand U9513 (N_9513,N_7191,N_7482);
nor U9514 (N_9514,N_5791,N_6185);
and U9515 (N_9515,N_6391,N_6496);
xor U9516 (N_9516,N_6548,N_5209);
and U9517 (N_9517,N_6984,N_6987);
or U9518 (N_9518,N_6313,N_5506);
or U9519 (N_9519,N_5326,N_6823);
and U9520 (N_9520,N_6278,N_5383);
nand U9521 (N_9521,N_6214,N_7353);
or U9522 (N_9522,N_5674,N_5956);
nor U9523 (N_9523,N_7095,N_6471);
nor U9524 (N_9524,N_6728,N_5091);
and U9525 (N_9525,N_5674,N_6691);
and U9526 (N_9526,N_5319,N_6522);
xor U9527 (N_9527,N_6435,N_7324);
nand U9528 (N_9528,N_5055,N_6404);
xnor U9529 (N_9529,N_6638,N_6215);
and U9530 (N_9530,N_6748,N_6848);
xor U9531 (N_9531,N_5437,N_5999);
nand U9532 (N_9532,N_5232,N_5039);
nand U9533 (N_9533,N_6632,N_5479);
xor U9534 (N_9534,N_7140,N_5315);
and U9535 (N_9535,N_5366,N_7377);
xnor U9536 (N_9536,N_6341,N_5336);
or U9537 (N_9537,N_7071,N_7390);
or U9538 (N_9538,N_6835,N_5504);
and U9539 (N_9539,N_6499,N_6166);
and U9540 (N_9540,N_5739,N_6020);
xor U9541 (N_9541,N_6908,N_6334);
xnor U9542 (N_9542,N_6605,N_5155);
xnor U9543 (N_9543,N_7069,N_5573);
xnor U9544 (N_9544,N_6573,N_6533);
nand U9545 (N_9545,N_5141,N_5278);
and U9546 (N_9546,N_5518,N_6316);
or U9547 (N_9547,N_7423,N_6028);
nand U9548 (N_9548,N_6162,N_7011);
nor U9549 (N_9549,N_6275,N_6117);
nand U9550 (N_9550,N_7309,N_5776);
or U9551 (N_9551,N_5798,N_7462);
nand U9552 (N_9552,N_7070,N_6443);
nand U9553 (N_9553,N_5521,N_7151);
and U9554 (N_9554,N_7326,N_6570);
nand U9555 (N_9555,N_5715,N_5164);
or U9556 (N_9556,N_7101,N_7146);
or U9557 (N_9557,N_7263,N_5127);
xor U9558 (N_9558,N_6862,N_6599);
or U9559 (N_9559,N_5025,N_7172);
xnor U9560 (N_9560,N_5601,N_7239);
and U9561 (N_9561,N_5247,N_7462);
xor U9562 (N_9562,N_5247,N_5276);
and U9563 (N_9563,N_6131,N_5032);
nor U9564 (N_9564,N_6200,N_5373);
xor U9565 (N_9565,N_5839,N_6480);
nand U9566 (N_9566,N_6328,N_7296);
nor U9567 (N_9567,N_6204,N_5491);
xnor U9568 (N_9568,N_5882,N_5613);
nor U9569 (N_9569,N_7048,N_6867);
nand U9570 (N_9570,N_6079,N_5052);
xnor U9571 (N_9571,N_5701,N_5735);
xnor U9572 (N_9572,N_6940,N_7127);
or U9573 (N_9573,N_5278,N_6694);
or U9574 (N_9574,N_5159,N_6726);
nand U9575 (N_9575,N_5806,N_6282);
nand U9576 (N_9576,N_6929,N_6903);
nand U9577 (N_9577,N_6548,N_6846);
nand U9578 (N_9578,N_7204,N_5954);
nand U9579 (N_9579,N_7339,N_6651);
xnor U9580 (N_9580,N_6841,N_6474);
or U9581 (N_9581,N_5730,N_6662);
and U9582 (N_9582,N_6706,N_5294);
xnor U9583 (N_9583,N_6293,N_5379);
or U9584 (N_9584,N_7265,N_6027);
xnor U9585 (N_9585,N_6677,N_7485);
nand U9586 (N_9586,N_5835,N_5936);
or U9587 (N_9587,N_6790,N_5335);
and U9588 (N_9588,N_6905,N_6267);
xnor U9589 (N_9589,N_6608,N_5282);
nand U9590 (N_9590,N_6315,N_6499);
xnor U9591 (N_9591,N_6692,N_5693);
or U9592 (N_9592,N_6382,N_6332);
and U9593 (N_9593,N_5932,N_5881);
or U9594 (N_9594,N_5761,N_5319);
or U9595 (N_9595,N_6417,N_6807);
nor U9596 (N_9596,N_5434,N_5901);
xnor U9597 (N_9597,N_5541,N_6507);
nor U9598 (N_9598,N_6462,N_6492);
xnor U9599 (N_9599,N_6357,N_7309);
or U9600 (N_9600,N_5381,N_6871);
and U9601 (N_9601,N_6805,N_6282);
xnor U9602 (N_9602,N_5835,N_5883);
nor U9603 (N_9603,N_5737,N_5626);
nor U9604 (N_9604,N_6787,N_5623);
or U9605 (N_9605,N_6972,N_5894);
nor U9606 (N_9606,N_5276,N_7156);
xor U9607 (N_9607,N_5480,N_5979);
or U9608 (N_9608,N_6393,N_5568);
nor U9609 (N_9609,N_6613,N_5976);
or U9610 (N_9610,N_6188,N_5189);
nor U9611 (N_9611,N_6467,N_5699);
xnor U9612 (N_9612,N_5378,N_6376);
xnor U9613 (N_9613,N_7235,N_6906);
nor U9614 (N_9614,N_6044,N_5888);
nand U9615 (N_9615,N_6382,N_7330);
nand U9616 (N_9616,N_5475,N_7007);
nor U9617 (N_9617,N_6845,N_6834);
xnor U9618 (N_9618,N_5119,N_7371);
xor U9619 (N_9619,N_6173,N_5746);
and U9620 (N_9620,N_5102,N_5124);
and U9621 (N_9621,N_6432,N_7413);
or U9622 (N_9622,N_7341,N_7012);
and U9623 (N_9623,N_6492,N_7022);
or U9624 (N_9624,N_7013,N_7270);
or U9625 (N_9625,N_7343,N_5670);
and U9626 (N_9626,N_5124,N_6256);
xor U9627 (N_9627,N_6198,N_5647);
xor U9628 (N_9628,N_5796,N_6575);
nand U9629 (N_9629,N_6384,N_7458);
xnor U9630 (N_9630,N_5210,N_7277);
or U9631 (N_9631,N_6814,N_6919);
and U9632 (N_9632,N_6608,N_5368);
and U9633 (N_9633,N_5571,N_5966);
nor U9634 (N_9634,N_5894,N_6214);
nor U9635 (N_9635,N_7016,N_6154);
or U9636 (N_9636,N_6599,N_5694);
nand U9637 (N_9637,N_7366,N_5562);
nor U9638 (N_9638,N_7180,N_6689);
nand U9639 (N_9639,N_5832,N_5463);
or U9640 (N_9640,N_7229,N_6315);
or U9641 (N_9641,N_5022,N_6662);
or U9642 (N_9642,N_5102,N_7081);
nor U9643 (N_9643,N_5025,N_5747);
nor U9644 (N_9644,N_6936,N_6140);
or U9645 (N_9645,N_6827,N_5918);
nor U9646 (N_9646,N_5108,N_7130);
nand U9647 (N_9647,N_5797,N_5156);
xnor U9648 (N_9648,N_5110,N_5364);
xnor U9649 (N_9649,N_7326,N_6223);
and U9650 (N_9650,N_7208,N_6444);
xor U9651 (N_9651,N_5468,N_5188);
and U9652 (N_9652,N_6612,N_6096);
nand U9653 (N_9653,N_6018,N_6712);
nor U9654 (N_9654,N_5259,N_7451);
or U9655 (N_9655,N_6327,N_5066);
or U9656 (N_9656,N_5682,N_5256);
nand U9657 (N_9657,N_5320,N_5648);
and U9658 (N_9658,N_5023,N_7291);
nor U9659 (N_9659,N_5848,N_7008);
nor U9660 (N_9660,N_7048,N_6143);
nand U9661 (N_9661,N_5836,N_7203);
or U9662 (N_9662,N_5608,N_6074);
and U9663 (N_9663,N_5667,N_5258);
or U9664 (N_9664,N_7350,N_6475);
xnor U9665 (N_9665,N_7154,N_7222);
nor U9666 (N_9666,N_5579,N_5807);
nor U9667 (N_9667,N_7291,N_5633);
or U9668 (N_9668,N_6657,N_6972);
or U9669 (N_9669,N_6014,N_6022);
and U9670 (N_9670,N_6354,N_5932);
xor U9671 (N_9671,N_7133,N_5222);
nand U9672 (N_9672,N_6073,N_5873);
nor U9673 (N_9673,N_7198,N_7460);
nand U9674 (N_9674,N_5851,N_7142);
and U9675 (N_9675,N_7038,N_5032);
nand U9676 (N_9676,N_5482,N_5034);
nand U9677 (N_9677,N_6955,N_7488);
xnor U9678 (N_9678,N_5797,N_5020);
and U9679 (N_9679,N_7043,N_5972);
xor U9680 (N_9680,N_6760,N_6366);
nand U9681 (N_9681,N_5228,N_7420);
nor U9682 (N_9682,N_6110,N_6057);
xor U9683 (N_9683,N_5424,N_5546);
xor U9684 (N_9684,N_6046,N_5663);
xnor U9685 (N_9685,N_6054,N_7203);
nand U9686 (N_9686,N_6773,N_7123);
xnor U9687 (N_9687,N_6323,N_6837);
or U9688 (N_9688,N_5358,N_5972);
xnor U9689 (N_9689,N_6249,N_5468);
xnor U9690 (N_9690,N_6073,N_5309);
xor U9691 (N_9691,N_6143,N_5672);
xor U9692 (N_9692,N_6419,N_5530);
xor U9693 (N_9693,N_6184,N_6674);
xnor U9694 (N_9694,N_7091,N_7344);
xor U9695 (N_9695,N_5200,N_7002);
nand U9696 (N_9696,N_5831,N_6022);
nor U9697 (N_9697,N_6383,N_7464);
or U9698 (N_9698,N_6040,N_6500);
nor U9699 (N_9699,N_5457,N_6488);
and U9700 (N_9700,N_5454,N_5892);
and U9701 (N_9701,N_5508,N_6318);
or U9702 (N_9702,N_6816,N_5881);
xnor U9703 (N_9703,N_5141,N_5169);
nand U9704 (N_9704,N_6842,N_6598);
nor U9705 (N_9705,N_6991,N_6416);
nor U9706 (N_9706,N_7356,N_6283);
nor U9707 (N_9707,N_6915,N_5802);
nand U9708 (N_9708,N_5850,N_7038);
or U9709 (N_9709,N_5969,N_6155);
and U9710 (N_9710,N_6143,N_7414);
xnor U9711 (N_9711,N_7303,N_7143);
xnor U9712 (N_9712,N_7284,N_5105);
nor U9713 (N_9713,N_5093,N_7425);
nand U9714 (N_9714,N_6435,N_6634);
xor U9715 (N_9715,N_6580,N_6731);
nand U9716 (N_9716,N_5154,N_5522);
or U9717 (N_9717,N_6168,N_5018);
nor U9718 (N_9718,N_6153,N_5806);
nand U9719 (N_9719,N_6272,N_7330);
nor U9720 (N_9720,N_5439,N_7200);
xnor U9721 (N_9721,N_6000,N_5682);
xnor U9722 (N_9722,N_6168,N_5769);
nor U9723 (N_9723,N_6999,N_6575);
and U9724 (N_9724,N_5865,N_5490);
and U9725 (N_9725,N_7441,N_7020);
or U9726 (N_9726,N_6950,N_6592);
or U9727 (N_9727,N_5811,N_6270);
nor U9728 (N_9728,N_5859,N_7097);
nor U9729 (N_9729,N_6974,N_6988);
and U9730 (N_9730,N_7303,N_5282);
nand U9731 (N_9731,N_5095,N_6466);
and U9732 (N_9732,N_7411,N_5150);
or U9733 (N_9733,N_6339,N_5660);
nand U9734 (N_9734,N_5687,N_5464);
and U9735 (N_9735,N_5884,N_6557);
xnor U9736 (N_9736,N_7042,N_7285);
or U9737 (N_9737,N_5871,N_7284);
nand U9738 (N_9738,N_7174,N_6847);
xnor U9739 (N_9739,N_6288,N_6525);
nand U9740 (N_9740,N_7339,N_5281);
or U9741 (N_9741,N_6552,N_6748);
or U9742 (N_9742,N_6951,N_5594);
xnor U9743 (N_9743,N_5315,N_5249);
and U9744 (N_9744,N_7441,N_6244);
xnor U9745 (N_9745,N_6640,N_6670);
xor U9746 (N_9746,N_7330,N_5477);
and U9747 (N_9747,N_7345,N_6485);
and U9748 (N_9748,N_6135,N_5579);
nor U9749 (N_9749,N_5667,N_6575);
and U9750 (N_9750,N_6524,N_6345);
xnor U9751 (N_9751,N_5924,N_6328);
and U9752 (N_9752,N_5919,N_6011);
nor U9753 (N_9753,N_5707,N_6966);
and U9754 (N_9754,N_7098,N_6957);
nor U9755 (N_9755,N_6560,N_5247);
xnor U9756 (N_9756,N_7060,N_6908);
and U9757 (N_9757,N_5394,N_5429);
or U9758 (N_9758,N_6398,N_7022);
nor U9759 (N_9759,N_5874,N_6264);
or U9760 (N_9760,N_5956,N_5201);
and U9761 (N_9761,N_5036,N_5677);
and U9762 (N_9762,N_7154,N_6535);
or U9763 (N_9763,N_5546,N_5818);
nand U9764 (N_9764,N_7393,N_7032);
xor U9765 (N_9765,N_5085,N_6455);
nand U9766 (N_9766,N_6019,N_5497);
nor U9767 (N_9767,N_5332,N_6291);
or U9768 (N_9768,N_5020,N_5041);
nor U9769 (N_9769,N_5263,N_7364);
xor U9770 (N_9770,N_5897,N_6685);
nand U9771 (N_9771,N_6651,N_5108);
xor U9772 (N_9772,N_6276,N_5689);
and U9773 (N_9773,N_6563,N_6499);
xnor U9774 (N_9774,N_5869,N_6405);
and U9775 (N_9775,N_5225,N_5766);
nand U9776 (N_9776,N_5461,N_7435);
nand U9777 (N_9777,N_6412,N_5076);
nand U9778 (N_9778,N_7079,N_5883);
nor U9779 (N_9779,N_6792,N_5980);
nor U9780 (N_9780,N_6046,N_5019);
and U9781 (N_9781,N_6602,N_6537);
nor U9782 (N_9782,N_6708,N_5655);
and U9783 (N_9783,N_5765,N_7388);
nand U9784 (N_9784,N_6228,N_7397);
nand U9785 (N_9785,N_6647,N_5171);
nor U9786 (N_9786,N_7171,N_5074);
or U9787 (N_9787,N_5569,N_6954);
or U9788 (N_9788,N_6996,N_6367);
or U9789 (N_9789,N_6688,N_5019);
xnor U9790 (N_9790,N_5868,N_5029);
nor U9791 (N_9791,N_7312,N_7439);
nand U9792 (N_9792,N_7230,N_6972);
xor U9793 (N_9793,N_6992,N_6209);
nand U9794 (N_9794,N_7053,N_6662);
and U9795 (N_9795,N_6255,N_7036);
or U9796 (N_9796,N_5869,N_6312);
or U9797 (N_9797,N_6144,N_7119);
xor U9798 (N_9798,N_6947,N_5946);
or U9799 (N_9799,N_6768,N_5190);
or U9800 (N_9800,N_5069,N_5464);
or U9801 (N_9801,N_6854,N_7095);
nor U9802 (N_9802,N_5488,N_7107);
nand U9803 (N_9803,N_5045,N_5627);
nor U9804 (N_9804,N_5313,N_7089);
nand U9805 (N_9805,N_5754,N_5661);
xor U9806 (N_9806,N_5020,N_6326);
and U9807 (N_9807,N_5860,N_6231);
and U9808 (N_9808,N_5516,N_5313);
nor U9809 (N_9809,N_5668,N_7443);
and U9810 (N_9810,N_6838,N_6878);
or U9811 (N_9811,N_7495,N_6087);
xnor U9812 (N_9812,N_5097,N_5982);
or U9813 (N_9813,N_5355,N_5609);
or U9814 (N_9814,N_5072,N_7177);
xor U9815 (N_9815,N_5128,N_7199);
or U9816 (N_9816,N_7008,N_6500);
nand U9817 (N_9817,N_5629,N_6345);
xor U9818 (N_9818,N_5061,N_5693);
or U9819 (N_9819,N_6463,N_5461);
or U9820 (N_9820,N_5286,N_7424);
nor U9821 (N_9821,N_6897,N_5600);
xnor U9822 (N_9822,N_6174,N_6348);
and U9823 (N_9823,N_5264,N_6118);
nand U9824 (N_9824,N_6718,N_6956);
nor U9825 (N_9825,N_5765,N_5922);
or U9826 (N_9826,N_5674,N_7230);
or U9827 (N_9827,N_7186,N_7358);
or U9828 (N_9828,N_5464,N_7014);
nor U9829 (N_9829,N_5953,N_7309);
xnor U9830 (N_9830,N_5039,N_6647);
xnor U9831 (N_9831,N_6735,N_5218);
and U9832 (N_9832,N_6056,N_7259);
nand U9833 (N_9833,N_6827,N_6856);
and U9834 (N_9834,N_5842,N_6500);
nand U9835 (N_9835,N_6299,N_5208);
xnor U9836 (N_9836,N_6898,N_7451);
and U9837 (N_9837,N_5087,N_7300);
or U9838 (N_9838,N_6704,N_5507);
nor U9839 (N_9839,N_6314,N_5197);
and U9840 (N_9840,N_5550,N_6842);
or U9841 (N_9841,N_6656,N_6601);
nor U9842 (N_9842,N_6291,N_6340);
xnor U9843 (N_9843,N_6494,N_7356);
and U9844 (N_9844,N_7194,N_6979);
xor U9845 (N_9845,N_6768,N_5024);
and U9846 (N_9846,N_7084,N_5941);
or U9847 (N_9847,N_7153,N_7170);
or U9848 (N_9848,N_7319,N_5103);
and U9849 (N_9849,N_5675,N_6097);
or U9850 (N_9850,N_7205,N_5474);
or U9851 (N_9851,N_6436,N_7003);
and U9852 (N_9852,N_6656,N_5716);
xnor U9853 (N_9853,N_6965,N_5707);
xor U9854 (N_9854,N_6494,N_6859);
nor U9855 (N_9855,N_5212,N_5263);
or U9856 (N_9856,N_7452,N_6606);
nor U9857 (N_9857,N_7174,N_6737);
nor U9858 (N_9858,N_5925,N_6709);
or U9859 (N_9859,N_6022,N_5720);
or U9860 (N_9860,N_6588,N_6967);
or U9861 (N_9861,N_6660,N_5467);
or U9862 (N_9862,N_6207,N_5855);
xnor U9863 (N_9863,N_5817,N_6163);
nand U9864 (N_9864,N_6621,N_7181);
or U9865 (N_9865,N_6127,N_5099);
and U9866 (N_9866,N_7088,N_5849);
nor U9867 (N_9867,N_6000,N_6491);
and U9868 (N_9868,N_7457,N_7139);
and U9869 (N_9869,N_5422,N_6503);
xnor U9870 (N_9870,N_5762,N_5928);
nand U9871 (N_9871,N_6532,N_6146);
or U9872 (N_9872,N_5883,N_6721);
xnor U9873 (N_9873,N_6603,N_5945);
or U9874 (N_9874,N_7025,N_6084);
nand U9875 (N_9875,N_6272,N_7136);
and U9876 (N_9876,N_5168,N_6429);
nor U9877 (N_9877,N_6109,N_6833);
xor U9878 (N_9878,N_5428,N_6779);
xor U9879 (N_9879,N_6691,N_5994);
and U9880 (N_9880,N_5187,N_6392);
or U9881 (N_9881,N_5815,N_5796);
nor U9882 (N_9882,N_5517,N_6866);
xor U9883 (N_9883,N_5490,N_7098);
and U9884 (N_9884,N_6667,N_6171);
or U9885 (N_9885,N_5675,N_6901);
and U9886 (N_9886,N_7098,N_7114);
nand U9887 (N_9887,N_7238,N_5771);
xnor U9888 (N_9888,N_6671,N_5261);
xnor U9889 (N_9889,N_6732,N_7021);
and U9890 (N_9890,N_6348,N_6949);
nand U9891 (N_9891,N_5042,N_6775);
xor U9892 (N_9892,N_6240,N_6697);
nand U9893 (N_9893,N_5511,N_6573);
and U9894 (N_9894,N_5574,N_5295);
xor U9895 (N_9895,N_6268,N_5354);
or U9896 (N_9896,N_6366,N_7115);
and U9897 (N_9897,N_5034,N_6953);
and U9898 (N_9898,N_6624,N_6659);
nand U9899 (N_9899,N_5688,N_5002);
and U9900 (N_9900,N_6636,N_5446);
or U9901 (N_9901,N_6367,N_5727);
and U9902 (N_9902,N_7133,N_5284);
nor U9903 (N_9903,N_6208,N_6869);
and U9904 (N_9904,N_6759,N_6888);
xor U9905 (N_9905,N_5006,N_5385);
xor U9906 (N_9906,N_6957,N_5214);
xor U9907 (N_9907,N_7261,N_7494);
nor U9908 (N_9908,N_7334,N_6055);
xnor U9909 (N_9909,N_7209,N_5464);
or U9910 (N_9910,N_6843,N_6686);
nand U9911 (N_9911,N_6040,N_5016);
or U9912 (N_9912,N_6719,N_6204);
xor U9913 (N_9913,N_7191,N_5702);
nand U9914 (N_9914,N_6272,N_6097);
nor U9915 (N_9915,N_6645,N_7180);
or U9916 (N_9916,N_5813,N_6838);
nand U9917 (N_9917,N_5309,N_6761);
xnor U9918 (N_9918,N_7495,N_7490);
xnor U9919 (N_9919,N_5464,N_7017);
and U9920 (N_9920,N_5817,N_5315);
and U9921 (N_9921,N_5179,N_6245);
and U9922 (N_9922,N_6516,N_6142);
nand U9923 (N_9923,N_5884,N_6667);
nor U9924 (N_9924,N_5906,N_5302);
nor U9925 (N_9925,N_5376,N_5758);
xor U9926 (N_9926,N_6235,N_6256);
and U9927 (N_9927,N_6583,N_6185);
and U9928 (N_9928,N_6344,N_7238);
or U9929 (N_9929,N_7078,N_5245);
nand U9930 (N_9930,N_6510,N_5891);
nor U9931 (N_9931,N_6353,N_5147);
or U9932 (N_9932,N_6241,N_5683);
nor U9933 (N_9933,N_6005,N_5464);
nor U9934 (N_9934,N_5504,N_5431);
or U9935 (N_9935,N_5380,N_6609);
and U9936 (N_9936,N_6199,N_7479);
nand U9937 (N_9937,N_6094,N_7412);
or U9938 (N_9938,N_7031,N_5457);
xnor U9939 (N_9939,N_7379,N_6603);
and U9940 (N_9940,N_5255,N_5623);
nand U9941 (N_9941,N_6759,N_6564);
and U9942 (N_9942,N_5970,N_6108);
xor U9943 (N_9943,N_7016,N_6233);
nand U9944 (N_9944,N_7169,N_5414);
xor U9945 (N_9945,N_5692,N_6886);
nand U9946 (N_9946,N_6899,N_6424);
xnor U9947 (N_9947,N_5789,N_6694);
and U9948 (N_9948,N_7456,N_5477);
xor U9949 (N_9949,N_5734,N_5745);
or U9950 (N_9950,N_7412,N_5407);
and U9951 (N_9951,N_5300,N_5130);
nand U9952 (N_9952,N_7378,N_6233);
or U9953 (N_9953,N_7286,N_5192);
and U9954 (N_9954,N_6248,N_5290);
nor U9955 (N_9955,N_7279,N_5788);
and U9956 (N_9956,N_7167,N_5813);
nand U9957 (N_9957,N_6688,N_7393);
or U9958 (N_9958,N_5611,N_6119);
or U9959 (N_9959,N_6935,N_6223);
xor U9960 (N_9960,N_7063,N_6318);
xor U9961 (N_9961,N_5051,N_6311);
and U9962 (N_9962,N_7111,N_6795);
xnor U9963 (N_9963,N_5526,N_6838);
nand U9964 (N_9964,N_5220,N_6448);
nand U9965 (N_9965,N_6290,N_5632);
and U9966 (N_9966,N_6759,N_5249);
and U9967 (N_9967,N_5203,N_6472);
nor U9968 (N_9968,N_5886,N_6997);
nand U9969 (N_9969,N_6886,N_6870);
and U9970 (N_9970,N_5941,N_5209);
nand U9971 (N_9971,N_6699,N_6440);
xor U9972 (N_9972,N_7034,N_6580);
and U9973 (N_9973,N_5966,N_7386);
xor U9974 (N_9974,N_5887,N_5902);
nand U9975 (N_9975,N_6650,N_6501);
nor U9976 (N_9976,N_6028,N_5725);
xnor U9977 (N_9977,N_5879,N_6091);
xnor U9978 (N_9978,N_5181,N_7052);
and U9979 (N_9979,N_6189,N_7243);
and U9980 (N_9980,N_5692,N_5487);
nand U9981 (N_9981,N_5907,N_5222);
nand U9982 (N_9982,N_7470,N_7417);
nor U9983 (N_9983,N_6385,N_6588);
and U9984 (N_9984,N_5846,N_6770);
and U9985 (N_9985,N_5715,N_6897);
and U9986 (N_9986,N_6480,N_7184);
nand U9987 (N_9987,N_6081,N_5353);
xor U9988 (N_9988,N_7001,N_5432);
or U9989 (N_9989,N_5829,N_6523);
and U9990 (N_9990,N_5061,N_5959);
nor U9991 (N_9991,N_5575,N_7461);
or U9992 (N_9992,N_5851,N_5109);
nor U9993 (N_9993,N_5169,N_7192);
xor U9994 (N_9994,N_6254,N_5131);
and U9995 (N_9995,N_6727,N_5743);
nand U9996 (N_9996,N_6423,N_6130);
nand U9997 (N_9997,N_5266,N_6131);
xnor U9998 (N_9998,N_5734,N_5830);
or U9999 (N_9999,N_5534,N_6698);
xnor U10000 (N_10000,N_8292,N_8263);
and U10001 (N_10001,N_9686,N_9266);
or U10002 (N_10002,N_9366,N_8844);
and U10003 (N_10003,N_8120,N_8702);
nor U10004 (N_10004,N_9554,N_8175);
or U10005 (N_10005,N_9903,N_7568);
and U10006 (N_10006,N_9828,N_8149);
nor U10007 (N_10007,N_9205,N_9852);
xnor U10008 (N_10008,N_9272,N_8726);
nand U10009 (N_10009,N_9467,N_9453);
nor U10010 (N_10010,N_8070,N_8199);
xor U10011 (N_10011,N_8687,N_9536);
xor U10012 (N_10012,N_9214,N_8434);
nand U10013 (N_10013,N_9660,N_8742);
xnor U10014 (N_10014,N_9392,N_8576);
nand U10015 (N_10015,N_8140,N_8237);
xor U10016 (N_10016,N_7585,N_9018);
xor U10017 (N_10017,N_9268,N_8316);
nor U10018 (N_10018,N_9324,N_8753);
and U10019 (N_10019,N_9327,N_8048);
and U10020 (N_10020,N_8606,N_8691);
xor U10021 (N_10021,N_9757,N_7762);
xor U10022 (N_10022,N_9808,N_7711);
nor U10023 (N_10023,N_7592,N_9121);
and U10024 (N_10024,N_8559,N_8022);
nand U10025 (N_10025,N_8283,N_8957);
nand U10026 (N_10026,N_7562,N_8129);
and U10027 (N_10027,N_9666,N_9241);
nand U10028 (N_10028,N_8697,N_8333);
xor U10029 (N_10029,N_9956,N_8666);
nor U10030 (N_10030,N_8570,N_9074);
nand U10031 (N_10031,N_9284,N_9551);
and U10032 (N_10032,N_8207,N_9661);
nor U10033 (N_10033,N_8342,N_9151);
nor U10034 (N_10034,N_7643,N_7725);
and U10035 (N_10035,N_7987,N_8154);
and U10036 (N_10036,N_7607,N_9306);
xnor U10037 (N_10037,N_9441,N_9002);
nand U10038 (N_10038,N_8472,N_8257);
nor U10039 (N_10039,N_8637,N_7552);
nor U10040 (N_10040,N_9581,N_7890);
nor U10041 (N_10041,N_7809,N_7814);
nand U10042 (N_10042,N_8698,N_9138);
and U10043 (N_10043,N_8716,N_7795);
or U10044 (N_10044,N_9457,N_9842);
or U10045 (N_10045,N_8216,N_8478);
xnor U10046 (N_10046,N_8229,N_7985);
nor U10047 (N_10047,N_8094,N_9297);
or U10048 (N_10048,N_9418,N_7615);
xor U10049 (N_10049,N_9647,N_8227);
xor U10050 (N_10050,N_9455,N_8176);
and U10051 (N_10051,N_9343,N_8302);
nor U10052 (N_10052,N_8276,N_8265);
nor U10053 (N_10053,N_8055,N_8830);
or U10054 (N_10054,N_9402,N_9899);
or U10055 (N_10055,N_9329,N_8778);
or U10056 (N_10056,N_9533,N_8101);
and U10057 (N_10057,N_8032,N_8117);
nor U10058 (N_10058,N_9375,N_8161);
and U10059 (N_10059,N_8714,N_7939);
or U10060 (N_10060,N_8690,N_9620);
and U10061 (N_10061,N_8718,N_8883);
or U10062 (N_10062,N_9696,N_7570);
or U10063 (N_10063,N_8505,N_9871);
xor U10064 (N_10064,N_9063,N_7571);
nor U10065 (N_10065,N_7750,N_9680);
xor U10066 (N_10066,N_8143,N_8988);
and U10067 (N_10067,N_8787,N_9942);
xor U10068 (N_10068,N_8616,N_8201);
nor U10069 (N_10069,N_7927,N_7652);
nand U10070 (N_10070,N_8410,N_9727);
and U10071 (N_10071,N_9722,N_7692);
or U10072 (N_10072,N_9090,N_9817);
xnor U10073 (N_10073,N_9712,N_7801);
or U10074 (N_10074,N_8943,N_9785);
nand U10075 (N_10075,N_9486,N_8673);
nor U10076 (N_10076,N_7875,N_8562);
or U10077 (N_10077,N_8496,N_9797);
nor U10078 (N_10078,N_8053,N_7966);
nand U10079 (N_10079,N_7885,N_9221);
nand U10080 (N_10080,N_9947,N_9333);
nand U10081 (N_10081,N_9251,N_8869);
or U10082 (N_10082,N_9195,N_9475);
and U10083 (N_10083,N_9381,N_7722);
or U10084 (N_10084,N_9881,N_9779);
nand U10085 (N_10085,N_9201,N_8851);
and U10086 (N_10086,N_9033,N_9364);
and U10087 (N_10087,N_9812,N_7908);
xor U10088 (N_10088,N_7907,N_8599);
or U10089 (N_10089,N_9978,N_8730);
or U10090 (N_10090,N_7926,N_9294);
nand U10091 (N_10091,N_8577,N_8605);
nor U10092 (N_10092,N_8008,N_8768);
nand U10093 (N_10093,N_7602,N_9060);
nand U10094 (N_10094,N_7586,N_7753);
or U10095 (N_10095,N_9986,N_8045);
and U10096 (N_10096,N_9580,N_8819);
or U10097 (N_10097,N_8274,N_8037);
nand U10098 (N_10098,N_7821,N_8332);
nor U10099 (N_10099,N_9636,N_8703);
xor U10100 (N_10100,N_9283,N_8223);
and U10101 (N_10101,N_8555,N_9851);
or U10102 (N_10102,N_9055,N_9365);
xnor U10103 (N_10103,N_8266,N_7740);
xnor U10104 (N_10104,N_9880,N_8195);
xor U10105 (N_10105,N_9111,N_9326);
nand U10106 (N_10106,N_9875,N_7746);
or U10107 (N_10107,N_7515,N_7895);
xnor U10108 (N_10108,N_8111,N_8717);
xor U10109 (N_10109,N_8650,N_8311);
nand U10110 (N_10110,N_9449,N_9385);
xor U10111 (N_10111,N_9070,N_9293);
xnor U10112 (N_10112,N_9827,N_8862);
nor U10113 (N_10113,N_9206,N_8738);
nand U10114 (N_10114,N_8466,N_9801);
nand U10115 (N_10115,N_8063,N_9612);
xor U10116 (N_10116,N_9788,N_8894);
or U10117 (N_10117,N_9445,N_8909);
nand U10118 (N_10118,N_8402,N_8928);
and U10119 (N_10119,N_9010,N_9425);
nand U10120 (N_10120,N_8281,N_7525);
xnor U10121 (N_10121,N_9292,N_9527);
or U10122 (N_10122,N_8357,N_8633);
nor U10123 (N_10123,N_9535,N_9637);
or U10124 (N_10124,N_8680,N_8362);
nand U10125 (N_10125,N_8388,N_8481);
xor U10126 (N_10126,N_8081,N_9725);
and U10127 (N_10127,N_9176,N_8829);
nand U10128 (N_10128,N_9480,N_8611);
nor U10129 (N_10129,N_9254,N_8471);
or U10130 (N_10130,N_8871,N_7680);
xor U10131 (N_10131,N_8099,N_8234);
and U10132 (N_10132,N_9006,N_8930);
and U10133 (N_10133,N_7797,N_9933);
or U10134 (N_10134,N_7835,N_9549);
and U10135 (N_10135,N_9314,N_7947);
nand U10136 (N_10136,N_9093,N_7655);
and U10137 (N_10137,N_8169,N_8556);
nand U10138 (N_10138,N_8743,N_8926);
and U10139 (N_10139,N_8961,N_8672);
and U10140 (N_10140,N_7911,N_8076);
or U10141 (N_10141,N_8712,N_7864);
nor U10142 (N_10142,N_9415,N_8312);
nand U10143 (N_10143,N_7697,N_9166);
nor U10144 (N_10144,N_9207,N_8425);
nor U10145 (N_10145,N_7812,N_9500);
nand U10146 (N_10146,N_8901,N_8809);
xor U10147 (N_10147,N_8021,N_9991);
and U10148 (N_10148,N_9879,N_8912);
and U10149 (N_10149,N_9622,N_8654);
xor U10150 (N_10150,N_8522,N_8214);
and U10151 (N_10151,N_7599,N_9945);
or U10152 (N_10152,N_9047,N_9731);
nor U10153 (N_10153,N_9965,N_8838);
or U10154 (N_10154,N_8763,N_7943);
or U10155 (N_10155,N_9191,N_9435);
xor U10156 (N_10156,N_8807,N_7806);
xor U10157 (N_10157,N_7535,N_8189);
or U10158 (N_10158,N_8891,N_9930);
nor U10159 (N_10159,N_8459,N_9180);
nor U10160 (N_10160,N_8122,N_7736);
or U10161 (N_10161,N_7855,N_9917);
and U10162 (N_10162,N_9038,N_9550);
or U10163 (N_10163,N_8791,N_7820);
and U10164 (N_10164,N_7636,N_8532);
nor U10165 (N_10165,N_9170,N_8074);
and U10166 (N_10166,N_7832,N_8011);
nand U10167 (N_10167,N_8774,N_9609);
xnor U10168 (N_10168,N_9753,N_8231);
and U10169 (N_10169,N_7671,N_9347);
xor U10170 (N_10170,N_9673,N_8446);
nand U10171 (N_10171,N_7548,N_8420);
and U10172 (N_10172,N_7970,N_8377);
and U10173 (N_10173,N_8136,N_8747);
nand U10174 (N_10174,N_7743,N_8879);
or U10175 (N_10175,N_7948,N_8550);
or U10176 (N_10176,N_8762,N_7900);
nand U10177 (N_10177,N_8445,N_9745);
or U10178 (N_10178,N_8956,N_8116);
nor U10179 (N_10179,N_9106,N_8013);
nand U10180 (N_10180,N_9037,N_8507);
or U10181 (N_10181,N_9939,N_9398);
xnor U10182 (N_10182,N_7617,N_9123);
and U10183 (N_10183,N_9743,N_7677);
nor U10184 (N_10184,N_8695,N_7506);
and U10185 (N_10185,N_7977,N_9977);
or U10186 (N_10186,N_8304,N_7935);
or U10187 (N_10187,N_9910,N_8275);
xor U10188 (N_10188,N_7681,N_9183);
nand U10189 (N_10189,N_9607,N_9579);
nand U10190 (N_10190,N_8877,N_7732);
nor U10191 (N_10191,N_8501,N_8392);
nand U10192 (N_10192,N_7955,N_8724);
or U10193 (N_10193,N_8942,N_9213);
nand U10194 (N_10194,N_9764,N_9127);
xor U10195 (N_10195,N_9429,N_9531);
nor U10196 (N_10196,N_8419,N_7557);
xnor U10197 (N_10197,N_8927,N_8024);
and U10198 (N_10198,N_7699,N_9937);
nor U10199 (N_10199,N_8187,N_8391);
and U10200 (N_10200,N_9859,N_7544);
or U10201 (N_10201,N_7919,N_9857);
and U10202 (N_10202,N_9136,N_9732);
nand U10203 (N_10203,N_7884,N_8315);
xor U10204 (N_10204,N_9290,N_8219);
xor U10205 (N_10205,N_8679,N_9529);
nand U10206 (N_10206,N_9845,N_9925);
nor U10207 (N_10207,N_9987,N_7789);
nand U10208 (N_10208,N_9586,N_9943);
or U10209 (N_10209,N_9525,N_9865);
or U10210 (N_10210,N_9331,N_8394);
nand U10211 (N_10211,N_9307,N_8360);
and U10212 (N_10212,N_9747,N_8084);
nor U10213 (N_10213,N_7594,N_7724);
and U10214 (N_10214,N_8424,N_8511);
and U10215 (N_10215,N_8861,N_8797);
nand U10216 (N_10216,N_7507,N_8153);
nor U10217 (N_10217,N_7794,N_9147);
nand U10218 (N_10218,N_8370,N_7800);
nand U10219 (N_10219,N_9724,N_8051);
or U10220 (N_10220,N_8247,N_8831);
nor U10221 (N_10221,N_9169,N_8164);
xnor U10222 (N_10222,N_9082,N_7577);
and U10223 (N_10223,N_8191,N_8645);
nor U10224 (N_10224,N_7971,N_8100);
nor U10225 (N_10225,N_8541,N_9019);
nand U10226 (N_10226,N_9589,N_7816);
or U10227 (N_10227,N_9892,N_9460);
nand U10228 (N_10228,N_8824,N_8594);
nor U10229 (N_10229,N_8454,N_9485);
xor U10230 (N_10230,N_9081,N_9838);
or U10231 (N_10231,N_7857,N_8764);
nand U10232 (N_10232,N_9472,N_7849);
or U10233 (N_10233,N_9878,N_7945);
or U10234 (N_10234,N_8069,N_9999);
nor U10235 (N_10235,N_7766,N_9354);
and U10236 (N_10236,N_9915,N_8465);
nor U10237 (N_10237,N_8089,N_9565);
nor U10238 (N_10238,N_9493,N_8442);
nand U10239 (N_10239,N_7742,N_9863);
nand U10240 (N_10240,N_8160,N_7940);
nor U10241 (N_10241,N_7865,N_9356);
or U10242 (N_10242,N_8749,N_7936);
nand U10243 (N_10243,N_7640,N_9440);
or U10244 (N_10244,N_8026,N_8364);
nor U10245 (N_10245,N_8427,N_7879);
and U10246 (N_10246,N_9746,N_7780);
and U10247 (N_10247,N_7771,N_8352);
xnor U10248 (N_10248,N_8506,N_9157);
nand U10249 (N_10249,N_7996,N_9796);
nor U10250 (N_10250,N_9172,N_9259);
or U10251 (N_10251,N_9739,N_9640);
and U10252 (N_10252,N_8924,N_9212);
and U10253 (N_10253,N_9015,N_9601);
or U10254 (N_10254,N_8765,N_8080);
nand U10255 (N_10255,N_9174,N_8498);
or U10256 (N_10256,N_9748,N_8363);
xor U10257 (N_10257,N_9644,N_9104);
or U10258 (N_10258,N_9322,N_9976);
and U10259 (N_10259,N_9576,N_8035);
and U10260 (N_10260,N_7872,N_9985);
nand U10261 (N_10261,N_7547,N_9377);
and U10262 (N_10262,N_8970,N_8182);
nand U10263 (N_10263,N_9328,N_7623);
nor U10264 (N_10264,N_9776,N_8233);
xor U10265 (N_10265,N_8918,N_8323);
nand U10266 (N_10266,N_9321,N_8018);
nor U10267 (N_10267,N_8638,N_7601);
and U10268 (N_10268,N_7739,N_8306);
and U10269 (N_10269,N_9907,N_9540);
nand U10270 (N_10270,N_8936,N_8582);
xor U10271 (N_10271,N_9846,N_9959);
xnor U10272 (N_10272,N_9787,N_9256);
or U10273 (N_10273,N_9962,N_9036);
or U10274 (N_10274,N_9419,N_9122);
nand U10275 (N_10275,N_9913,N_8287);
nand U10276 (N_10276,N_9594,N_8810);
nand U10277 (N_10277,N_9783,N_8401);
nor U10278 (N_10278,N_7756,N_7566);
xnor U10279 (N_10279,N_9583,N_7706);
nor U10280 (N_10280,N_8412,N_8158);
nand U10281 (N_10281,N_8553,N_9974);
nand U10282 (N_10282,N_9113,N_8657);
nand U10283 (N_10283,N_7824,N_8945);
and U10284 (N_10284,N_9416,N_9626);
or U10285 (N_10285,N_8317,N_8196);
nor U10286 (N_10286,N_9308,N_7880);
xnor U10287 (N_10287,N_8808,N_9394);
xor U10288 (N_10288,N_7504,N_8515);
xnor U10289 (N_10289,N_9720,N_8248);
xnor U10290 (N_10290,N_7963,N_8755);
or U10291 (N_10291,N_7641,N_8091);
xnor U10292 (N_10292,N_9901,N_7503);
or U10293 (N_10293,N_9459,N_9932);
xor U10294 (N_10294,N_8186,N_9678);
nor U10295 (N_10295,N_8845,N_8882);
nor U10296 (N_10296,N_7558,N_9571);
nand U10297 (N_10297,N_8905,N_9515);
and U10298 (N_10298,N_9345,N_8060);
or U10299 (N_10299,N_9239,N_8781);
xnor U10300 (N_10300,N_8676,N_9617);
xnor U10301 (N_10301,N_8353,N_9923);
and U10302 (N_10302,N_8139,N_9387);
xor U10303 (N_10303,N_8236,N_7997);
or U10304 (N_10304,N_9502,N_9654);
or U10305 (N_10305,N_7583,N_9026);
or U10306 (N_10306,N_8001,N_8795);
nor U10307 (N_10307,N_8150,N_8141);
xor U10308 (N_10308,N_7654,N_9649);
nand U10309 (N_10309,N_9013,N_9164);
xor U10310 (N_10310,N_8056,N_8581);
xnor U10311 (N_10311,N_7632,N_7944);
nand U10312 (N_10312,N_8623,N_9714);
nand U10313 (N_10313,N_9920,N_9688);
or U10314 (N_10314,N_9483,N_8524);
xor U10315 (N_10315,N_7679,N_9588);
or U10316 (N_10316,N_9008,N_8962);
or U10317 (N_10317,N_9229,N_8152);
nand U10318 (N_10318,N_7682,N_9894);
nand U10319 (N_10319,N_8497,N_8873);
or U10320 (N_10320,N_9426,N_8414);
and U10321 (N_10321,N_8652,N_7606);
xnor U10322 (N_10322,N_9924,N_8536);
and U10323 (N_10323,N_8888,N_7894);
nand U10324 (N_10324,N_8239,N_7634);
nor U10325 (N_10325,N_8895,N_7590);
nor U10326 (N_10326,N_8293,N_9633);
nor U10327 (N_10327,N_9064,N_8295);
nor U10328 (N_10328,N_9456,N_9162);
or U10329 (N_10329,N_7647,N_7836);
xor U10330 (N_10330,N_9603,N_9028);
and U10331 (N_10331,N_7973,N_9372);
and U10332 (N_10332,N_7658,N_9995);
or U10333 (N_10333,N_8321,N_9902);
nor U10334 (N_10334,N_9302,N_8502);
nand U10335 (N_10335,N_7694,N_8610);
nand U10336 (N_10336,N_8899,N_8359);
and U10337 (N_10337,N_7691,N_8543);
xor U10338 (N_10338,N_7912,N_8254);
and U10339 (N_10339,N_9181,N_7834);
or U10340 (N_10340,N_9866,N_7698);
and U10341 (N_10341,N_9975,N_7823);
nand U10342 (N_10342,N_9705,N_8782);
nand U10343 (N_10343,N_9885,N_9477);
nor U10344 (N_10344,N_9309,N_8426);
nand U10345 (N_10345,N_9476,N_9427);
and U10346 (N_10346,N_9560,N_7883);
or U10347 (N_10347,N_8917,N_9046);
and U10348 (N_10348,N_8416,N_9397);
nor U10349 (N_10349,N_8908,N_8017);
xnor U10350 (N_10350,N_7862,N_9348);
nor U10351 (N_10351,N_9790,N_9886);
nand U10352 (N_10352,N_8925,N_9918);
or U10353 (N_10353,N_8270,N_7953);
nand U10354 (N_10354,N_9573,N_9171);
nor U10355 (N_10355,N_8386,N_8000);
xor U10356 (N_10356,N_8615,N_8727);
or U10357 (N_10357,N_7892,N_7538);
and U10358 (N_10358,N_9780,N_7888);
nor U10359 (N_10359,N_7576,N_8735);
nand U10360 (N_10360,N_8959,N_8533);
nor U10361 (N_10361,N_9646,N_8826);
or U10362 (N_10362,N_8566,N_9811);
and U10363 (N_10363,N_7745,N_8110);
nand U10364 (N_10364,N_7610,N_8480);
nor U10365 (N_10365,N_9786,N_9358);
and U10366 (N_10366,N_9534,N_8846);
or U10367 (N_10367,N_8713,N_8612);
nand U10368 (N_10368,N_7887,N_9778);
xor U10369 (N_10369,N_8955,N_9856);
nand U10370 (N_10370,N_8996,N_9446);
xnor U10371 (N_10371,N_8334,N_9411);
nor U10372 (N_10372,N_7564,N_7511);
nand U10373 (N_10373,N_7501,N_9247);
or U10374 (N_10374,N_7786,N_7828);
or U10375 (N_10375,N_9657,N_8272);
xnor U10376 (N_10376,N_8458,N_8843);
nor U10377 (N_10377,N_9103,N_9717);
xor U10378 (N_10378,N_9401,N_8546);
or U10379 (N_10379,N_8054,N_8689);
nor U10380 (N_10380,N_7803,N_8664);
nand U10381 (N_10381,N_7891,N_9927);
and U10382 (N_10382,N_8429,N_8356);
xnor U10383 (N_10383,N_9631,N_8519);
and U10384 (N_10384,N_8126,N_7755);
or U10385 (N_10385,N_9393,N_9088);
nor U10386 (N_10386,N_7702,N_9216);
and U10387 (N_10387,N_9862,N_7877);
nand U10388 (N_10388,N_9623,N_7534);
or U10389 (N_10389,N_7550,N_9210);
nand U10390 (N_10390,N_7841,N_9775);
nor U10391 (N_10391,N_8318,N_7792);
and U10392 (N_10392,N_9628,N_9044);
nor U10393 (N_10393,N_9056,N_8213);
nor U10394 (N_10394,N_7931,N_8107);
nor U10395 (N_10395,N_8596,N_9854);
and U10396 (N_10396,N_7509,N_8322);
nand U10397 (N_10397,N_7998,N_8548);
and U10398 (N_10398,N_7642,N_9009);
nor U10399 (N_10399,N_7512,N_9955);
and U10400 (N_10400,N_8721,N_9001);
and U10401 (N_10401,N_9248,N_9156);
nor U10402 (N_10402,N_9043,N_7720);
nor U10403 (N_10403,N_8834,N_8104);
nor U10404 (N_10404,N_9729,N_9570);
and U10405 (N_10405,N_8818,N_9726);
nand U10406 (N_10406,N_8887,N_8284);
xor U10407 (N_10407,N_8208,N_9921);
nor U10408 (N_10408,N_7782,N_8732);
nand U10409 (N_10409,N_8619,N_9243);
or U10410 (N_10410,N_9552,N_8545);
xnor U10411 (N_10411,N_7840,N_8508);
nand U10412 (N_10412,N_9412,N_8435);
or U10413 (N_10413,N_8404,N_8984);
or U10414 (N_10414,N_9518,N_9360);
xnor U10415 (N_10415,N_9610,N_8969);
xnor U10416 (N_10416,N_9815,N_8397);
or U10417 (N_10417,N_8681,N_8889);
nand U10418 (N_10418,N_9627,N_9887);
and U10419 (N_10419,N_8975,N_7685);
nor U10420 (N_10420,N_8893,N_7733);
nand U10421 (N_10421,N_9490,N_7580);
nor U10422 (N_10422,N_8244,N_9514);
and U10423 (N_10423,N_9114,N_8340);
and U10424 (N_10424,N_8047,N_8057);
nor U10425 (N_10425,N_9185,N_8850);
or U10426 (N_10426,N_9754,N_9330);
and U10427 (N_10427,N_7545,N_8935);
xnor U10428 (N_10428,N_9900,N_9316);
nand U10429 (N_10429,N_8789,N_9512);
xor U10430 (N_10430,N_9810,N_8137);
and U10431 (N_10431,N_8800,N_8347);
nand U10432 (N_10432,N_8669,N_7696);
xnor U10433 (N_10433,N_9964,N_9703);
xnor U10434 (N_10434,N_7833,N_9682);
xor U10435 (N_10435,N_7729,N_9155);
nand U10436 (N_10436,N_8963,N_7916);
xor U10437 (N_10437,N_7761,N_9813);
xor U10438 (N_10438,N_9509,N_9339);
nor U10439 (N_10439,N_9882,N_8568);
xnor U10440 (N_10440,N_8285,N_8407);
or U10441 (N_10441,N_8422,N_8603);
and U10442 (N_10442,N_8171,N_9774);
or U10443 (N_10443,N_8618,N_8853);
and U10444 (N_10444,N_8897,N_7593);
nand U10445 (N_10445,N_7981,N_8190);
xor U10446 (N_10446,N_8484,N_9130);
nor U10447 (N_10447,N_9034,N_9906);
nand U10448 (N_10448,N_9697,N_9370);
or U10449 (N_10449,N_8031,N_8595);
and U10450 (N_10450,N_8804,N_8486);
xnor U10451 (N_10451,N_8470,N_9767);
and U10452 (N_10452,N_8162,N_7644);
and U10453 (N_10453,N_8954,N_9843);
xor U10454 (N_10454,N_8335,N_8865);
nor U10455 (N_10455,N_7903,N_8210);
nor U10456 (N_10456,N_8088,N_9116);
xor U10457 (N_10457,N_7728,N_8997);
and U10458 (N_10458,N_7510,N_8518);
xnor U10459 (N_10459,N_9458,N_7744);
nand U10460 (N_10460,N_7645,N_8464);
nand U10461 (N_10461,N_9198,N_9659);
or U10462 (N_10462,N_8477,N_9606);
xnor U10463 (N_10463,N_9532,N_9369);
and U10464 (N_10464,N_8251,N_8977);
xor U10465 (N_10465,N_7560,N_9542);
xnor U10466 (N_10466,N_8500,N_9406);
and U10467 (N_10467,N_9728,N_8597);
or U10468 (N_10468,N_9281,N_9340);
and U10469 (N_10469,N_9410,N_8439);
and U10470 (N_10470,N_8232,N_9639);
and U10471 (N_10471,N_9698,N_9668);
xnor U10472 (N_10472,N_9223,N_7710);
nand U10473 (N_10473,N_8794,N_7650);
and U10474 (N_10474,N_8715,N_7920);
xor U10475 (N_10475,N_7822,N_9545);
and U10476 (N_10476,N_9877,N_9471);
and U10477 (N_10477,N_8798,N_7791);
nand U10478 (N_10478,N_8866,N_8181);
nor U10479 (N_10479,N_7873,N_9249);
and U10480 (N_10480,N_9215,N_8857);
or U10481 (N_10481,N_8142,N_8042);
xnor U10482 (N_10482,N_8677,N_7529);
and U10483 (N_10483,N_9112,N_8282);
xnor U10484 (N_10484,N_9662,N_9708);
or U10485 (N_10485,N_8268,N_9635);
and U10486 (N_10486,N_9177,N_9618);
and U10487 (N_10487,N_8994,N_9519);
nor U10488 (N_10488,N_8780,N_9966);
nor U10489 (N_10489,N_7866,N_8542);
and U10490 (N_10490,N_7964,N_8303);
nor U10491 (N_10491,N_9798,N_7850);
nand U10492 (N_10492,N_8922,N_9675);
nand U10493 (N_10493,N_8561,N_8253);
nand U10494 (N_10494,N_8156,N_8646);
nand U10495 (N_10495,N_9858,N_8197);
nor U10496 (N_10496,N_8572,N_8365);
or U10497 (N_10497,N_8444,N_9593);
or U10498 (N_10498,N_9814,N_7752);
nor U10499 (N_10499,N_8479,N_8025);
nand U10500 (N_10500,N_9602,N_7969);
nand U10501 (N_10501,N_8813,N_8408);
or U10502 (N_10502,N_9874,N_9848);
and U10503 (N_10503,N_7867,N_8958);
xor U10504 (N_10504,N_9099,N_8348);
nor U10505 (N_10505,N_9718,N_9648);
nor U10506 (N_10506,N_9832,N_9758);
and U10507 (N_10507,N_9756,N_8504);
and U10508 (N_10508,N_8886,N_9988);
or U10509 (N_10509,N_7874,N_8934);
nand U10510 (N_10510,N_8371,N_7613);
and U10511 (N_10511,N_8939,N_8784);
nor U10512 (N_10512,N_8124,N_9335);
nor U10513 (N_10513,N_8978,N_8447);
or U10514 (N_10514,N_7608,N_8510);
nand U10515 (N_10515,N_9624,N_7713);
and U10516 (N_10516,N_7889,N_8567);
or U10517 (N_10517,N_7735,N_8585);
nor U10518 (N_10518,N_8225,N_9761);
or U10519 (N_10519,N_8146,N_8170);
xnor U10520 (N_10520,N_7561,N_9474);
nand U10521 (N_10521,N_9679,N_9141);
nand U10522 (N_10522,N_9496,N_9528);
or U10523 (N_10523,N_7952,N_8584);
and U10524 (N_10524,N_8355,N_8050);
and U10525 (N_10525,N_9694,N_9653);
nand U10526 (N_10526,N_9065,N_8709);
xor U10527 (N_10527,N_7785,N_9847);
nor U10528 (N_10528,N_9444,N_9833);
and U10529 (N_10529,N_9834,N_9053);
and U10530 (N_10530,N_8805,N_9323);
or U10531 (N_10531,N_9341,N_8168);
and U10532 (N_10532,N_9400,N_7757);
nand U10533 (N_10533,N_8923,N_8684);
and U10534 (N_10534,N_9944,N_8399);
xor U10535 (N_10535,N_8417,N_8551);
or U10536 (N_10536,N_9704,N_7553);
and U10537 (N_10537,N_8868,N_9396);
nor U10538 (N_10538,N_8569,N_8766);
xor U10539 (N_10539,N_9431,N_7901);
nor U10540 (N_10540,N_7995,N_7520);
nor U10541 (N_10541,N_9860,N_8754);
nor U10542 (N_10542,N_7628,N_7881);
nor U10543 (N_10543,N_7959,N_9693);
and U10544 (N_10544,N_7633,N_7773);
nor U10545 (N_10545,N_8406,N_8185);
nor U10546 (N_10546,N_9363,N_7991);
nor U10547 (N_10547,N_7618,N_8858);
nor U10548 (N_10548,N_7788,N_8493);
nor U10549 (N_10549,N_9039,N_7626);
nor U10550 (N_10550,N_9572,N_9524);
or U10551 (N_10551,N_7878,N_7818);
or U10552 (N_10552,N_9523,N_8589);
xor U10553 (N_10553,N_9017,N_9409);
and U10554 (N_10554,N_9012,N_8779);
nand U10555 (N_10555,N_9124,N_9506);
nor U10556 (N_10556,N_8995,N_8108);
and U10557 (N_10557,N_8114,N_8375);
or U10558 (N_10558,N_9296,N_9650);
nor U10559 (N_10559,N_8913,N_8876);
nor U10560 (N_10560,N_8704,N_8243);
nand U10561 (N_10561,N_8972,N_7845);
or U10562 (N_10562,N_7717,N_9107);
and U10563 (N_10563,N_9094,N_8106);
xor U10564 (N_10564,N_7767,N_9751);
or U10565 (N_10565,N_9547,N_9226);
nand U10566 (N_10566,N_7775,N_9569);
nor U10567 (N_10567,N_7559,N_9789);
or U10568 (N_10568,N_9526,N_8448);
xor U10569 (N_10569,N_8639,N_9159);
nor U10570 (N_10570,N_9605,N_9663);
or U10571 (N_10571,N_8395,N_8489);
or U10572 (N_10572,N_8198,N_8644);
or U10573 (N_10573,N_9041,N_8613);
or U10574 (N_10574,N_9766,N_9084);
and U10575 (N_10575,N_7869,N_8558);
nand U10576 (N_10576,N_8267,N_7581);
and U10577 (N_10577,N_9148,N_7539);
xor U10578 (N_10578,N_8771,N_9802);
nor U10579 (N_10579,N_8062,N_7530);
nor U10580 (N_10580,N_8313,N_9125);
nor U10581 (N_10581,N_8630,N_9218);
nor U10582 (N_10582,N_9931,N_8590);
xor U10583 (N_10583,N_9299,N_7846);
nor U10584 (N_10584,N_7829,N_9664);
or U10585 (N_10585,N_9303,N_7635);
xor U10586 (N_10586,N_9119,N_9643);
nand U10587 (N_10587,N_7531,N_9282);
nor U10588 (N_10588,N_7831,N_8855);
xnor U10589 (N_10589,N_9338,N_7505);
nand U10590 (N_10590,N_9765,N_9548);
or U10591 (N_10591,N_9199,N_8938);
or U10592 (N_10592,N_8421,N_8430);
nand U10593 (N_10593,N_9342,N_7604);
xnor U10594 (N_10594,N_9516,N_8092);
nor U10595 (N_10595,N_8940,N_7960);
nand U10596 (N_10596,N_7573,N_8872);
or U10597 (N_10597,N_7651,N_9521);
nor U10598 (N_10598,N_9577,N_9539);
and U10599 (N_10599,N_7619,N_9355);
xor U10600 (N_10600,N_8604,N_9443);
nor U10601 (N_10601,N_7993,N_9799);
and U10602 (N_10602,N_8686,N_8989);
nor U10603 (N_10603,N_9888,N_9240);
xor U10604 (N_10604,N_8212,N_7899);
nand U10605 (N_10605,N_8226,N_8678);
and U10606 (N_10606,N_7582,N_9128);
nand U10607 (N_10607,N_8600,N_9153);
and U10608 (N_10608,N_9231,N_8077);
nor U10609 (N_10609,N_8256,N_9481);
nor U10610 (N_10610,N_9278,N_8663);
nand U10611 (N_10611,N_7625,N_9464);
xnor U10612 (N_10612,N_8300,N_9793);
and U10613 (N_10613,N_8628,N_8368);
nand U10614 (N_10614,N_9186,N_8565);
and U10615 (N_10615,N_9803,N_7827);
xor U10616 (N_10616,N_9567,N_9839);
nor U10617 (N_10617,N_7638,N_8919);
and U10618 (N_10618,N_8965,N_8815);
xnor U10619 (N_10619,N_9408,N_9837);
xnor U10620 (N_10620,N_8286,N_9211);
and U10621 (N_10621,N_8202,N_9928);
xor U10622 (N_10622,N_8786,N_8029);
nand U10623 (N_10623,N_8517,N_8006);
and U10624 (N_10624,N_7826,N_7676);
nor U10625 (N_10625,N_7675,N_7662);
or U10626 (N_10626,N_9439,N_8674);
xnor U10627 (N_10627,N_8783,N_8220);
xor U10628 (N_10628,N_9651,N_8647);
nand U10629 (N_10629,N_9741,N_8526);
nor U10630 (N_10630,N_9513,N_8987);
or U10631 (N_10631,N_9820,N_9204);
or U10632 (N_10632,N_9451,N_9263);
xor U10633 (N_10633,N_8005,N_8291);
nand U10634 (N_10634,N_8067,N_7781);
nand U10635 (N_10635,N_7502,N_7783);
xnor U10636 (N_10636,N_8750,N_9996);
and U10637 (N_10637,N_8528,N_8799);
nand U10638 (N_10638,N_9940,N_7913);
xnor U10639 (N_10639,N_9792,N_8661);
nor U10640 (N_10640,N_8583,N_8163);
xor U10641 (N_10641,N_8587,N_7584);
or U10642 (N_10642,N_8588,N_8580);
and U10643 (N_10643,N_8289,N_9244);
and U10644 (N_10644,N_9404,N_9831);
xor U10645 (N_10645,N_7990,N_8651);
nor U10646 (N_10646,N_8722,N_9075);
nand U10647 (N_10647,N_8003,N_8881);
xor U10648 (N_10648,N_8981,N_7543);
nand U10649 (N_10649,N_8044,N_7763);
xnor U10650 (N_10650,N_8564,N_8937);
nor U10651 (N_10651,N_9684,N_8211);
nand U10652 (N_10652,N_7897,N_9491);
and U10653 (N_10653,N_8949,N_9829);
nor U10654 (N_10654,N_9970,N_9736);
or U10655 (N_10655,N_7851,N_9884);
nor U10656 (N_10656,N_8903,N_8350);
nor U10657 (N_10657,N_9257,N_9466);
nand U10658 (N_10658,N_9578,N_7716);
nor U10659 (N_10659,N_8832,N_9553);
xor U10660 (N_10660,N_9655,N_8344);
nand U10661 (N_10661,N_7666,N_8443);
xor U10662 (N_10662,N_8041,N_8953);
nor U10663 (N_10663,N_9187,N_8330);
nand U10664 (N_10664,N_8354,N_9992);
nand U10665 (N_10665,N_8915,N_8217);
and U10666 (N_10666,N_7631,N_8761);
nand U10667 (N_10667,N_9699,N_8892);
and U10668 (N_10668,N_8411,N_8135);
nor U10669 (N_10669,N_9224,N_7804);
nand U10670 (N_10670,N_9770,N_8167);
nand U10671 (N_10671,N_8552,N_9421);
or U10672 (N_10672,N_7978,N_9641);
xor U10673 (N_10673,N_7726,N_9738);
nand U10674 (N_10674,N_8878,N_8811);
xnor U10675 (N_10675,N_7688,N_9035);
nor U10676 (N_10676,N_9997,N_9737);
and U10677 (N_10677,N_7779,N_9024);
and U10678 (N_10678,N_9361,N_9344);
or U10679 (N_10679,N_7853,N_9687);
or U10680 (N_10680,N_9824,N_8710);
nand U10681 (N_10681,N_7989,N_9032);
and U10682 (N_10682,N_8733,N_7704);
or U10683 (N_10683,N_8173,N_7589);
nand U10684 (N_10684,N_9709,N_8061);
nor U10685 (N_10685,N_9178,N_9971);
or U10686 (N_10686,N_8290,N_7917);
nor U10687 (N_10687,N_8491,N_8387);
or U10688 (N_10688,N_8971,N_8776);
nor U10689 (N_10689,N_9165,N_9083);
or U10690 (N_10690,N_9870,N_9543);
nor U10691 (N_10691,N_9690,N_8848);
nor U10692 (N_10692,N_7802,N_8720);
xor U10693 (N_10693,N_9537,N_8485);
nand U10694 (N_10694,N_9574,N_8549);
or U10695 (N_10695,N_7693,N_8601);
or U10696 (N_10696,N_8906,N_7915);
and U10697 (N_10697,N_9557,N_8308);
xor U10698 (N_10698,N_9969,N_8261);
nor U10699 (N_10699,N_8102,N_7612);
xor U10700 (N_10700,N_8640,N_8269);
nor U10701 (N_10701,N_8516,N_9597);
or U10702 (N_10702,N_9559,N_8675);
or U10703 (N_10703,N_8773,N_8941);
or U10704 (N_10704,N_8902,N_9671);
nor U10705 (N_10705,N_8598,N_7522);
nor U10706 (N_10706,N_8205,N_9235);
xor U10707 (N_10707,N_8383,N_7627);
xor U10708 (N_10708,N_8288,N_8023);
or U10709 (N_10709,N_9163,N_9118);
or U10710 (N_10710,N_9073,N_9100);
nor U10711 (N_10711,N_9794,N_9983);
xor U10712 (N_10712,N_9488,N_7738);
nand U10713 (N_10713,N_7578,N_7709);
and U10714 (N_10714,N_9929,N_9246);
xor U10715 (N_10715,N_8240,N_8259);
and U10716 (N_10716,N_7813,N_8854);
xnor U10717 (N_10717,N_7871,N_8885);
or U10718 (N_10718,N_9953,N_9040);
xor U10719 (N_10719,N_7563,N_7830);
and U10720 (N_10720,N_8499,N_8736);
nor U10721 (N_10721,N_8728,N_8707);
and U10722 (N_10722,N_8560,N_9442);
xnor U10723 (N_10723,N_7979,N_9069);
nand U10724 (N_10724,N_9585,N_7624);
nand U10725 (N_10725,N_8494,N_8817);
nor U10726 (N_10726,N_8297,N_9473);
xnor U10727 (N_10727,N_9101,N_9707);
and U10728 (N_10728,N_9981,N_9368);
nor U10729 (N_10729,N_8235,N_9998);
nor U10730 (N_10730,N_9479,N_8010);
and U10731 (N_10731,N_7657,N_8453);
xnor U10732 (N_10732,N_9295,N_8823);
nand U10733 (N_10733,N_8653,N_9030);
nand U10734 (N_10734,N_9301,N_9079);
and U10735 (N_10735,N_7870,N_8767);
or U10736 (N_10736,N_9777,N_8144);
or U10737 (N_10737,N_9716,N_9197);
nand U10738 (N_10738,N_8193,N_8592);
nor U10739 (N_10739,N_8538,N_8803);
or U10740 (N_10740,N_9949,N_8482);
xnor U10741 (N_10741,N_8151,N_9298);
xor U10742 (N_10742,N_9505,N_9462);
nand U10743 (N_10743,N_9071,N_9098);
nand U10744 (N_10744,N_8842,N_7528);
and U10745 (N_10745,N_7852,N_9371);
nand U10746 (N_10746,N_9700,N_9872);
nand U10747 (N_10747,N_9004,N_9667);
or U10748 (N_10748,N_9300,N_8130);
xor U10749 (N_10749,N_9386,N_9658);
nand U10750 (N_10750,N_8324,N_7541);
nand U10751 (N_10751,N_9271,N_8574);
or U10752 (N_10752,N_8020,N_7760);
or U10753 (N_10753,N_7967,N_9556);
xor U10754 (N_10754,N_9706,N_9274);
or U10755 (N_10755,N_7549,N_9461);
nor U10756 (N_10756,N_8449,N_8078);
or U10757 (N_10757,N_9227,N_8900);
or U10758 (N_10758,N_9482,N_8166);
xnor U10759 (N_10759,N_8921,N_8827);
or U10760 (N_10760,N_7609,N_7734);
and U10761 (N_10761,N_8758,N_8875);
and U10762 (N_10762,N_9105,N_8474);
nand U10763 (N_10763,N_8951,N_8932);
xor U10764 (N_10764,N_7567,N_7790);
xor U10765 (N_10765,N_9132,N_7741);
nand U10766 (N_10766,N_9634,N_7986);
or U10767 (N_10767,N_8336,N_7918);
and U10768 (N_10768,N_9468,N_9423);
or U10769 (N_10769,N_8525,N_9253);
xor U10770 (N_10770,N_7708,N_8097);
and U10771 (N_10771,N_7938,N_8535);
nand U10772 (N_10772,N_9422,N_8822);
nand U10773 (N_10773,N_9267,N_9584);
or U10774 (N_10774,N_9334,N_9511);
or U10775 (N_10775,N_8621,N_9614);
nor U10776 (N_10776,N_8415,N_8573);
and U10777 (N_10777,N_7648,N_7957);
or U10778 (N_10778,N_9555,N_8660);
nand U10779 (N_10779,N_9864,N_8490);
or U10780 (N_10780,N_7574,N_9723);
nor U10781 (N_10781,N_8775,N_9389);
nand U10782 (N_10782,N_8856,N_9568);
or U10783 (N_10783,N_9742,N_8015);
and U10784 (N_10784,N_9311,N_9265);
and U10785 (N_10785,N_8820,N_9869);
and U10786 (N_10786,N_9430,N_8351);
or U10787 (N_10787,N_8228,N_9599);
xnor U10788 (N_10788,N_7975,N_8338);
or U10789 (N_10789,N_8503,N_8626);
or U10790 (N_10790,N_9438,N_9189);
nand U10791 (N_10791,N_8475,N_8495);
nand U10792 (N_10792,N_9867,N_9003);
nor U10793 (N_10793,N_9095,N_9049);
xor U10794 (N_10794,N_9150,N_8757);
nor U10795 (N_10795,N_7579,N_8487);
xor U10796 (N_10796,N_9109,N_9450);
or U10797 (N_10797,N_8301,N_8469);
nand U10798 (N_10798,N_7837,N_8165);
or U10799 (N_10799,N_9200,N_8874);
and U10800 (N_10800,N_9582,N_8440);
and U10801 (N_10801,N_9131,N_9642);
nor U10802 (N_10802,N_7811,N_9711);
or U10803 (N_10803,N_9285,N_7784);
nor U10804 (N_10804,N_8400,N_8960);
xor U10805 (N_10805,N_7683,N_8920);
nand U10806 (N_10806,N_8133,N_8575);
nor U10807 (N_10807,N_7956,N_8983);
nand U10808 (N_10808,N_9424,N_9390);
nand U10809 (N_10809,N_9021,N_9926);
xnor U10810 (N_10810,N_8701,N_8999);
and U10811 (N_10811,N_8931,N_7819);
or U10812 (N_10812,N_8904,N_9129);
nor U10813 (N_10813,N_9562,N_8483);
xor U10814 (N_10814,N_9142,N_9674);
or U10815 (N_10815,N_7514,N_9273);
nand U10816 (N_10816,N_8539,N_9315);
or U10817 (N_10817,N_9275,N_8343);
nand U10818 (N_10818,N_9052,N_9317);
nand U10819 (N_10819,N_8328,N_7933);
nand U10820 (N_10820,N_8346,N_8086);
and U10821 (N_10821,N_8314,N_8683);
nand U10822 (N_10822,N_8118,N_9805);
or U10823 (N_10823,N_8770,N_8148);
or U10824 (N_10824,N_8307,N_7843);
or U10825 (N_10825,N_8529,N_7700);
nor U10826 (N_10826,N_9914,N_9558);
xor U10827 (N_10827,N_8534,N_9484);
nor U10828 (N_10828,N_9149,N_8523);
nor U10829 (N_10829,N_9517,N_8438);
and U10830 (N_10830,N_8299,N_8172);
or U10831 (N_10831,N_9849,N_8521);
or U10832 (N_10832,N_7527,N_8772);
and U10833 (N_10833,N_9161,N_8706);
or U10834 (N_10834,N_8852,N_9608);
and U10835 (N_10835,N_7695,N_7893);
or U10836 (N_10836,N_9225,N_9332);
nand U10837 (N_10837,N_8252,N_8369);
xor U10838 (N_10838,N_9508,N_8944);
nor U10839 (N_10839,N_8933,N_7860);
or U10840 (N_10840,N_9896,N_8947);
xnor U10841 (N_10841,N_8096,N_9209);
nor U10842 (N_10842,N_8870,N_8095);
nand U10843 (N_10843,N_7614,N_8034);
nand U10844 (N_10844,N_8729,N_7925);
nor U10845 (N_10845,N_9380,N_9379);
or U10846 (N_10846,N_9217,N_8224);
nand U10847 (N_10847,N_7923,N_8514);
and U10848 (N_10848,N_7906,N_8682);
and U10849 (N_10849,N_9252,N_7669);
nor U10850 (N_10850,N_9670,N_9507);
nor U10851 (N_10851,N_8769,N_9382);
nor U10852 (N_10852,N_7863,N_9436);
nor U10853 (N_10853,N_8396,N_9951);
xnor U10854 (N_10854,N_9652,N_7542);
nand U10855 (N_10855,N_9269,N_9463);
nand U10856 (N_10856,N_8632,N_8741);
or U10857 (N_10857,N_8309,N_8467);
nand U10858 (N_10858,N_7810,N_9068);
nand U10859 (N_10859,N_9238,N_9014);
xnor U10860 (N_10860,N_9152,N_9208);
xnor U10861 (N_10861,N_7946,N_8009);
nor U10862 (N_10862,N_7656,N_8433);
nand U10863 (N_10863,N_9616,N_9110);
or U10864 (N_10864,N_8052,N_9134);
xor U10865 (N_10865,N_7886,N_8655);
nand U10866 (N_10866,N_8123,N_9665);
nor U10867 (N_10867,N_9823,N_8624);
nand U10868 (N_10868,N_8320,N_9994);
xnor U10869 (N_10869,N_8381,N_9057);
or U10870 (N_10870,N_7859,N_9196);
nand U10871 (N_10871,N_8071,N_7999);
and U10872 (N_10872,N_8264,N_8746);
nand U10873 (N_10873,N_9821,N_7523);
xnor U10874 (N_10874,N_9952,N_8178);
or U10875 (N_10875,N_9733,N_9936);
nand U10876 (N_10876,N_7569,N_8038);
nand U10877 (N_10877,N_8744,N_9054);
nor U10878 (N_10878,N_8218,N_7984);
xnor U10879 (N_10879,N_8085,N_9819);
or U10880 (N_10880,N_7754,N_7672);
nor U10881 (N_10881,N_9948,N_9395);
nand U10882 (N_10882,N_8456,N_7898);
nand U10883 (N_10883,N_8043,N_7748);
and U10884 (N_10884,N_9139,N_7924);
and U10885 (N_10885,N_9861,N_7941);
xnor U10886 (N_10886,N_9072,N_8756);
or U10887 (N_10887,N_8331,N_7731);
or U10888 (N_10888,N_8837,N_8468);
and U10889 (N_10889,N_8159,N_8668);
or U10890 (N_10890,N_9432,N_7670);
or U10891 (N_10891,N_8374,N_7847);
nor U10892 (N_10892,N_8579,N_8389);
nand U10893 (N_10893,N_9219,N_9374);
nor U10894 (N_10894,N_9781,N_8788);
nor U10895 (N_10895,N_9563,N_9889);
nand U10896 (N_10896,N_9522,N_9841);
and U10897 (N_10897,N_7516,N_9245);
or U10898 (N_10898,N_7730,N_9689);
xor U10899 (N_10899,N_8777,N_7705);
and U10900 (N_10900,N_9076,N_8833);
xnor U10901 (N_10901,N_9062,N_8473);
and U10902 (N_10902,N_9818,N_8296);
and U10903 (N_10903,N_8759,N_8859);
nand U10904 (N_10904,N_8463,N_7616);
xor U10905 (N_10905,N_8385,N_9855);
nand U10906 (N_10906,N_7793,N_8694);
nor U10907 (N_10907,N_7772,N_7942);
nand U10908 (N_10908,N_7737,N_7882);
nor U10909 (N_10909,N_9919,N_8155);
nor U10910 (N_10910,N_7749,N_9168);
nand U10911 (N_10911,N_9561,N_7532);
and U10912 (N_10912,N_9349,N_7572);
xor U10913 (N_10913,N_9120,N_8002);
nor U10914 (N_10914,N_9681,N_9184);
or U10915 (N_10915,N_7673,N_9433);
or U10916 (N_10916,N_9769,N_7714);
or U10917 (N_10917,N_9498,N_8298);
nor U10918 (N_10918,N_9469,N_8379);
or U10919 (N_10919,N_9182,N_7799);
nand U10920 (N_10920,N_9840,N_8277);
and U10921 (N_10921,N_8625,N_9192);
xnor U10922 (N_10922,N_8708,N_8209);
nand U10923 (N_10923,N_9312,N_8450);
or U10924 (N_10924,N_7661,N_9407);
nor U10925 (N_10925,N_8609,N_8914);
xor U10926 (N_10926,N_9089,N_8734);
or U10927 (N_10927,N_7949,N_7597);
xor U10928 (N_10928,N_8007,N_9625);
nor U10929 (N_10929,N_9173,N_7861);
nor U10930 (N_10930,N_9230,N_9715);
nor U10931 (N_10931,N_8806,N_9701);
nor U10932 (N_10932,N_8200,N_8667);
nor U10933 (N_10933,N_8260,N_9066);
nor U10934 (N_10934,N_9025,N_8230);
xor U10935 (N_10935,N_9320,N_7921);
and U10936 (N_10936,N_9319,N_7703);
nor U10937 (N_10937,N_9538,N_8194);
nor U10938 (N_10938,N_8083,N_7605);
xor U10939 (N_10939,N_8617,N_8985);
xnor U10940 (N_10940,N_7951,N_8622);
and U10941 (N_10941,N_8174,N_8245);
nor U10942 (N_10942,N_9806,N_7715);
nand U10943 (N_10943,N_7777,N_9905);
nand U10944 (N_10944,N_8816,N_8423);
nand U10945 (N_10945,N_8109,N_8372);
xor U10946 (N_10946,N_8390,N_8366);
xnor U10947 (N_10947,N_7965,N_9289);
nand U10948 (N_10948,N_9934,N_8093);
or U10949 (N_10949,N_8836,N_9279);
nor U10950 (N_10950,N_9384,N_8671);
nand U10951 (N_10951,N_7630,N_9993);
and U10952 (N_10952,N_9615,N_7930);
and U10953 (N_10953,N_9989,N_9611);
xnor U10954 (N_10954,N_8393,N_8250);
nand U10955 (N_10955,N_9980,N_8752);
nor U10956 (N_10956,N_7721,N_8183);
xnor U10957 (N_10957,N_8537,N_7817);
nor U10958 (N_10958,N_7660,N_7524);
xor U10959 (N_10959,N_9911,N_8968);
and U10960 (N_10960,N_8952,N_8221);
nand U10961 (N_10961,N_9188,N_7513);
xor U10962 (N_10962,N_9604,N_8271);
nor U10963 (N_10963,N_8132,N_8512);
xnor U10964 (N_10964,N_8373,N_8064);
and U10965 (N_10965,N_9954,N_9898);
nand U10966 (N_10966,N_8145,N_8188);
nand U10967 (N_10967,N_8027,N_9762);
xnor U10968 (N_10968,N_8241,N_9853);
nand U10969 (N_10969,N_9092,N_8636);
xor U10970 (N_10970,N_8796,N_7928);
or U10971 (N_10971,N_8740,N_7808);
nor U10972 (N_10972,N_7665,N_9973);
xnor U10973 (N_10973,N_7842,N_8635);
or U10974 (N_10974,N_7980,N_8068);
xnor U10975 (N_10975,N_9734,N_7758);
xnor U10976 (N_10976,N_8540,N_8884);
xor U10977 (N_10977,N_7974,N_8242);
and U10978 (N_10978,N_9672,N_8280);
xnor U10979 (N_10979,N_7914,N_8665);
xnor U10980 (N_10980,N_8310,N_8863);
xnor U10981 (N_10981,N_9117,N_7932);
xor U10982 (N_10982,N_8907,N_9541);
nand U10983 (N_10983,N_8403,N_7954);
and U10984 (N_10984,N_8890,N_8457);
xnor U10985 (N_10985,N_7540,N_8019);
and U10986 (N_10986,N_9097,N_9058);
nand U10987 (N_10987,N_7622,N_7668);
nand U10988 (N_10988,N_9876,N_8380);
xnor U10989 (N_10989,N_7896,N_8998);
xor U10990 (N_10990,N_7764,N_9050);
nand U10991 (N_10991,N_8896,N_8591);
and U10992 (N_10992,N_8705,N_9938);
or U10993 (N_10993,N_8693,N_8950);
or U10994 (N_10994,N_8488,N_7595);
and U10995 (N_10995,N_9530,N_7659);
or U10996 (N_10996,N_8910,N_8337);
nor U10997 (N_10997,N_9167,N_8075);
xor U10998 (N_10998,N_9359,N_8964);
nor U10999 (N_10999,N_7982,N_8557);
or U11000 (N_11000,N_9102,N_9494);
xor U11001 (N_11001,N_9749,N_8378);
nor U11002 (N_11002,N_7778,N_8692);
or U11003 (N_11003,N_8602,N_8204);
xnor U11004 (N_11004,N_9434,N_8059);
and U11005 (N_11005,N_7937,N_9763);
and U11006 (N_11006,N_9470,N_9304);
and U11007 (N_11007,N_8929,N_7854);
and U11008 (N_11008,N_8793,N_9000);
and U11009 (N_11009,N_7518,N_9750);
xnor U11010 (N_11010,N_9194,N_8409);
xor U11011 (N_11011,N_8476,N_8916);
nor U11012 (N_11012,N_7727,N_9804);
xnor U11013 (N_11013,N_8629,N_7637);
nand U11014 (N_11014,N_9826,N_8821);
nor U11015 (N_11015,N_9310,N_7825);
nand U11016 (N_11016,N_9016,N_8115);
nor U11017 (N_11017,N_8180,N_8992);
nand U11018 (N_11018,N_9487,N_7620);
and U11019 (N_11019,N_8329,N_9735);
or U11020 (N_11020,N_7876,N_7962);
or U11021 (N_11021,N_7551,N_7701);
nor U11022 (N_11022,N_8451,N_7621);
nor U11023 (N_11023,N_9264,N_7591);
nor U11024 (N_11024,N_9941,N_9772);
and U11025 (N_11025,N_8880,N_7910);
and U11026 (N_11026,N_9115,N_9760);
or U11027 (N_11027,N_9784,N_7687);
nor U11028 (N_11028,N_9236,N_9291);
and U11029 (N_11029,N_8979,N_9596);
or U11030 (N_11030,N_8432,N_9873);
nand U11031 (N_11031,N_9403,N_9771);
nand U11032 (N_11032,N_9984,N_9564);
xnor U11033 (N_11033,N_8405,N_7856);
or U11034 (N_11034,N_7537,N_9908);
xor U11035 (N_11035,N_8112,N_9020);
nand U11036 (N_11036,N_9600,N_7994);
and U11037 (N_11037,N_8014,N_9378);
xnor U11038 (N_11038,N_9143,N_8087);
or U11039 (N_11039,N_8258,N_9203);
or U11040 (N_11040,N_8711,N_7678);
nand U11041 (N_11041,N_7968,N_8898);
nor U11042 (N_11042,N_9544,N_9791);
nor U11043 (N_11043,N_9972,N_9935);
xor U11044 (N_11044,N_8367,N_8642);
xor U11045 (N_11045,N_8192,N_9782);
and U11046 (N_11046,N_9007,N_8688);
or U11047 (N_11047,N_8437,N_9313);
and U11048 (N_11048,N_9087,N_9702);
nor U11049 (N_11049,N_7719,N_8531);
and U11050 (N_11050,N_8460,N_8849);
nor U11051 (N_11051,N_8586,N_8492);
and U11052 (N_11052,N_9059,N_8036);
and U11053 (N_11053,N_9276,N_7674);
and U11054 (N_11054,N_9222,N_7667);
nand U11055 (N_11055,N_9904,N_9454);
or U11056 (N_11056,N_9960,N_7769);
xor U11057 (N_11057,N_9376,N_7554);
nor U11058 (N_11058,N_8441,N_8058);
and U11059 (N_11059,N_8222,N_9645);
nand U11060 (N_11060,N_9270,N_8382);
nand U11061 (N_11061,N_9499,N_8649);
xnor U11062 (N_11062,N_9795,N_9146);
or U11063 (N_11063,N_8016,N_8066);
xor U11064 (N_11064,N_8436,N_9383);
and U11065 (N_11065,N_8121,N_9405);
and U11066 (N_11066,N_9695,N_7988);
nor U11067 (N_11067,N_8049,N_8203);
and U11068 (N_11068,N_9413,N_7844);
nand U11069 (N_11069,N_9958,N_9575);
or U11070 (N_11070,N_9895,N_8341);
nand U11071 (N_11071,N_9957,N_8748);
nand U11072 (N_11072,N_9692,N_7664);
nor U11073 (N_11073,N_8841,N_9916);
xnor U11074 (N_11074,N_8571,N_8319);
xor U11075 (N_11075,N_7902,N_9260);
or U11076 (N_11076,N_9045,N_9133);
nand U11077 (N_11077,N_8127,N_8119);
or U11078 (N_11078,N_9807,N_8627);
or U11079 (N_11079,N_9137,N_9492);
nand U11080 (N_11080,N_7663,N_9890);
or U11081 (N_11081,N_8278,N_7649);
xnor U11082 (N_11082,N_8814,N_8131);
xor U11083 (N_11083,N_9280,N_9656);
nor U11084 (N_11084,N_9233,N_9503);
nor U11085 (N_11085,N_7868,N_8812);
nor U11086 (N_11086,N_9710,N_7774);
nand U11087 (N_11087,N_8413,N_7598);
or U11088 (N_11088,N_9825,N_8262);
nor U11089 (N_11089,N_9835,N_8847);
or U11090 (N_11090,N_9193,N_8376);
or U11091 (N_11091,N_8825,N_9912);
nor U11092 (N_11092,N_8138,N_8973);
and U11093 (N_11093,N_8279,N_9388);
or U11094 (N_11094,N_8530,N_9632);
and U11095 (N_11095,N_9286,N_9676);
or U11096 (N_11096,N_8751,N_8349);
nor U11097 (N_11097,N_9031,N_9126);
nor U11098 (N_11098,N_9414,N_9621);
and U11099 (N_11099,N_9968,N_7556);
or U11100 (N_11100,N_9768,N_9140);
nor U11101 (N_11101,N_8699,N_9202);
xnor U11102 (N_11102,N_9922,N_8828);
nand U11103 (N_11103,N_9085,N_8090);
nand U11104 (N_11104,N_9051,N_9891);
and U11105 (N_11105,N_7508,N_9613);
and U11106 (N_11106,N_8079,N_8643);
xor U11107 (N_11107,N_9288,N_8255);
nand U11108 (N_11108,N_7751,N_8739);
nand U11109 (N_11109,N_8113,N_8461);
or U11110 (N_11110,N_8065,N_7858);
nor U11111 (N_11111,N_8455,N_8040);
nor U11112 (N_11112,N_8662,N_8134);
nor U11113 (N_11113,N_8840,N_9362);
nor U11114 (N_11114,N_8685,N_9086);
and U11115 (N_11115,N_9809,N_8462);
or U11116 (N_11116,N_8593,N_9373);
and U11117 (N_11117,N_9220,N_8563);
nand U11118 (N_11118,N_9428,N_9029);
or U11119 (N_11119,N_8760,N_7684);
and U11120 (N_11120,N_8520,N_9108);
and U11121 (N_11121,N_9504,N_7546);
xor U11122 (N_11122,N_9242,N_8039);
nand U11123 (N_11123,N_9190,N_9318);
nor U11124 (N_11124,N_7653,N_8206);
nand U11125 (N_11125,N_8620,N_9669);
nor U11126 (N_11126,N_9452,N_7629);
xor U11127 (N_11127,N_9590,N_9816);
xnor U11128 (N_11128,N_7712,N_8246);
xnor U11129 (N_11129,N_9510,N_9713);
nor U11130 (N_11130,N_9255,N_8527);
nor U11131 (N_11131,N_8345,N_8976);
or U11132 (N_11132,N_8641,N_7929);
and U11133 (N_11133,N_9262,N_9495);
nand U11134 (N_11134,N_7961,N_9478);
or U11135 (N_11135,N_8967,N_8513);
nand U11136 (N_11136,N_8547,N_8648);
nand U11137 (N_11137,N_8725,N_8867);
nand U11138 (N_11138,N_9336,N_9258);
or U11139 (N_11139,N_9982,N_8790);
or U11140 (N_11140,N_9391,N_8509);
nor U11141 (N_11141,N_9740,N_7972);
nor U11142 (N_11142,N_9893,N_9237);
xor U11143 (N_11143,N_8384,N_8835);
or U11144 (N_11144,N_7787,N_9961);
xnor U11145 (N_11145,N_8802,N_7798);
or U11146 (N_11146,N_9752,N_8719);
nor U11147 (N_11147,N_9448,N_7805);
nor U11148 (N_11148,N_8428,N_9836);
xnor U11149 (N_11149,N_8696,N_9325);
nor U11150 (N_11150,N_7747,N_7526);
xor U11151 (N_11151,N_7815,N_8105);
xor U11152 (N_11152,N_9909,N_8554);
xnor U11153 (N_11153,N_7905,N_8157);
or U11154 (N_11154,N_9179,N_9154);
nand U11155 (N_11155,N_9629,N_9228);
or U11156 (N_11156,N_9967,N_9566);
nand U11157 (N_11157,N_7517,N_9067);
nand U11158 (N_11158,N_8658,N_9759);
nand U11159 (N_11159,N_7765,N_7759);
and U11160 (N_11160,N_7839,N_7536);
and U11161 (N_11161,N_9546,N_7796);
nand U11162 (N_11162,N_8737,N_9078);
nand U11163 (N_11163,N_9135,N_8305);
or U11164 (N_11164,N_8215,N_8358);
or U11165 (N_11165,N_8326,N_8839);
nor U11166 (N_11166,N_8082,N_9830);
and U11167 (N_11167,N_8578,N_7646);
or U11168 (N_11168,N_8238,N_8608);
nor U11169 (N_11169,N_7690,N_8864);
nor U11170 (N_11170,N_9683,N_9619);
xor U11171 (N_11171,N_9592,N_9744);
and U11172 (N_11172,N_7838,N_9234);
xnor U11173 (N_11173,N_8004,N_7600);
xnor U11174 (N_11174,N_7718,N_9844);
and U11175 (N_11175,N_9447,N_9011);
xor U11176 (N_11176,N_9868,N_9005);
nand U11177 (N_11177,N_9048,N_9489);
xor U11178 (N_11178,N_9022,N_9638);
or U11179 (N_11179,N_8072,N_7588);
xnor U11180 (N_11180,N_8103,N_8785);
or U11181 (N_11181,N_8700,N_8659);
or U11182 (N_11182,N_9351,N_9352);
and U11183 (N_11183,N_7521,N_7922);
xor U11184 (N_11184,N_9145,N_9587);
or U11185 (N_11185,N_7807,N_8946);
or U11186 (N_11186,N_9417,N_8273);
and U11187 (N_11187,N_9353,N_9077);
nand U11188 (N_11188,N_9346,N_9691);
nand U11189 (N_11189,N_8147,N_7770);
and U11190 (N_11190,N_9023,N_9175);
and U11191 (N_11191,N_8982,N_9979);
nand U11192 (N_11192,N_8431,N_9677);
nor U11193 (N_11193,N_9337,N_9950);
or U11194 (N_11194,N_7934,N_8544);
and U11195 (N_11195,N_9399,N_9287);
nand U11196 (N_11196,N_8249,N_8986);
and U11197 (N_11197,N_9497,N_9595);
xor U11198 (N_11198,N_7686,N_8801);
and U11199 (N_11199,N_9158,N_8656);
and U11200 (N_11200,N_8974,N_9367);
nand U11201 (N_11201,N_8398,N_8073);
or U11202 (N_11202,N_7500,N_9946);
xnor U11203 (N_11203,N_7575,N_7992);
or U11204 (N_11204,N_9719,N_9598);
nor U11205 (N_11205,N_8731,N_7603);
xnor U11206 (N_11206,N_9420,N_7611);
and U11207 (N_11207,N_7587,N_9261);
and U11208 (N_11208,N_9437,N_8033);
nor U11209 (N_11209,N_9144,N_8128);
nor U11210 (N_11210,N_7768,N_8948);
nand U11211 (N_11211,N_7904,N_8723);
nand U11212 (N_11212,N_8184,N_8179);
or U11213 (N_11213,N_9773,N_9501);
nor U11214 (N_11214,N_7639,N_8028);
xor U11215 (N_11215,N_7983,N_9591);
nand U11216 (N_11216,N_8452,N_7519);
and U11217 (N_11217,N_8993,N_9721);
xnor U11218 (N_11218,N_8990,N_8631);
nor U11219 (N_11219,N_9091,N_9465);
nor U11220 (N_11220,N_8980,N_9520);
or U11221 (N_11221,N_8125,N_8860);
xnor U11222 (N_11222,N_9027,N_7555);
nor U11223 (N_11223,N_9822,N_8327);
and U11224 (N_11224,N_7596,N_9350);
and U11225 (N_11225,N_9990,N_7976);
and U11226 (N_11226,N_8294,N_9305);
or U11227 (N_11227,N_9800,N_7950);
xnor U11228 (N_11228,N_8177,N_8325);
or U11229 (N_11229,N_8745,N_7707);
nor U11230 (N_11230,N_7909,N_9755);
nand U11231 (N_11231,N_9277,N_7776);
xnor U11232 (N_11232,N_7533,N_8030);
xor U11233 (N_11233,N_9080,N_8911);
xor U11234 (N_11234,N_8012,N_8991);
nand U11235 (N_11235,N_9096,N_9160);
xor U11236 (N_11236,N_8098,N_9357);
nand U11237 (N_11237,N_8634,N_8339);
nand U11238 (N_11238,N_9042,N_8418);
xnor U11239 (N_11239,N_8792,N_9250);
nand U11240 (N_11240,N_9850,N_9061);
nand U11241 (N_11241,N_7958,N_9897);
nand U11242 (N_11242,N_9730,N_7565);
and U11243 (N_11243,N_8614,N_8046);
xnor U11244 (N_11244,N_9963,N_8670);
xor U11245 (N_11245,N_7848,N_9630);
or U11246 (N_11246,N_8361,N_8966);
or U11247 (N_11247,N_7723,N_9883);
xnor U11248 (N_11248,N_7689,N_8607);
and U11249 (N_11249,N_9232,N_9685);
nor U11250 (N_11250,N_7741,N_9641);
nor U11251 (N_11251,N_7644,N_8560);
xor U11252 (N_11252,N_9871,N_7694);
or U11253 (N_11253,N_7906,N_8417);
or U11254 (N_11254,N_9046,N_9341);
or U11255 (N_11255,N_9786,N_9562);
nand U11256 (N_11256,N_8444,N_9465);
nand U11257 (N_11257,N_9622,N_8898);
xor U11258 (N_11258,N_9229,N_9971);
nor U11259 (N_11259,N_9531,N_8958);
and U11260 (N_11260,N_8247,N_9259);
nor U11261 (N_11261,N_7886,N_8658);
xnor U11262 (N_11262,N_7656,N_7741);
nor U11263 (N_11263,N_8600,N_8008);
nand U11264 (N_11264,N_8962,N_8711);
xor U11265 (N_11265,N_9601,N_8115);
nor U11266 (N_11266,N_9841,N_9445);
nand U11267 (N_11267,N_8803,N_9551);
nor U11268 (N_11268,N_7598,N_9766);
or U11269 (N_11269,N_9029,N_7732);
nand U11270 (N_11270,N_8961,N_9276);
nor U11271 (N_11271,N_8069,N_9452);
or U11272 (N_11272,N_9225,N_8980);
or U11273 (N_11273,N_9386,N_8624);
xor U11274 (N_11274,N_8946,N_9505);
nor U11275 (N_11275,N_7910,N_9316);
nand U11276 (N_11276,N_9869,N_9034);
xor U11277 (N_11277,N_9102,N_9089);
nor U11278 (N_11278,N_9521,N_8991);
xor U11279 (N_11279,N_8923,N_8232);
xnor U11280 (N_11280,N_9874,N_7743);
and U11281 (N_11281,N_7510,N_8350);
nand U11282 (N_11282,N_8751,N_9805);
xor U11283 (N_11283,N_9130,N_8400);
or U11284 (N_11284,N_7595,N_7693);
xor U11285 (N_11285,N_7913,N_8476);
nor U11286 (N_11286,N_8073,N_9285);
nor U11287 (N_11287,N_9850,N_8108);
nand U11288 (N_11288,N_9457,N_7771);
nor U11289 (N_11289,N_9974,N_9092);
and U11290 (N_11290,N_9629,N_8006);
xor U11291 (N_11291,N_8844,N_7593);
nor U11292 (N_11292,N_9287,N_7912);
xor U11293 (N_11293,N_9402,N_7673);
nor U11294 (N_11294,N_9776,N_9545);
nor U11295 (N_11295,N_9187,N_7531);
nand U11296 (N_11296,N_7520,N_7602);
or U11297 (N_11297,N_9108,N_7541);
nand U11298 (N_11298,N_9222,N_9175);
nor U11299 (N_11299,N_7863,N_8727);
nand U11300 (N_11300,N_8149,N_9330);
or U11301 (N_11301,N_8016,N_7608);
and U11302 (N_11302,N_7993,N_9899);
nand U11303 (N_11303,N_9222,N_8427);
and U11304 (N_11304,N_9291,N_9724);
nor U11305 (N_11305,N_7632,N_8098);
xor U11306 (N_11306,N_7590,N_9628);
nand U11307 (N_11307,N_8580,N_9318);
nand U11308 (N_11308,N_9775,N_7606);
xnor U11309 (N_11309,N_7826,N_8980);
nor U11310 (N_11310,N_9481,N_8060);
or U11311 (N_11311,N_8566,N_9537);
nand U11312 (N_11312,N_8237,N_9905);
xnor U11313 (N_11313,N_9832,N_9911);
nand U11314 (N_11314,N_8233,N_8466);
xnor U11315 (N_11315,N_9205,N_9061);
or U11316 (N_11316,N_9770,N_9361);
nand U11317 (N_11317,N_7887,N_7770);
or U11318 (N_11318,N_9645,N_9683);
nor U11319 (N_11319,N_9231,N_7631);
xor U11320 (N_11320,N_9186,N_8468);
nand U11321 (N_11321,N_7847,N_7986);
and U11322 (N_11322,N_9169,N_9008);
or U11323 (N_11323,N_8567,N_9952);
nand U11324 (N_11324,N_8102,N_9600);
nand U11325 (N_11325,N_7647,N_8979);
xnor U11326 (N_11326,N_8981,N_8616);
nand U11327 (N_11327,N_8907,N_8942);
nor U11328 (N_11328,N_8618,N_9112);
and U11329 (N_11329,N_8728,N_8765);
xnor U11330 (N_11330,N_7633,N_9396);
and U11331 (N_11331,N_9106,N_9176);
xor U11332 (N_11332,N_7615,N_9067);
xor U11333 (N_11333,N_9272,N_8923);
nand U11334 (N_11334,N_8452,N_8934);
nor U11335 (N_11335,N_9391,N_9477);
xor U11336 (N_11336,N_9600,N_9138);
nor U11337 (N_11337,N_7716,N_8628);
nor U11338 (N_11338,N_9620,N_7866);
xor U11339 (N_11339,N_8107,N_9883);
nor U11340 (N_11340,N_8210,N_9754);
xnor U11341 (N_11341,N_8579,N_9408);
and U11342 (N_11342,N_8185,N_8235);
nor U11343 (N_11343,N_7756,N_9128);
or U11344 (N_11344,N_9084,N_8198);
or U11345 (N_11345,N_8044,N_8380);
xor U11346 (N_11346,N_7923,N_8366);
nand U11347 (N_11347,N_9050,N_9127);
and U11348 (N_11348,N_8926,N_9898);
xnor U11349 (N_11349,N_7622,N_9701);
and U11350 (N_11350,N_9898,N_8094);
or U11351 (N_11351,N_9708,N_7649);
nor U11352 (N_11352,N_9608,N_9433);
nor U11353 (N_11353,N_9841,N_8632);
nand U11354 (N_11354,N_8126,N_9373);
and U11355 (N_11355,N_9782,N_7599);
xnor U11356 (N_11356,N_8632,N_9627);
and U11357 (N_11357,N_7850,N_7580);
and U11358 (N_11358,N_7872,N_7642);
and U11359 (N_11359,N_8347,N_8918);
nor U11360 (N_11360,N_8131,N_8439);
or U11361 (N_11361,N_8210,N_8432);
xor U11362 (N_11362,N_9948,N_8587);
and U11363 (N_11363,N_7708,N_8074);
nor U11364 (N_11364,N_9390,N_8096);
and U11365 (N_11365,N_8443,N_8999);
or U11366 (N_11366,N_7890,N_8345);
nor U11367 (N_11367,N_8356,N_9013);
and U11368 (N_11368,N_8317,N_9248);
xnor U11369 (N_11369,N_8851,N_8117);
xnor U11370 (N_11370,N_8024,N_7822);
and U11371 (N_11371,N_8201,N_9815);
xor U11372 (N_11372,N_7550,N_9823);
nor U11373 (N_11373,N_7684,N_8083);
nor U11374 (N_11374,N_8016,N_8756);
or U11375 (N_11375,N_9361,N_9211);
xnor U11376 (N_11376,N_9749,N_7687);
xor U11377 (N_11377,N_9566,N_7845);
and U11378 (N_11378,N_9562,N_9642);
and U11379 (N_11379,N_8420,N_8771);
and U11380 (N_11380,N_7547,N_9119);
nand U11381 (N_11381,N_8677,N_8870);
xor U11382 (N_11382,N_9414,N_7662);
xnor U11383 (N_11383,N_7716,N_9328);
xor U11384 (N_11384,N_8928,N_9397);
nor U11385 (N_11385,N_8884,N_8088);
nand U11386 (N_11386,N_8342,N_7569);
and U11387 (N_11387,N_9013,N_9196);
or U11388 (N_11388,N_8366,N_9424);
and U11389 (N_11389,N_9192,N_7867);
nor U11390 (N_11390,N_7670,N_9568);
or U11391 (N_11391,N_7962,N_9609);
xor U11392 (N_11392,N_9713,N_7667);
or U11393 (N_11393,N_9015,N_9246);
or U11394 (N_11394,N_8276,N_7845);
or U11395 (N_11395,N_8597,N_8646);
nor U11396 (N_11396,N_7736,N_9420);
nor U11397 (N_11397,N_9521,N_7976);
nand U11398 (N_11398,N_8034,N_7749);
xor U11399 (N_11399,N_8166,N_8522);
xor U11400 (N_11400,N_8564,N_8468);
or U11401 (N_11401,N_7863,N_9502);
and U11402 (N_11402,N_9637,N_8009);
xor U11403 (N_11403,N_8830,N_7956);
and U11404 (N_11404,N_8455,N_9171);
and U11405 (N_11405,N_7628,N_9634);
and U11406 (N_11406,N_7947,N_8280);
nor U11407 (N_11407,N_8474,N_9231);
nor U11408 (N_11408,N_9438,N_9085);
and U11409 (N_11409,N_9042,N_9791);
and U11410 (N_11410,N_9837,N_9106);
nand U11411 (N_11411,N_9515,N_8474);
nor U11412 (N_11412,N_8103,N_8352);
nand U11413 (N_11413,N_7683,N_9736);
xnor U11414 (N_11414,N_8891,N_9752);
nor U11415 (N_11415,N_9005,N_9296);
nand U11416 (N_11416,N_9749,N_9802);
and U11417 (N_11417,N_9370,N_9538);
nand U11418 (N_11418,N_8815,N_9389);
nand U11419 (N_11419,N_7942,N_9434);
and U11420 (N_11420,N_9493,N_7526);
xnor U11421 (N_11421,N_9733,N_9990);
xnor U11422 (N_11422,N_9815,N_8636);
nand U11423 (N_11423,N_7962,N_9117);
nand U11424 (N_11424,N_9731,N_9953);
nand U11425 (N_11425,N_9356,N_9247);
and U11426 (N_11426,N_8844,N_8806);
xnor U11427 (N_11427,N_8746,N_7950);
xor U11428 (N_11428,N_9571,N_8174);
nor U11429 (N_11429,N_8695,N_8000);
nand U11430 (N_11430,N_7587,N_9611);
or U11431 (N_11431,N_8177,N_8441);
or U11432 (N_11432,N_8516,N_9895);
nor U11433 (N_11433,N_7628,N_7813);
and U11434 (N_11434,N_8751,N_8974);
xor U11435 (N_11435,N_8550,N_8544);
or U11436 (N_11436,N_9184,N_8716);
and U11437 (N_11437,N_9805,N_7738);
xnor U11438 (N_11438,N_9738,N_9338);
or U11439 (N_11439,N_9092,N_9433);
xnor U11440 (N_11440,N_8991,N_9402);
xor U11441 (N_11441,N_9570,N_7689);
or U11442 (N_11442,N_8317,N_9885);
xor U11443 (N_11443,N_7701,N_9205);
or U11444 (N_11444,N_7743,N_8520);
nor U11445 (N_11445,N_7631,N_8254);
xor U11446 (N_11446,N_8336,N_8692);
nand U11447 (N_11447,N_8104,N_9706);
xor U11448 (N_11448,N_8106,N_9798);
or U11449 (N_11449,N_7886,N_8281);
and U11450 (N_11450,N_8825,N_9142);
xnor U11451 (N_11451,N_9892,N_8700);
and U11452 (N_11452,N_8595,N_9603);
nor U11453 (N_11453,N_7913,N_8438);
nand U11454 (N_11454,N_9587,N_9741);
nand U11455 (N_11455,N_9727,N_8114);
or U11456 (N_11456,N_7743,N_9465);
xor U11457 (N_11457,N_9733,N_8596);
nand U11458 (N_11458,N_9488,N_8507);
xnor U11459 (N_11459,N_7661,N_9682);
nand U11460 (N_11460,N_8242,N_8634);
and U11461 (N_11461,N_8033,N_8210);
nand U11462 (N_11462,N_9707,N_8328);
nor U11463 (N_11463,N_9834,N_7917);
or U11464 (N_11464,N_9282,N_7670);
xor U11465 (N_11465,N_7805,N_9611);
nor U11466 (N_11466,N_8182,N_7596);
or U11467 (N_11467,N_9683,N_7536);
nor U11468 (N_11468,N_9216,N_9466);
nand U11469 (N_11469,N_9343,N_9391);
and U11470 (N_11470,N_9771,N_9855);
or U11471 (N_11471,N_8370,N_8112);
or U11472 (N_11472,N_8800,N_9165);
xnor U11473 (N_11473,N_8474,N_9151);
nand U11474 (N_11474,N_9369,N_8681);
and U11475 (N_11475,N_8214,N_8326);
xnor U11476 (N_11476,N_7594,N_9143);
nand U11477 (N_11477,N_9787,N_9520);
nor U11478 (N_11478,N_8130,N_9812);
or U11479 (N_11479,N_8020,N_8127);
xor U11480 (N_11480,N_9738,N_8458);
nor U11481 (N_11481,N_8585,N_8766);
or U11482 (N_11482,N_8158,N_8977);
xnor U11483 (N_11483,N_8115,N_9194);
nor U11484 (N_11484,N_9481,N_9261);
or U11485 (N_11485,N_8098,N_8652);
and U11486 (N_11486,N_9134,N_8589);
nor U11487 (N_11487,N_8301,N_7522);
nor U11488 (N_11488,N_9149,N_8630);
xnor U11489 (N_11489,N_7589,N_8922);
xnor U11490 (N_11490,N_9487,N_8645);
xor U11491 (N_11491,N_9336,N_8147);
or U11492 (N_11492,N_9520,N_9583);
nor U11493 (N_11493,N_8522,N_9377);
nand U11494 (N_11494,N_7860,N_9681);
nand U11495 (N_11495,N_9978,N_7908);
nor U11496 (N_11496,N_9207,N_9773);
xnor U11497 (N_11497,N_7579,N_9623);
xor U11498 (N_11498,N_8844,N_9415);
or U11499 (N_11499,N_7848,N_9856);
nor U11500 (N_11500,N_7831,N_7506);
xnor U11501 (N_11501,N_9514,N_7690);
xor U11502 (N_11502,N_7605,N_7933);
or U11503 (N_11503,N_8837,N_7654);
nor U11504 (N_11504,N_9346,N_8790);
nand U11505 (N_11505,N_8735,N_9090);
nand U11506 (N_11506,N_8241,N_7712);
nor U11507 (N_11507,N_8571,N_8867);
or U11508 (N_11508,N_9060,N_8180);
nor U11509 (N_11509,N_8550,N_8092);
and U11510 (N_11510,N_8986,N_9945);
nand U11511 (N_11511,N_8042,N_8542);
nand U11512 (N_11512,N_9645,N_7588);
or U11513 (N_11513,N_8970,N_9199);
nand U11514 (N_11514,N_9339,N_7540);
xnor U11515 (N_11515,N_8599,N_8776);
or U11516 (N_11516,N_7696,N_7947);
and U11517 (N_11517,N_7621,N_8358);
and U11518 (N_11518,N_8287,N_8660);
and U11519 (N_11519,N_8310,N_9901);
or U11520 (N_11520,N_9028,N_9761);
nor U11521 (N_11521,N_8351,N_8249);
and U11522 (N_11522,N_9276,N_9705);
xor U11523 (N_11523,N_9958,N_8818);
nand U11524 (N_11524,N_7830,N_8533);
nor U11525 (N_11525,N_9676,N_9911);
nand U11526 (N_11526,N_9735,N_8681);
nand U11527 (N_11527,N_9914,N_9764);
or U11528 (N_11528,N_8245,N_9017);
and U11529 (N_11529,N_8953,N_9294);
nand U11530 (N_11530,N_8616,N_7778);
nor U11531 (N_11531,N_8107,N_8506);
nand U11532 (N_11532,N_9990,N_9022);
nor U11533 (N_11533,N_8125,N_8523);
nor U11534 (N_11534,N_9721,N_9754);
or U11535 (N_11535,N_9691,N_7988);
xor U11536 (N_11536,N_8229,N_9738);
nor U11537 (N_11537,N_8317,N_8675);
and U11538 (N_11538,N_7656,N_8287);
nor U11539 (N_11539,N_7905,N_7917);
or U11540 (N_11540,N_8074,N_8387);
and U11541 (N_11541,N_9954,N_8498);
nor U11542 (N_11542,N_9246,N_8959);
nor U11543 (N_11543,N_7508,N_9024);
or U11544 (N_11544,N_8092,N_9460);
nor U11545 (N_11545,N_9510,N_8387);
or U11546 (N_11546,N_8455,N_8980);
xnor U11547 (N_11547,N_8946,N_9219);
xnor U11548 (N_11548,N_8016,N_9838);
nand U11549 (N_11549,N_9993,N_8043);
and U11550 (N_11550,N_9984,N_8234);
nor U11551 (N_11551,N_8303,N_9168);
nor U11552 (N_11552,N_8896,N_8221);
nor U11553 (N_11553,N_7746,N_8294);
or U11554 (N_11554,N_8729,N_7971);
or U11555 (N_11555,N_8707,N_9732);
xor U11556 (N_11556,N_8705,N_9921);
nand U11557 (N_11557,N_8518,N_9163);
or U11558 (N_11558,N_8713,N_9502);
nor U11559 (N_11559,N_8602,N_9120);
nand U11560 (N_11560,N_9020,N_8543);
and U11561 (N_11561,N_9319,N_7634);
nor U11562 (N_11562,N_9668,N_8617);
nand U11563 (N_11563,N_8647,N_9092);
and U11564 (N_11564,N_7628,N_8594);
or U11565 (N_11565,N_8449,N_9663);
nor U11566 (N_11566,N_8359,N_8339);
or U11567 (N_11567,N_8872,N_7714);
nor U11568 (N_11568,N_9757,N_9800);
and U11569 (N_11569,N_8492,N_8727);
nor U11570 (N_11570,N_9530,N_8301);
xor U11571 (N_11571,N_8673,N_9974);
xnor U11572 (N_11572,N_9378,N_8369);
and U11573 (N_11573,N_8775,N_7822);
nor U11574 (N_11574,N_8877,N_9599);
and U11575 (N_11575,N_7993,N_9081);
nor U11576 (N_11576,N_8996,N_9240);
or U11577 (N_11577,N_9825,N_9386);
nor U11578 (N_11578,N_8329,N_7843);
xnor U11579 (N_11579,N_9556,N_7652);
or U11580 (N_11580,N_8995,N_9437);
and U11581 (N_11581,N_8851,N_7760);
or U11582 (N_11582,N_7856,N_7811);
and U11583 (N_11583,N_9292,N_9430);
or U11584 (N_11584,N_8482,N_9265);
and U11585 (N_11585,N_9145,N_9598);
xnor U11586 (N_11586,N_8429,N_9990);
and U11587 (N_11587,N_7934,N_8419);
nand U11588 (N_11588,N_9227,N_8557);
xnor U11589 (N_11589,N_8046,N_9354);
xor U11590 (N_11590,N_8893,N_8594);
and U11591 (N_11591,N_8076,N_8106);
nand U11592 (N_11592,N_9836,N_8277);
nor U11593 (N_11593,N_7525,N_8317);
nand U11594 (N_11594,N_9302,N_9404);
nand U11595 (N_11595,N_8168,N_9164);
xor U11596 (N_11596,N_8163,N_9812);
nand U11597 (N_11597,N_8009,N_7751);
nor U11598 (N_11598,N_8031,N_9771);
nand U11599 (N_11599,N_9635,N_8573);
xor U11600 (N_11600,N_9086,N_9073);
or U11601 (N_11601,N_8619,N_9760);
nor U11602 (N_11602,N_7884,N_8313);
nand U11603 (N_11603,N_7599,N_8860);
or U11604 (N_11604,N_8987,N_8594);
and U11605 (N_11605,N_7910,N_9575);
nor U11606 (N_11606,N_7990,N_8507);
nand U11607 (N_11607,N_8013,N_8375);
nand U11608 (N_11608,N_8909,N_8367);
nand U11609 (N_11609,N_9714,N_9738);
or U11610 (N_11610,N_7657,N_8325);
and U11611 (N_11611,N_9420,N_8022);
or U11612 (N_11612,N_8444,N_9104);
nor U11613 (N_11613,N_7976,N_9712);
or U11614 (N_11614,N_7735,N_7714);
nor U11615 (N_11615,N_9582,N_9995);
and U11616 (N_11616,N_8091,N_9619);
or U11617 (N_11617,N_9931,N_7500);
or U11618 (N_11618,N_9964,N_8942);
xor U11619 (N_11619,N_7864,N_8204);
nor U11620 (N_11620,N_9626,N_8744);
nand U11621 (N_11621,N_8781,N_8300);
nand U11622 (N_11622,N_9884,N_9414);
nor U11623 (N_11623,N_7595,N_7601);
nor U11624 (N_11624,N_8122,N_8283);
nor U11625 (N_11625,N_9968,N_8670);
and U11626 (N_11626,N_9014,N_7684);
xor U11627 (N_11627,N_9515,N_9527);
xor U11628 (N_11628,N_9776,N_9827);
xnor U11629 (N_11629,N_7649,N_8808);
nor U11630 (N_11630,N_9364,N_8996);
or U11631 (N_11631,N_9505,N_9328);
nor U11632 (N_11632,N_7905,N_7801);
nand U11633 (N_11633,N_8022,N_9928);
nor U11634 (N_11634,N_8033,N_9142);
or U11635 (N_11635,N_8485,N_8812);
nor U11636 (N_11636,N_8774,N_9220);
and U11637 (N_11637,N_8448,N_8405);
xnor U11638 (N_11638,N_8990,N_9605);
xor U11639 (N_11639,N_9638,N_7590);
and U11640 (N_11640,N_8926,N_8281);
nor U11641 (N_11641,N_7524,N_9669);
xnor U11642 (N_11642,N_9618,N_7693);
xnor U11643 (N_11643,N_7568,N_8189);
or U11644 (N_11644,N_8646,N_9107);
xor U11645 (N_11645,N_9599,N_8773);
and U11646 (N_11646,N_8742,N_8232);
or U11647 (N_11647,N_8514,N_7555);
xnor U11648 (N_11648,N_7883,N_7640);
nor U11649 (N_11649,N_9846,N_9039);
or U11650 (N_11650,N_9070,N_8291);
nand U11651 (N_11651,N_9311,N_7748);
and U11652 (N_11652,N_7979,N_8096);
nor U11653 (N_11653,N_9070,N_9036);
or U11654 (N_11654,N_8856,N_9055);
xor U11655 (N_11655,N_8933,N_8388);
or U11656 (N_11656,N_8290,N_8450);
nor U11657 (N_11657,N_9475,N_7996);
or U11658 (N_11658,N_8279,N_8244);
and U11659 (N_11659,N_8933,N_9803);
nand U11660 (N_11660,N_9580,N_8840);
nor U11661 (N_11661,N_9339,N_9568);
nor U11662 (N_11662,N_8547,N_7760);
or U11663 (N_11663,N_7650,N_7734);
nand U11664 (N_11664,N_9134,N_8277);
and U11665 (N_11665,N_8097,N_9977);
and U11666 (N_11666,N_8303,N_7541);
nand U11667 (N_11667,N_8841,N_9774);
or U11668 (N_11668,N_8624,N_9293);
nand U11669 (N_11669,N_8898,N_8389);
or U11670 (N_11670,N_8202,N_9489);
nor U11671 (N_11671,N_7996,N_9740);
nor U11672 (N_11672,N_9816,N_9524);
or U11673 (N_11673,N_8062,N_9531);
nand U11674 (N_11674,N_9110,N_8850);
or U11675 (N_11675,N_9816,N_9527);
nand U11676 (N_11676,N_7785,N_8827);
nor U11677 (N_11677,N_9691,N_9096);
or U11678 (N_11678,N_9753,N_8728);
nor U11679 (N_11679,N_8039,N_9574);
nor U11680 (N_11680,N_7924,N_8711);
nand U11681 (N_11681,N_9587,N_9325);
nor U11682 (N_11682,N_9379,N_7670);
xnor U11683 (N_11683,N_7958,N_9281);
or U11684 (N_11684,N_8912,N_8177);
nand U11685 (N_11685,N_8423,N_9854);
xnor U11686 (N_11686,N_7585,N_9321);
xor U11687 (N_11687,N_8095,N_8538);
nand U11688 (N_11688,N_9007,N_8752);
nand U11689 (N_11689,N_8080,N_7719);
nand U11690 (N_11690,N_8843,N_7952);
nor U11691 (N_11691,N_7928,N_9031);
or U11692 (N_11692,N_9618,N_9488);
nand U11693 (N_11693,N_7512,N_9682);
nor U11694 (N_11694,N_8331,N_8724);
and U11695 (N_11695,N_9024,N_7994);
nor U11696 (N_11696,N_7552,N_7716);
nand U11697 (N_11697,N_9256,N_9193);
nand U11698 (N_11698,N_7517,N_9090);
and U11699 (N_11699,N_9126,N_7716);
nor U11700 (N_11700,N_9103,N_8742);
and U11701 (N_11701,N_7598,N_8426);
and U11702 (N_11702,N_8516,N_8256);
xnor U11703 (N_11703,N_7512,N_9159);
or U11704 (N_11704,N_9636,N_9884);
and U11705 (N_11705,N_9713,N_9586);
nor U11706 (N_11706,N_9057,N_7601);
or U11707 (N_11707,N_9943,N_8081);
nand U11708 (N_11708,N_8883,N_9899);
nand U11709 (N_11709,N_9685,N_9322);
nor U11710 (N_11710,N_8560,N_9100);
xor U11711 (N_11711,N_9979,N_9676);
or U11712 (N_11712,N_9792,N_7586);
and U11713 (N_11713,N_8600,N_7641);
and U11714 (N_11714,N_8672,N_8063);
nor U11715 (N_11715,N_7922,N_9723);
and U11716 (N_11716,N_8318,N_9244);
or U11717 (N_11717,N_7541,N_8530);
nand U11718 (N_11718,N_9377,N_8217);
and U11719 (N_11719,N_8560,N_7943);
or U11720 (N_11720,N_8572,N_8979);
nor U11721 (N_11721,N_7692,N_7509);
xnor U11722 (N_11722,N_9290,N_8331);
and U11723 (N_11723,N_8562,N_8345);
and U11724 (N_11724,N_9412,N_9856);
xnor U11725 (N_11725,N_7895,N_8419);
xnor U11726 (N_11726,N_8732,N_9477);
xor U11727 (N_11727,N_7530,N_9651);
and U11728 (N_11728,N_8432,N_8053);
nor U11729 (N_11729,N_9970,N_8015);
xnor U11730 (N_11730,N_8340,N_9073);
and U11731 (N_11731,N_7600,N_8994);
xor U11732 (N_11732,N_9393,N_8128);
or U11733 (N_11733,N_8083,N_8928);
and U11734 (N_11734,N_8868,N_9095);
and U11735 (N_11735,N_8910,N_8496);
nand U11736 (N_11736,N_8744,N_9926);
or U11737 (N_11737,N_8495,N_7799);
and U11738 (N_11738,N_8404,N_7990);
or U11739 (N_11739,N_8749,N_9005);
xnor U11740 (N_11740,N_8184,N_8684);
xor U11741 (N_11741,N_8874,N_9176);
xnor U11742 (N_11742,N_8754,N_9907);
and U11743 (N_11743,N_8494,N_8591);
nand U11744 (N_11744,N_8410,N_7789);
xnor U11745 (N_11745,N_9530,N_7821);
nand U11746 (N_11746,N_7966,N_9856);
xor U11747 (N_11747,N_9485,N_9058);
xor U11748 (N_11748,N_7578,N_7819);
and U11749 (N_11749,N_8160,N_9115);
or U11750 (N_11750,N_9308,N_9643);
and U11751 (N_11751,N_9979,N_8431);
nor U11752 (N_11752,N_8393,N_7890);
xor U11753 (N_11753,N_7516,N_8500);
and U11754 (N_11754,N_8478,N_8686);
or U11755 (N_11755,N_7742,N_8375);
and U11756 (N_11756,N_9636,N_9158);
and U11757 (N_11757,N_8209,N_8428);
nor U11758 (N_11758,N_7525,N_8959);
and U11759 (N_11759,N_8756,N_9379);
nand U11760 (N_11760,N_9523,N_7986);
xor U11761 (N_11761,N_7745,N_8204);
nand U11762 (N_11762,N_9404,N_7670);
nor U11763 (N_11763,N_8712,N_7574);
and U11764 (N_11764,N_7945,N_8672);
or U11765 (N_11765,N_9982,N_9516);
or U11766 (N_11766,N_9844,N_9920);
xor U11767 (N_11767,N_9465,N_9661);
nor U11768 (N_11768,N_7658,N_9933);
nand U11769 (N_11769,N_7575,N_9690);
xnor U11770 (N_11770,N_8199,N_7614);
and U11771 (N_11771,N_9595,N_9677);
or U11772 (N_11772,N_7923,N_9531);
xnor U11773 (N_11773,N_9104,N_7540);
or U11774 (N_11774,N_7581,N_9178);
nor U11775 (N_11775,N_9188,N_8851);
or U11776 (N_11776,N_7549,N_7890);
and U11777 (N_11777,N_8322,N_9994);
nand U11778 (N_11778,N_8414,N_8196);
nor U11779 (N_11779,N_7664,N_8262);
and U11780 (N_11780,N_8436,N_7669);
or U11781 (N_11781,N_8198,N_9611);
nand U11782 (N_11782,N_8151,N_8536);
or U11783 (N_11783,N_8900,N_7641);
or U11784 (N_11784,N_9419,N_9885);
and U11785 (N_11785,N_7561,N_7519);
or U11786 (N_11786,N_9976,N_8523);
or U11787 (N_11787,N_8354,N_9972);
or U11788 (N_11788,N_9528,N_7693);
nand U11789 (N_11789,N_9707,N_8702);
and U11790 (N_11790,N_7627,N_7658);
xnor U11791 (N_11791,N_7609,N_9231);
or U11792 (N_11792,N_8021,N_9853);
nor U11793 (N_11793,N_8182,N_9561);
nand U11794 (N_11794,N_8771,N_7930);
and U11795 (N_11795,N_7807,N_7721);
nand U11796 (N_11796,N_8889,N_9996);
nor U11797 (N_11797,N_8781,N_9185);
or U11798 (N_11798,N_8073,N_7602);
xnor U11799 (N_11799,N_9993,N_9275);
and U11800 (N_11800,N_7551,N_8034);
nor U11801 (N_11801,N_8247,N_8762);
nor U11802 (N_11802,N_7519,N_9570);
nand U11803 (N_11803,N_9627,N_9797);
nand U11804 (N_11804,N_9733,N_9824);
nor U11805 (N_11805,N_7637,N_9351);
or U11806 (N_11806,N_8025,N_9754);
nand U11807 (N_11807,N_8677,N_7756);
xnor U11808 (N_11808,N_9143,N_7824);
or U11809 (N_11809,N_9009,N_8021);
nand U11810 (N_11810,N_9111,N_7605);
xor U11811 (N_11811,N_8469,N_9764);
nor U11812 (N_11812,N_9146,N_9038);
or U11813 (N_11813,N_8487,N_9003);
or U11814 (N_11814,N_8360,N_8636);
nor U11815 (N_11815,N_9589,N_9666);
xnor U11816 (N_11816,N_9018,N_7625);
or U11817 (N_11817,N_8006,N_7738);
nor U11818 (N_11818,N_7858,N_9588);
or U11819 (N_11819,N_9628,N_8614);
xor U11820 (N_11820,N_8620,N_9802);
and U11821 (N_11821,N_9065,N_7858);
and U11822 (N_11822,N_9967,N_8941);
nand U11823 (N_11823,N_9140,N_7980);
nand U11824 (N_11824,N_8148,N_8900);
or U11825 (N_11825,N_7501,N_8738);
xor U11826 (N_11826,N_8077,N_9437);
and U11827 (N_11827,N_9449,N_9073);
nor U11828 (N_11828,N_8469,N_9069);
or U11829 (N_11829,N_7943,N_8572);
xor U11830 (N_11830,N_9224,N_9822);
nor U11831 (N_11831,N_9995,N_9873);
or U11832 (N_11832,N_8574,N_9931);
or U11833 (N_11833,N_8328,N_9304);
xor U11834 (N_11834,N_8312,N_9685);
nor U11835 (N_11835,N_9471,N_9519);
or U11836 (N_11836,N_9750,N_9330);
xnor U11837 (N_11837,N_7741,N_8020);
and U11838 (N_11838,N_9136,N_7717);
nand U11839 (N_11839,N_7616,N_8429);
or U11840 (N_11840,N_9367,N_9441);
nor U11841 (N_11841,N_7755,N_9152);
nand U11842 (N_11842,N_7680,N_8994);
or U11843 (N_11843,N_8933,N_8493);
xnor U11844 (N_11844,N_8022,N_7935);
xor U11845 (N_11845,N_9719,N_8995);
and U11846 (N_11846,N_9929,N_8092);
and U11847 (N_11847,N_8479,N_8333);
nand U11848 (N_11848,N_8411,N_8829);
nor U11849 (N_11849,N_8847,N_9443);
xor U11850 (N_11850,N_9208,N_8731);
and U11851 (N_11851,N_8165,N_9389);
xnor U11852 (N_11852,N_7594,N_8907);
nor U11853 (N_11853,N_9318,N_8186);
nor U11854 (N_11854,N_7615,N_7925);
nor U11855 (N_11855,N_8232,N_9174);
or U11856 (N_11856,N_9452,N_8654);
or U11857 (N_11857,N_9242,N_8148);
nand U11858 (N_11858,N_9596,N_8890);
nand U11859 (N_11859,N_8679,N_8116);
or U11860 (N_11860,N_8088,N_8765);
nand U11861 (N_11861,N_9490,N_7638);
nand U11862 (N_11862,N_7680,N_8026);
nor U11863 (N_11863,N_8052,N_9687);
nand U11864 (N_11864,N_7726,N_8526);
and U11865 (N_11865,N_9997,N_8380);
nor U11866 (N_11866,N_8289,N_7827);
xor U11867 (N_11867,N_9096,N_9045);
nor U11868 (N_11868,N_7507,N_8635);
nand U11869 (N_11869,N_8951,N_8440);
or U11870 (N_11870,N_8155,N_9100);
xor U11871 (N_11871,N_7978,N_9938);
or U11872 (N_11872,N_8626,N_9244);
xor U11873 (N_11873,N_9003,N_8981);
and U11874 (N_11874,N_9160,N_8121);
or U11875 (N_11875,N_9675,N_8440);
or U11876 (N_11876,N_8823,N_7944);
nand U11877 (N_11877,N_8608,N_9390);
nor U11878 (N_11878,N_8842,N_8243);
or U11879 (N_11879,N_7705,N_7979);
or U11880 (N_11880,N_9074,N_7761);
and U11881 (N_11881,N_8116,N_7522);
xor U11882 (N_11882,N_8344,N_8637);
nand U11883 (N_11883,N_8133,N_7620);
or U11884 (N_11884,N_7567,N_8610);
and U11885 (N_11885,N_9196,N_9771);
and U11886 (N_11886,N_9220,N_8298);
nor U11887 (N_11887,N_7745,N_7613);
nand U11888 (N_11888,N_7698,N_9458);
nand U11889 (N_11889,N_9807,N_8477);
xor U11890 (N_11890,N_9489,N_8793);
nand U11891 (N_11891,N_7512,N_8428);
and U11892 (N_11892,N_8999,N_8080);
and U11893 (N_11893,N_9964,N_8618);
xnor U11894 (N_11894,N_7966,N_8319);
or U11895 (N_11895,N_7664,N_7527);
and U11896 (N_11896,N_8252,N_8210);
nor U11897 (N_11897,N_8770,N_9979);
nor U11898 (N_11898,N_7847,N_9493);
and U11899 (N_11899,N_9215,N_9084);
nor U11900 (N_11900,N_7541,N_9136);
nand U11901 (N_11901,N_8041,N_8871);
and U11902 (N_11902,N_9391,N_9956);
nor U11903 (N_11903,N_9751,N_9068);
or U11904 (N_11904,N_8840,N_9259);
nand U11905 (N_11905,N_9496,N_8692);
and U11906 (N_11906,N_7534,N_9585);
nand U11907 (N_11907,N_9476,N_7953);
or U11908 (N_11908,N_8809,N_9249);
or U11909 (N_11909,N_8810,N_9933);
nor U11910 (N_11910,N_9952,N_8279);
xor U11911 (N_11911,N_9749,N_8866);
and U11912 (N_11912,N_9831,N_8691);
xor U11913 (N_11913,N_9584,N_8412);
or U11914 (N_11914,N_9073,N_9203);
or U11915 (N_11915,N_8875,N_8616);
or U11916 (N_11916,N_9398,N_8229);
or U11917 (N_11917,N_9978,N_9715);
nand U11918 (N_11918,N_9160,N_9452);
and U11919 (N_11919,N_7760,N_7522);
and U11920 (N_11920,N_7841,N_8422);
or U11921 (N_11921,N_9221,N_9347);
and U11922 (N_11922,N_9423,N_8229);
and U11923 (N_11923,N_8221,N_9063);
nor U11924 (N_11924,N_8232,N_8225);
xnor U11925 (N_11925,N_8323,N_9873);
or U11926 (N_11926,N_8808,N_9285);
nor U11927 (N_11927,N_9186,N_8820);
and U11928 (N_11928,N_8491,N_9763);
and U11929 (N_11929,N_8726,N_9523);
or U11930 (N_11930,N_8667,N_8313);
nand U11931 (N_11931,N_7503,N_9390);
nor U11932 (N_11932,N_7510,N_8130);
xor U11933 (N_11933,N_7819,N_8517);
nor U11934 (N_11934,N_7666,N_7710);
and U11935 (N_11935,N_9893,N_7837);
and U11936 (N_11936,N_7980,N_7916);
and U11937 (N_11937,N_8833,N_9907);
nor U11938 (N_11938,N_8195,N_7674);
nand U11939 (N_11939,N_9201,N_8635);
and U11940 (N_11940,N_8579,N_8924);
or U11941 (N_11941,N_9501,N_7910);
xor U11942 (N_11942,N_9529,N_8535);
xnor U11943 (N_11943,N_9643,N_8438);
nand U11944 (N_11944,N_8772,N_8233);
nor U11945 (N_11945,N_7583,N_9698);
xnor U11946 (N_11946,N_8710,N_7755);
nand U11947 (N_11947,N_8240,N_8269);
or U11948 (N_11948,N_8998,N_9504);
or U11949 (N_11949,N_9640,N_7941);
nand U11950 (N_11950,N_8716,N_7931);
or U11951 (N_11951,N_8352,N_8050);
nand U11952 (N_11952,N_7540,N_8186);
xnor U11953 (N_11953,N_8709,N_7661);
and U11954 (N_11954,N_9791,N_8334);
nor U11955 (N_11955,N_9216,N_8553);
nor U11956 (N_11956,N_9788,N_7867);
xor U11957 (N_11957,N_9008,N_8325);
and U11958 (N_11958,N_8787,N_8769);
xor U11959 (N_11959,N_9072,N_9867);
xor U11960 (N_11960,N_9162,N_9580);
and U11961 (N_11961,N_9372,N_8739);
nor U11962 (N_11962,N_8163,N_8570);
xor U11963 (N_11963,N_9523,N_7623);
and U11964 (N_11964,N_9134,N_8485);
nand U11965 (N_11965,N_7773,N_8172);
nor U11966 (N_11966,N_7545,N_9501);
and U11967 (N_11967,N_9996,N_8152);
nor U11968 (N_11968,N_8628,N_8553);
xnor U11969 (N_11969,N_9055,N_7742);
nand U11970 (N_11970,N_7546,N_9587);
xnor U11971 (N_11971,N_9111,N_9188);
xnor U11972 (N_11972,N_7618,N_7541);
xnor U11973 (N_11973,N_9637,N_7581);
nand U11974 (N_11974,N_9090,N_9693);
xnor U11975 (N_11975,N_9464,N_9076);
and U11976 (N_11976,N_8941,N_7738);
and U11977 (N_11977,N_9823,N_8760);
nand U11978 (N_11978,N_8670,N_7864);
and U11979 (N_11979,N_8243,N_9078);
nand U11980 (N_11980,N_8650,N_8519);
and U11981 (N_11981,N_8999,N_9209);
xor U11982 (N_11982,N_7570,N_9648);
or U11983 (N_11983,N_7828,N_7820);
and U11984 (N_11984,N_8732,N_9134);
or U11985 (N_11985,N_7546,N_7648);
or U11986 (N_11986,N_8725,N_9618);
nor U11987 (N_11987,N_7726,N_9558);
xnor U11988 (N_11988,N_9023,N_9127);
nor U11989 (N_11989,N_7687,N_9062);
nand U11990 (N_11990,N_7999,N_7781);
or U11991 (N_11991,N_8423,N_9435);
and U11992 (N_11992,N_7607,N_8883);
nand U11993 (N_11993,N_8998,N_7828);
nor U11994 (N_11994,N_8988,N_8668);
or U11995 (N_11995,N_9346,N_8772);
or U11996 (N_11996,N_9469,N_9082);
and U11997 (N_11997,N_8757,N_8134);
and U11998 (N_11998,N_8586,N_7766);
and U11999 (N_11999,N_7551,N_8371);
nand U12000 (N_12000,N_9508,N_8647);
and U12001 (N_12001,N_9756,N_9659);
nor U12002 (N_12002,N_8613,N_9860);
or U12003 (N_12003,N_8081,N_9843);
xnor U12004 (N_12004,N_8835,N_9769);
or U12005 (N_12005,N_7617,N_8779);
nand U12006 (N_12006,N_8309,N_8178);
and U12007 (N_12007,N_9694,N_9016);
and U12008 (N_12008,N_8199,N_8092);
nand U12009 (N_12009,N_8184,N_8647);
or U12010 (N_12010,N_7617,N_7698);
or U12011 (N_12011,N_9083,N_9103);
nor U12012 (N_12012,N_9240,N_8958);
xnor U12013 (N_12013,N_9603,N_7740);
or U12014 (N_12014,N_8214,N_8061);
or U12015 (N_12015,N_8518,N_9851);
or U12016 (N_12016,N_7508,N_9996);
nor U12017 (N_12017,N_7720,N_8060);
xor U12018 (N_12018,N_9547,N_8199);
xor U12019 (N_12019,N_8674,N_9448);
and U12020 (N_12020,N_8762,N_8700);
and U12021 (N_12021,N_8531,N_8139);
xnor U12022 (N_12022,N_7772,N_9756);
and U12023 (N_12023,N_8675,N_9585);
or U12024 (N_12024,N_8212,N_8691);
xor U12025 (N_12025,N_8369,N_9414);
nand U12026 (N_12026,N_8824,N_7824);
or U12027 (N_12027,N_9404,N_9760);
nor U12028 (N_12028,N_7661,N_9658);
nand U12029 (N_12029,N_9951,N_8155);
or U12030 (N_12030,N_8451,N_9962);
nand U12031 (N_12031,N_9390,N_9555);
or U12032 (N_12032,N_7924,N_9733);
nand U12033 (N_12033,N_7757,N_9560);
xor U12034 (N_12034,N_8888,N_8366);
xnor U12035 (N_12035,N_9202,N_8974);
xor U12036 (N_12036,N_7925,N_8546);
nor U12037 (N_12037,N_9438,N_9398);
and U12038 (N_12038,N_9050,N_9191);
xor U12039 (N_12039,N_7838,N_7707);
nand U12040 (N_12040,N_9100,N_9442);
or U12041 (N_12041,N_7876,N_8950);
nand U12042 (N_12042,N_9332,N_7979);
and U12043 (N_12043,N_7821,N_9827);
nand U12044 (N_12044,N_9753,N_7934);
xor U12045 (N_12045,N_8745,N_7529);
nand U12046 (N_12046,N_9764,N_8694);
or U12047 (N_12047,N_9444,N_9794);
nand U12048 (N_12048,N_7907,N_7715);
nor U12049 (N_12049,N_8819,N_8357);
nand U12050 (N_12050,N_8948,N_9509);
nand U12051 (N_12051,N_8275,N_8767);
and U12052 (N_12052,N_8080,N_7592);
nand U12053 (N_12053,N_8823,N_9782);
or U12054 (N_12054,N_8061,N_9901);
xnor U12055 (N_12055,N_7952,N_9187);
or U12056 (N_12056,N_8289,N_8414);
or U12057 (N_12057,N_8803,N_7617);
and U12058 (N_12058,N_8207,N_9955);
or U12059 (N_12059,N_7679,N_9377);
or U12060 (N_12060,N_8925,N_9807);
nand U12061 (N_12061,N_9056,N_8453);
or U12062 (N_12062,N_9640,N_9546);
nor U12063 (N_12063,N_9780,N_7574);
nor U12064 (N_12064,N_8150,N_8056);
xnor U12065 (N_12065,N_8433,N_9328);
and U12066 (N_12066,N_9293,N_8765);
nor U12067 (N_12067,N_9713,N_7897);
and U12068 (N_12068,N_8246,N_7949);
nor U12069 (N_12069,N_8306,N_9710);
xnor U12070 (N_12070,N_8263,N_9007);
nor U12071 (N_12071,N_7549,N_8776);
or U12072 (N_12072,N_8807,N_7824);
and U12073 (N_12073,N_8573,N_8597);
and U12074 (N_12074,N_9878,N_9880);
or U12075 (N_12075,N_9058,N_7810);
or U12076 (N_12076,N_9588,N_9160);
xnor U12077 (N_12077,N_9970,N_8510);
xor U12078 (N_12078,N_9455,N_9217);
xor U12079 (N_12079,N_9198,N_7566);
nand U12080 (N_12080,N_8335,N_9068);
and U12081 (N_12081,N_9910,N_8368);
or U12082 (N_12082,N_7526,N_7690);
xnor U12083 (N_12083,N_9880,N_7982);
nor U12084 (N_12084,N_8418,N_8743);
and U12085 (N_12085,N_7963,N_8658);
or U12086 (N_12086,N_9965,N_9681);
or U12087 (N_12087,N_8677,N_8054);
and U12088 (N_12088,N_8526,N_7621);
nand U12089 (N_12089,N_8583,N_8534);
nand U12090 (N_12090,N_8280,N_8930);
or U12091 (N_12091,N_9701,N_8249);
nor U12092 (N_12092,N_8587,N_8035);
or U12093 (N_12093,N_8216,N_8461);
and U12094 (N_12094,N_7690,N_9816);
or U12095 (N_12095,N_8344,N_8584);
and U12096 (N_12096,N_8037,N_9336);
xnor U12097 (N_12097,N_9848,N_8834);
nand U12098 (N_12098,N_9321,N_8204);
or U12099 (N_12099,N_9048,N_8329);
xor U12100 (N_12100,N_8572,N_7788);
nand U12101 (N_12101,N_7732,N_8633);
nand U12102 (N_12102,N_7651,N_9069);
nand U12103 (N_12103,N_9257,N_9598);
xor U12104 (N_12104,N_7900,N_9674);
nor U12105 (N_12105,N_7965,N_7896);
xor U12106 (N_12106,N_8485,N_9264);
or U12107 (N_12107,N_9442,N_8422);
xor U12108 (N_12108,N_8636,N_9034);
nor U12109 (N_12109,N_9791,N_8223);
or U12110 (N_12110,N_8018,N_7560);
nor U12111 (N_12111,N_9093,N_8432);
nor U12112 (N_12112,N_9203,N_8598);
or U12113 (N_12113,N_7706,N_9905);
nor U12114 (N_12114,N_7682,N_9926);
or U12115 (N_12115,N_9838,N_9890);
xnor U12116 (N_12116,N_9820,N_8024);
and U12117 (N_12117,N_8848,N_8301);
nor U12118 (N_12118,N_9642,N_7681);
nor U12119 (N_12119,N_9841,N_8507);
xor U12120 (N_12120,N_8015,N_8500);
nor U12121 (N_12121,N_8973,N_7565);
and U12122 (N_12122,N_9884,N_8554);
xnor U12123 (N_12123,N_9505,N_8820);
and U12124 (N_12124,N_7515,N_9524);
xnor U12125 (N_12125,N_8539,N_9610);
nor U12126 (N_12126,N_9643,N_9317);
xor U12127 (N_12127,N_8104,N_7775);
and U12128 (N_12128,N_9782,N_8839);
xor U12129 (N_12129,N_7532,N_9480);
nand U12130 (N_12130,N_9678,N_8625);
or U12131 (N_12131,N_9101,N_7874);
xnor U12132 (N_12132,N_8340,N_9750);
or U12133 (N_12133,N_8658,N_8741);
xor U12134 (N_12134,N_9529,N_8523);
or U12135 (N_12135,N_8548,N_9661);
or U12136 (N_12136,N_8995,N_7897);
xor U12137 (N_12137,N_8145,N_7907);
nor U12138 (N_12138,N_9594,N_9775);
or U12139 (N_12139,N_9092,N_9025);
nor U12140 (N_12140,N_9518,N_8031);
and U12141 (N_12141,N_9140,N_9872);
and U12142 (N_12142,N_7676,N_9797);
and U12143 (N_12143,N_8837,N_9637);
nand U12144 (N_12144,N_9160,N_7512);
nor U12145 (N_12145,N_7946,N_7673);
and U12146 (N_12146,N_8578,N_8695);
xnor U12147 (N_12147,N_9026,N_7703);
and U12148 (N_12148,N_8533,N_9051);
xnor U12149 (N_12149,N_8041,N_9444);
nor U12150 (N_12150,N_7693,N_9933);
and U12151 (N_12151,N_9649,N_8509);
nand U12152 (N_12152,N_8273,N_8724);
xor U12153 (N_12153,N_9192,N_9901);
nand U12154 (N_12154,N_9473,N_9635);
xnor U12155 (N_12155,N_8117,N_8726);
or U12156 (N_12156,N_7515,N_8864);
nand U12157 (N_12157,N_9968,N_9022);
or U12158 (N_12158,N_8101,N_8145);
nand U12159 (N_12159,N_8264,N_8806);
nand U12160 (N_12160,N_7684,N_7814);
and U12161 (N_12161,N_9821,N_8826);
or U12162 (N_12162,N_9474,N_9473);
xor U12163 (N_12163,N_8162,N_9087);
nand U12164 (N_12164,N_9186,N_9884);
and U12165 (N_12165,N_8085,N_8478);
xnor U12166 (N_12166,N_8603,N_8659);
and U12167 (N_12167,N_9328,N_8575);
nand U12168 (N_12168,N_8089,N_9984);
nand U12169 (N_12169,N_8618,N_8337);
nand U12170 (N_12170,N_8850,N_8436);
or U12171 (N_12171,N_8971,N_9435);
or U12172 (N_12172,N_8872,N_9027);
and U12173 (N_12173,N_9191,N_8169);
nor U12174 (N_12174,N_9469,N_8649);
or U12175 (N_12175,N_9195,N_7919);
nor U12176 (N_12176,N_9354,N_9083);
xor U12177 (N_12177,N_8846,N_7778);
or U12178 (N_12178,N_8600,N_9850);
nor U12179 (N_12179,N_7633,N_9243);
or U12180 (N_12180,N_9060,N_7524);
and U12181 (N_12181,N_8128,N_9175);
nand U12182 (N_12182,N_9031,N_8831);
nand U12183 (N_12183,N_8876,N_7955);
nor U12184 (N_12184,N_8777,N_8672);
or U12185 (N_12185,N_7832,N_8359);
and U12186 (N_12186,N_9556,N_8003);
nor U12187 (N_12187,N_9969,N_8173);
nand U12188 (N_12188,N_7724,N_9645);
nor U12189 (N_12189,N_8584,N_7991);
or U12190 (N_12190,N_8838,N_9540);
or U12191 (N_12191,N_9999,N_8425);
nor U12192 (N_12192,N_9723,N_8214);
nor U12193 (N_12193,N_9375,N_8653);
nor U12194 (N_12194,N_8318,N_9141);
and U12195 (N_12195,N_9340,N_9616);
nor U12196 (N_12196,N_9213,N_9145);
or U12197 (N_12197,N_9530,N_9337);
xor U12198 (N_12198,N_9727,N_7863);
and U12199 (N_12199,N_8954,N_7889);
or U12200 (N_12200,N_8826,N_7806);
or U12201 (N_12201,N_9656,N_7813);
nand U12202 (N_12202,N_9205,N_8812);
nand U12203 (N_12203,N_8789,N_8644);
nand U12204 (N_12204,N_9368,N_9500);
nor U12205 (N_12205,N_9672,N_8245);
or U12206 (N_12206,N_8005,N_7622);
nor U12207 (N_12207,N_8730,N_8465);
nand U12208 (N_12208,N_8005,N_9755);
xor U12209 (N_12209,N_7722,N_9725);
nor U12210 (N_12210,N_8190,N_7590);
nor U12211 (N_12211,N_9057,N_9683);
nor U12212 (N_12212,N_8352,N_8524);
nor U12213 (N_12213,N_7921,N_9673);
or U12214 (N_12214,N_9408,N_9558);
nor U12215 (N_12215,N_8620,N_8348);
nand U12216 (N_12216,N_9266,N_8550);
nand U12217 (N_12217,N_8794,N_8643);
and U12218 (N_12218,N_8345,N_9967);
and U12219 (N_12219,N_9051,N_9967);
and U12220 (N_12220,N_9573,N_9601);
xnor U12221 (N_12221,N_9461,N_9029);
or U12222 (N_12222,N_7590,N_8560);
nand U12223 (N_12223,N_8595,N_9133);
nand U12224 (N_12224,N_8785,N_8585);
and U12225 (N_12225,N_8133,N_7911);
nor U12226 (N_12226,N_7986,N_7502);
xnor U12227 (N_12227,N_8716,N_8125);
nor U12228 (N_12228,N_7814,N_8821);
xnor U12229 (N_12229,N_8469,N_8361);
and U12230 (N_12230,N_9998,N_9258);
nor U12231 (N_12231,N_9726,N_8305);
and U12232 (N_12232,N_8070,N_9530);
nor U12233 (N_12233,N_9807,N_7537);
nand U12234 (N_12234,N_8676,N_8766);
nor U12235 (N_12235,N_9535,N_9174);
and U12236 (N_12236,N_9792,N_7953);
nor U12237 (N_12237,N_8069,N_8984);
nand U12238 (N_12238,N_7873,N_7851);
and U12239 (N_12239,N_9997,N_8071);
and U12240 (N_12240,N_9924,N_9668);
xnor U12241 (N_12241,N_9295,N_9289);
and U12242 (N_12242,N_8806,N_8122);
xor U12243 (N_12243,N_7737,N_9578);
nand U12244 (N_12244,N_9022,N_7768);
and U12245 (N_12245,N_8294,N_8884);
or U12246 (N_12246,N_9322,N_9084);
nand U12247 (N_12247,N_7694,N_8236);
and U12248 (N_12248,N_9815,N_9376);
nor U12249 (N_12249,N_8834,N_9638);
or U12250 (N_12250,N_7534,N_9986);
xnor U12251 (N_12251,N_9816,N_8257);
or U12252 (N_12252,N_9815,N_9620);
and U12253 (N_12253,N_7926,N_8779);
or U12254 (N_12254,N_8709,N_7618);
nand U12255 (N_12255,N_8501,N_9899);
or U12256 (N_12256,N_9558,N_8181);
xnor U12257 (N_12257,N_9424,N_8324);
xnor U12258 (N_12258,N_7709,N_7614);
nand U12259 (N_12259,N_7731,N_7633);
nor U12260 (N_12260,N_9175,N_9331);
or U12261 (N_12261,N_9763,N_8029);
or U12262 (N_12262,N_8192,N_8660);
xor U12263 (N_12263,N_8547,N_8501);
xor U12264 (N_12264,N_9529,N_9677);
nand U12265 (N_12265,N_8510,N_9069);
and U12266 (N_12266,N_7971,N_9354);
xor U12267 (N_12267,N_9242,N_9128);
nor U12268 (N_12268,N_9916,N_9862);
nor U12269 (N_12269,N_7754,N_8847);
nand U12270 (N_12270,N_7957,N_8351);
nand U12271 (N_12271,N_8259,N_9963);
or U12272 (N_12272,N_8035,N_7960);
nor U12273 (N_12273,N_8960,N_9885);
or U12274 (N_12274,N_8082,N_8097);
nor U12275 (N_12275,N_8913,N_9617);
xnor U12276 (N_12276,N_8524,N_9794);
nor U12277 (N_12277,N_7835,N_9580);
and U12278 (N_12278,N_9922,N_8849);
nor U12279 (N_12279,N_8556,N_8526);
xnor U12280 (N_12280,N_9893,N_8296);
xor U12281 (N_12281,N_8923,N_8490);
nor U12282 (N_12282,N_8790,N_8864);
nand U12283 (N_12283,N_8983,N_8854);
nor U12284 (N_12284,N_8384,N_9852);
or U12285 (N_12285,N_7931,N_7820);
and U12286 (N_12286,N_9573,N_7760);
xnor U12287 (N_12287,N_9849,N_9543);
or U12288 (N_12288,N_9801,N_8137);
nor U12289 (N_12289,N_8147,N_8154);
xor U12290 (N_12290,N_8611,N_8928);
xor U12291 (N_12291,N_8865,N_8742);
or U12292 (N_12292,N_9588,N_9364);
nand U12293 (N_12293,N_9066,N_9147);
or U12294 (N_12294,N_9952,N_9963);
nand U12295 (N_12295,N_7767,N_7631);
nor U12296 (N_12296,N_8615,N_9250);
nor U12297 (N_12297,N_8504,N_9854);
nor U12298 (N_12298,N_8823,N_8203);
nand U12299 (N_12299,N_9138,N_9346);
nand U12300 (N_12300,N_8241,N_9573);
and U12301 (N_12301,N_9219,N_9026);
or U12302 (N_12302,N_9052,N_9304);
or U12303 (N_12303,N_9331,N_9949);
xor U12304 (N_12304,N_8115,N_9685);
xor U12305 (N_12305,N_9724,N_9875);
xor U12306 (N_12306,N_9060,N_9558);
or U12307 (N_12307,N_8554,N_8095);
or U12308 (N_12308,N_7504,N_7661);
or U12309 (N_12309,N_8891,N_9115);
nor U12310 (N_12310,N_7982,N_9903);
nand U12311 (N_12311,N_9012,N_8588);
nand U12312 (N_12312,N_7522,N_8285);
nor U12313 (N_12313,N_9999,N_9380);
or U12314 (N_12314,N_9560,N_8476);
nor U12315 (N_12315,N_9989,N_8752);
nor U12316 (N_12316,N_8584,N_9218);
and U12317 (N_12317,N_7649,N_9160);
xnor U12318 (N_12318,N_8145,N_8046);
nor U12319 (N_12319,N_8319,N_7594);
nand U12320 (N_12320,N_9293,N_8047);
nor U12321 (N_12321,N_9294,N_8141);
xor U12322 (N_12322,N_8102,N_7726);
and U12323 (N_12323,N_9072,N_9539);
or U12324 (N_12324,N_7750,N_7948);
xor U12325 (N_12325,N_9939,N_8644);
nor U12326 (N_12326,N_8253,N_7977);
nor U12327 (N_12327,N_9033,N_9955);
and U12328 (N_12328,N_8990,N_7513);
nand U12329 (N_12329,N_7690,N_7792);
and U12330 (N_12330,N_9930,N_8999);
nor U12331 (N_12331,N_8415,N_8910);
or U12332 (N_12332,N_9062,N_7716);
nand U12333 (N_12333,N_8603,N_9749);
and U12334 (N_12334,N_9010,N_7659);
and U12335 (N_12335,N_9960,N_7848);
xnor U12336 (N_12336,N_8095,N_7622);
nand U12337 (N_12337,N_8090,N_8143);
or U12338 (N_12338,N_9073,N_9436);
xnor U12339 (N_12339,N_8433,N_9013);
nand U12340 (N_12340,N_9062,N_9598);
and U12341 (N_12341,N_9956,N_8254);
and U12342 (N_12342,N_8359,N_9550);
or U12343 (N_12343,N_8469,N_9915);
or U12344 (N_12344,N_7953,N_9481);
and U12345 (N_12345,N_8087,N_9988);
nand U12346 (N_12346,N_9029,N_7736);
nor U12347 (N_12347,N_8365,N_8110);
nor U12348 (N_12348,N_9123,N_8881);
xnor U12349 (N_12349,N_9876,N_8073);
and U12350 (N_12350,N_7948,N_8313);
xor U12351 (N_12351,N_9476,N_8931);
xnor U12352 (N_12352,N_9020,N_9265);
or U12353 (N_12353,N_9429,N_9603);
nor U12354 (N_12354,N_9745,N_9529);
nand U12355 (N_12355,N_7543,N_8693);
nand U12356 (N_12356,N_9174,N_7595);
xor U12357 (N_12357,N_8904,N_8295);
or U12358 (N_12358,N_9227,N_8253);
or U12359 (N_12359,N_8829,N_7915);
or U12360 (N_12360,N_8945,N_9591);
and U12361 (N_12361,N_7584,N_8925);
nor U12362 (N_12362,N_9437,N_9194);
and U12363 (N_12363,N_9676,N_7541);
nor U12364 (N_12364,N_9845,N_9580);
nand U12365 (N_12365,N_9500,N_7586);
or U12366 (N_12366,N_8023,N_8085);
or U12367 (N_12367,N_9105,N_7666);
or U12368 (N_12368,N_7956,N_8416);
and U12369 (N_12369,N_8655,N_8914);
or U12370 (N_12370,N_8785,N_8712);
nand U12371 (N_12371,N_7899,N_9524);
nand U12372 (N_12372,N_8478,N_8289);
or U12373 (N_12373,N_9956,N_8142);
or U12374 (N_12374,N_8055,N_7516);
nand U12375 (N_12375,N_8377,N_9322);
xnor U12376 (N_12376,N_8185,N_8064);
nor U12377 (N_12377,N_8564,N_7592);
and U12378 (N_12378,N_9608,N_7601);
or U12379 (N_12379,N_8913,N_7965);
nor U12380 (N_12380,N_8148,N_9160);
and U12381 (N_12381,N_9874,N_8316);
xnor U12382 (N_12382,N_7839,N_9209);
and U12383 (N_12383,N_8467,N_9108);
nor U12384 (N_12384,N_9103,N_9670);
and U12385 (N_12385,N_8362,N_8188);
and U12386 (N_12386,N_7681,N_9694);
xnor U12387 (N_12387,N_7648,N_8931);
and U12388 (N_12388,N_8325,N_8499);
nand U12389 (N_12389,N_8849,N_7870);
nor U12390 (N_12390,N_8868,N_9364);
and U12391 (N_12391,N_8399,N_7693);
and U12392 (N_12392,N_9236,N_9587);
and U12393 (N_12393,N_8742,N_9643);
nor U12394 (N_12394,N_9231,N_9053);
xor U12395 (N_12395,N_8767,N_7709);
xor U12396 (N_12396,N_7698,N_7963);
nand U12397 (N_12397,N_9971,N_7637);
nand U12398 (N_12398,N_8112,N_9267);
or U12399 (N_12399,N_7602,N_8742);
nor U12400 (N_12400,N_8335,N_7721);
nand U12401 (N_12401,N_9724,N_9701);
nor U12402 (N_12402,N_9199,N_7535);
and U12403 (N_12403,N_9860,N_8149);
or U12404 (N_12404,N_8958,N_8876);
xnor U12405 (N_12405,N_9507,N_9285);
and U12406 (N_12406,N_7600,N_7792);
and U12407 (N_12407,N_8162,N_8896);
nor U12408 (N_12408,N_8442,N_8480);
xor U12409 (N_12409,N_8013,N_8316);
and U12410 (N_12410,N_9041,N_9147);
and U12411 (N_12411,N_8087,N_8541);
and U12412 (N_12412,N_7592,N_8366);
or U12413 (N_12413,N_9646,N_7878);
and U12414 (N_12414,N_8445,N_8754);
xnor U12415 (N_12415,N_8239,N_9885);
nor U12416 (N_12416,N_8472,N_7729);
and U12417 (N_12417,N_7863,N_7848);
nand U12418 (N_12418,N_7782,N_8974);
and U12419 (N_12419,N_9391,N_8138);
and U12420 (N_12420,N_7974,N_7741);
or U12421 (N_12421,N_8428,N_8004);
or U12422 (N_12422,N_9720,N_9953);
xor U12423 (N_12423,N_7870,N_8191);
and U12424 (N_12424,N_8797,N_8450);
nor U12425 (N_12425,N_8737,N_7744);
and U12426 (N_12426,N_8640,N_7987);
nor U12427 (N_12427,N_7985,N_9024);
or U12428 (N_12428,N_9082,N_7971);
or U12429 (N_12429,N_8278,N_7871);
or U12430 (N_12430,N_8387,N_9272);
nand U12431 (N_12431,N_8891,N_8086);
and U12432 (N_12432,N_9879,N_8733);
nor U12433 (N_12433,N_8975,N_8195);
xor U12434 (N_12434,N_7689,N_8173);
or U12435 (N_12435,N_9580,N_9276);
nor U12436 (N_12436,N_7778,N_8529);
nor U12437 (N_12437,N_7974,N_7641);
xnor U12438 (N_12438,N_9236,N_8729);
nand U12439 (N_12439,N_9410,N_7503);
or U12440 (N_12440,N_9257,N_8351);
or U12441 (N_12441,N_9094,N_7509);
nor U12442 (N_12442,N_7926,N_8642);
or U12443 (N_12443,N_8518,N_9858);
nand U12444 (N_12444,N_8231,N_8227);
and U12445 (N_12445,N_8403,N_7693);
or U12446 (N_12446,N_9035,N_9014);
or U12447 (N_12447,N_8610,N_8059);
nor U12448 (N_12448,N_9307,N_7535);
xnor U12449 (N_12449,N_9175,N_9028);
nor U12450 (N_12450,N_9673,N_9737);
nand U12451 (N_12451,N_9892,N_9024);
nand U12452 (N_12452,N_8468,N_8642);
nor U12453 (N_12453,N_7849,N_8198);
nor U12454 (N_12454,N_8847,N_7710);
nor U12455 (N_12455,N_7677,N_7812);
or U12456 (N_12456,N_7998,N_7636);
or U12457 (N_12457,N_7959,N_9976);
nand U12458 (N_12458,N_9613,N_9345);
or U12459 (N_12459,N_7991,N_9588);
nor U12460 (N_12460,N_9459,N_8630);
nor U12461 (N_12461,N_9944,N_8298);
or U12462 (N_12462,N_9126,N_7535);
nand U12463 (N_12463,N_9288,N_9227);
nor U12464 (N_12464,N_8171,N_9384);
or U12465 (N_12465,N_8103,N_8227);
or U12466 (N_12466,N_8341,N_8296);
nand U12467 (N_12467,N_9874,N_7976);
nor U12468 (N_12468,N_7948,N_7752);
nor U12469 (N_12469,N_8166,N_8899);
nor U12470 (N_12470,N_8379,N_9029);
and U12471 (N_12471,N_8653,N_8691);
xnor U12472 (N_12472,N_9454,N_8497);
nor U12473 (N_12473,N_8456,N_7677);
or U12474 (N_12474,N_8352,N_9679);
nor U12475 (N_12475,N_9269,N_9230);
and U12476 (N_12476,N_9611,N_8567);
nor U12477 (N_12477,N_7932,N_8467);
nor U12478 (N_12478,N_7829,N_9743);
nand U12479 (N_12479,N_9625,N_8779);
and U12480 (N_12480,N_8240,N_9890);
and U12481 (N_12481,N_8396,N_8035);
nand U12482 (N_12482,N_9365,N_8824);
or U12483 (N_12483,N_8119,N_9193);
and U12484 (N_12484,N_9748,N_7628);
nor U12485 (N_12485,N_8986,N_8940);
nand U12486 (N_12486,N_9271,N_8535);
and U12487 (N_12487,N_8934,N_8536);
nand U12488 (N_12488,N_9752,N_9993);
or U12489 (N_12489,N_9611,N_9202);
nor U12490 (N_12490,N_8131,N_8531);
or U12491 (N_12491,N_7556,N_9131);
and U12492 (N_12492,N_9625,N_7522);
nand U12493 (N_12493,N_8815,N_9139);
and U12494 (N_12494,N_8498,N_8934);
nand U12495 (N_12495,N_7748,N_8795);
xor U12496 (N_12496,N_7544,N_8006);
xnor U12497 (N_12497,N_9074,N_8267);
nor U12498 (N_12498,N_9895,N_7800);
xnor U12499 (N_12499,N_9384,N_8397);
and U12500 (N_12500,N_11763,N_11775);
nand U12501 (N_12501,N_10197,N_11268);
nor U12502 (N_12502,N_11559,N_10876);
nor U12503 (N_12503,N_10454,N_11525);
nand U12504 (N_12504,N_12402,N_10935);
or U12505 (N_12505,N_11243,N_10016);
nand U12506 (N_12506,N_11776,N_10635);
nand U12507 (N_12507,N_11847,N_10201);
nor U12508 (N_12508,N_10772,N_11265);
or U12509 (N_12509,N_12266,N_11089);
nor U12510 (N_12510,N_12497,N_10920);
xnor U12511 (N_12511,N_12324,N_11537);
and U12512 (N_12512,N_10571,N_10256);
and U12513 (N_12513,N_11557,N_10470);
and U12514 (N_12514,N_10659,N_10701);
or U12515 (N_12515,N_10729,N_11068);
nor U12516 (N_12516,N_10594,N_11083);
xnor U12517 (N_12517,N_11027,N_10037);
xor U12518 (N_12518,N_10789,N_10123);
nor U12519 (N_12519,N_11182,N_11153);
or U12520 (N_12520,N_10409,N_10181);
nand U12521 (N_12521,N_11056,N_12140);
nand U12522 (N_12522,N_11953,N_10033);
nor U12523 (N_12523,N_11780,N_10687);
nor U12524 (N_12524,N_10620,N_10485);
or U12525 (N_12525,N_11736,N_11959);
and U12526 (N_12526,N_10452,N_10413);
or U12527 (N_12527,N_12086,N_10491);
or U12528 (N_12528,N_11290,N_10686);
xor U12529 (N_12529,N_11261,N_11766);
and U12530 (N_12530,N_11555,N_11839);
and U12531 (N_12531,N_10255,N_10711);
xor U12532 (N_12532,N_12187,N_11721);
or U12533 (N_12533,N_10272,N_11573);
nand U12534 (N_12534,N_10805,N_10154);
or U12535 (N_12535,N_10679,N_10046);
or U12536 (N_12536,N_10088,N_12428);
nand U12537 (N_12537,N_10095,N_11779);
nand U12538 (N_12538,N_10008,N_12348);
and U12539 (N_12539,N_12453,N_11408);
and U12540 (N_12540,N_12117,N_11515);
and U12541 (N_12541,N_10105,N_11693);
or U12542 (N_12542,N_10036,N_11064);
and U12543 (N_12543,N_12470,N_12265);
nand U12544 (N_12544,N_11589,N_11458);
nand U12545 (N_12545,N_10050,N_10195);
nand U12546 (N_12546,N_11772,N_12025);
nor U12547 (N_12547,N_11065,N_11548);
and U12548 (N_12548,N_11575,N_12109);
or U12549 (N_12549,N_12092,N_11394);
nand U12550 (N_12550,N_10278,N_11412);
and U12551 (N_12551,N_10150,N_11560);
or U12552 (N_12552,N_12474,N_12476);
and U12553 (N_12553,N_10192,N_10247);
and U12554 (N_12554,N_11577,N_12085);
nand U12555 (N_12555,N_12492,N_10137);
nor U12556 (N_12556,N_11747,N_12175);
nor U12557 (N_12557,N_11163,N_10652);
nor U12558 (N_12558,N_10482,N_10784);
nor U12559 (N_12559,N_12316,N_10610);
nor U12560 (N_12560,N_10458,N_10641);
xnor U12561 (N_12561,N_10143,N_12421);
xnor U12562 (N_12562,N_12046,N_12131);
and U12563 (N_12563,N_12264,N_11624);
nand U12564 (N_12564,N_10078,N_12256);
nor U12565 (N_12565,N_10827,N_10063);
or U12566 (N_12566,N_11255,N_11278);
and U12567 (N_12567,N_10169,N_11718);
xnor U12568 (N_12568,N_12398,N_10795);
nand U12569 (N_12569,N_11994,N_12242);
nor U12570 (N_12570,N_10138,N_10629);
nand U12571 (N_12571,N_11415,N_10263);
or U12572 (N_12572,N_10324,N_10584);
xor U12573 (N_12573,N_11605,N_11485);
or U12574 (N_12574,N_10486,N_11761);
and U12575 (N_12575,N_12258,N_12125);
or U12576 (N_12576,N_11621,N_12107);
or U12577 (N_12577,N_11285,N_12279);
and U12578 (N_12578,N_11087,N_10356);
and U12579 (N_12579,N_11025,N_10998);
or U12580 (N_12580,N_11383,N_11347);
or U12581 (N_12581,N_10184,N_10307);
nand U12582 (N_12582,N_10999,N_10311);
or U12583 (N_12583,N_10791,N_11364);
nand U12584 (N_12584,N_10733,N_12208);
xnor U12585 (N_12585,N_10100,N_10070);
nand U12586 (N_12586,N_10394,N_11316);
or U12587 (N_12587,N_10222,N_12103);
nand U12588 (N_12588,N_11096,N_12020);
nand U12589 (N_12589,N_12192,N_11220);
nor U12590 (N_12590,N_12004,N_10021);
nor U12591 (N_12591,N_12200,N_11990);
and U12592 (N_12592,N_10799,N_11053);
and U12593 (N_12593,N_11774,N_10187);
xnor U12594 (N_12594,N_11727,N_10212);
nor U12595 (N_12595,N_10749,N_11300);
and U12596 (N_12596,N_11864,N_12496);
xor U12597 (N_12597,N_10329,N_10358);
or U12598 (N_12598,N_11158,N_11622);
xor U12599 (N_12599,N_11791,N_10564);
nor U12600 (N_12600,N_11417,N_12405);
and U12601 (N_12601,N_11162,N_11317);
and U12602 (N_12602,N_11295,N_11030);
nand U12603 (N_12603,N_10650,N_10258);
nor U12604 (N_12604,N_10414,N_10405);
nand U12605 (N_12605,N_11494,N_10821);
or U12606 (N_12606,N_11778,N_11699);
or U12607 (N_12607,N_12159,N_11737);
xor U12608 (N_12608,N_11218,N_11665);
or U12609 (N_12609,N_10605,N_11429);
nand U12610 (N_12610,N_10481,N_10198);
nor U12611 (N_12611,N_11368,N_10883);
or U12612 (N_12612,N_10094,N_10699);
nor U12613 (N_12613,N_10541,N_12024);
nand U12614 (N_12614,N_11873,N_12328);
and U12615 (N_12615,N_11487,N_10320);
or U12616 (N_12616,N_10846,N_10044);
nor U12617 (N_12617,N_10524,N_11574);
nor U12618 (N_12618,N_10609,N_10042);
and U12619 (N_12619,N_12194,N_12077);
and U12620 (N_12620,N_11860,N_10980);
nand U12621 (N_12621,N_10200,N_11912);
nand U12622 (N_12622,N_11880,N_10755);
nor U12623 (N_12623,N_12041,N_11156);
nor U12624 (N_12624,N_11660,N_10534);
nand U12625 (N_12625,N_10732,N_12010);
or U12626 (N_12626,N_10336,N_11437);
nand U12627 (N_12627,N_12036,N_10644);
nand U12628 (N_12628,N_11824,N_11044);
nand U12629 (N_12629,N_10569,N_11113);
or U12630 (N_12630,N_10497,N_11854);
and U12631 (N_12631,N_11657,N_10292);
nand U12632 (N_12632,N_12227,N_10345);
xnor U12633 (N_12633,N_12263,N_10553);
nand U12634 (N_12634,N_12346,N_11564);
nor U12635 (N_12635,N_12207,N_11687);
xnor U12636 (N_12636,N_12183,N_11572);
nor U12637 (N_12637,N_11932,N_10575);
and U12638 (N_12638,N_11263,N_10382);
nand U12639 (N_12639,N_11334,N_12053);
or U12640 (N_12640,N_11998,N_11277);
xor U12641 (N_12641,N_12147,N_11512);
and U12642 (N_12642,N_10508,N_10365);
and U12643 (N_12643,N_10996,N_12271);
or U12644 (N_12644,N_11129,N_12411);
nand U12645 (N_12645,N_11611,N_10376);
nand U12646 (N_12646,N_10933,N_10781);
nand U12647 (N_12647,N_11333,N_10713);
or U12648 (N_12648,N_12312,N_11318);
and U12649 (N_12649,N_12409,N_10052);
and U12650 (N_12650,N_11844,N_12199);
nor U12651 (N_12651,N_11244,N_11945);
and U12652 (N_12652,N_10602,N_11093);
and U12653 (N_12653,N_10489,N_10472);
nor U12654 (N_12654,N_10591,N_10640);
and U12655 (N_12655,N_11911,N_11418);
nand U12656 (N_12656,N_10587,N_10364);
nor U12657 (N_12657,N_10165,N_12285);
xor U12658 (N_12658,N_11730,N_12116);
nand U12659 (N_12659,N_10374,N_11058);
nand U12660 (N_12660,N_11444,N_12093);
nor U12661 (N_12661,N_12127,N_10000);
nor U12662 (N_12662,N_11592,N_11389);
nor U12663 (N_12663,N_11731,N_10361);
xor U12664 (N_12664,N_11118,N_10588);
or U12665 (N_12665,N_10825,N_10461);
xnor U12666 (N_12666,N_10990,N_10303);
nor U12667 (N_12667,N_10438,N_12365);
or U12668 (N_12668,N_10202,N_10054);
nor U12669 (N_12669,N_11608,N_12274);
nand U12670 (N_12670,N_11652,N_10455);
and U12671 (N_12671,N_12394,N_10969);
nand U12672 (N_12672,N_11099,N_11190);
xnor U12673 (N_12673,N_11997,N_10873);
xor U12674 (N_12674,N_11471,N_10225);
and U12675 (N_12675,N_10199,N_10972);
xor U12676 (N_12676,N_11985,N_12165);
or U12677 (N_12677,N_12099,N_10214);
xor U12678 (N_12678,N_11395,N_10538);
and U12679 (N_12679,N_10496,N_12225);
or U12680 (N_12680,N_10331,N_10203);
nor U12681 (N_12681,N_11014,N_10228);
nand U12682 (N_12682,N_10899,N_10817);
nand U12683 (N_12683,N_11170,N_10312);
nand U12684 (N_12684,N_10774,N_11746);
nand U12685 (N_12685,N_10257,N_12074);
nor U12686 (N_12686,N_11576,N_10060);
and U12687 (N_12687,N_10171,N_12172);
or U12688 (N_12688,N_11786,N_11594);
and U12689 (N_12689,N_11326,N_11151);
nor U12690 (N_12690,N_12370,N_11958);
nand U12691 (N_12691,N_10991,N_11180);
and U12692 (N_12692,N_12157,N_11069);
nor U12693 (N_12693,N_10707,N_11940);
nand U12694 (N_12694,N_10279,N_11668);
or U12695 (N_12695,N_12115,N_10872);
and U12696 (N_12696,N_12221,N_10466);
nand U12697 (N_12697,N_10527,N_10062);
or U12698 (N_12698,N_10338,N_11047);
nor U12699 (N_12699,N_11764,N_10695);
and U12700 (N_12700,N_12069,N_10007);
nand U12701 (N_12701,N_11691,N_11253);
or U12702 (N_12702,N_11989,N_11527);
or U12703 (N_12703,N_11528,N_10589);
nor U12704 (N_12704,N_12050,N_10163);
xnor U12705 (N_12705,N_10006,N_11688);
nor U12706 (N_12706,N_11116,N_10389);
and U12707 (N_12707,N_12252,N_11451);
and U12708 (N_12708,N_10617,N_11358);
xor U12709 (N_12709,N_11236,N_11449);
and U12710 (N_12710,N_10537,N_10089);
nor U12711 (N_12711,N_11125,N_10921);
or U12712 (N_12712,N_10932,N_10581);
nand U12713 (N_12713,N_11714,N_10528);
xnor U12714 (N_12714,N_11461,N_10959);
or U12715 (N_12715,N_11877,N_12180);
nor U12716 (N_12716,N_12422,N_11882);
nand U12717 (N_12717,N_11583,N_11428);
nand U12718 (N_12718,N_12123,N_10579);
and U12719 (N_12719,N_12206,N_12397);
nor U12720 (N_12720,N_10747,N_10009);
xor U12721 (N_12721,N_11967,N_11739);
and U12722 (N_12722,N_11770,N_10299);
xnor U12723 (N_12723,N_12215,N_10313);
or U12724 (N_12724,N_11452,N_11550);
nand U12725 (N_12725,N_10140,N_11910);
nor U12726 (N_12726,N_11393,N_10759);
or U12727 (N_12727,N_11946,N_11705);
xor U12728 (N_12728,N_10210,N_11876);
nor U12729 (N_12729,N_12419,N_12446);
or U12730 (N_12730,N_10884,N_12095);
xnor U12731 (N_12731,N_11225,N_10977);
xor U12732 (N_12732,N_10211,N_10683);
nor U12733 (N_12733,N_11674,N_10310);
nand U12734 (N_12734,N_10855,N_12467);
nor U12735 (N_12735,N_12204,N_10107);
xnor U12736 (N_12736,N_12073,N_11052);
or U12737 (N_12737,N_12190,N_12436);
nand U12738 (N_12738,N_10194,N_11907);
or U12739 (N_12739,N_10549,N_12401);
and U12740 (N_12740,N_10113,N_11003);
and U12741 (N_12741,N_11149,N_10393);
nor U12742 (N_12742,N_11883,N_11787);
or U12743 (N_12743,N_10362,N_12356);
or U12744 (N_12744,N_11916,N_11918);
nor U12745 (N_12745,N_11508,N_10535);
nand U12746 (N_12746,N_10432,N_10412);
xor U12747 (N_12747,N_11411,N_11063);
or U12748 (N_12748,N_10974,N_10055);
xnor U12749 (N_12749,N_11045,N_12425);
nand U12750 (N_12750,N_12361,N_12321);
nand U12751 (N_12751,N_10282,N_11728);
or U12752 (N_12752,N_10468,N_12112);
nand U12753 (N_12753,N_10475,N_12217);
or U12754 (N_12754,N_12484,N_11987);
xor U12755 (N_12755,N_11901,N_11552);
and U12756 (N_12756,N_11034,N_11595);
nand U12757 (N_12757,N_11330,N_11524);
nand U12758 (N_12758,N_10106,N_10810);
nand U12759 (N_12759,N_10543,N_11273);
nand U12760 (N_12760,N_12473,N_10844);
and U12761 (N_12761,N_10819,N_11857);
or U12762 (N_12762,N_10566,N_11321);
nor U12763 (N_12763,N_10041,N_10047);
xor U12764 (N_12764,N_10295,N_10596);
nand U12765 (N_12765,N_10845,N_10580);
or U12766 (N_12766,N_10155,N_10536);
xor U12767 (N_12767,N_10419,N_11986);
nor U12768 (N_12768,N_10500,N_11861);
and U12769 (N_12769,N_10387,N_11019);
xnor U12770 (N_12770,N_12284,N_12008);
nor U12771 (N_12771,N_10424,N_11545);
or U12772 (N_12772,N_10829,N_10624);
or U12773 (N_12773,N_11425,N_12337);
nand U12774 (N_12774,N_10631,N_11782);
xor U12775 (N_12775,N_12403,N_11396);
nor U12776 (N_12776,N_12006,N_11909);
or U12777 (N_12777,N_10418,N_11613);
xor U12778 (N_12778,N_12291,N_10077);
xor U12779 (N_12779,N_12045,N_10838);
nor U12780 (N_12780,N_11349,N_10168);
or U12781 (N_12781,N_10868,N_10334);
nand U12782 (N_12782,N_12426,N_10885);
and U12783 (N_12783,N_11536,N_11309);
or U12784 (N_12784,N_10728,N_11335);
nand U12785 (N_12785,N_10141,N_12283);
and U12786 (N_12786,N_11815,N_11260);
and U12787 (N_12787,N_10476,N_12210);
xor U12788 (N_12788,N_10297,N_11896);
xor U12789 (N_12789,N_11547,N_11284);
or U12790 (N_12790,N_10120,N_11441);
xnor U12791 (N_12791,N_11091,N_12261);
nand U12792 (N_12792,N_10018,N_11222);
nand U12793 (N_12793,N_10778,N_11154);
and U12794 (N_12794,N_10011,N_12448);
or U12795 (N_12795,N_10191,N_11055);
and U12796 (N_12796,N_12414,N_12173);
nand U12797 (N_12797,N_12150,N_10383);
nand U12798 (N_12798,N_12044,N_11313);
or U12799 (N_12799,N_11629,N_10801);
nand U12800 (N_12800,N_11305,N_11686);
nand U12801 (N_12801,N_11212,N_10121);
and U12802 (N_12802,N_10862,N_10665);
and U12803 (N_12803,N_10045,N_10286);
or U12804 (N_12804,N_11700,N_11371);
or U12805 (N_12805,N_11571,N_10722);
nor U12806 (N_12806,N_10246,N_11177);
xnor U12807 (N_12807,N_12386,N_10632);
or U12808 (N_12808,N_10606,N_11105);
and U12809 (N_12809,N_12384,N_10682);
nor U12810 (N_12810,N_10558,N_11210);
and U12811 (N_12811,N_11460,N_11308);
nor U12812 (N_12812,N_10407,N_10850);
nand U12813 (N_12813,N_10226,N_10207);
or U12814 (N_12814,N_10131,N_11826);
or U12815 (N_12815,N_11040,N_11757);
nand U12816 (N_12816,N_11399,N_10953);
nand U12817 (N_12817,N_11216,N_11832);
xnor U12818 (N_12818,N_12331,N_10448);
nand U12819 (N_12819,N_12481,N_11507);
xnor U12820 (N_12820,N_10645,N_10762);
or U12821 (N_12821,N_10798,N_10942);
and U12822 (N_12822,N_11521,N_12267);
xor U12823 (N_12823,N_11167,N_11634);
and U12824 (N_12824,N_11711,N_11797);
nand U12825 (N_12825,N_12042,N_10578);
nand U12826 (N_12826,N_10354,N_11000);
or U12827 (N_12827,N_11311,N_10309);
or U12828 (N_12828,N_12021,N_12495);
nand U12829 (N_12829,N_10786,N_10291);
xor U12830 (N_12830,N_11495,N_12105);
or U12831 (N_12831,N_10988,N_11601);
and U12832 (N_12832,N_11898,N_11327);
or U12833 (N_12833,N_10704,N_10048);
xor U12834 (N_12834,N_12219,N_12243);
and U12835 (N_12835,N_11203,N_11375);
and U12836 (N_12836,N_11293,N_10188);
nor U12837 (N_12837,N_12390,N_10469);
and U12838 (N_12838,N_10901,N_12491);
or U12839 (N_12839,N_10236,N_11565);
and U12840 (N_12840,N_10714,N_10480);
nand U12841 (N_12841,N_12434,N_10938);
xor U12842 (N_12842,N_10718,N_10928);
and U12843 (N_12843,N_11174,N_10305);
and U12844 (N_12844,N_11410,N_10135);
xnor U12845 (N_12845,N_11843,N_11971);
and U12846 (N_12846,N_10675,N_11783);
or U12847 (N_12847,N_10937,N_12315);
xor U12848 (N_12848,N_11023,N_10895);
nor U12849 (N_12849,N_11179,N_10435);
and U12850 (N_12850,N_10170,N_11707);
xor U12851 (N_12851,N_11017,N_11459);
xor U12852 (N_12852,N_12415,N_11233);
nor U12853 (N_12853,N_12152,N_10902);
or U12854 (N_12854,N_10029,N_11175);
or U12855 (N_12855,N_11892,N_11221);
or U12856 (N_12856,N_10989,N_11596);
nor U12857 (N_12857,N_11920,N_12134);
nand U12858 (N_12858,N_11900,N_10751);
and U12859 (N_12859,N_10341,N_12160);
nand U12860 (N_12860,N_10750,N_12454);
xnor U12861 (N_12861,N_10615,N_10881);
xnor U12862 (N_12862,N_11132,N_12121);
or U12863 (N_12863,N_10693,N_10067);
nor U12864 (N_12864,N_10290,N_10287);
or U12865 (N_12865,N_11540,N_10814);
and U12866 (N_12866,N_12114,N_10132);
nor U12867 (N_12867,N_12369,N_11473);
xor U12868 (N_12868,N_11365,N_11343);
nand U12869 (N_12869,N_11569,N_10146);
nor U12870 (N_12870,N_12489,N_11369);
and U12871 (N_12871,N_11504,N_10443);
xnor U12872 (N_12872,N_12342,N_10560);
or U12873 (N_12873,N_10325,N_10522);
xnor U12874 (N_12874,N_11913,N_10218);
and U12875 (N_12875,N_10125,N_10849);
or U12876 (N_12876,N_12354,N_12241);
and U12877 (N_12877,N_11223,N_10093);
nand U12878 (N_12878,N_11204,N_11035);
and U12879 (N_12879,N_11743,N_11704);
nand U12880 (N_12880,N_10372,N_10944);
or U12881 (N_12881,N_10806,N_10219);
or U12882 (N_12882,N_10385,N_11381);
nor U12883 (N_12883,N_12000,N_12177);
and U12884 (N_12884,N_12334,N_11871);
xor U12885 (N_12885,N_12238,N_11534);
nor U12886 (N_12886,N_11819,N_12013);
nand U12887 (N_12887,N_10671,N_11879);
xor U12888 (N_12888,N_10080,N_10182);
or U12889 (N_12889,N_10504,N_11114);
or U12890 (N_12890,N_11570,N_12332);
nor U12891 (N_12891,N_10843,N_12360);
or U12892 (N_12892,N_12406,N_11109);
xnor U12893 (N_12893,N_11983,N_12326);
nand U12894 (N_12894,N_11367,N_12335);
nand U12895 (N_12895,N_12358,N_11587);
xnor U12896 (N_12896,N_12087,N_10919);
or U12897 (N_12897,N_11713,N_10208);
and U12898 (N_12898,N_10501,N_10516);
nor U12899 (N_12899,N_10532,N_11046);
or U12900 (N_12900,N_11443,N_10488);
nand U12901 (N_12901,N_10744,N_10517);
or U12902 (N_12902,N_10076,N_11039);
and U12903 (N_12903,N_12143,N_10353);
nor U12904 (N_12904,N_11538,N_10963);
nor U12905 (N_12905,N_11081,N_12288);
nor U12906 (N_12906,N_12465,N_11600);
xor U12907 (N_12907,N_10807,N_11789);
nand U12908 (N_12908,N_10017,N_10661);
nor U12909 (N_12909,N_12230,N_12417);
xor U12910 (N_12910,N_10451,N_11478);
xor U12911 (N_12911,N_10540,N_10178);
nor U12912 (N_12912,N_11562,N_10521);
and U12913 (N_12913,N_10498,N_11188);
xnor U12914 (N_12914,N_12433,N_11931);
xnor U12915 (N_12915,N_12477,N_10262);
nor U12916 (N_12916,N_10916,N_11211);
or U12917 (N_12917,N_11933,N_10509);
nor U12918 (N_12918,N_11407,N_10043);
nand U12919 (N_12919,N_10294,N_12378);
nor U12920 (N_12920,N_11868,N_10927);
nor U12921 (N_12921,N_11127,N_10975);
nor U12922 (N_12922,N_11532,N_11673);
nor U12923 (N_12923,N_11191,N_11742);
xor U12924 (N_12924,N_11430,N_10127);
xor U12925 (N_12925,N_10585,N_12003);
nand U12926 (N_12926,N_10072,N_12383);
nand U12927 (N_12927,N_12202,N_12336);
nor U12928 (N_12928,N_12387,N_10563);
or U12929 (N_12929,N_10764,N_10788);
or U12930 (N_12930,N_11974,N_12244);
or U12931 (N_12931,N_10839,N_10217);
and U12932 (N_12932,N_10028,N_12028);
and U12933 (N_12933,N_11831,N_12188);
xnor U12934 (N_12934,N_12389,N_12056);
nor U12935 (N_12935,N_10274,N_12393);
nand U12936 (N_12936,N_11602,N_11376);
or U12937 (N_12937,N_11921,N_10343);
nor U12938 (N_12938,N_11890,N_12171);
or U12939 (N_12939,N_12063,N_11620);
or U12940 (N_12940,N_11799,N_10657);
nand U12941 (N_12941,N_12254,N_11497);
or U12942 (N_12942,N_11006,N_11062);
nor U12943 (N_12943,N_11362,N_12431);
nand U12944 (N_12944,N_10276,N_12246);
xor U12945 (N_12945,N_12349,N_12163);
xnor U12946 (N_12946,N_11630,N_11950);
or U12947 (N_12947,N_11276,N_12060);
xnor U12948 (N_12948,N_10719,N_12270);
and U12949 (N_12949,N_10865,N_12449);
and U12950 (N_12950,N_10275,N_11853);
nand U12951 (N_12951,N_11667,N_10431);
xnor U12952 (N_12952,N_11298,N_11659);
and U12953 (N_12953,N_12048,N_10705);
or U12954 (N_12954,N_11924,N_11715);
xor U12955 (N_12955,N_10337,N_10812);
nand U12956 (N_12956,N_11446,N_11701);
nor U12957 (N_12957,N_10685,N_10625);
nand U12958 (N_12958,N_11760,N_12323);
xnor U12959 (N_12959,N_11199,N_10244);
xor U12960 (N_12960,N_10880,N_10993);
and U12961 (N_12961,N_11914,N_10375);
nor U12962 (N_12962,N_11496,N_10956);
or U12963 (N_12963,N_10743,N_10633);
nor U12964 (N_12964,N_12438,N_12019);
or U12965 (N_12965,N_11245,N_10677);
xor U12966 (N_12966,N_11505,N_11484);
xor U12967 (N_12967,N_10097,N_11848);
nor U12968 (N_12968,N_11102,N_11681);
nand U12969 (N_12969,N_12359,N_10623);
xor U12970 (N_12970,N_10450,N_11670);
or U12971 (N_12971,N_11838,N_12237);
nand U12972 (N_12972,N_11533,N_12343);
nand U12973 (N_12973,N_10024,N_11208);
nand U12974 (N_12974,N_10666,N_11226);
nand U12975 (N_12975,N_11121,N_10058);
or U12976 (N_12976,N_10092,N_10149);
xnor U12977 (N_12977,N_12007,N_12404);
xnor U12978 (N_12978,N_10315,N_11609);
or U12979 (N_12979,N_11426,N_11092);
nor U12980 (N_12980,N_11173,N_12377);
xor U12981 (N_12981,N_11716,N_10440);
xor U12982 (N_12982,N_12460,N_10185);
or U12983 (N_12983,N_11481,N_10979);
and U12984 (N_12984,N_11954,N_10117);
and U12985 (N_12985,N_11798,N_12026);
or U12986 (N_12986,N_11623,N_10530);
or U12987 (N_12987,N_10227,N_11227);
and U12988 (N_12988,N_10694,N_10056);
and U12989 (N_12989,N_12305,N_11676);
nand U12990 (N_12990,N_12303,N_12196);
or U12991 (N_12991,N_11283,N_11171);
nor U12992 (N_12992,N_11689,N_11568);
nor U12993 (N_12993,N_11827,N_11751);
nand U12994 (N_12994,N_12374,N_12493);
nand U12995 (N_12995,N_10483,N_10724);
xnor U12996 (N_12996,N_12466,N_11526);
or U12997 (N_12997,N_11520,N_11784);
or U12998 (N_12998,N_10936,N_10505);
and U12999 (N_12999,N_11627,N_12385);
or U13000 (N_13000,N_10022,N_10032);
and U13001 (N_13001,N_11082,N_12122);
nor U13002 (N_13002,N_11679,N_10391);
and U13003 (N_13003,N_11115,N_10399);
nand U13004 (N_13004,N_11345,N_12412);
xnor U13005 (N_13005,N_10720,N_11131);
xor U13006 (N_13006,N_12313,N_10688);
or U13007 (N_13007,N_12338,N_12130);
and U13008 (N_13008,N_11957,N_10739);
and U13009 (N_13009,N_10952,N_11262);
and U13010 (N_13010,N_10301,N_11808);
nand U13011 (N_13011,N_11462,N_10869);
nor U13012 (N_13012,N_12487,N_12068);
nor U13013 (N_13013,N_11097,N_10355);
xnor U13014 (N_13014,N_11556,N_12286);
and U13015 (N_13015,N_12424,N_11554);
xnor U13016 (N_13016,N_12480,N_12032);
nand U13017 (N_13017,N_12164,N_11447);
xor U13018 (N_13018,N_11685,N_10847);
and U13019 (N_13019,N_10152,N_10968);
or U13020 (N_13020,N_10085,N_11250);
nand U13021 (N_13021,N_11465,N_11071);
and U13022 (N_13022,N_10648,N_11755);
or U13023 (N_13023,N_11740,N_12135);
or U13024 (N_13024,N_11328,N_11392);
xor U13025 (N_13025,N_10235,N_12220);
nor U13026 (N_13026,N_11166,N_11982);
nand U13027 (N_13027,N_12295,N_11207);
and U13028 (N_13028,N_10074,N_12307);
nor U13029 (N_13029,N_11561,N_12399);
nor U13030 (N_13030,N_11943,N_10283);
or U13031 (N_13031,N_10684,N_12213);
or U13032 (N_13032,N_10215,N_10231);
xor U13033 (N_13033,N_10453,N_10164);
xnor U13034 (N_13034,N_11357,N_12325);
or U13035 (N_13035,N_10518,N_10690);
nor U13036 (N_13036,N_11279,N_10660);
nand U13037 (N_13037,N_10793,N_10441);
nand U13038 (N_13038,N_11722,N_10860);
xnor U13039 (N_13039,N_12138,N_11294);
and U13040 (N_13040,N_11022,N_10422);
and U13041 (N_13041,N_10561,N_10119);
and U13042 (N_13042,N_11650,N_11979);
or U13043 (N_13043,N_11869,N_11809);
nand U13044 (N_13044,N_11938,N_11988);
nor U13045 (N_13045,N_10940,N_11406);
or U13046 (N_13046,N_11683,N_10269);
nand U13047 (N_13047,N_11617,N_10866);
or U13048 (N_13048,N_10408,N_11581);
nor U13049 (N_13049,N_11269,N_10248);
or U13050 (N_13050,N_11135,N_10867);
and U13051 (N_13051,N_11214,N_10878);
xnor U13052 (N_13052,N_11029,N_10233);
nand U13053 (N_13053,N_10012,N_12094);
and U13054 (N_13054,N_11331,N_12445);
and U13055 (N_13055,N_12066,N_11654);
or U13056 (N_13056,N_11563,N_11996);
and U13057 (N_13057,N_12249,N_11106);
xnor U13058 (N_13058,N_10700,N_12352);
nor U13059 (N_13059,N_11354,N_11015);
and U13060 (N_13060,N_11432,N_11010);
or U13061 (N_13061,N_10401,N_11863);
xor U13062 (N_13062,N_11834,N_11500);
nand U13063 (N_13063,N_11889,N_10319);
nand U13064 (N_13064,N_10363,N_12102);
or U13065 (N_13065,N_10388,N_11427);
xor U13066 (N_13066,N_12088,N_11257);
nor U13067 (N_13067,N_10573,N_12193);
nand U13068 (N_13068,N_10582,N_10698);
or U13069 (N_13069,N_11104,N_11964);
or U13070 (N_13070,N_11256,N_12300);
xor U13071 (N_13071,N_11516,N_11599);
xor U13072 (N_13072,N_12118,N_10966);
nand U13073 (N_13073,N_10603,N_12486);
nand U13074 (N_13074,N_12071,N_11433);
xor U13075 (N_13075,N_10708,N_11598);
and U13076 (N_13076,N_11694,N_10333);
and U13077 (N_13077,N_12442,N_10040);
nand U13078 (N_13078,N_11531,N_11682);
nand U13079 (N_13079,N_11553,N_11192);
xnor U13080 (N_13080,N_10861,N_11514);
nand U13081 (N_13081,N_12057,N_11975);
xor U13082 (N_13082,N_11140,N_11805);
and U13083 (N_13083,N_11024,N_11150);
nand U13084 (N_13084,N_12292,N_10053);
nand U13085 (N_13085,N_10555,N_12278);
nor U13086 (N_13086,N_10223,N_11641);
nand U13087 (N_13087,N_11165,N_10831);
nand U13088 (N_13088,N_11806,N_10349);
and U13089 (N_13089,N_11384,N_10434);
xnor U13090 (N_13090,N_10782,N_12141);
xor U13091 (N_13091,N_12472,N_11830);
xor U13092 (N_13092,N_10780,N_11796);
nand U13093 (N_13093,N_10709,N_11315);
and U13094 (N_13094,N_10678,N_11419);
nor U13095 (N_13095,N_11899,N_10725);
nand U13096 (N_13096,N_10061,N_10129);
nor U13097 (N_13097,N_10945,N_11678);
or U13098 (N_13098,N_10655,N_12098);
nor U13099 (N_13099,N_12039,N_10766);
and U13100 (N_13100,N_10706,N_12214);
and U13101 (N_13101,N_11137,N_11511);
nor U13102 (N_13102,N_10479,N_10917);
nor U13103 (N_13103,N_11157,N_11342);
or U13104 (N_13104,N_10071,N_10264);
and U13105 (N_13105,N_11235,N_11607);
nand U13106 (N_13106,N_10160,N_10176);
xnor U13107 (N_13107,N_12078,N_11382);
xnor U13108 (N_13108,N_12185,N_11733);
nand U13109 (N_13109,N_12233,N_10392);
xor U13110 (N_13110,N_10104,N_11038);
and U13111 (N_13111,N_12381,N_11965);
nand U13112 (N_13112,N_12396,N_10525);
and U13113 (N_13113,N_11870,N_11973);
and U13114 (N_13114,N_11671,N_11509);
nand U13115 (N_13115,N_11292,N_10811);
and U13116 (N_13116,N_10462,N_12153);
or U13117 (N_13117,N_11631,N_11636);
nand U13118 (N_13118,N_11963,N_10417);
nor U13119 (N_13119,N_10371,N_10108);
xor U13120 (N_13120,N_11304,N_12051);
or U13121 (N_13121,N_11597,N_11401);
and U13122 (N_13122,N_12260,N_12392);
nor U13123 (N_13123,N_10904,N_10915);
nor U13124 (N_13124,N_10614,N_12120);
nor U13125 (N_13125,N_11404,N_11881);
or U13126 (N_13126,N_11781,N_11440);
and U13127 (N_13127,N_11002,N_11080);
nor U13128 (N_13128,N_10096,N_11662);
and U13129 (N_13129,N_11661,N_11992);
and U13130 (N_13130,N_10205,N_11301);
nand U13131 (N_13131,N_11201,N_11200);
xor U13132 (N_13132,N_11995,N_12176);
nand U13133 (N_13133,N_10397,N_11351);
xor U13134 (N_13134,N_11146,N_11859);
and U13135 (N_13135,N_10600,N_10403);
and U13136 (N_13136,N_10754,N_11578);
or U13137 (N_13137,N_11142,N_11119);
or U13138 (N_13138,N_10503,N_10001);
or U13139 (N_13139,N_11398,N_10740);
nor U13140 (N_13140,N_11271,N_11615);
and U13141 (N_13141,N_12070,N_10960);
nand U13142 (N_13142,N_10949,N_10510);
nor U13143 (N_13143,N_11625,N_11072);
and U13144 (N_13144,N_11147,N_10158);
and U13145 (N_13145,N_11841,N_11810);
nand U13146 (N_13146,N_12327,N_10014);
xor U13147 (N_13147,N_10647,N_11246);
or U13148 (N_13148,N_11604,N_11632);
or U13149 (N_13149,N_10837,N_12298);
nand U13150 (N_13150,N_11855,N_11626);
nand U13151 (N_13151,N_12301,N_11468);
nor U13152 (N_13152,N_10221,N_12273);
xor U13153 (N_13153,N_11152,N_11066);
or U13154 (N_13154,N_11852,N_10025);
xnor U13155 (N_13155,N_10406,N_12110);
or U13156 (N_13156,N_12250,N_12097);
and U13157 (N_13157,N_11111,N_10068);
nand U13158 (N_13158,N_12084,N_10691);
and U13159 (N_13159,N_10241,N_11197);
xor U13160 (N_13160,N_11340,N_10820);
and U13161 (N_13161,N_10249,N_10395);
nor U13162 (N_13162,N_11028,N_11803);
or U13163 (N_13163,N_11457,N_11346);
and U13164 (N_13164,N_12395,N_10368);
or U13165 (N_13165,N_12224,N_10069);
xnor U13166 (N_13166,N_10946,N_11048);
or U13167 (N_13167,N_11241,N_10459);
and U13168 (N_13168,N_10144,N_10857);
and U13169 (N_13169,N_11544,N_10598);
nor U13170 (N_13170,N_12310,N_11231);
nor U13171 (N_13171,N_12280,N_11923);
or U13172 (N_13172,N_12209,N_11926);
and U13173 (N_13173,N_10981,N_10285);
xnor U13174 (N_13174,N_10663,N_10520);
xor U13175 (N_13175,N_11475,N_12104);
or U13176 (N_13176,N_11423,N_12136);
nor U13177 (N_13177,N_11436,N_11619);
xor U13178 (N_13178,N_10083,N_12052);
xor U13179 (N_13179,N_10970,N_10662);
or U13180 (N_13180,N_11373,N_10351);
nand U13181 (N_13181,N_11108,N_10396);
nand U13182 (N_13182,N_11785,N_12174);
or U13183 (N_13183,N_12216,N_10172);
xor U13184 (N_13184,N_10823,N_10546);
or U13185 (N_13185,N_10444,N_11377);
nand U13186 (N_13186,N_11732,N_12255);
nand U13187 (N_13187,N_11925,N_11530);
nand U13188 (N_13188,N_11720,N_10193);
nand U13189 (N_13189,N_11112,N_11274);
nand U13190 (N_13190,N_11323,N_11546);
and U13191 (N_13191,N_10523,N_11818);
or U13192 (N_13192,N_10656,N_10442);
or U13193 (N_13193,N_11252,N_10010);
or U13194 (N_13194,N_11130,N_10941);
xnor U13195 (N_13195,N_10853,N_12170);
or U13196 (N_13196,N_12282,N_10870);
xnor U13197 (N_13197,N_10384,N_12471);
nor U13198 (N_13198,N_10828,N_11310);
nand U13199 (N_13199,N_11051,N_10493);
xnor U13200 (N_13200,N_10487,N_10122);
nand U13201 (N_13201,N_11939,N_12049);
xnor U13202 (N_13202,N_10057,N_11275);
nand U13203 (N_13203,N_11588,N_10326);
nor U13204 (N_13204,N_11498,N_10346);
nor U13205 (N_13205,N_12076,N_12309);
and U13206 (N_13206,N_11948,N_12031);
nor U13207 (N_13207,N_11719,N_12340);
nand U13208 (N_13208,N_10910,N_10787);
xor U13209 (N_13209,N_10891,N_12353);
and U13210 (N_13210,N_10271,N_10289);
and U13211 (N_13211,N_12231,N_11822);
nor U13212 (N_13212,N_10971,N_11400);
nand U13213 (N_13213,N_11117,N_11126);
or U13214 (N_13214,N_12124,N_11289);
nor U13215 (N_13215,N_10402,N_10906);
xnor U13216 (N_13216,N_11363,N_11438);
xnor U13217 (N_13217,N_11800,N_10209);
or U13218 (N_13218,N_11181,N_10586);
and U13219 (N_13219,N_11647,N_12034);
and U13220 (N_13220,N_11237,N_11833);
nor U13221 (N_13221,N_10756,N_10268);
nor U13222 (N_13222,N_11143,N_12455);
nand U13223 (N_13223,N_10929,N_10421);
nand U13224 (N_13224,N_10304,N_11648);
xnor U13225 (N_13225,N_11049,N_11205);
and U13226 (N_13226,N_11741,N_11710);
xor U13227 (N_13227,N_10833,N_10091);
xnor U13228 (N_13228,N_10410,N_12373);
and U13229 (N_13229,N_10890,N_10892);
and U13230 (N_13230,N_12144,N_10515);
nor U13231 (N_13231,N_10595,N_12423);
xor U13232 (N_13232,N_11885,N_12128);
and U13233 (N_13233,N_10183,N_10177);
nand U13234 (N_13234,N_10983,N_11008);
and U13235 (N_13235,N_11489,N_11264);
or U13236 (N_13236,N_11232,N_12211);
nand U13237 (N_13237,N_10513,N_11603);
xor U13238 (N_13238,N_10809,N_11480);
nand U13239 (N_13239,N_11016,N_11302);
and U13240 (N_13240,N_12362,N_10133);
or U13241 (N_13241,N_11139,N_10710);
and U13242 (N_13242,N_10035,N_11807);
or U13243 (N_13243,N_10887,N_11355);
and U13244 (N_13244,N_11060,N_11420);
or U13245 (N_13245,N_10982,N_11193);
nand U13246 (N_13246,N_12368,N_11007);
and U13247 (N_13247,N_10703,N_10726);
or U13248 (N_13248,N_10544,N_10259);
xnor U13249 (N_13249,N_11771,N_10692);
nand U13250 (N_13250,N_12444,N_10038);
and U13251 (N_13251,N_11501,N_12139);
xnor U13252 (N_13252,N_11765,N_10565);
nand U13253 (N_13253,N_10931,N_10757);
xor U13254 (N_13254,N_11936,N_10626);
or U13255 (N_13255,N_11878,N_10502);
nand U13256 (N_13256,N_10005,N_12137);
nor U13257 (N_13257,N_10745,N_10552);
xnor U13258 (N_13258,N_10049,N_11314);
xor U13259 (N_13259,N_11836,N_10347);
or U13260 (N_13260,N_10689,N_10474);
and U13261 (N_13261,N_11729,N_10712);
xor U13262 (N_13262,N_10465,N_10914);
nand U13263 (N_13263,N_10322,N_11350);
xnor U13264 (N_13264,N_11133,N_10548);
nor U13265 (N_13265,N_11209,N_10604);
and U13266 (N_13266,N_11299,N_11078);
nor U13267 (N_13267,N_11070,N_10109);
nand U13268 (N_13268,N_10273,N_10567);
or U13269 (N_13269,N_12228,N_10216);
nand U13270 (N_13270,N_10761,N_11927);
nand U13271 (N_13271,N_11840,N_10267);
nor U13272 (N_13272,N_11435,N_10934);
nand U13273 (N_13273,N_10110,N_11353);
or U13274 (N_13274,N_11697,N_10116);
and U13275 (N_13275,N_10196,N_11238);
nand U13276 (N_13276,N_10894,N_11455);
and U13277 (N_13277,N_12450,N_11886);
and U13278 (N_13278,N_11677,N_10542);
nor U13279 (N_13279,N_10797,N_10545);
xor U13280 (N_13280,N_11952,N_11306);
nand U13281 (N_13281,N_12413,N_12457);
and U13282 (N_13282,N_12079,N_10175);
and U13283 (N_13283,N_10619,N_10075);
xor U13284 (N_13284,N_10649,N_12005);
nor U13285 (N_13285,N_12205,N_10316);
nor U13286 (N_13286,N_10955,N_10340);
xor U13287 (N_13287,N_11829,N_11884);
and U13288 (N_13288,N_10871,N_10463);
xor U13289 (N_13289,N_12289,N_10590);
xor U13290 (N_13290,N_10237,N_11385);
nor U13291 (N_13291,N_11872,N_10015);
xnor U13292 (N_13292,N_10717,N_10676);
and U13293 (N_13293,N_10308,N_11145);
nand U13294 (N_13294,N_11874,N_11768);
xnor U13295 (N_13295,N_11084,N_11037);
nor U13296 (N_13296,N_10879,N_11178);
or U13297 (N_13297,N_10557,N_11134);
and U13298 (N_13298,N_11185,N_10987);
nor U13299 (N_13299,N_12379,N_10531);
nand U13300 (N_13300,N_10909,N_10568);
and U13301 (N_13301,N_10180,N_10327);
xnor U13302 (N_13302,N_11409,N_12113);
or U13303 (N_13303,N_12058,N_11414);
or U13304 (N_13304,N_10783,N_10852);
nand U13305 (N_13305,N_10875,N_10746);
nand U13306 (N_13306,N_10512,N_11380);
or U13307 (N_13307,N_10254,N_10494);
nand U13308 (N_13308,N_11324,N_10098);
nor U13309 (N_13309,N_10922,N_12132);
and U13310 (N_13310,N_11591,N_10103);
xor U13311 (N_13311,N_11054,N_11230);
xor U13312 (N_13312,N_10019,N_11095);
nand U13313 (N_13313,N_12482,N_11813);
or U13314 (N_13314,N_12226,N_11424);
nor U13315 (N_13315,N_10457,N_10826);
nor U13316 (N_13316,N_12311,N_11195);
or U13317 (N_13317,N_10293,N_12023);
xnor U13318 (N_13318,N_11219,N_11692);
nand U13319 (N_13319,N_10266,N_11640);
and U13320 (N_13320,N_10723,N_11013);
xor U13321 (N_13321,N_10467,N_12029);
or U13322 (N_13322,N_12146,N_11032);
nand U13323 (N_13323,N_12375,N_10352);
nor U13324 (N_13324,N_11593,N_12475);
nor U13325 (N_13325,N_11675,N_11894);
nand U13326 (N_13326,N_11176,N_10767);
nor U13327 (N_13327,N_10769,N_11821);
and U13328 (N_13328,N_10926,N_11769);
nor U13329 (N_13329,N_11442,N_11240);
nor U13330 (N_13330,N_11762,N_11138);
nor U13331 (N_13331,N_11286,N_12464);
or U13332 (N_13332,N_10059,N_11703);
xnor U13333 (N_13333,N_10378,N_10986);
xnor U13334 (N_13334,N_12075,N_10529);
xnor U13335 (N_13335,N_12240,N_11075);
nand U13336 (N_13336,N_10943,N_10366);
or U13337 (N_13337,N_10484,N_12483);
xor U13338 (N_13338,N_11476,N_11332);
nand U13339 (N_13339,N_11107,N_11811);
xor U13340 (N_13340,N_11748,N_11845);
and U13341 (N_13341,N_11325,N_10574);
nand U13342 (N_13342,N_11266,N_10350);
or U13343 (N_13343,N_10836,N_11352);
and U13344 (N_13344,N_10288,N_11666);
nand U13345 (N_13345,N_11434,N_12065);
xnor U13346 (N_13346,N_10253,N_11043);
and U13347 (N_13347,N_11773,N_10539);
xnor U13348 (N_13348,N_11795,N_10903);
nand U13349 (N_13349,N_10673,N_11041);
or U13350 (N_13350,N_11402,N_10335);
or U13351 (N_13351,N_10668,N_12468);
nand U13352 (N_13352,N_12089,N_11767);
nor U13353 (N_13353,N_12257,N_10206);
nor U13354 (N_13354,N_10818,N_12443);
or U13355 (N_13355,N_10882,N_10697);
or U13356 (N_13356,N_11969,N_11103);
nor U13357 (N_13357,N_10607,N_12429);
and U13358 (N_13358,N_12407,N_11999);
and U13359 (N_13359,N_10420,N_10147);
nor U13360 (N_13360,N_11794,N_11649);
nand U13361 (N_13361,N_11968,N_10101);
xor U13362 (N_13362,N_10284,N_11942);
or U13363 (N_13363,N_10066,N_10734);
nor U13364 (N_13364,N_11031,N_12363);
xnor U13365 (N_13365,N_10930,N_12232);
nor U13366 (N_13366,N_11539,N_10957);
nand U13367 (N_13367,N_10775,N_10426);
xor U13368 (N_13368,N_11930,N_10962);
xor U13369 (N_13369,N_10186,N_12145);
xnor U13370 (N_13370,N_10898,N_10251);
nor U13371 (N_13371,N_11849,N_10925);
nand U13372 (N_13372,N_10148,N_10994);
and U13373 (N_13373,N_11663,N_12372);
and U13374 (N_13374,N_11169,N_12191);
nand U13375 (N_13375,N_11633,N_12350);
nor U13376 (N_13376,N_11506,N_11217);
nor U13377 (N_13377,N_11919,N_11148);
nor U13378 (N_13378,N_10554,N_11307);
nor U13379 (N_13379,N_10667,N_11291);
nand U13380 (N_13380,N_11823,N_11628);
or U13381 (N_13381,N_11984,N_10859);
nand U13382 (N_13382,N_12357,N_10840);
nor U13383 (N_13383,N_12440,N_10612);
xnor U13384 (N_13384,N_11726,N_12318);
and U13385 (N_13385,N_11493,N_10064);
nor U13386 (N_13386,N_10507,N_12236);
nor U13387 (N_13387,N_10976,N_11817);
and U13388 (N_13388,N_11754,N_10576);
nor U13389 (N_13389,N_12494,N_10339);
xor U13390 (N_13390,N_11472,N_11858);
nand U13391 (N_13391,N_12380,N_11492);
nand U13392 (N_13392,N_10130,N_12420);
xnor U13393 (N_13393,N_11403,N_10954);
xnor U13394 (N_13394,N_10593,N_10913);
nor U13395 (N_13395,N_11584,N_11922);
and U13396 (N_13396,N_12371,N_12179);
and U13397 (N_13397,N_11837,N_12400);
nor U13398 (N_13398,N_12490,N_11360);
or U13399 (N_13399,N_10034,N_12080);
nor U13400 (N_13400,N_12033,N_12447);
and U13401 (N_13401,N_10252,N_11464);
nand U13402 (N_13402,N_10822,N_11866);
xnor U13403 (N_13403,N_10145,N_10967);
or U13404 (N_13404,N_11690,N_11606);
nand U13405 (N_13405,N_11033,N_10437);
nor U13406 (N_13406,N_11397,N_11944);
xor U13407 (N_13407,N_11224,N_11610);
nor U13408 (N_13408,N_11431,N_11288);
nor U13409 (N_13409,N_12302,N_11061);
and U13410 (N_13410,N_11144,N_12451);
xor U13411 (N_13411,N_11655,N_12151);
and U13412 (N_13412,N_11474,N_10670);
or U13413 (N_13413,N_10157,N_10912);
xor U13414 (N_13414,N_12017,N_12364);
nand U13415 (N_13415,N_12022,N_11036);
nand U13416 (N_13416,N_11888,N_10429);
nand U13417 (N_13417,N_10583,N_11651);
xnor U13418 (N_13418,N_12320,N_10134);
nor U13419 (N_13419,N_10302,N_10330);
or U13420 (N_13420,N_11580,N_10893);
nand U13421 (N_13421,N_11749,N_12427);
or U13422 (N_13422,N_11164,N_10863);
and U13423 (N_13423,N_10918,N_10984);
or U13424 (N_13424,N_11820,N_11073);
nor U13425 (N_13425,N_11960,N_12441);
or U13426 (N_13426,N_10794,N_11356);
xnor U13427 (N_13427,N_10240,N_10082);
and U13428 (N_13428,N_12330,N_11696);
nor U13429 (N_13429,N_12293,N_11076);
or U13430 (N_13430,N_10179,N_12351);
and U13431 (N_13431,N_10115,N_12297);
nand U13432 (N_13432,N_12418,N_12203);
and U13433 (N_13433,N_11788,N_10473);
xor U13434 (N_13434,N_11312,N_11186);
and U13435 (N_13435,N_11215,N_11001);
and U13436 (N_13436,N_10306,N_11519);
nor U13437 (N_13437,N_12015,N_12154);
and U13438 (N_13438,N_10298,N_10173);
nor U13439 (N_13439,N_11280,N_12035);
and U13440 (N_13440,N_11009,N_10622);
nand U13441 (N_13441,N_11790,N_12218);
xor U13442 (N_13442,N_11725,N_10716);
or U13443 (N_13443,N_10947,N_12061);
or U13444 (N_13444,N_11951,N_11902);
xnor U13445 (N_13445,N_11672,N_11386);
nand U13446 (N_13446,N_11366,N_10166);
nor U13447 (N_13447,N_11281,N_11196);
or U13448 (N_13448,N_11792,N_10802);
and U13449 (N_13449,N_11978,N_11270);
nor U13450 (N_13450,N_12090,N_10114);
or U13451 (N_13451,N_12142,N_11011);
and U13452 (N_13452,N_12339,N_12347);
or U13453 (N_13453,N_10735,N_12072);
nand U13454 (N_13454,N_10900,N_11329);
nor U13455 (N_13455,N_11793,N_10445);
and U13456 (N_13456,N_12382,N_10785);
and U13457 (N_13457,N_12009,N_11961);
nand U13458 (N_13458,N_10189,N_10250);
and U13459 (N_13459,N_10950,N_11698);
nand U13460 (N_13460,N_11582,N_12294);
xnor U13461 (N_13461,N_10813,N_12189);
or U13462 (N_13462,N_11247,N_11499);
or U13463 (N_13463,N_12037,N_12166);
or U13464 (N_13464,N_12247,N_11825);
or U13465 (N_13465,N_12100,N_11862);
and U13466 (N_13466,N_11467,N_10321);
nor U13467 (N_13467,N_11439,N_12197);
or U13468 (N_13468,N_11490,N_11454);
nor U13469 (N_13469,N_10051,N_11867);
and U13470 (N_13470,N_11510,N_10213);
and U13471 (N_13471,N_12223,N_10239);
nor U13472 (N_13472,N_10630,N_11503);
nand U13473 (N_13473,N_11251,N_11935);
nand U13474 (N_13474,N_10317,N_10995);
and U13475 (N_13475,N_11374,N_12111);
or U13476 (N_13476,N_10816,N_10658);
nor U13477 (N_13477,N_10079,N_12317);
and U13478 (N_13478,N_10611,N_12212);
nor U13479 (N_13479,N_11734,N_10471);
nor U13480 (N_13480,N_11272,N_10416);
or U13481 (N_13481,N_12054,N_10680);
nor U13482 (N_13482,N_10702,N_11450);
xnor U13483 (N_13483,N_12277,N_11549);
and U13484 (N_13484,N_11387,N_10436);
nand U13485 (N_13485,N_12245,N_10460);
nand U13486 (N_13486,N_11344,N_10526);
xor U13487 (N_13487,N_10519,N_12251);
and U13488 (N_13488,N_10477,N_11228);
nor U13489 (N_13489,N_11486,N_12435);
and U13490 (N_13490,N_10731,N_11456);
nand U13491 (N_13491,N_12059,N_11777);
and U13492 (N_13492,N_10423,N_11851);
xor U13493 (N_13493,N_10907,N_10084);
nor U13494 (N_13494,N_11322,N_10777);
nor U13495 (N_13495,N_11477,N_10499);
xor U13496 (N_13496,N_10495,N_11172);
and U13497 (N_13497,N_11724,N_10715);
nor U13498 (N_13498,N_10627,N_10506);
and U13499 (N_13499,N_12067,N_11421);
nor U13500 (N_13500,N_10851,N_11669);
nand U13501 (N_13501,N_12235,N_10370);
and U13502 (N_13502,N_10765,N_11348);
nor U13503 (N_13503,N_11491,N_11229);
nor U13504 (N_13504,N_10748,N_11723);
or U13505 (N_13505,N_11664,N_12275);
nand U13506 (N_13506,N_11258,N_11296);
or U13507 (N_13507,N_11120,N_12158);
nand U13508 (N_13508,N_10357,N_12366);
nor U13509 (N_13509,N_10741,N_11067);
nor U13510 (N_13510,N_12038,N_11956);
xor U13511 (N_13511,N_11445,N_11586);
or U13512 (N_13512,N_12479,N_11695);
xnor U13513 (N_13513,N_10803,N_10923);
nand U13514 (N_13514,N_10415,N_10280);
nand U13515 (N_13515,N_11717,N_10628);
nand U13516 (N_13516,N_10961,N_11816);
and U13517 (N_13517,N_10300,N_10270);
nor U13518 (N_13518,N_10642,N_11937);
and U13519 (N_13519,N_10854,N_11018);
xnor U13520 (N_13520,N_10834,N_10242);
or U13521 (N_13521,N_11012,N_10559);
nor U13522 (N_13522,N_12178,N_12222);
xor U13523 (N_13523,N_11558,N_10492);
xor U13524 (N_13524,N_10874,N_11947);
nand U13525 (N_13525,N_10379,N_11523);
and U13526 (N_13526,N_12306,N_11887);
nor U13527 (N_13527,N_11642,N_10323);
and U13528 (N_13528,N_12126,N_11529);
xnor U13529 (N_13529,N_10013,N_10551);
and U13530 (N_13530,N_12064,N_11542);
nand U13531 (N_13531,N_10948,N_10841);
xnor U13532 (N_13532,N_11712,N_11966);
and U13533 (N_13533,N_10550,N_10664);
nand U13534 (N_13534,N_11198,N_11812);
nor U13535 (N_13535,N_12016,N_11124);
nand U13536 (N_13536,N_12101,N_10896);
or U13537 (N_13537,N_10597,N_12416);
xor U13538 (N_13538,N_10102,N_11413);
nand U13539 (N_13539,N_10779,N_12469);
nor U13540 (N_13540,N_11955,N_10428);
xor U13541 (N_13541,N_11339,N_10634);
and U13542 (N_13542,N_10314,N_11802);
xor U13543 (N_13543,N_11059,N_10639);
and U13544 (N_13544,N_12162,N_10696);
nor U13545 (N_13545,N_12459,N_12014);
or U13546 (N_13546,N_11359,N_11042);
or U13547 (N_13547,N_11579,N_11482);
or U13548 (N_13548,N_10136,N_10997);
nand U13549 (N_13549,N_12055,N_10533);
and U13550 (N_13550,N_11585,N_12439);
or U13551 (N_13551,N_10427,N_10449);
nor U13552 (N_13552,N_10277,N_10889);
and U13553 (N_13553,N_10864,N_11470);
or U13554 (N_13554,N_11735,N_10111);
xnor U13555 (N_13555,N_11756,N_12001);
and U13556 (N_13556,N_12432,N_11897);
nand U13557 (N_13557,N_10570,N_11020);
and U13558 (N_13558,N_11202,N_11234);
xor U13559 (N_13559,N_12239,N_11567);
xnor U13560 (N_13560,N_10646,N_12322);
xnor U13561 (N_13561,N_12186,N_10328);
or U13562 (N_13562,N_10577,N_10601);
nor U13563 (N_13563,N_11110,N_10238);
xnor U13564 (N_13564,N_12408,N_10128);
xnor U13565 (N_13565,N_10939,N_12319);
xnor U13566 (N_13566,N_11390,N_10964);
nand U13567 (N_13567,N_10190,N_10672);
xnor U13568 (N_13568,N_11098,N_10373);
nor U13569 (N_13569,N_11259,N_10830);
and U13570 (N_13570,N_12262,N_12461);
and U13571 (N_13571,N_10118,N_11391);
xor U13572 (N_13572,N_12410,N_10592);
and U13573 (N_13573,N_11422,N_11645);
nand U13574 (N_13574,N_10162,N_10230);
or U13575 (N_13575,N_10877,N_11535);
and U13576 (N_13576,N_11287,N_11337);
xor U13577 (N_13577,N_11846,N_10464);
nor U13578 (N_13578,N_11448,N_11745);
nand U13579 (N_13579,N_11865,N_11977);
xor U13580 (N_13580,N_10808,N_11094);
nand U13581 (N_13581,N_12452,N_10386);
nand U13582 (N_13582,N_10367,N_11303);
nand U13583 (N_13583,N_10490,N_12030);
or U13584 (N_13584,N_11469,N_11388);
xnor U13585 (N_13585,N_10651,N_11242);
xnor U13586 (N_13586,N_12287,N_10245);
nor U13587 (N_13587,N_10281,N_12018);
or U13588 (N_13588,N_11050,N_12462);
xnor U13589 (N_13589,N_11155,N_10572);
or U13590 (N_13590,N_10771,N_10348);
nor U13591 (N_13591,N_12269,N_11488);
nand U13592 (N_13592,N_12248,N_11183);
xor U13593 (N_13593,N_10456,N_11644);
or U13594 (N_13594,N_10514,N_12156);
nor U13595 (N_13595,N_12082,N_10637);
or U13596 (N_13596,N_11338,N_10790);
nand U13597 (N_13597,N_11744,N_10776);
or U13598 (N_13598,N_11522,N_10911);
xor U13599 (N_13599,N_11949,N_11502);
xor U13600 (N_13600,N_10404,N_11708);
and U13601 (N_13601,N_10161,N_11706);
xnor U13602 (N_13602,N_10973,N_11074);
nand U13603 (N_13603,N_10433,N_10721);
or U13604 (N_13604,N_11122,N_11513);
nand U13605 (N_13605,N_12129,N_11801);
or U13606 (N_13606,N_10026,N_11517);
and U13607 (N_13607,N_11814,N_10562);
nand U13608 (N_13608,N_12463,N_10381);
nor U13609 (N_13609,N_12201,N_12488);
nand U13610 (N_13610,N_11090,N_11206);
nor U13611 (N_13611,N_12391,N_11566);
nor U13612 (N_13612,N_12355,N_11026);
nand U13613 (N_13613,N_10430,N_10858);
nor U13614 (N_13614,N_10167,N_12182);
nor U13615 (N_13615,N_11004,N_11738);
xor U13616 (N_13616,N_10768,N_11934);
or U13617 (N_13617,N_11972,N_10204);
nor U13618 (N_13618,N_12304,N_11917);
nand U13619 (N_13619,N_10003,N_12281);
nand U13620 (N_13620,N_12276,N_10737);
nor U13621 (N_13621,N_12043,N_10804);
nor U13622 (N_13622,N_11160,N_10296);
and U13623 (N_13623,N_11684,N_10951);
nand U13624 (N_13624,N_10073,N_11213);
and U13625 (N_13625,N_10842,N_10669);
nor U13626 (N_13626,N_11184,N_12253);
nor U13627 (N_13627,N_10081,N_11905);
and U13628 (N_13628,N_11638,N_12108);
and U13629 (N_13629,N_10174,N_12167);
xnor U13630 (N_13630,N_10439,N_11835);
nand U13631 (N_13631,N_11646,N_12096);
and U13632 (N_13632,N_12149,N_10800);
nor U13633 (N_13633,N_11618,N_11361);
xor U13634 (N_13634,N_12184,N_12333);
nand U13635 (N_13635,N_10425,N_10599);
nand U13636 (N_13636,N_10065,N_12195);
or U13637 (N_13637,N_11551,N_11466);
xnor U13638 (N_13638,N_12341,N_10447);
nor U13639 (N_13639,N_10992,N_10030);
xnor U13640 (N_13640,N_12345,N_11702);
and U13641 (N_13641,N_12458,N_12081);
xor U13642 (N_13642,N_10232,N_11319);
nor U13643 (N_13643,N_10985,N_10770);
and U13644 (N_13644,N_12168,N_12314);
nor U13645 (N_13645,N_11416,N_10359);
or U13646 (N_13646,N_10897,N_11980);
and U13647 (N_13647,N_11612,N_10344);
nand U13648 (N_13648,N_12498,N_10086);
xor U13649 (N_13649,N_12376,N_10618);
xnor U13650 (N_13650,N_10224,N_12181);
or U13651 (N_13651,N_11981,N_12329);
and U13652 (N_13652,N_11750,N_10260);
or U13653 (N_13653,N_11908,N_11079);
nand U13654 (N_13654,N_12091,N_11378);
nand U13655 (N_13655,N_10478,N_12478);
xnor U13656 (N_13656,N_11941,N_11875);
xnor U13657 (N_13657,N_11976,N_10727);
or U13658 (N_13658,N_11249,N_10020);
xnor U13659 (N_13659,N_10832,N_11005);
xor U13660 (N_13660,N_10151,N_10446);
xnor U13661 (N_13661,N_11895,N_11085);
and U13662 (N_13662,N_10234,N_12083);
or U13663 (N_13663,N_12198,N_10265);
and U13664 (N_13664,N_11453,N_11194);
xor U13665 (N_13665,N_10139,N_12268);
xor U13666 (N_13666,N_12456,N_11804);
nand U13667 (N_13667,N_10773,N_11906);
xor U13668 (N_13668,N_12437,N_10908);
nor U13669 (N_13669,N_12002,N_10087);
or U13670 (N_13670,N_11962,N_10556);
nand U13671 (N_13671,N_11248,N_12485);
nor U13672 (N_13672,N_12430,N_11993);
or U13673 (N_13673,N_11590,N_10511);
nor U13674 (N_13674,N_11086,N_10681);
and U13675 (N_13675,N_10039,N_10220);
nand U13676 (N_13676,N_11637,N_10736);
nor U13677 (N_13677,N_12290,N_12169);
nand U13678 (N_13678,N_11929,N_12062);
xor U13679 (N_13679,N_10888,N_11282);
or U13680 (N_13680,N_11893,N_10924);
and U13681 (N_13681,N_10380,N_10856);
and U13682 (N_13682,N_12308,N_10360);
and U13683 (N_13683,N_11341,N_10643);
xor U13684 (N_13684,N_11758,N_11159);
or U13685 (N_13685,N_11842,N_10090);
xor U13686 (N_13686,N_10653,N_11616);
nand U13687 (N_13687,N_11463,N_11267);
and U13688 (N_13688,N_12388,N_10730);
nand U13689 (N_13689,N_10332,N_11483);
or U13690 (N_13690,N_10835,N_11656);
and U13691 (N_13691,N_11370,N_10390);
xnor U13692 (N_13692,N_10738,N_10002);
xnor U13693 (N_13693,N_11168,N_12234);
nor U13694 (N_13694,N_11856,N_12229);
nand U13695 (N_13695,N_10608,N_11635);
nand U13696 (N_13696,N_11658,N_12344);
nand U13697 (N_13697,N_10796,N_11123);
and U13698 (N_13698,N_12047,N_10613);
nor U13699 (N_13699,N_11991,N_11320);
nand U13700 (N_13700,N_12012,N_11639);
and U13701 (N_13701,N_12027,N_10752);
and U13702 (N_13702,N_10159,N_11709);
nor U13703 (N_13703,N_11828,N_11405);
xnor U13704 (N_13704,N_11077,N_10318);
nand U13705 (N_13705,N_10112,N_10229);
nor U13706 (N_13706,N_11543,N_12106);
xor U13707 (N_13707,N_12133,N_11057);
and U13708 (N_13708,N_11101,N_10636);
xor U13709 (N_13709,N_11891,N_10621);
xor U13710 (N_13710,N_11680,N_10958);
nor U13711 (N_13711,N_11753,N_10616);
and U13712 (N_13712,N_11915,N_11372);
and U13713 (N_13713,N_10547,N_10824);
nor U13714 (N_13714,N_11643,N_10978);
and U13715 (N_13715,N_10763,N_12499);
nand U13716 (N_13716,N_10400,N_11128);
xor U13717 (N_13717,N_11752,N_10023);
nor U13718 (N_13718,N_10153,N_11970);
xnor U13719 (N_13719,N_11088,N_11136);
nand U13720 (N_13720,N_12296,N_11479);
xor U13721 (N_13721,N_11189,N_12259);
and U13722 (N_13722,N_12119,N_11239);
nand U13723 (N_13723,N_10243,N_11141);
or U13724 (N_13724,N_12011,N_12272);
nand U13725 (N_13725,N_10398,N_12155);
nand U13726 (N_13726,N_11850,N_12148);
nand U13727 (N_13727,N_10126,N_11904);
xnor U13728 (N_13728,N_11759,N_10369);
nor U13729 (N_13729,N_11187,N_11254);
or U13730 (N_13730,N_11297,N_11541);
and U13731 (N_13731,N_10654,N_10377);
nand U13732 (N_13732,N_11903,N_12367);
nor U13733 (N_13733,N_10027,N_10848);
nand U13734 (N_13734,N_11928,N_10815);
nand U13735 (N_13735,N_10124,N_11161);
and U13736 (N_13736,N_10099,N_10760);
nand U13737 (N_13737,N_11653,N_10674);
nor U13738 (N_13738,N_10758,N_11379);
or U13739 (N_13739,N_10004,N_10742);
xnor U13740 (N_13740,N_10142,N_10792);
xnor U13741 (N_13741,N_12040,N_10342);
nor U13742 (N_13742,N_11100,N_10261);
xor U13743 (N_13743,N_10031,N_11518);
nor U13744 (N_13744,N_11614,N_10411);
nor U13745 (N_13745,N_10753,N_10965);
nand U13746 (N_13746,N_10156,N_10905);
or U13747 (N_13747,N_11336,N_11021);
and U13748 (N_13748,N_10886,N_12299);
and U13749 (N_13749,N_10638,N_12161);
and U13750 (N_13750,N_10112,N_10893);
nand U13751 (N_13751,N_10697,N_11059);
nor U13752 (N_13752,N_12202,N_12499);
and U13753 (N_13753,N_12070,N_12379);
xor U13754 (N_13754,N_10671,N_11274);
or U13755 (N_13755,N_11574,N_12279);
xnor U13756 (N_13756,N_12331,N_12036);
xnor U13757 (N_13757,N_12101,N_11961);
nand U13758 (N_13758,N_12365,N_10503);
or U13759 (N_13759,N_10453,N_11864);
or U13760 (N_13760,N_12275,N_10107);
or U13761 (N_13761,N_11597,N_11520);
xnor U13762 (N_13762,N_10533,N_11433);
nor U13763 (N_13763,N_11625,N_11622);
nor U13764 (N_13764,N_10582,N_11500);
nor U13765 (N_13765,N_10086,N_10858);
nand U13766 (N_13766,N_11172,N_12301);
nor U13767 (N_13767,N_10658,N_10042);
nand U13768 (N_13768,N_10802,N_10704);
xor U13769 (N_13769,N_10798,N_11855);
xnor U13770 (N_13770,N_11819,N_11378);
and U13771 (N_13771,N_10977,N_10499);
xor U13772 (N_13772,N_11474,N_12172);
nor U13773 (N_13773,N_12395,N_12449);
xor U13774 (N_13774,N_10971,N_12458);
and U13775 (N_13775,N_11605,N_10159);
nor U13776 (N_13776,N_10004,N_10613);
xnor U13777 (N_13777,N_10732,N_10671);
nor U13778 (N_13778,N_10581,N_11010);
and U13779 (N_13779,N_10238,N_10255);
xor U13780 (N_13780,N_10223,N_10396);
nor U13781 (N_13781,N_10775,N_10552);
or U13782 (N_13782,N_11178,N_10119);
or U13783 (N_13783,N_10755,N_10329);
and U13784 (N_13784,N_12032,N_12349);
xor U13785 (N_13785,N_11611,N_11860);
and U13786 (N_13786,N_10118,N_10591);
nor U13787 (N_13787,N_10992,N_11306);
xor U13788 (N_13788,N_10419,N_11803);
and U13789 (N_13789,N_10156,N_12377);
and U13790 (N_13790,N_11281,N_12012);
and U13791 (N_13791,N_11237,N_10911);
nor U13792 (N_13792,N_11146,N_12119);
and U13793 (N_13793,N_10329,N_11945);
nand U13794 (N_13794,N_10696,N_10389);
xnor U13795 (N_13795,N_11374,N_12435);
nor U13796 (N_13796,N_12309,N_12255);
or U13797 (N_13797,N_11081,N_10285);
and U13798 (N_13798,N_10047,N_11042);
and U13799 (N_13799,N_12375,N_10416);
and U13800 (N_13800,N_10452,N_10643);
or U13801 (N_13801,N_12414,N_10093);
and U13802 (N_13802,N_10317,N_10347);
nor U13803 (N_13803,N_11952,N_10108);
xnor U13804 (N_13804,N_10284,N_11637);
xor U13805 (N_13805,N_11073,N_11530);
and U13806 (N_13806,N_10902,N_12137);
and U13807 (N_13807,N_11270,N_10025);
nor U13808 (N_13808,N_10974,N_11568);
and U13809 (N_13809,N_11255,N_10857);
or U13810 (N_13810,N_11019,N_11463);
xnor U13811 (N_13811,N_11735,N_10517);
xnor U13812 (N_13812,N_10963,N_12487);
or U13813 (N_13813,N_11044,N_10836);
xor U13814 (N_13814,N_10093,N_11153);
or U13815 (N_13815,N_11459,N_12328);
or U13816 (N_13816,N_10118,N_11437);
and U13817 (N_13817,N_11173,N_10230);
or U13818 (N_13818,N_11300,N_11696);
nand U13819 (N_13819,N_11063,N_10148);
or U13820 (N_13820,N_12407,N_11028);
nor U13821 (N_13821,N_12347,N_12243);
xnor U13822 (N_13822,N_11798,N_10371);
nor U13823 (N_13823,N_11176,N_11949);
or U13824 (N_13824,N_10921,N_10932);
nand U13825 (N_13825,N_12216,N_10897);
nand U13826 (N_13826,N_10086,N_11359);
or U13827 (N_13827,N_12230,N_11049);
and U13828 (N_13828,N_10194,N_11560);
or U13829 (N_13829,N_11694,N_10739);
xnor U13830 (N_13830,N_10157,N_10324);
nor U13831 (N_13831,N_10178,N_11430);
xor U13832 (N_13832,N_10183,N_12009);
nand U13833 (N_13833,N_12065,N_12252);
nor U13834 (N_13834,N_10016,N_10480);
nand U13835 (N_13835,N_10469,N_11694);
nor U13836 (N_13836,N_10841,N_12387);
nand U13837 (N_13837,N_12105,N_11071);
xnor U13838 (N_13838,N_11974,N_11470);
nor U13839 (N_13839,N_10985,N_11832);
nand U13840 (N_13840,N_11811,N_11093);
xor U13841 (N_13841,N_10904,N_11734);
xor U13842 (N_13842,N_11186,N_12259);
xnor U13843 (N_13843,N_10973,N_11003);
or U13844 (N_13844,N_12325,N_10193);
xnor U13845 (N_13845,N_11206,N_12323);
xnor U13846 (N_13846,N_11205,N_11395);
or U13847 (N_13847,N_10290,N_10118);
xnor U13848 (N_13848,N_11867,N_11647);
or U13849 (N_13849,N_12380,N_11862);
nand U13850 (N_13850,N_11687,N_10582);
and U13851 (N_13851,N_10996,N_11460);
or U13852 (N_13852,N_11027,N_11398);
or U13853 (N_13853,N_10352,N_11719);
and U13854 (N_13854,N_10570,N_12156);
or U13855 (N_13855,N_12162,N_10216);
nand U13856 (N_13856,N_11673,N_11970);
nor U13857 (N_13857,N_10029,N_12139);
or U13858 (N_13858,N_10502,N_12194);
nand U13859 (N_13859,N_10896,N_11179);
nor U13860 (N_13860,N_12431,N_12130);
nor U13861 (N_13861,N_11370,N_11865);
xnor U13862 (N_13862,N_10965,N_11287);
and U13863 (N_13863,N_11965,N_11613);
or U13864 (N_13864,N_10681,N_11222);
or U13865 (N_13865,N_11525,N_11575);
or U13866 (N_13866,N_12415,N_11780);
xor U13867 (N_13867,N_11804,N_12140);
xnor U13868 (N_13868,N_11699,N_11369);
or U13869 (N_13869,N_11714,N_11544);
xnor U13870 (N_13870,N_10357,N_12177);
and U13871 (N_13871,N_11036,N_11354);
nand U13872 (N_13872,N_10808,N_12389);
or U13873 (N_13873,N_12102,N_10199);
xor U13874 (N_13874,N_11482,N_11266);
and U13875 (N_13875,N_12052,N_10311);
xor U13876 (N_13876,N_10745,N_12064);
and U13877 (N_13877,N_10156,N_12056);
and U13878 (N_13878,N_11112,N_12129);
nor U13879 (N_13879,N_11004,N_10255);
nor U13880 (N_13880,N_11725,N_11406);
or U13881 (N_13881,N_11970,N_10145);
or U13882 (N_13882,N_11449,N_10124);
nand U13883 (N_13883,N_12098,N_11965);
and U13884 (N_13884,N_10471,N_12193);
and U13885 (N_13885,N_10499,N_10315);
nor U13886 (N_13886,N_11494,N_11986);
xor U13887 (N_13887,N_10117,N_12089);
or U13888 (N_13888,N_11523,N_11231);
and U13889 (N_13889,N_10719,N_11822);
nor U13890 (N_13890,N_10004,N_11150);
or U13891 (N_13891,N_10128,N_11550);
and U13892 (N_13892,N_11990,N_12107);
nand U13893 (N_13893,N_10874,N_11008);
or U13894 (N_13894,N_11155,N_11671);
or U13895 (N_13895,N_10586,N_11680);
nor U13896 (N_13896,N_11495,N_11061);
nor U13897 (N_13897,N_11766,N_10462);
or U13898 (N_13898,N_10492,N_11663);
xnor U13899 (N_13899,N_11078,N_10986);
nand U13900 (N_13900,N_10619,N_10411);
and U13901 (N_13901,N_10839,N_10004);
nand U13902 (N_13902,N_10331,N_11536);
nand U13903 (N_13903,N_10115,N_12444);
and U13904 (N_13904,N_12133,N_12044);
nand U13905 (N_13905,N_10436,N_12115);
and U13906 (N_13906,N_10744,N_11288);
or U13907 (N_13907,N_11788,N_11343);
nor U13908 (N_13908,N_10007,N_11830);
or U13909 (N_13909,N_11364,N_10381);
and U13910 (N_13910,N_12171,N_10430);
xor U13911 (N_13911,N_11257,N_11544);
nand U13912 (N_13912,N_11595,N_10827);
nor U13913 (N_13913,N_11852,N_11762);
xnor U13914 (N_13914,N_12470,N_10761);
nand U13915 (N_13915,N_12451,N_10274);
xor U13916 (N_13916,N_11892,N_11294);
or U13917 (N_13917,N_10528,N_10481);
and U13918 (N_13918,N_10554,N_12352);
nand U13919 (N_13919,N_10021,N_10580);
xor U13920 (N_13920,N_10060,N_11838);
nor U13921 (N_13921,N_11782,N_10664);
nand U13922 (N_13922,N_12113,N_10772);
nor U13923 (N_13923,N_11270,N_10832);
or U13924 (N_13924,N_11309,N_11510);
nor U13925 (N_13925,N_12459,N_12095);
and U13926 (N_13926,N_10431,N_12462);
nand U13927 (N_13927,N_10257,N_10869);
or U13928 (N_13928,N_11519,N_10005);
xnor U13929 (N_13929,N_11130,N_12279);
nor U13930 (N_13930,N_10837,N_10069);
or U13931 (N_13931,N_11154,N_11639);
xnor U13932 (N_13932,N_10108,N_11560);
xnor U13933 (N_13933,N_10364,N_10110);
nand U13934 (N_13934,N_11427,N_10000);
nand U13935 (N_13935,N_10782,N_11202);
nor U13936 (N_13936,N_12158,N_11727);
and U13937 (N_13937,N_11564,N_12332);
nand U13938 (N_13938,N_10202,N_12436);
nor U13939 (N_13939,N_11891,N_10394);
and U13940 (N_13940,N_10381,N_12292);
xnor U13941 (N_13941,N_11650,N_10614);
nand U13942 (N_13942,N_12429,N_11172);
xor U13943 (N_13943,N_12185,N_11996);
or U13944 (N_13944,N_12401,N_11161);
and U13945 (N_13945,N_11072,N_10011);
and U13946 (N_13946,N_10692,N_11533);
xnor U13947 (N_13947,N_10729,N_11270);
and U13948 (N_13948,N_11814,N_12069);
nor U13949 (N_13949,N_11796,N_11684);
nand U13950 (N_13950,N_11238,N_11631);
nand U13951 (N_13951,N_10396,N_11975);
or U13952 (N_13952,N_10614,N_12357);
or U13953 (N_13953,N_11459,N_12181);
and U13954 (N_13954,N_11424,N_12453);
nor U13955 (N_13955,N_12119,N_10436);
nand U13956 (N_13956,N_12365,N_11627);
and U13957 (N_13957,N_10173,N_10774);
and U13958 (N_13958,N_12402,N_10180);
nor U13959 (N_13959,N_11701,N_12195);
nor U13960 (N_13960,N_11497,N_11413);
xor U13961 (N_13961,N_10359,N_12084);
and U13962 (N_13962,N_10059,N_11739);
xnor U13963 (N_13963,N_11590,N_12207);
and U13964 (N_13964,N_10944,N_12074);
nand U13965 (N_13965,N_10695,N_10564);
and U13966 (N_13966,N_10901,N_11414);
nor U13967 (N_13967,N_10781,N_11647);
nor U13968 (N_13968,N_11538,N_12105);
or U13969 (N_13969,N_12379,N_12095);
xor U13970 (N_13970,N_12034,N_12338);
nand U13971 (N_13971,N_10337,N_10987);
and U13972 (N_13972,N_10463,N_12091);
nor U13973 (N_13973,N_11098,N_10157);
nand U13974 (N_13974,N_11851,N_12341);
nand U13975 (N_13975,N_10710,N_10905);
nand U13976 (N_13976,N_11050,N_12238);
or U13977 (N_13977,N_10180,N_10235);
nor U13978 (N_13978,N_12178,N_12302);
nor U13979 (N_13979,N_10708,N_10351);
and U13980 (N_13980,N_11566,N_12496);
nand U13981 (N_13981,N_11201,N_11048);
nand U13982 (N_13982,N_11902,N_12154);
nor U13983 (N_13983,N_11934,N_11069);
nand U13984 (N_13984,N_12003,N_11215);
and U13985 (N_13985,N_10521,N_11801);
and U13986 (N_13986,N_10394,N_11493);
nand U13987 (N_13987,N_11109,N_11517);
or U13988 (N_13988,N_11594,N_10576);
and U13989 (N_13989,N_11458,N_10995);
and U13990 (N_13990,N_10103,N_10065);
xor U13991 (N_13991,N_11541,N_12080);
and U13992 (N_13992,N_10860,N_10805);
and U13993 (N_13993,N_10258,N_12490);
xnor U13994 (N_13994,N_12062,N_11973);
and U13995 (N_13995,N_10582,N_10779);
nor U13996 (N_13996,N_10558,N_11573);
and U13997 (N_13997,N_11453,N_10483);
nand U13998 (N_13998,N_12034,N_10582);
and U13999 (N_13999,N_11790,N_12202);
or U14000 (N_14000,N_11783,N_10248);
nand U14001 (N_14001,N_10475,N_10319);
xor U14002 (N_14002,N_11345,N_12280);
xor U14003 (N_14003,N_11028,N_10056);
nand U14004 (N_14004,N_10570,N_11944);
and U14005 (N_14005,N_10460,N_11242);
and U14006 (N_14006,N_11774,N_10763);
nor U14007 (N_14007,N_12218,N_12135);
nand U14008 (N_14008,N_11490,N_11427);
and U14009 (N_14009,N_10013,N_10626);
nand U14010 (N_14010,N_11578,N_12087);
nand U14011 (N_14011,N_11029,N_10671);
nor U14012 (N_14012,N_10498,N_11671);
and U14013 (N_14013,N_10876,N_10444);
xor U14014 (N_14014,N_10389,N_11492);
or U14015 (N_14015,N_12497,N_11252);
or U14016 (N_14016,N_10000,N_11068);
nand U14017 (N_14017,N_10049,N_11919);
nor U14018 (N_14018,N_12461,N_12090);
nor U14019 (N_14019,N_10546,N_12321);
nor U14020 (N_14020,N_12394,N_11263);
or U14021 (N_14021,N_11019,N_10000);
and U14022 (N_14022,N_12459,N_11610);
or U14023 (N_14023,N_11235,N_11751);
or U14024 (N_14024,N_10996,N_10066);
or U14025 (N_14025,N_10080,N_10317);
xor U14026 (N_14026,N_10161,N_12270);
nand U14027 (N_14027,N_11715,N_10132);
xnor U14028 (N_14028,N_11736,N_12169);
nand U14029 (N_14029,N_10372,N_11323);
nand U14030 (N_14030,N_10981,N_10493);
nor U14031 (N_14031,N_12032,N_10472);
or U14032 (N_14032,N_11167,N_10768);
xor U14033 (N_14033,N_11993,N_10253);
and U14034 (N_14034,N_12412,N_10726);
and U14035 (N_14035,N_11101,N_12119);
nor U14036 (N_14036,N_12397,N_11734);
or U14037 (N_14037,N_11793,N_10604);
xor U14038 (N_14038,N_10235,N_11928);
nand U14039 (N_14039,N_10079,N_11061);
xor U14040 (N_14040,N_11194,N_12040);
nand U14041 (N_14041,N_11106,N_11450);
xor U14042 (N_14042,N_10339,N_10688);
nand U14043 (N_14043,N_11194,N_10699);
nor U14044 (N_14044,N_10005,N_11283);
nor U14045 (N_14045,N_11121,N_11751);
and U14046 (N_14046,N_12280,N_11778);
nand U14047 (N_14047,N_11315,N_12061);
nor U14048 (N_14048,N_10630,N_11190);
nand U14049 (N_14049,N_12208,N_12021);
nand U14050 (N_14050,N_12275,N_10373);
or U14051 (N_14051,N_10432,N_11298);
nand U14052 (N_14052,N_10679,N_10091);
or U14053 (N_14053,N_10628,N_11103);
and U14054 (N_14054,N_10761,N_11940);
xnor U14055 (N_14055,N_10685,N_12042);
nand U14056 (N_14056,N_12462,N_10689);
or U14057 (N_14057,N_12466,N_12303);
or U14058 (N_14058,N_10363,N_12304);
xnor U14059 (N_14059,N_12429,N_12462);
or U14060 (N_14060,N_11151,N_11111);
xnor U14061 (N_14061,N_12447,N_12392);
or U14062 (N_14062,N_11072,N_10682);
and U14063 (N_14063,N_10428,N_11194);
xnor U14064 (N_14064,N_10513,N_10218);
nand U14065 (N_14065,N_11364,N_10121);
and U14066 (N_14066,N_11412,N_11186);
and U14067 (N_14067,N_11763,N_11797);
and U14068 (N_14068,N_10778,N_10265);
xor U14069 (N_14069,N_10884,N_10026);
and U14070 (N_14070,N_12489,N_10616);
xnor U14071 (N_14071,N_10542,N_10259);
or U14072 (N_14072,N_11947,N_11268);
xor U14073 (N_14073,N_12482,N_11871);
xnor U14074 (N_14074,N_11004,N_10836);
nor U14075 (N_14075,N_10347,N_10172);
nor U14076 (N_14076,N_10883,N_12011);
nor U14077 (N_14077,N_10493,N_10343);
nand U14078 (N_14078,N_10320,N_11838);
xnor U14079 (N_14079,N_11269,N_12017);
nor U14080 (N_14080,N_11624,N_11831);
or U14081 (N_14081,N_10238,N_10684);
or U14082 (N_14082,N_11189,N_10521);
nand U14083 (N_14083,N_11613,N_12068);
xor U14084 (N_14084,N_11239,N_10428);
nor U14085 (N_14085,N_10037,N_10481);
or U14086 (N_14086,N_10032,N_10212);
xor U14087 (N_14087,N_11454,N_12244);
or U14088 (N_14088,N_10651,N_10577);
and U14089 (N_14089,N_10262,N_12323);
nand U14090 (N_14090,N_11155,N_12075);
xor U14091 (N_14091,N_11211,N_11405);
and U14092 (N_14092,N_10408,N_10926);
nand U14093 (N_14093,N_12179,N_10953);
or U14094 (N_14094,N_11780,N_11292);
and U14095 (N_14095,N_11648,N_12496);
xnor U14096 (N_14096,N_11803,N_11886);
xnor U14097 (N_14097,N_11342,N_11186);
nand U14098 (N_14098,N_10825,N_11210);
or U14099 (N_14099,N_11004,N_10403);
and U14100 (N_14100,N_12029,N_10991);
nor U14101 (N_14101,N_10487,N_11237);
and U14102 (N_14102,N_11295,N_11081);
or U14103 (N_14103,N_10077,N_10341);
and U14104 (N_14104,N_10427,N_12398);
nor U14105 (N_14105,N_12202,N_12177);
and U14106 (N_14106,N_10068,N_10098);
nor U14107 (N_14107,N_10784,N_12016);
nand U14108 (N_14108,N_11904,N_10894);
nand U14109 (N_14109,N_11712,N_11443);
nand U14110 (N_14110,N_11592,N_12094);
xor U14111 (N_14111,N_12260,N_12014);
or U14112 (N_14112,N_11950,N_11245);
nand U14113 (N_14113,N_10721,N_11958);
nand U14114 (N_14114,N_11571,N_11267);
xor U14115 (N_14115,N_11243,N_10679);
and U14116 (N_14116,N_10391,N_11666);
or U14117 (N_14117,N_10062,N_12321);
nand U14118 (N_14118,N_10536,N_11524);
or U14119 (N_14119,N_12243,N_11767);
and U14120 (N_14120,N_10425,N_12222);
and U14121 (N_14121,N_12380,N_10943);
xor U14122 (N_14122,N_11352,N_11800);
xnor U14123 (N_14123,N_10264,N_10717);
nand U14124 (N_14124,N_12422,N_11391);
nand U14125 (N_14125,N_10725,N_12231);
nand U14126 (N_14126,N_11692,N_10438);
nor U14127 (N_14127,N_11350,N_10805);
nand U14128 (N_14128,N_12416,N_12473);
and U14129 (N_14129,N_11135,N_10479);
nor U14130 (N_14130,N_11533,N_11325);
and U14131 (N_14131,N_12270,N_10585);
and U14132 (N_14132,N_11267,N_10754);
nand U14133 (N_14133,N_11188,N_12390);
nand U14134 (N_14134,N_10555,N_12070);
nand U14135 (N_14135,N_10534,N_10684);
nor U14136 (N_14136,N_10699,N_10143);
or U14137 (N_14137,N_10420,N_10135);
nor U14138 (N_14138,N_10688,N_11870);
nor U14139 (N_14139,N_11838,N_10407);
nor U14140 (N_14140,N_10411,N_12166);
nor U14141 (N_14141,N_11300,N_10641);
nand U14142 (N_14142,N_11244,N_11106);
or U14143 (N_14143,N_11973,N_10769);
and U14144 (N_14144,N_12037,N_12183);
nor U14145 (N_14145,N_12338,N_12026);
nor U14146 (N_14146,N_10366,N_10670);
or U14147 (N_14147,N_11682,N_10048);
nor U14148 (N_14148,N_12495,N_10052);
or U14149 (N_14149,N_12486,N_12442);
and U14150 (N_14150,N_11515,N_10581);
or U14151 (N_14151,N_11178,N_10914);
and U14152 (N_14152,N_10660,N_10878);
nor U14153 (N_14153,N_11215,N_11672);
xor U14154 (N_14154,N_10708,N_10094);
nor U14155 (N_14155,N_11136,N_10247);
and U14156 (N_14156,N_11561,N_11259);
or U14157 (N_14157,N_10905,N_11226);
xor U14158 (N_14158,N_11548,N_12486);
xnor U14159 (N_14159,N_12441,N_10441);
xor U14160 (N_14160,N_11689,N_12228);
nand U14161 (N_14161,N_10981,N_11455);
and U14162 (N_14162,N_10043,N_10706);
xor U14163 (N_14163,N_12020,N_11639);
xnor U14164 (N_14164,N_11838,N_10489);
or U14165 (N_14165,N_10992,N_11309);
xnor U14166 (N_14166,N_10989,N_10626);
or U14167 (N_14167,N_11366,N_11008);
or U14168 (N_14168,N_10567,N_12416);
nand U14169 (N_14169,N_10002,N_10313);
nor U14170 (N_14170,N_11516,N_12460);
nor U14171 (N_14171,N_10488,N_11737);
nor U14172 (N_14172,N_11298,N_12246);
nor U14173 (N_14173,N_10073,N_12020);
nand U14174 (N_14174,N_11482,N_10502);
and U14175 (N_14175,N_10275,N_10517);
and U14176 (N_14176,N_10447,N_10879);
nor U14177 (N_14177,N_10392,N_11476);
nand U14178 (N_14178,N_10134,N_10219);
xnor U14179 (N_14179,N_11406,N_11224);
or U14180 (N_14180,N_12161,N_12219);
nor U14181 (N_14181,N_10594,N_11263);
and U14182 (N_14182,N_10091,N_10235);
and U14183 (N_14183,N_12148,N_10554);
and U14184 (N_14184,N_10324,N_10665);
xor U14185 (N_14185,N_10369,N_12411);
xor U14186 (N_14186,N_12495,N_10297);
xnor U14187 (N_14187,N_11468,N_12446);
and U14188 (N_14188,N_11852,N_10353);
or U14189 (N_14189,N_11755,N_11889);
nand U14190 (N_14190,N_11968,N_12288);
or U14191 (N_14191,N_12198,N_11466);
nand U14192 (N_14192,N_10863,N_11018);
and U14193 (N_14193,N_11864,N_10029);
nor U14194 (N_14194,N_12024,N_12311);
and U14195 (N_14195,N_12044,N_11599);
nand U14196 (N_14196,N_10356,N_12418);
or U14197 (N_14197,N_11269,N_10792);
or U14198 (N_14198,N_11023,N_10890);
nand U14199 (N_14199,N_10534,N_12454);
nor U14200 (N_14200,N_12276,N_12282);
and U14201 (N_14201,N_11618,N_11839);
and U14202 (N_14202,N_12029,N_11678);
nor U14203 (N_14203,N_10271,N_12126);
nand U14204 (N_14204,N_11655,N_10251);
and U14205 (N_14205,N_11527,N_10934);
nand U14206 (N_14206,N_11163,N_12269);
nand U14207 (N_14207,N_10526,N_12139);
nand U14208 (N_14208,N_11990,N_12015);
or U14209 (N_14209,N_11364,N_12471);
or U14210 (N_14210,N_11288,N_10251);
nor U14211 (N_14211,N_11856,N_12129);
nand U14212 (N_14212,N_10302,N_10570);
xnor U14213 (N_14213,N_10974,N_12447);
nor U14214 (N_14214,N_11700,N_10147);
or U14215 (N_14215,N_10441,N_11955);
nand U14216 (N_14216,N_11715,N_11518);
nor U14217 (N_14217,N_11849,N_10619);
nand U14218 (N_14218,N_11433,N_11003);
nor U14219 (N_14219,N_12434,N_10750);
nor U14220 (N_14220,N_10262,N_10375);
or U14221 (N_14221,N_10708,N_11715);
or U14222 (N_14222,N_11523,N_12194);
nand U14223 (N_14223,N_12003,N_10948);
nor U14224 (N_14224,N_11382,N_11183);
nor U14225 (N_14225,N_10773,N_11950);
nand U14226 (N_14226,N_11822,N_10382);
xnor U14227 (N_14227,N_10127,N_12447);
or U14228 (N_14228,N_11419,N_10193);
or U14229 (N_14229,N_11244,N_10721);
nand U14230 (N_14230,N_12480,N_11911);
nand U14231 (N_14231,N_12266,N_12022);
nand U14232 (N_14232,N_11826,N_11960);
nand U14233 (N_14233,N_12148,N_11135);
nand U14234 (N_14234,N_11704,N_10596);
nand U14235 (N_14235,N_11050,N_10747);
and U14236 (N_14236,N_11953,N_11464);
nor U14237 (N_14237,N_10966,N_11579);
and U14238 (N_14238,N_11702,N_11846);
xnor U14239 (N_14239,N_11129,N_12265);
xnor U14240 (N_14240,N_10226,N_11572);
nand U14241 (N_14241,N_11971,N_10806);
or U14242 (N_14242,N_11622,N_11708);
xnor U14243 (N_14243,N_10869,N_11869);
nor U14244 (N_14244,N_10776,N_11448);
nor U14245 (N_14245,N_11565,N_11610);
xnor U14246 (N_14246,N_11050,N_11153);
or U14247 (N_14247,N_12230,N_10866);
and U14248 (N_14248,N_10622,N_10653);
xnor U14249 (N_14249,N_11964,N_11050);
nand U14250 (N_14250,N_10500,N_10139);
or U14251 (N_14251,N_12310,N_11040);
or U14252 (N_14252,N_10398,N_11642);
and U14253 (N_14253,N_11572,N_10531);
nor U14254 (N_14254,N_11802,N_11081);
or U14255 (N_14255,N_11722,N_11200);
xnor U14256 (N_14256,N_10310,N_11310);
or U14257 (N_14257,N_11341,N_10970);
xnor U14258 (N_14258,N_10008,N_11693);
nor U14259 (N_14259,N_11059,N_11458);
xnor U14260 (N_14260,N_12474,N_12487);
nand U14261 (N_14261,N_11802,N_11666);
or U14262 (N_14262,N_10800,N_10258);
and U14263 (N_14263,N_11241,N_11532);
nand U14264 (N_14264,N_10544,N_10025);
xor U14265 (N_14265,N_10184,N_11475);
and U14266 (N_14266,N_11311,N_11457);
nor U14267 (N_14267,N_10641,N_10590);
nor U14268 (N_14268,N_11241,N_10489);
nand U14269 (N_14269,N_11495,N_12223);
or U14270 (N_14270,N_11005,N_12015);
xnor U14271 (N_14271,N_12168,N_10936);
and U14272 (N_14272,N_11142,N_10461);
or U14273 (N_14273,N_10782,N_11414);
nand U14274 (N_14274,N_10515,N_10556);
or U14275 (N_14275,N_12423,N_10587);
nand U14276 (N_14276,N_12241,N_11807);
nor U14277 (N_14277,N_10506,N_11929);
or U14278 (N_14278,N_11740,N_10783);
xnor U14279 (N_14279,N_11211,N_10955);
and U14280 (N_14280,N_11611,N_11614);
xor U14281 (N_14281,N_10834,N_12170);
and U14282 (N_14282,N_10655,N_10612);
xor U14283 (N_14283,N_11481,N_10499);
xor U14284 (N_14284,N_12320,N_11883);
or U14285 (N_14285,N_12253,N_10894);
or U14286 (N_14286,N_10102,N_10313);
and U14287 (N_14287,N_11452,N_11753);
and U14288 (N_14288,N_10813,N_12145);
xnor U14289 (N_14289,N_10457,N_12010);
and U14290 (N_14290,N_10778,N_11360);
nor U14291 (N_14291,N_11351,N_10820);
nor U14292 (N_14292,N_11146,N_11104);
or U14293 (N_14293,N_11923,N_10342);
xor U14294 (N_14294,N_10342,N_10411);
nand U14295 (N_14295,N_12464,N_11667);
xnor U14296 (N_14296,N_10522,N_10102);
nor U14297 (N_14297,N_11247,N_10719);
xnor U14298 (N_14298,N_11968,N_10664);
nor U14299 (N_14299,N_10101,N_12448);
nand U14300 (N_14300,N_10942,N_10581);
nand U14301 (N_14301,N_12339,N_10914);
and U14302 (N_14302,N_12383,N_11096);
xnor U14303 (N_14303,N_10343,N_12387);
or U14304 (N_14304,N_11084,N_12276);
xor U14305 (N_14305,N_11643,N_11326);
xnor U14306 (N_14306,N_10653,N_11770);
xor U14307 (N_14307,N_12082,N_10125);
xor U14308 (N_14308,N_10473,N_12476);
nand U14309 (N_14309,N_10764,N_12166);
nor U14310 (N_14310,N_10940,N_10462);
xnor U14311 (N_14311,N_11587,N_11438);
nor U14312 (N_14312,N_10073,N_10245);
or U14313 (N_14313,N_12299,N_11050);
or U14314 (N_14314,N_10141,N_12458);
and U14315 (N_14315,N_10197,N_11417);
and U14316 (N_14316,N_10650,N_10163);
xnor U14317 (N_14317,N_10130,N_11141);
and U14318 (N_14318,N_10568,N_10445);
nand U14319 (N_14319,N_10004,N_12107);
nor U14320 (N_14320,N_12053,N_10324);
nand U14321 (N_14321,N_11389,N_12111);
nor U14322 (N_14322,N_11154,N_10638);
xnor U14323 (N_14323,N_11505,N_11337);
and U14324 (N_14324,N_12171,N_10791);
and U14325 (N_14325,N_11233,N_11945);
nor U14326 (N_14326,N_10757,N_10493);
and U14327 (N_14327,N_11730,N_12194);
or U14328 (N_14328,N_12436,N_12340);
and U14329 (N_14329,N_10298,N_11354);
xor U14330 (N_14330,N_10006,N_10654);
nor U14331 (N_14331,N_10236,N_12060);
nand U14332 (N_14332,N_10518,N_12465);
and U14333 (N_14333,N_11502,N_10191);
nand U14334 (N_14334,N_10644,N_11771);
nand U14335 (N_14335,N_10750,N_11207);
and U14336 (N_14336,N_12193,N_11171);
and U14337 (N_14337,N_12410,N_11444);
and U14338 (N_14338,N_12430,N_11721);
nand U14339 (N_14339,N_12434,N_12392);
and U14340 (N_14340,N_12373,N_11902);
nand U14341 (N_14341,N_12193,N_11973);
or U14342 (N_14342,N_10291,N_11540);
or U14343 (N_14343,N_10088,N_11562);
xnor U14344 (N_14344,N_10619,N_11769);
nand U14345 (N_14345,N_10900,N_11576);
and U14346 (N_14346,N_10269,N_10288);
or U14347 (N_14347,N_11958,N_12304);
and U14348 (N_14348,N_10000,N_10720);
or U14349 (N_14349,N_12385,N_12168);
and U14350 (N_14350,N_11287,N_10599);
xnor U14351 (N_14351,N_10108,N_10208);
and U14352 (N_14352,N_10683,N_12060);
nor U14353 (N_14353,N_12042,N_12356);
or U14354 (N_14354,N_11244,N_10863);
or U14355 (N_14355,N_11758,N_12339);
or U14356 (N_14356,N_12421,N_11504);
nor U14357 (N_14357,N_12157,N_11138);
xor U14358 (N_14358,N_11468,N_12215);
xor U14359 (N_14359,N_10409,N_11117);
xor U14360 (N_14360,N_11982,N_11854);
xnor U14361 (N_14361,N_11234,N_11211);
or U14362 (N_14362,N_10421,N_11072);
and U14363 (N_14363,N_11673,N_11988);
xor U14364 (N_14364,N_10128,N_12413);
xor U14365 (N_14365,N_11541,N_12142);
nor U14366 (N_14366,N_12463,N_10057);
and U14367 (N_14367,N_11670,N_11895);
and U14368 (N_14368,N_12374,N_11684);
or U14369 (N_14369,N_10792,N_11611);
or U14370 (N_14370,N_11207,N_11320);
nor U14371 (N_14371,N_11335,N_12446);
nor U14372 (N_14372,N_12046,N_11161);
xor U14373 (N_14373,N_11092,N_10891);
nand U14374 (N_14374,N_12156,N_10268);
xnor U14375 (N_14375,N_10998,N_11882);
nand U14376 (N_14376,N_10543,N_11922);
xnor U14377 (N_14377,N_11352,N_11556);
nand U14378 (N_14378,N_11908,N_10470);
nand U14379 (N_14379,N_10350,N_10749);
or U14380 (N_14380,N_10475,N_11781);
nand U14381 (N_14381,N_11944,N_10023);
or U14382 (N_14382,N_11110,N_10851);
nor U14383 (N_14383,N_10723,N_11922);
nand U14384 (N_14384,N_11232,N_10220);
or U14385 (N_14385,N_10788,N_10414);
xnor U14386 (N_14386,N_11895,N_12082);
or U14387 (N_14387,N_10651,N_10521);
nand U14388 (N_14388,N_12022,N_11736);
nand U14389 (N_14389,N_12306,N_10018);
nor U14390 (N_14390,N_12261,N_12223);
nand U14391 (N_14391,N_11287,N_11974);
xor U14392 (N_14392,N_11944,N_11603);
nand U14393 (N_14393,N_11444,N_10836);
xor U14394 (N_14394,N_11275,N_12143);
nand U14395 (N_14395,N_11525,N_12471);
xnor U14396 (N_14396,N_11837,N_12484);
nand U14397 (N_14397,N_10471,N_11681);
nand U14398 (N_14398,N_11788,N_11725);
or U14399 (N_14399,N_10637,N_12105);
nor U14400 (N_14400,N_10433,N_10913);
and U14401 (N_14401,N_11002,N_10195);
xnor U14402 (N_14402,N_11542,N_12300);
and U14403 (N_14403,N_11105,N_11903);
xor U14404 (N_14404,N_11988,N_10148);
nor U14405 (N_14405,N_10092,N_11909);
nand U14406 (N_14406,N_12488,N_12486);
and U14407 (N_14407,N_12321,N_12385);
or U14408 (N_14408,N_11417,N_12283);
nand U14409 (N_14409,N_11615,N_11917);
and U14410 (N_14410,N_10074,N_10838);
and U14411 (N_14411,N_11282,N_10823);
xnor U14412 (N_14412,N_10855,N_10585);
or U14413 (N_14413,N_10081,N_10341);
nor U14414 (N_14414,N_11460,N_11245);
and U14415 (N_14415,N_12289,N_11124);
or U14416 (N_14416,N_10217,N_12081);
nand U14417 (N_14417,N_12017,N_10319);
xor U14418 (N_14418,N_10544,N_10224);
nor U14419 (N_14419,N_12478,N_10606);
nand U14420 (N_14420,N_12385,N_12423);
nand U14421 (N_14421,N_11041,N_10620);
xnor U14422 (N_14422,N_12026,N_11026);
nand U14423 (N_14423,N_11230,N_12344);
nand U14424 (N_14424,N_11790,N_10595);
or U14425 (N_14425,N_10697,N_12133);
and U14426 (N_14426,N_11274,N_11513);
xnor U14427 (N_14427,N_10902,N_10327);
xnor U14428 (N_14428,N_11798,N_10834);
nor U14429 (N_14429,N_12285,N_11347);
or U14430 (N_14430,N_12433,N_10755);
and U14431 (N_14431,N_10255,N_10174);
xnor U14432 (N_14432,N_11153,N_11973);
or U14433 (N_14433,N_11685,N_10543);
and U14434 (N_14434,N_11289,N_10463);
nand U14435 (N_14435,N_11208,N_12350);
xnor U14436 (N_14436,N_10466,N_10684);
xor U14437 (N_14437,N_11664,N_10481);
xnor U14438 (N_14438,N_11856,N_11328);
and U14439 (N_14439,N_11878,N_11270);
nor U14440 (N_14440,N_10947,N_10569);
nand U14441 (N_14441,N_10016,N_10042);
and U14442 (N_14442,N_12043,N_12293);
nor U14443 (N_14443,N_10800,N_11420);
or U14444 (N_14444,N_11051,N_12289);
nand U14445 (N_14445,N_10768,N_11119);
xor U14446 (N_14446,N_12022,N_11537);
xor U14447 (N_14447,N_11494,N_10381);
nor U14448 (N_14448,N_12276,N_12114);
nor U14449 (N_14449,N_11988,N_11607);
nand U14450 (N_14450,N_10703,N_10098);
or U14451 (N_14451,N_12165,N_10227);
nor U14452 (N_14452,N_11640,N_11688);
or U14453 (N_14453,N_10918,N_10233);
and U14454 (N_14454,N_10701,N_11343);
xnor U14455 (N_14455,N_11120,N_11178);
nand U14456 (N_14456,N_10791,N_10542);
nor U14457 (N_14457,N_11271,N_10833);
or U14458 (N_14458,N_11407,N_10311);
or U14459 (N_14459,N_11181,N_12443);
nand U14460 (N_14460,N_12329,N_10282);
nand U14461 (N_14461,N_10650,N_10125);
and U14462 (N_14462,N_11863,N_10517);
and U14463 (N_14463,N_11962,N_10726);
and U14464 (N_14464,N_12257,N_11296);
nor U14465 (N_14465,N_10947,N_11593);
nor U14466 (N_14466,N_10654,N_11452);
nor U14467 (N_14467,N_10272,N_12230);
nand U14468 (N_14468,N_11602,N_10768);
and U14469 (N_14469,N_12000,N_10956);
nand U14470 (N_14470,N_10746,N_10266);
xor U14471 (N_14471,N_10679,N_11803);
and U14472 (N_14472,N_10302,N_11687);
or U14473 (N_14473,N_10204,N_12139);
xnor U14474 (N_14474,N_11391,N_10411);
and U14475 (N_14475,N_10474,N_10804);
or U14476 (N_14476,N_11715,N_10037);
nand U14477 (N_14477,N_11322,N_10606);
or U14478 (N_14478,N_11003,N_12441);
or U14479 (N_14479,N_10467,N_11728);
nand U14480 (N_14480,N_11110,N_10065);
or U14481 (N_14481,N_10966,N_11785);
nor U14482 (N_14482,N_11568,N_10431);
and U14483 (N_14483,N_11964,N_11809);
nand U14484 (N_14484,N_12210,N_12131);
xnor U14485 (N_14485,N_11745,N_11365);
xor U14486 (N_14486,N_10016,N_11267);
and U14487 (N_14487,N_12407,N_12277);
or U14488 (N_14488,N_12394,N_10497);
and U14489 (N_14489,N_10042,N_11538);
xor U14490 (N_14490,N_10409,N_10114);
nor U14491 (N_14491,N_11249,N_10494);
nor U14492 (N_14492,N_11600,N_10815);
and U14493 (N_14493,N_10021,N_11301);
nor U14494 (N_14494,N_11834,N_11818);
or U14495 (N_14495,N_11924,N_10627);
xor U14496 (N_14496,N_10632,N_10306);
nand U14497 (N_14497,N_12221,N_11499);
or U14498 (N_14498,N_11802,N_10998);
nand U14499 (N_14499,N_10557,N_11771);
or U14500 (N_14500,N_11003,N_10846);
xnor U14501 (N_14501,N_11799,N_12083);
nand U14502 (N_14502,N_10597,N_12042);
nand U14503 (N_14503,N_11846,N_11837);
and U14504 (N_14504,N_10214,N_10595);
nand U14505 (N_14505,N_11098,N_11818);
or U14506 (N_14506,N_12307,N_11552);
nand U14507 (N_14507,N_10291,N_12315);
or U14508 (N_14508,N_10621,N_11725);
nor U14509 (N_14509,N_10996,N_10633);
nor U14510 (N_14510,N_11720,N_10949);
xor U14511 (N_14511,N_12185,N_10866);
xor U14512 (N_14512,N_10203,N_10024);
xor U14513 (N_14513,N_11219,N_10701);
nor U14514 (N_14514,N_10987,N_10264);
or U14515 (N_14515,N_12220,N_10681);
or U14516 (N_14516,N_10503,N_12344);
nor U14517 (N_14517,N_11280,N_12129);
xnor U14518 (N_14518,N_10791,N_10955);
and U14519 (N_14519,N_10761,N_10529);
and U14520 (N_14520,N_10914,N_11433);
nand U14521 (N_14521,N_10711,N_12386);
nor U14522 (N_14522,N_11409,N_10788);
and U14523 (N_14523,N_10550,N_12276);
nor U14524 (N_14524,N_11298,N_10678);
nand U14525 (N_14525,N_12245,N_10191);
xnor U14526 (N_14526,N_10459,N_10545);
or U14527 (N_14527,N_10714,N_11796);
nor U14528 (N_14528,N_12271,N_11753);
nor U14529 (N_14529,N_10847,N_11412);
or U14530 (N_14530,N_10139,N_10172);
nand U14531 (N_14531,N_11415,N_11879);
nor U14532 (N_14532,N_11022,N_11216);
xor U14533 (N_14533,N_10290,N_11269);
or U14534 (N_14534,N_11437,N_10786);
and U14535 (N_14535,N_12222,N_11169);
and U14536 (N_14536,N_10213,N_12431);
nand U14537 (N_14537,N_10611,N_12395);
xnor U14538 (N_14538,N_11915,N_12359);
or U14539 (N_14539,N_10162,N_11974);
or U14540 (N_14540,N_11210,N_11346);
or U14541 (N_14541,N_10290,N_11209);
and U14542 (N_14542,N_12191,N_10544);
xor U14543 (N_14543,N_11134,N_10230);
or U14544 (N_14544,N_11019,N_10578);
nor U14545 (N_14545,N_10820,N_12025);
or U14546 (N_14546,N_10594,N_10885);
nand U14547 (N_14547,N_10698,N_12251);
and U14548 (N_14548,N_12332,N_10065);
nor U14549 (N_14549,N_11203,N_10243);
nor U14550 (N_14550,N_11575,N_10603);
nor U14551 (N_14551,N_10752,N_10233);
or U14552 (N_14552,N_11751,N_11036);
xnor U14553 (N_14553,N_11873,N_10491);
xor U14554 (N_14554,N_10775,N_10698);
xor U14555 (N_14555,N_12171,N_12433);
xor U14556 (N_14556,N_10821,N_11200);
nand U14557 (N_14557,N_11397,N_11094);
nand U14558 (N_14558,N_12235,N_10144);
xnor U14559 (N_14559,N_10170,N_12023);
and U14560 (N_14560,N_11736,N_12143);
and U14561 (N_14561,N_12443,N_10638);
xnor U14562 (N_14562,N_10568,N_12360);
and U14563 (N_14563,N_12111,N_12431);
nand U14564 (N_14564,N_10753,N_12315);
nand U14565 (N_14565,N_11348,N_11063);
and U14566 (N_14566,N_11911,N_12370);
nand U14567 (N_14567,N_11670,N_11950);
and U14568 (N_14568,N_11529,N_11800);
nor U14569 (N_14569,N_12191,N_12188);
and U14570 (N_14570,N_10155,N_10265);
and U14571 (N_14571,N_11784,N_11388);
or U14572 (N_14572,N_10890,N_11391);
and U14573 (N_14573,N_11847,N_12349);
xnor U14574 (N_14574,N_10554,N_10131);
nand U14575 (N_14575,N_11632,N_11534);
xor U14576 (N_14576,N_12411,N_11608);
nand U14577 (N_14577,N_10903,N_10218);
or U14578 (N_14578,N_11438,N_10977);
nor U14579 (N_14579,N_11295,N_11721);
xnor U14580 (N_14580,N_11640,N_11254);
nand U14581 (N_14581,N_12004,N_11401);
and U14582 (N_14582,N_11499,N_10563);
or U14583 (N_14583,N_10618,N_10927);
xnor U14584 (N_14584,N_11726,N_10404);
nand U14585 (N_14585,N_12255,N_11161);
xor U14586 (N_14586,N_10075,N_10708);
and U14587 (N_14587,N_10716,N_11719);
xor U14588 (N_14588,N_10171,N_12226);
and U14589 (N_14589,N_12430,N_10077);
nor U14590 (N_14590,N_11309,N_10560);
nor U14591 (N_14591,N_11307,N_12162);
nor U14592 (N_14592,N_10996,N_10924);
nor U14593 (N_14593,N_10340,N_11536);
and U14594 (N_14594,N_10932,N_10656);
nor U14595 (N_14595,N_12266,N_11609);
nor U14596 (N_14596,N_10116,N_12019);
nand U14597 (N_14597,N_10720,N_11480);
xor U14598 (N_14598,N_12467,N_10430);
nor U14599 (N_14599,N_11353,N_11924);
nand U14600 (N_14600,N_10444,N_10182);
xnor U14601 (N_14601,N_10669,N_11995);
and U14602 (N_14602,N_12272,N_10578);
nand U14603 (N_14603,N_12113,N_10257);
nor U14604 (N_14604,N_12338,N_12306);
and U14605 (N_14605,N_11177,N_10948);
xor U14606 (N_14606,N_11541,N_10179);
nor U14607 (N_14607,N_11696,N_10417);
xor U14608 (N_14608,N_12295,N_10699);
xor U14609 (N_14609,N_11493,N_12155);
nor U14610 (N_14610,N_11468,N_10966);
xnor U14611 (N_14611,N_12431,N_10091);
or U14612 (N_14612,N_10229,N_11344);
nor U14613 (N_14613,N_12288,N_11617);
xnor U14614 (N_14614,N_10252,N_10375);
nor U14615 (N_14615,N_10011,N_10802);
xor U14616 (N_14616,N_12189,N_12332);
nand U14617 (N_14617,N_11097,N_10128);
and U14618 (N_14618,N_11654,N_10122);
and U14619 (N_14619,N_12082,N_10485);
xnor U14620 (N_14620,N_10068,N_10793);
nand U14621 (N_14621,N_11068,N_11821);
and U14622 (N_14622,N_11492,N_10561);
nand U14623 (N_14623,N_11548,N_10843);
nand U14624 (N_14624,N_10553,N_10450);
nor U14625 (N_14625,N_10010,N_12262);
or U14626 (N_14626,N_12205,N_10958);
xnor U14627 (N_14627,N_10388,N_10864);
or U14628 (N_14628,N_11570,N_11072);
or U14629 (N_14629,N_12101,N_11171);
nand U14630 (N_14630,N_11279,N_11506);
and U14631 (N_14631,N_11049,N_11687);
nor U14632 (N_14632,N_11034,N_12021);
xnor U14633 (N_14633,N_11171,N_11320);
nor U14634 (N_14634,N_11718,N_10335);
nor U14635 (N_14635,N_10159,N_11071);
nand U14636 (N_14636,N_12199,N_12321);
nand U14637 (N_14637,N_12486,N_11188);
nand U14638 (N_14638,N_11491,N_12065);
and U14639 (N_14639,N_10321,N_12187);
nor U14640 (N_14640,N_11126,N_10789);
or U14641 (N_14641,N_10065,N_10437);
xor U14642 (N_14642,N_10889,N_11613);
nand U14643 (N_14643,N_12415,N_11801);
xnor U14644 (N_14644,N_11489,N_12276);
xnor U14645 (N_14645,N_11211,N_12339);
nor U14646 (N_14646,N_10050,N_12406);
xor U14647 (N_14647,N_10343,N_10626);
xnor U14648 (N_14648,N_10279,N_11658);
nand U14649 (N_14649,N_10648,N_10915);
nand U14650 (N_14650,N_10269,N_10849);
nand U14651 (N_14651,N_10210,N_11244);
nand U14652 (N_14652,N_10870,N_10734);
nor U14653 (N_14653,N_11004,N_12498);
xor U14654 (N_14654,N_12306,N_10381);
and U14655 (N_14655,N_11448,N_11591);
and U14656 (N_14656,N_10601,N_10980);
and U14657 (N_14657,N_10959,N_11415);
nand U14658 (N_14658,N_11648,N_11692);
nand U14659 (N_14659,N_12075,N_11645);
or U14660 (N_14660,N_11715,N_10179);
nor U14661 (N_14661,N_11027,N_12456);
nor U14662 (N_14662,N_12429,N_12181);
xor U14663 (N_14663,N_11623,N_12462);
xnor U14664 (N_14664,N_12402,N_11612);
and U14665 (N_14665,N_11120,N_10216);
xnor U14666 (N_14666,N_12406,N_12119);
nand U14667 (N_14667,N_10233,N_11355);
nor U14668 (N_14668,N_12052,N_10865);
and U14669 (N_14669,N_10843,N_11437);
nor U14670 (N_14670,N_11305,N_11155);
and U14671 (N_14671,N_11087,N_11173);
or U14672 (N_14672,N_10870,N_12290);
and U14673 (N_14673,N_10523,N_11552);
xnor U14674 (N_14674,N_10592,N_10181);
or U14675 (N_14675,N_11135,N_12018);
nand U14676 (N_14676,N_11761,N_10675);
xor U14677 (N_14677,N_11972,N_10058);
nor U14678 (N_14678,N_10169,N_10910);
or U14679 (N_14679,N_10937,N_12180);
xnor U14680 (N_14680,N_12184,N_10840);
and U14681 (N_14681,N_12394,N_11341);
and U14682 (N_14682,N_12123,N_12107);
nor U14683 (N_14683,N_10256,N_10025);
or U14684 (N_14684,N_11896,N_11169);
xnor U14685 (N_14685,N_12056,N_11289);
nand U14686 (N_14686,N_11826,N_10711);
and U14687 (N_14687,N_11065,N_11885);
nand U14688 (N_14688,N_11437,N_11356);
nand U14689 (N_14689,N_10981,N_11498);
nor U14690 (N_14690,N_10515,N_11171);
and U14691 (N_14691,N_11572,N_12172);
xor U14692 (N_14692,N_10926,N_12256);
and U14693 (N_14693,N_11008,N_12252);
xnor U14694 (N_14694,N_11775,N_11989);
or U14695 (N_14695,N_10558,N_12482);
nor U14696 (N_14696,N_12034,N_12215);
xor U14697 (N_14697,N_10018,N_10293);
nor U14698 (N_14698,N_10903,N_12392);
nor U14699 (N_14699,N_10748,N_12065);
xor U14700 (N_14700,N_11672,N_10336);
nor U14701 (N_14701,N_10039,N_10703);
nand U14702 (N_14702,N_12026,N_11437);
or U14703 (N_14703,N_10363,N_11062);
or U14704 (N_14704,N_11995,N_12247);
xor U14705 (N_14705,N_12219,N_11353);
or U14706 (N_14706,N_12389,N_12047);
xor U14707 (N_14707,N_10075,N_11962);
xnor U14708 (N_14708,N_11018,N_11843);
or U14709 (N_14709,N_12299,N_10744);
nor U14710 (N_14710,N_12483,N_11904);
nor U14711 (N_14711,N_10469,N_12367);
or U14712 (N_14712,N_11731,N_11446);
or U14713 (N_14713,N_10143,N_10257);
and U14714 (N_14714,N_10248,N_10153);
and U14715 (N_14715,N_12077,N_12246);
or U14716 (N_14716,N_10741,N_11792);
nor U14717 (N_14717,N_11990,N_10921);
nor U14718 (N_14718,N_11115,N_10786);
and U14719 (N_14719,N_11393,N_10581);
or U14720 (N_14720,N_11114,N_10241);
and U14721 (N_14721,N_11220,N_11895);
and U14722 (N_14722,N_10002,N_10913);
xor U14723 (N_14723,N_10774,N_12303);
nand U14724 (N_14724,N_12055,N_11099);
xnor U14725 (N_14725,N_10853,N_11635);
nor U14726 (N_14726,N_11130,N_10147);
or U14727 (N_14727,N_12217,N_10140);
and U14728 (N_14728,N_11650,N_12223);
nor U14729 (N_14729,N_10318,N_10555);
and U14730 (N_14730,N_10704,N_12160);
nor U14731 (N_14731,N_10059,N_11616);
xnor U14732 (N_14732,N_12356,N_10416);
and U14733 (N_14733,N_10147,N_12436);
or U14734 (N_14734,N_11703,N_10525);
or U14735 (N_14735,N_10881,N_10431);
nor U14736 (N_14736,N_11247,N_10666);
nor U14737 (N_14737,N_12268,N_12155);
and U14738 (N_14738,N_12399,N_10700);
nand U14739 (N_14739,N_11969,N_11578);
or U14740 (N_14740,N_11324,N_12261);
and U14741 (N_14741,N_10136,N_10457);
nor U14742 (N_14742,N_11088,N_10730);
nor U14743 (N_14743,N_11607,N_12392);
and U14744 (N_14744,N_11534,N_11018);
or U14745 (N_14745,N_12141,N_10801);
and U14746 (N_14746,N_11002,N_10683);
and U14747 (N_14747,N_12021,N_10725);
nor U14748 (N_14748,N_12315,N_11979);
xnor U14749 (N_14749,N_10935,N_11663);
nor U14750 (N_14750,N_10110,N_12023);
and U14751 (N_14751,N_11945,N_10967);
nor U14752 (N_14752,N_11231,N_10985);
xnor U14753 (N_14753,N_11027,N_12239);
nor U14754 (N_14754,N_12473,N_10872);
xnor U14755 (N_14755,N_10164,N_11497);
and U14756 (N_14756,N_10629,N_11266);
nand U14757 (N_14757,N_11056,N_10197);
xor U14758 (N_14758,N_12236,N_11414);
and U14759 (N_14759,N_11850,N_10201);
nor U14760 (N_14760,N_12190,N_10682);
or U14761 (N_14761,N_12328,N_12253);
and U14762 (N_14762,N_12309,N_10019);
nand U14763 (N_14763,N_12096,N_10807);
or U14764 (N_14764,N_12032,N_11713);
and U14765 (N_14765,N_11567,N_11296);
or U14766 (N_14766,N_11913,N_12004);
and U14767 (N_14767,N_11928,N_11590);
nor U14768 (N_14768,N_11841,N_10158);
and U14769 (N_14769,N_10522,N_11148);
and U14770 (N_14770,N_11012,N_12116);
nor U14771 (N_14771,N_10223,N_11420);
and U14772 (N_14772,N_10531,N_12087);
or U14773 (N_14773,N_11347,N_11610);
xnor U14774 (N_14774,N_11189,N_11415);
or U14775 (N_14775,N_11053,N_10924);
nor U14776 (N_14776,N_10450,N_10245);
xnor U14777 (N_14777,N_12406,N_11388);
or U14778 (N_14778,N_10342,N_12260);
nor U14779 (N_14779,N_12498,N_11256);
and U14780 (N_14780,N_11749,N_10208);
nor U14781 (N_14781,N_12262,N_11723);
nor U14782 (N_14782,N_10168,N_10613);
or U14783 (N_14783,N_11639,N_11959);
or U14784 (N_14784,N_11320,N_11692);
nor U14785 (N_14785,N_11501,N_10321);
xnor U14786 (N_14786,N_10586,N_11294);
or U14787 (N_14787,N_10371,N_12391);
nor U14788 (N_14788,N_11570,N_11800);
and U14789 (N_14789,N_10144,N_11965);
or U14790 (N_14790,N_10094,N_10732);
xor U14791 (N_14791,N_12157,N_10532);
xor U14792 (N_14792,N_10541,N_10869);
nand U14793 (N_14793,N_10556,N_11207);
nor U14794 (N_14794,N_10198,N_10147);
xnor U14795 (N_14795,N_11022,N_10434);
xnor U14796 (N_14796,N_11137,N_11105);
nand U14797 (N_14797,N_11551,N_11519);
nand U14798 (N_14798,N_10046,N_11923);
or U14799 (N_14799,N_10698,N_12015);
xor U14800 (N_14800,N_12298,N_11764);
and U14801 (N_14801,N_10616,N_11016);
xnor U14802 (N_14802,N_11997,N_10358);
nand U14803 (N_14803,N_12235,N_10179);
nor U14804 (N_14804,N_11716,N_11631);
xor U14805 (N_14805,N_10463,N_11877);
xor U14806 (N_14806,N_12369,N_11128);
and U14807 (N_14807,N_11539,N_10203);
and U14808 (N_14808,N_11402,N_11878);
and U14809 (N_14809,N_10172,N_10160);
and U14810 (N_14810,N_10314,N_10894);
and U14811 (N_14811,N_12419,N_11052);
nor U14812 (N_14812,N_10172,N_11499);
or U14813 (N_14813,N_11825,N_10984);
nor U14814 (N_14814,N_10654,N_10821);
xnor U14815 (N_14815,N_10991,N_11256);
nor U14816 (N_14816,N_11160,N_11282);
nand U14817 (N_14817,N_11783,N_11132);
or U14818 (N_14818,N_11716,N_10296);
xor U14819 (N_14819,N_11181,N_10203);
and U14820 (N_14820,N_11265,N_12258);
xor U14821 (N_14821,N_11877,N_11259);
xor U14822 (N_14822,N_11254,N_12179);
xnor U14823 (N_14823,N_10239,N_11556);
nor U14824 (N_14824,N_10839,N_12465);
and U14825 (N_14825,N_11295,N_10212);
xor U14826 (N_14826,N_10235,N_10631);
nor U14827 (N_14827,N_10776,N_11048);
nand U14828 (N_14828,N_10338,N_11804);
nand U14829 (N_14829,N_12315,N_11122);
nor U14830 (N_14830,N_11549,N_10531);
xor U14831 (N_14831,N_10722,N_10530);
and U14832 (N_14832,N_11485,N_11777);
and U14833 (N_14833,N_10519,N_11034);
and U14834 (N_14834,N_11722,N_12462);
nand U14835 (N_14835,N_11225,N_12049);
xnor U14836 (N_14836,N_11368,N_11528);
and U14837 (N_14837,N_10039,N_12072);
and U14838 (N_14838,N_11097,N_10620);
nor U14839 (N_14839,N_11919,N_10989);
xnor U14840 (N_14840,N_12258,N_12160);
or U14841 (N_14841,N_11157,N_10113);
and U14842 (N_14842,N_11754,N_11211);
or U14843 (N_14843,N_10517,N_10418);
nand U14844 (N_14844,N_11287,N_11549);
nand U14845 (N_14845,N_10826,N_10057);
or U14846 (N_14846,N_11134,N_11998);
or U14847 (N_14847,N_10112,N_11631);
nand U14848 (N_14848,N_11108,N_11876);
or U14849 (N_14849,N_11643,N_11942);
xor U14850 (N_14850,N_10231,N_10311);
nor U14851 (N_14851,N_10008,N_11190);
nand U14852 (N_14852,N_11919,N_10436);
and U14853 (N_14853,N_10249,N_10421);
or U14854 (N_14854,N_10100,N_11403);
nor U14855 (N_14855,N_11163,N_11041);
nand U14856 (N_14856,N_12496,N_10696);
nor U14857 (N_14857,N_10416,N_10514);
xnor U14858 (N_14858,N_10897,N_12290);
or U14859 (N_14859,N_10505,N_11641);
and U14860 (N_14860,N_12349,N_10346);
nand U14861 (N_14861,N_11326,N_11093);
xnor U14862 (N_14862,N_12327,N_12297);
and U14863 (N_14863,N_12083,N_12306);
xor U14864 (N_14864,N_10382,N_10906);
or U14865 (N_14865,N_11270,N_11926);
xnor U14866 (N_14866,N_11813,N_10690);
nor U14867 (N_14867,N_11898,N_12100);
nand U14868 (N_14868,N_10892,N_11741);
or U14869 (N_14869,N_10900,N_11625);
or U14870 (N_14870,N_10137,N_11901);
nand U14871 (N_14871,N_12143,N_10303);
or U14872 (N_14872,N_10701,N_11699);
or U14873 (N_14873,N_11731,N_10025);
xor U14874 (N_14874,N_10549,N_12428);
nand U14875 (N_14875,N_11152,N_10247);
xnor U14876 (N_14876,N_10666,N_12053);
or U14877 (N_14877,N_11513,N_11479);
nand U14878 (N_14878,N_10299,N_10132);
or U14879 (N_14879,N_12382,N_12049);
or U14880 (N_14880,N_10415,N_10146);
or U14881 (N_14881,N_11244,N_11971);
nor U14882 (N_14882,N_10853,N_11999);
or U14883 (N_14883,N_10585,N_11228);
nor U14884 (N_14884,N_10000,N_10789);
xnor U14885 (N_14885,N_10145,N_12361);
nor U14886 (N_14886,N_10215,N_10571);
xnor U14887 (N_14887,N_10678,N_11903);
nor U14888 (N_14888,N_12454,N_12447);
and U14889 (N_14889,N_10171,N_12483);
nand U14890 (N_14890,N_11557,N_12061);
and U14891 (N_14891,N_10215,N_10612);
nor U14892 (N_14892,N_11851,N_11555);
or U14893 (N_14893,N_10000,N_12262);
and U14894 (N_14894,N_11066,N_10131);
xor U14895 (N_14895,N_12149,N_12240);
nand U14896 (N_14896,N_12227,N_11498);
xor U14897 (N_14897,N_12426,N_10183);
nor U14898 (N_14898,N_10649,N_10150);
nor U14899 (N_14899,N_11746,N_12356);
xor U14900 (N_14900,N_10967,N_12470);
and U14901 (N_14901,N_10118,N_10657);
xor U14902 (N_14902,N_10514,N_10451);
or U14903 (N_14903,N_11408,N_11268);
xnor U14904 (N_14904,N_12140,N_11066);
nor U14905 (N_14905,N_10203,N_10378);
and U14906 (N_14906,N_11766,N_11456);
nor U14907 (N_14907,N_12017,N_10468);
and U14908 (N_14908,N_11496,N_12218);
nor U14909 (N_14909,N_11878,N_10331);
nor U14910 (N_14910,N_12007,N_10494);
nand U14911 (N_14911,N_11021,N_11767);
nor U14912 (N_14912,N_11471,N_10928);
xnor U14913 (N_14913,N_10602,N_10546);
nand U14914 (N_14914,N_11351,N_10205);
nor U14915 (N_14915,N_10012,N_11492);
nand U14916 (N_14916,N_10770,N_10847);
nor U14917 (N_14917,N_11275,N_10751);
xor U14918 (N_14918,N_10708,N_10321);
xor U14919 (N_14919,N_10558,N_10523);
nand U14920 (N_14920,N_10924,N_11303);
xnor U14921 (N_14921,N_11402,N_10902);
nor U14922 (N_14922,N_12184,N_12201);
and U14923 (N_14923,N_12475,N_11987);
xor U14924 (N_14924,N_11890,N_11955);
nor U14925 (N_14925,N_10079,N_11460);
and U14926 (N_14926,N_11625,N_12185);
and U14927 (N_14927,N_12333,N_10780);
and U14928 (N_14928,N_11065,N_10614);
nand U14929 (N_14929,N_10269,N_10952);
nor U14930 (N_14930,N_11338,N_11540);
nor U14931 (N_14931,N_10680,N_11406);
and U14932 (N_14932,N_11362,N_10035);
and U14933 (N_14933,N_11117,N_12178);
or U14934 (N_14934,N_11843,N_10251);
and U14935 (N_14935,N_10606,N_11441);
xnor U14936 (N_14936,N_12050,N_12094);
xor U14937 (N_14937,N_12272,N_10782);
nand U14938 (N_14938,N_11252,N_10330);
xnor U14939 (N_14939,N_11994,N_11266);
nand U14940 (N_14940,N_12131,N_11195);
and U14941 (N_14941,N_10299,N_11633);
and U14942 (N_14942,N_11169,N_11665);
and U14943 (N_14943,N_12485,N_12122);
xor U14944 (N_14944,N_11799,N_12056);
and U14945 (N_14945,N_10693,N_10638);
nand U14946 (N_14946,N_10812,N_11469);
nor U14947 (N_14947,N_10317,N_10748);
nand U14948 (N_14948,N_10409,N_11341);
xor U14949 (N_14949,N_10528,N_12013);
nand U14950 (N_14950,N_12185,N_11146);
xnor U14951 (N_14951,N_11750,N_10929);
and U14952 (N_14952,N_10899,N_10963);
nand U14953 (N_14953,N_10910,N_11970);
nand U14954 (N_14954,N_11103,N_10257);
or U14955 (N_14955,N_11753,N_11631);
nand U14956 (N_14956,N_11653,N_11505);
nor U14957 (N_14957,N_12027,N_10146);
nor U14958 (N_14958,N_11475,N_11454);
nor U14959 (N_14959,N_10279,N_12148);
xnor U14960 (N_14960,N_10359,N_12157);
nand U14961 (N_14961,N_10646,N_12242);
nand U14962 (N_14962,N_11661,N_11197);
nor U14963 (N_14963,N_12032,N_12197);
nand U14964 (N_14964,N_11837,N_12284);
nor U14965 (N_14965,N_10617,N_10726);
nand U14966 (N_14966,N_12094,N_10299);
or U14967 (N_14967,N_11524,N_10667);
and U14968 (N_14968,N_12117,N_10970);
or U14969 (N_14969,N_11126,N_10447);
nand U14970 (N_14970,N_10306,N_11916);
nor U14971 (N_14971,N_11120,N_10342);
or U14972 (N_14972,N_10733,N_12209);
nor U14973 (N_14973,N_10824,N_12364);
and U14974 (N_14974,N_11341,N_12296);
nor U14975 (N_14975,N_11612,N_11322);
nor U14976 (N_14976,N_10158,N_11758);
xor U14977 (N_14977,N_12484,N_10425);
or U14978 (N_14978,N_12138,N_11066);
nor U14979 (N_14979,N_10253,N_10967);
nor U14980 (N_14980,N_10333,N_10151);
xnor U14981 (N_14981,N_10722,N_10493);
and U14982 (N_14982,N_11338,N_10257);
or U14983 (N_14983,N_12165,N_11467);
nor U14984 (N_14984,N_11488,N_10619);
and U14985 (N_14985,N_12010,N_12292);
nor U14986 (N_14986,N_11986,N_11456);
nand U14987 (N_14987,N_10846,N_10069);
nand U14988 (N_14988,N_11013,N_10512);
and U14989 (N_14989,N_10397,N_11716);
nand U14990 (N_14990,N_10235,N_11293);
xor U14991 (N_14991,N_10801,N_11998);
nand U14992 (N_14992,N_11648,N_12199);
or U14993 (N_14993,N_10326,N_11018);
and U14994 (N_14994,N_11472,N_12321);
or U14995 (N_14995,N_11866,N_11553);
xnor U14996 (N_14996,N_11363,N_11070);
or U14997 (N_14997,N_10264,N_11129);
xnor U14998 (N_14998,N_11983,N_11901);
nor U14999 (N_14999,N_10276,N_10615);
or U15000 (N_15000,N_14138,N_13358);
or U15001 (N_15001,N_14928,N_13866);
nor U15002 (N_15002,N_14437,N_14370);
nor U15003 (N_15003,N_14399,N_12919);
or U15004 (N_15004,N_13256,N_13251);
nand U15005 (N_15005,N_14111,N_14285);
nand U15006 (N_15006,N_13466,N_14359);
nand U15007 (N_15007,N_12784,N_14702);
xor U15008 (N_15008,N_14470,N_14409);
and U15009 (N_15009,N_13956,N_14292);
nor U15010 (N_15010,N_13116,N_14110);
nor U15011 (N_15011,N_12933,N_12538);
and U15012 (N_15012,N_13492,N_14451);
or U15013 (N_15013,N_13984,N_14654);
nor U15014 (N_15014,N_12521,N_13662);
xnor U15015 (N_15015,N_13094,N_13913);
nor U15016 (N_15016,N_12858,N_13874);
or U15017 (N_15017,N_14068,N_14097);
nor U15018 (N_15018,N_12861,N_12949);
nand U15019 (N_15019,N_12757,N_12745);
or U15020 (N_15020,N_13709,N_12659);
nand U15021 (N_15021,N_12721,N_12500);
nand U15022 (N_15022,N_14326,N_13652);
nor U15023 (N_15023,N_12536,N_14173);
or U15024 (N_15024,N_12711,N_13851);
nor U15025 (N_15025,N_14759,N_14710);
nand U15026 (N_15026,N_12585,N_14338);
xnor U15027 (N_15027,N_13828,N_12629);
and U15028 (N_15028,N_13494,N_12887);
or U15029 (N_15029,N_13462,N_13957);
nand U15030 (N_15030,N_12916,N_14739);
xor U15031 (N_15031,N_14044,N_12756);
nor U15032 (N_15032,N_14170,N_13777);
nor U15033 (N_15033,N_13380,N_12881);
and U15034 (N_15034,N_13742,N_13496);
and U15035 (N_15035,N_14055,N_13520);
and U15036 (N_15036,N_14941,N_13562);
and U15037 (N_15037,N_12733,N_14210);
nor U15038 (N_15038,N_13598,N_14954);
and U15039 (N_15039,N_12886,N_14865);
xor U15040 (N_15040,N_13924,N_13650);
nor U15041 (N_15041,N_12559,N_13590);
and U15042 (N_15042,N_12786,N_12912);
nand U15043 (N_15043,N_12951,N_13185);
nand U15044 (N_15044,N_14414,N_12618);
xnor U15045 (N_15045,N_13345,N_14423);
and U15046 (N_15046,N_12569,N_13350);
or U15047 (N_15047,N_13940,N_13182);
or U15048 (N_15048,N_14099,N_13565);
xnor U15049 (N_15049,N_13075,N_12883);
nor U15050 (N_15050,N_14386,N_13689);
or U15051 (N_15051,N_14971,N_13810);
or U15052 (N_15052,N_12915,N_13581);
and U15053 (N_15053,N_14936,N_13306);
nand U15054 (N_15054,N_14150,N_14488);
and U15055 (N_15055,N_14814,N_14938);
xnor U15056 (N_15056,N_13656,N_14464);
and U15057 (N_15057,N_12955,N_13629);
xnor U15058 (N_15058,N_12766,N_12667);
nand U15059 (N_15059,N_14331,N_13384);
nand U15060 (N_15060,N_14351,N_12654);
xor U15061 (N_15061,N_13275,N_12616);
xnor U15062 (N_15062,N_13136,N_12987);
or U15063 (N_15063,N_13600,N_14366);
or U15064 (N_15064,N_14268,N_14295);
nor U15065 (N_15065,N_14144,N_14393);
xnor U15066 (N_15066,N_12526,N_12888);
or U15067 (N_15067,N_14993,N_13544);
or U15068 (N_15068,N_13511,N_13531);
nor U15069 (N_15069,N_13425,N_14013);
and U15070 (N_15070,N_13242,N_14568);
nand U15071 (N_15071,N_13174,N_13090);
or U15072 (N_15072,N_14195,N_14644);
nor U15073 (N_15073,N_12741,N_13120);
xnor U15074 (N_15074,N_13213,N_14005);
xnor U15075 (N_15075,N_12508,N_13607);
nor U15076 (N_15076,N_13336,N_14255);
nand U15077 (N_15077,N_12787,N_14070);
nand U15078 (N_15078,N_14037,N_13694);
xor U15079 (N_15079,N_12907,N_12801);
xor U15080 (N_15080,N_13687,N_12825);
and U15081 (N_15081,N_14107,N_12964);
xor U15082 (N_15082,N_13692,N_14518);
nand U15083 (N_15083,N_13325,N_13859);
nor U15084 (N_15084,N_13161,N_14826);
or U15085 (N_15085,N_14406,N_14240);
xor U15086 (N_15086,N_12931,N_12587);
xor U15087 (N_15087,N_13611,N_13084);
or U15088 (N_15088,N_13180,N_14157);
or U15089 (N_15089,N_14973,N_14340);
nor U15090 (N_15090,N_13767,N_14582);
and U15091 (N_15091,N_12792,N_13197);
nand U15092 (N_15092,N_12665,N_12655);
and U15093 (N_15093,N_12657,N_14322);
nand U15094 (N_15094,N_12829,N_12793);
or U15095 (N_15095,N_13034,N_13809);
nor U15096 (N_15096,N_13606,N_14707);
and U15097 (N_15097,N_13241,N_13470);
or U15098 (N_15098,N_12905,N_14842);
and U15099 (N_15099,N_14611,N_14453);
nor U15100 (N_15100,N_14232,N_14856);
or U15101 (N_15101,N_13451,N_14774);
nand U15102 (N_15102,N_14927,N_14081);
or U15103 (N_15103,N_14897,N_14565);
nand U15104 (N_15104,N_14363,N_14324);
nor U15105 (N_15105,N_12978,N_12947);
xnor U15106 (N_15106,N_13898,N_14425);
nor U15107 (N_15107,N_14229,N_13103);
and U15108 (N_15108,N_13745,N_13098);
nand U15109 (N_15109,N_12533,N_14188);
and U15110 (N_15110,N_14302,N_14696);
nand U15111 (N_15111,N_13784,N_14925);
and U15112 (N_15112,N_13623,N_13093);
or U15113 (N_15113,N_13664,N_12639);
or U15114 (N_15114,N_14521,N_13764);
nand U15115 (N_15115,N_13168,N_14580);
or U15116 (N_15116,N_14102,N_13026);
nand U15117 (N_15117,N_13554,N_14402);
nand U15118 (N_15118,N_13058,N_13686);
nor U15119 (N_15119,N_13817,N_13181);
xor U15120 (N_15120,N_13835,N_14633);
and U15121 (N_15121,N_14329,N_14801);
and U15122 (N_15122,N_14078,N_14282);
xor U15123 (N_15123,N_13928,N_14764);
nand U15124 (N_15124,N_14498,N_14713);
and U15125 (N_15125,N_13557,N_13348);
or U15126 (N_15126,N_13079,N_13677);
or U15127 (N_15127,N_14638,N_14598);
nand U15128 (N_15128,N_13647,N_13782);
xnor U15129 (N_15129,N_13801,N_14738);
and U15130 (N_15130,N_13149,N_14827);
nor U15131 (N_15131,N_13618,N_14203);
and U15132 (N_15132,N_14678,N_13108);
xor U15133 (N_15133,N_13726,N_14587);
nand U15134 (N_15134,N_14500,N_13019);
xor U15135 (N_15135,N_14442,N_13294);
or U15136 (N_15136,N_13163,N_14661);
and U15137 (N_15137,N_14923,N_14477);
nand U15138 (N_15138,N_13884,N_14804);
and U15139 (N_15139,N_12682,N_13787);
or U15140 (N_15140,N_13264,N_14251);
and U15141 (N_15141,N_14450,N_12610);
or U15142 (N_15142,N_13445,N_14259);
nor U15143 (N_15143,N_13569,N_14847);
xor U15144 (N_15144,N_13398,N_14028);
or U15145 (N_15145,N_13006,N_12518);
or U15146 (N_15146,N_13698,N_13203);
or U15147 (N_15147,N_13449,N_13602);
nor U15148 (N_15148,N_13482,N_13527);
xnor U15149 (N_15149,N_13340,N_13892);
nor U15150 (N_15150,N_14373,N_14825);
xnor U15151 (N_15151,N_12504,N_14432);
and U15152 (N_15152,N_14625,N_12572);
or U15153 (N_15153,N_13959,N_14602);
nand U15154 (N_15154,N_13137,N_13043);
and U15155 (N_15155,N_13349,N_13986);
and U15156 (N_15156,N_14960,N_12830);
nor U15157 (N_15157,N_12561,N_13328);
and U15158 (N_15158,N_12838,N_14357);
or U15159 (N_15159,N_13521,N_13808);
or U15160 (N_15160,N_13238,N_14610);
or U15161 (N_15161,N_14628,N_12890);
xor U15162 (N_15162,N_12531,N_14887);
xor U15163 (N_15163,N_13639,N_13134);
and U15164 (N_15164,N_13863,N_12516);
or U15165 (N_15165,N_14216,N_13070);
and U15166 (N_15166,N_14433,N_14986);
xnor U15167 (N_15167,N_12902,N_14378);
nor U15168 (N_15168,N_12621,N_13452);
and U15169 (N_15169,N_14548,N_13690);
and U15170 (N_15170,N_14014,N_13009);
xor U15171 (N_15171,N_14069,N_13469);
or U15172 (N_15172,N_13036,N_12926);
nand U15173 (N_15173,N_13700,N_13681);
and U15174 (N_15174,N_12970,N_14485);
and U15175 (N_15175,N_14265,N_14141);
or U15176 (N_15176,N_13286,N_13024);
or U15177 (N_15177,N_13123,N_12724);
or U15178 (N_15178,N_14073,N_14832);
and U15179 (N_15179,N_14946,N_14218);
or U15180 (N_15180,N_14164,N_12627);
and U15181 (N_15181,N_13030,N_14679);
or U15182 (N_15182,N_13505,N_14920);
nor U15183 (N_15183,N_13910,N_13312);
xnor U15184 (N_15184,N_13483,N_13974);
or U15185 (N_15185,N_13891,N_13985);
nand U15186 (N_15186,N_13798,N_14056);
nor U15187 (N_15187,N_13593,N_14116);
nand U15188 (N_15188,N_13438,N_13184);
or U15189 (N_15189,N_13517,N_12702);
or U15190 (N_15190,N_14356,N_14163);
or U15191 (N_15191,N_13839,N_13113);
and U15192 (N_15192,N_13735,N_14647);
xor U15193 (N_15193,N_13240,N_14523);
nor U15194 (N_15194,N_14919,N_14151);
xor U15195 (N_15195,N_14271,N_13697);
xnor U15196 (N_15196,N_13570,N_13508);
xnor U15197 (N_15197,N_13774,N_14571);
nor U15198 (N_15198,N_13969,N_14724);
and U15199 (N_15199,N_13287,N_13622);
xor U15200 (N_15200,N_14176,N_12591);
nor U15201 (N_15201,N_13323,N_13150);
xnor U15202 (N_15202,N_13805,N_14117);
nand U15203 (N_15203,N_14597,N_13538);
nand U15204 (N_15204,N_14039,N_14996);
and U15205 (N_15205,N_13245,N_14276);
nand U15206 (N_15206,N_13410,N_13230);
nand U15207 (N_15207,N_12864,N_14940);
and U15208 (N_15208,N_13359,N_14063);
nor U15209 (N_15209,N_14554,N_12982);
nor U15210 (N_15210,N_13591,N_13951);
or U15211 (N_15211,N_14040,N_13715);
and U15212 (N_15212,N_13279,N_14193);
xnor U15213 (N_15213,N_13704,N_14031);
or U15214 (N_15214,N_14420,N_13977);
nand U15215 (N_15215,N_14362,N_13608);
and U15216 (N_15216,N_12980,N_12775);
nor U15217 (N_15217,N_14112,N_14454);
or U15218 (N_15218,N_13243,N_14857);
or U15219 (N_15219,N_13276,N_14918);
nand U15220 (N_15220,N_14088,N_13971);
nand U15221 (N_15221,N_14152,N_13816);
xor U15222 (N_15222,N_14410,N_13731);
nand U15223 (N_15223,N_12619,N_14656);
nor U15224 (N_15224,N_14058,N_14632);
or U15225 (N_15225,N_13751,N_13566);
nor U15226 (N_15226,N_12804,N_14030);
nand U15227 (N_15227,N_14562,N_13057);
or U15228 (N_15228,N_12515,N_14226);
nor U15229 (N_15229,N_14036,N_14660);
xor U15230 (N_15230,N_13446,N_13615);
xor U15231 (N_15231,N_14280,N_13394);
or U15232 (N_15232,N_13574,N_13781);
nor U15233 (N_15233,N_13176,N_14299);
and U15234 (N_15234,N_14023,N_12633);
and U15235 (N_15235,N_14360,N_14049);
nand U15236 (N_15236,N_12545,N_13405);
or U15237 (N_15237,N_12773,N_12566);
nor U15238 (N_15238,N_14736,N_14428);
nor U15239 (N_15239,N_12811,N_13175);
nor U15240 (N_15240,N_14156,N_14743);
or U15241 (N_15241,N_13304,N_14038);
and U15242 (N_15242,N_13732,N_12769);
xor U15243 (N_15243,N_13377,N_14675);
and U15244 (N_15244,N_12731,N_14966);
and U15245 (N_15245,N_14215,N_12755);
nand U15246 (N_15246,N_14802,N_14520);
nor U15247 (N_15247,N_14581,N_14260);
nor U15248 (N_15248,N_13290,N_13993);
nor U15249 (N_15249,N_13053,N_14975);
nand U15250 (N_15250,N_12750,N_13818);
nor U15251 (N_15251,N_13645,N_14950);
or U15252 (N_15252,N_13119,N_14981);
nor U15253 (N_15253,N_14583,N_14594);
or U15254 (N_15254,N_14977,N_14318);
xnor U15255 (N_15255,N_14435,N_12712);
xnor U15256 (N_15256,N_14025,N_13560);
or U15257 (N_15257,N_14881,N_13747);
xnor U15258 (N_15258,N_14926,N_13025);
xnor U15259 (N_15259,N_13640,N_13041);
nor U15260 (N_15260,N_14573,N_12794);
nor U15261 (N_15261,N_14962,N_12567);
nand U15262 (N_15262,N_13865,N_13016);
and U15263 (N_15263,N_13779,N_14389);
xor U15264 (N_15264,N_12513,N_13771);
nor U15265 (N_15265,N_12939,N_14001);
nor U15266 (N_15266,N_13044,N_14061);
nand U15267 (N_15267,N_12672,N_13049);
nor U15268 (N_15268,N_13837,N_12590);
xor U15269 (N_15269,N_14830,N_12839);
xor U15270 (N_15270,N_13217,N_14643);
nor U15271 (N_15271,N_13867,N_14325);
nand U15272 (N_15272,N_13671,N_13792);
and U15273 (N_15273,N_13729,N_12581);
nor U15274 (N_15274,N_12602,N_14480);
nor U15275 (N_15275,N_14662,N_14264);
nand U15276 (N_15276,N_14642,N_14531);
and U15277 (N_15277,N_13198,N_14145);
xnor U15278 (N_15278,N_14648,N_12634);
xor U15279 (N_15279,N_14512,N_12891);
nor U15280 (N_15280,N_12800,N_12683);
or U15281 (N_15281,N_13225,N_12743);
or U15282 (N_15282,N_13210,N_14524);
or U15283 (N_15283,N_13786,N_13341);
xor U15284 (N_15284,N_13497,N_13983);
nor U15285 (N_15285,N_13135,N_12934);
xnor U15286 (N_15286,N_14692,N_14646);
nand U15287 (N_15287,N_13847,N_14806);
or U15288 (N_15288,N_12870,N_14430);
nor U15289 (N_15289,N_13007,N_13518);
xnor U15290 (N_15290,N_13834,N_13015);
and U15291 (N_15291,N_14365,N_14294);
or U15292 (N_15292,N_12880,N_14388);
nor U15293 (N_15293,N_12502,N_13435);
xnor U15294 (N_15294,N_13526,N_14734);
and U15295 (N_15295,N_12529,N_14822);
nor U15296 (N_15296,N_12971,N_13540);
xor U15297 (N_15297,N_13826,N_13332);
nand U15298 (N_15298,N_13223,N_13717);
xor U15299 (N_15299,N_14538,N_12999);
xor U15300 (N_15300,N_12664,N_14530);
nor U15301 (N_15301,N_12514,N_12828);
nor U15302 (N_15302,N_13799,N_14397);
nand U15303 (N_15303,N_13580,N_13261);
nand U15304 (N_15304,N_13357,N_13923);
xor U15305 (N_15305,N_13945,N_13486);
and U15306 (N_15306,N_14411,N_14737);
or U15307 (N_15307,N_12668,N_14328);
xor U15308 (N_15308,N_13942,N_14659);
and U15309 (N_15309,N_13107,N_13250);
nor U15310 (N_15310,N_13080,N_12645);
nor U15311 (N_15311,N_14903,N_13564);
xor U15312 (N_15312,N_14653,N_14348);
xor U15313 (N_15313,N_12661,N_14899);
nand U15314 (N_15314,N_13067,N_13088);
nor U15315 (N_15315,N_13551,N_14385);
nand U15316 (N_15316,N_13424,N_12898);
and U15317 (N_15317,N_14048,N_13988);
and U15318 (N_15318,N_14283,N_14933);
nand U15319 (N_15319,N_13141,N_12944);
or U15320 (N_15320,N_12795,N_13824);
or U15321 (N_15321,N_12681,N_12930);
nor U15322 (N_15322,N_14391,N_13651);
nand U15323 (N_15323,N_13973,N_14481);
nor U15324 (N_15324,N_13227,N_13762);
and U15325 (N_15325,N_14862,N_12985);
xnor U15326 (N_15326,N_13588,N_14335);
or U15327 (N_15327,N_12640,N_14727);
and U15328 (N_15328,N_14426,N_13352);
nand U15329 (N_15329,N_13793,N_13008);
nand U15330 (N_15330,N_13413,N_12807);
or U15331 (N_15331,N_14236,N_14935);
nor U15332 (N_15332,N_14017,N_13720);
xor U15333 (N_15333,N_14060,N_13712);
nor U15334 (N_15334,N_14020,N_14553);
xnor U15335 (N_15335,N_14509,N_14071);
or U15336 (N_15336,N_14600,N_12688);
nand U15337 (N_15337,N_14834,N_13794);
nand U15338 (N_15338,N_13914,N_13087);
nor U15339 (N_15339,N_13760,N_13682);
and U15340 (N_15340,N_13125,N_14693);
nand U15341 (N_15341,N_14452,N_13173);
nor U15342 (N_15342,N_13236,N_13547);
nor U15343 (N_15343,N_14382,N_14390);
nand U15344 (N_15344,N_12760,N_13515);
and U15345 (N_15345,N_12856,N_13953);
and U15346 (N_15346,N_13365,N_12753);
and U15347 (N_15347,N_13274,N_13096);
and U15348 (N_15348,N_13430,N_13795);
nand U15349 (N_15349,N_14718,N_14957);
nand U15350 (N_15350,N_14533,N_13244);
xnor U15351 (N_15351,N_14368,N_13536);
nand U15352 (N_15352,N_12563,N_13829);
xnor U15353 (N_15353,N_13699,N_12601);
nor U15354 (N_15354,N_13807,N_13339);
and U15355 (N_15355,N_14135,N_13374);
or U15356 (N_15356,N_12981,N_13537);
nand U15357 (N_15357,N_13832,N_14939);
or U15358 (N_15358,N_13595,N_13917);
nand U15359 (N_15359,N_13159,N_14345);
and U15360 (N_15360,N_14082,N_14160);
and U15361 (N_15361,N_14243,N_13548);
or U15362 (N_15362,N_12726,N_14494);
or U15363 (N_15363,N_13933,N_13936);
nand U15364 (N_15364,N_14891,N_14012);
xnor U15365 (N_15365,N_13632,N_13734);
and U15366 (N_15366,N_14904,N_12878);
nor U15367 (N_15367,N_13576,N_12606);
or U15368 (N_15368,N_14209,N_14616);
xor U15369 (N_15369,N_13975,N_13129);
xnor U15370 (N_15370,N_13321,N_14279);
nand U15371 (N_15371,N_14242,N_14085);
or U15372 (N_15372,N_14290,N_14846);
xor U15373 (N_15373,N_14510,N_12577);
nand U15374 (N_15374,N_13237,N_13167);
xor U15375 (N_15375,N_14945,N_13707);
and U15376 (N_15376,N_13603,N_14998);
nand U15377 (N_15377,N_14109,N_14009);
xor U15378 (N_15378,N_14779,N_13232);
or U15379 (N_15379,N_13759,N_13376);
nand U15380 (N_15380,N_12613,N_13468);
or U15381 (N_15381,N_14871,N_14408);
xnor U15382 (N_15382,N_12853,N_14343);
nor U15383 (N_15383,N_13702,N_14606);
nand U15384 (N_15384,N_12727,N_13802);
xnor U15385 (N_15385,N_14191,N_13364);
xnor U15386 (N_15386,N_14793,N_12836);
nor U15387 (N_15387,N_14791,N_12805);
xor U15388 (N_15388,N_14221,N_14888);
or U15389 (N_15389,N_12802,N_14495);
and U15390 (N_15390,N_13385,N_13806);
and U15391 (N_15391,N_13389,N_13485);
xor U15392 (N_15392,N_14608,N_12942);
and U15393 (N_15393,N_13463,N_13897);
or U15394 (N_15394,N_14204,N_12604);
and U15395 (N_15395,N_14709,N_14394);
or U15396 (N_15396,N_14412,N_12770);
and U15397 (N_15397,N_12691,N_14851);
and U15398 (N_15398,N_13642,N_12894);
nand U15399 (N_15399,N_12908,N_13431);
nand U15400 (N_15400,N_14353,N_13931);
nor U15401 (N_15401,N_14697,N_13937);
nand U15402 (N_15402,N_14064,N_12777);
nand U15403 (N_15403,N_14721,N_13559);
and U15404 (N_15404,N_13653,N_14262);
nor U15405 (N_15405,N_13991,N_14944);
nor U15406 (N_15406,N_14369,N_14785);
and U15407 (N_15407,N_12698,N_13789);
nand U15408 (N_15408,N_13018,N_14835);
nor U15409 (N_15409,N_12859,N_13005);
or U15410 (N_15410,N_13379,N_14747);
and U15411 (N_15411,N_14824,N_13318);
xnor U15412 (N_15412,N_12656,N_12670);
and U15413 (N_15413,N_13625,N_14569);
xnor U15414 (N_15414,N_12710,N_14788);
xnor U15415 (N_15415,N_14244,N_12865);
and U15416 (N_15416,N_14441,N_13319);
nand U15417 (N_15417,N_14869,N_14168);
and U15418 (N_15418,N_13730,N_14916);
or U15419 (N_15419,N_14893,N_12582);
or U15420 (N_15420,N_14008,N_12625);
nand U15421 (N_15421,N_13401,N_14455);
and U15422 (N_15422,N_12628,N_13819);
or U15423 (N_15423,N_13719,N_14550);
nor U15424 (N_15424,N_13032,N_12693);
or U15425 (N_15425,N_14046,N_12872);
nand U15426 (N_15426,N_12764,N_13990);
and U15427 (N_15427,N_12967,N_14732);
and U15428 (N_15428,N_13214,N_14689);
nor U15429 (N_15429,N_13219,N_13965);
nand U15430 (N_15430,N_14900,N_14978);
nand U15431 (N_15431,N_13477,N_12718);
xor U15432 (N_15432,N_12783,N_13800);
nor U15433 (N_15433,N_13474,N_14468);
nand U15434 (N_15434,N_13077,N_14970);
nand U15435 (N_15435,N_13711,N_13278);
or U15436 (N_15436,N_13571,N_12954);
and U15437 (N_15437,N_13033,N_12692);
xor U15438 (N_15438,N_13420,N_13233);
nor U15439 (N_15439,N_14029,N_13128);
xor U15440 (N_15440,N_12637,N_13169);
nand U15441 (N_15441,N_14974,N_13327);
nor U15442 (N_15442,N_14703,N_14798);
and U15443 (N_15443,N_12810,N_12622);
and U15444 (N_15444,N_12984,N_12744);
nor U15445 (N_15445,N_13130,N_14377);
or U15446 (N_15446,N_12534,N_13894);
nand U15447 (N_15447,N_13654,N_12523);
or U15448 (N_15448,N_13387,N_13627);
nand U15449 (N_15449,N_14021,N_13020);
and U15450 (N_15450,N_14987,N_14748);
nor U15451 (N_15451,N_13481,N_13281);
xor U15452 (N_15452,N_14560,N_14605);
nand U15453 (N_15453,N_13165,N_14120);
nor U15454 (N_15454,N_12507,N_14472);
nor U15455 (N_15455,N_13490,N_14557);
nor U15456 (N_15456,N_13621,N_13029);
or U15457 (N_15457,N_14577,N_14400);
nor U15458 (N_15458,N_14407,N_14622);
or U15459 (N_15459,N_14740,N_12568);
and U15460 (N_15460,N_12706,N_13706);
and U15461 (N_15461,N_13102,N_12740);
and U15462 (N_15462,N_14317,N_13218);
or U15463 (N_15463,N_14549,N_12528);
nor U15464 (N_15464,N_13186,N_13701);
or U15465 (N_15465,N_14127,N_12676);
and U15466 (N_15466,N_13981,N_14090);
nand U15467 (N_15467,N_13427,N_13000);
nand U15468 (N_15468,N_13335,N_14769);
and U15469 (N_15469,N_13331,N_12960);
or U15470 (N_15470,N_14235,N_13407);
nand U15471 (N_15471,N_12713,N_14883);
and U15472 (N_15472,N_12584,N_12700);
or U15473 (N_15473,N_13888,N_13912);
xor U15474 (N_15474,N_13860,N_12684);
nor U15475 (N_15475,N_14123,N_13882);
xor U15476 (N_15476,N_12993,N_14607);
nand U15477 (N_15477,N_14489,N_14951);
nor U15478 (N_15478,N_12834,N_13060);
nor U15479 (N_15479,N_14416,N_14716);
nand U15480 (N_15480,N_13825,N_13941);
or U15481 (N_15481,N_14287,N_13397);
nand U15482 (N_15482,N_13226,N_14757);
or U15483 (N_15483,N_14256,N_12956);
nor U15484 (N_15484,N_13613,N_13585);
nor U15485 (N_15485,N_14131,N_14541);
xnor U15486 (N_15486,N_13151,N_13929);
nor U15487 (N_15487,N_13146,N_13599);
xor U15488 (N_15488,N_14006,N_13001);
nand U15489 (N_15489,N_13309,N_13523);
and U15490 (N_15490,N_12849,N_13143);
or U15491 (N_15491,N_12644,N_14617);
or U15492 (N_15492,N_14228,N_13282);
or U15493 (N_15493,N_14231,N_12928);
and U15494 (N_15494,N_13416,N_14114);
xor U15495 (N_15495,N_12547,N_14821);
nand U15496 (N_15496,N_14701,N_14527);
nor U15497 (N_15497,N_12535,N_14080);
nor U15498 (N_15498,N_14665,N_13519);
xor U15499 (N_15499,N_14760,N_12806);
xor U15500 (N_15500,N_14418,N_13199);
nor U15501 (N_15501,N_13708,N_12882);
or U15502 (N_15502,N_12937,N_13408);
xnor U15503 (N_15503,N_13052,N_12565);
and U15504 (N_15504,N_13178,N_14969);
and U15505 (N_15505,N_14961,N_13231);
or U15506 (N_15506,N_14041,N_13065);
nor U15507 (N_15507,N_14537,N_12917);
nor U15508 (N_15508,N_13507,N_14161);
xnor U15509 (N_15509,N_13194,N_13062);
nor U15510 (N_15510,N_12943,N_14576);
and U15511 (N_15511,N_12948,N_14908);
nand U15512 (N_15512,N_13283,N_14086);
nand U15513 (N_15513,N_14198,N_13118);
nand U15514 (N_15514,N_14682,N_14301);
or U15515 (N_15515,N_14735,N_12738);
and U15516 (N_15516,N_14750,N_12748);
and U15517 (N_15517,N_13317,N_14860);
nand U15518 (N_15518,N_13678,N_13943);
nand U15519 (N_15519,N_12714,N_14965);
or U15520 (N_15520,N_12695,N_12852);
xnor U15521 (N_15521,N_14487,N_13890);
nand U15522 (N_15522,N_14267,N_13908);
xor U15523 (N_15523,N_13674,N_13628);
nor U15524 (N_15524,N_14202,N_14010);
nand U15525 (N_15525,N_13351,N_13976);
and U15526 (N_15526,N_12532,N_13864);
and U15527 (N_15527,N_12658,N_12735);
and U15528 (N_15528,N_13703,N_13710);
and U15529 (N_15529,N_13516,N_13872);
nand U15530 (N_15530,N_12586,N_13121);
nand U15531 (N_15531,N_13665,N_14492);
xor U15532 (N_15532,N_14474,N_13797);
xnor U15533 (N_15533,N_14536,N_14705);
nor U15534 (N_15534,N_12752,N_13960);
xnor U15535 (N_15535,N_13458,N_13450);
or U15536 (N_15536,N_13447,N_13746);
or U15537 (N_15537,N_14823,N_13259);
nor U15538 (N_15538,N_13982,N_13368);
or U15539 (N_15539,N_14415,N_14953);
xnor U15540 (N_15540,N_14314,N_12790);
nand U15541 (N_15541,N_14190,N_14811);
or U15542 (N_15542,N_13780,N_12910);
nor U15543 (N_15543,N_13191,N_14354);
nand U15544 (N_15544,N_12961,N_12571);
xor U15545 (N_15545,N_12686,N_13224);
nand U15546 (N_15546,N_14711,N_12778);
and U15547 (N_15547,N_13371,N_14796);
and U15548 (N_15548,N_14332,N_13428);
xor U15549 (N_15549,N_13946,N_14140);
nand U15550 (N_15550,N_12599,N_13017);
nor U15551 (N_15551,N_14208,N_12774);
and U15552 (N_15552,N_12952,N_12819);
nand U15553 (N_15553,N_13947,N_12509);
nor U15554 (N_15554,N_14684,N_14934);
nor U15555 (N_15555,N_14629,N_14189);
nor U15556 (N_15556,N_14912,N_14446);
xnor U15557 (N_15557,N_14277,N_12990);
or U15558 (N_15558,N_13578,N_13761);
or U15559 (N_15559,N_13220,N_12958);
nor U15560 (N_15560,N_13395,N_14578);
or U15561 (N_15561,N_14753,N_12719);
and U15562 (N_15562,N_14310,N_14004);
nor U15563 (N_15563,N_14890,N_13263);
or U15564 (N_15564,N_14274,N_13392);
and U15565 (N_15565,N_14752,N_14503);
xnor U15566 (N_15566,N_12573,N_13756);
nor U15567 (N_15567,N_14434,N_12651);
nor U15568 (N_15568,N_14507,N_14057);
nand U15569 (N_15569,N_13297,N_12583);
nand U15570 (N_15570,N_14902,N_13723);
nor U15571 (N_15571,N_14540,N_12868);
and U15572 (N_15572,N_13111,N_13743);
nor U15573 (N_15573,N_14575,N_13644);
xnor U15574 (N_15574,N_13610,N_13970);
or U15575 (N_15575,N_13586,N_14207);
xor U15576 (N_15576,N_13858,N_13919);
nand U15577 (N_15577,N_14905,N_13004);
or U15578 (N_15578,N_13267,N_13343);
and U15579 (N_15579,N_14631,N_12772);
nor U15580 (N_15580,N_14761,N_13534);
or U15581 (N_15581,N_14379,N_13346);
nand U15582 (N_15582,N_13272,N_14375);
and U15583 (N_15583,N_14618,N_14513);
xor U15584 (N_15584,N_13310,N_13737);
nor U15585 (N_15585,N_13201,N_12844);
nor U15586 (N_15586,N_12593,N_14884);
nor U15587 (N_15587,N_12742,N_12552);
nor U15588 (N_15588,N_13370,N_14914);
nor U15589 (N_15589,N_13054,N_13669);
and U15590 (N_15590,N_13848,N_13383);
or U15591 (N_15591,N_13616,N_13273);
and U15592 (N_15592,N_14858,N_14197);
and U15593 (N_15593,N_14273,N_14850);
nand U15594 (N_15594,N_14948,N_13905);
and U15595 (N_15595,N_12510,N_12678);
nand U15596 (N_15596,N_12636,N_14723);
xor U15597 (N_15597,N_13691,N_14075);
nand U15598 (N_15598,N_13010,N_12873);
nand U15599 (N_15599,N_13510,N_13964);
nor U15600 (N_15600,N_13879,N_14181);
or U15601 (N_15601,N_14800,N_14475);
or U15602 (N_15602,N_13280,N_14213);
or U15603 (N_15603,N_13772,N_13594);
xnor U15604 (N_15604,N_14065,N_14989);
or U15605 (N_15605,N_12694,N_14700);
xor U15606 (N_15606,N_14516,N_13266);
and U15607 (N_15607,N_13495,N_13889);
xnor U15608 (N_15608,N_14298,N_12953);
nor U15609 (N_15609,N_14398,N_13337);
nor U15610 (N_15610,N_13028,N_13739);
nand U15611 (N_15611,N_14591,N_13292);
nor U15612 (N_15612,N_13360,N_13736);
and U15613 (N_15613,N_12903,N_13157);
and U15614 (N_15614,N_12867,N_14671);
xnor U15615 (N_15615,N_12959,N_12550);
nand U15616 (N_15616,N_14991,N_13039);
xnor U15617 (N_15617,N_13902,N_13162);
or U15618 (N_15618,N_14346,N_13915);
nand U15619 (N_15619,N_13553,N_12605);
nor U15620 (N_15620,N_12570,N_14148);
nor U15621 (N_15621,N_12963,N_14054);
nand U15622 (N_15622,N_12986,N_12722);
or U15623 (N_15623,N_13073,N_13893);
nand U15624 (N_15624,N_13400,N_13785);
xor U15625 (N_15625,N_12729,N_12871);
xnor U15626 (N_15626,N_14122,N_13042);
xor U15627 (N_15627,N_13269,N_13432);
or U15628 (N_15628,N_13439,N_13453);
nor U15629 (N_15629,N_13850,N_13436);
and U15630 (N_15630,N_13166,N_14763);
nor U15631 (N_15631,N_12904,N_12595);
and U15632 (N_15632,N_14288,N_13992);
nor U15633 (N_15633,N_14187,N_12546);
or U15634 (N_15634,N_14755,N_13156);
and U15635 (N_15635,N_13877,N_13666);
xnor U15636 (N_15636,N_14364,N_14084);
and U15637 (N_15637,N_13814,N_13952);
nor U15638 (N_15638,N_12648,N_14669);
and U15639 (N_15639,N_14108,N_13744);
and U15640 (N_15640,N_13811,N_13106);
nand U15641 (N_15641,N_12701,N_14932);
xor U15642 (N_15642,N_13633,N_14924);
and U15643 (N_15643,N_12669,N_13247);
nor U15644 (N_15644,N_13758,N_13133);
or U15645 (N_15645,N_13499,N_14812);
nand U15646 (N_15646,N_13308,N_13680);
xnor U15647 (N_15647,N_14483,N_13443);
xnor U15648 (N_15648,N_12716,N_13855);
xnor U15649 (N_15649,N_12708,N_13542);
nand U15650 (N_15650,N_14493,N_14154);
or U15651 (N_15651,N_13949,N_12992);
and U15652 (N_15652,N_12615,N_13967);
or U15653 (N_15653,N_14270,N_12715);
nor U15654 (N_15654,N_13672,N_13841);
or U15655 (N_15655,N_14690,N_13448);
nand U15656 (N_15656,N_12997,N_13880);
xor U15657 (N_15657,N_14535,N_12703);
nor U15658 (N_15658,N_13461,N_13770);
nand U15659 (N_15659,N_14119,N_13649);
or U15660 (N_15660,N_14601,N_13980);
or U15661 (N_15661,N_13301,N_14741);
nand U15662 (N_15662,N_14639,N_14992);
nand U15663 (N_15663,N_13260,N_14999);
or U15664 (N_15664,N_14125,N_14680);
xor U15665 (N_15665,N_14349,N_14342);
xor U15666 (N_15666,N_14956,N_14526);
xnor U15667 (N_15667,N_14034,N_13568);
xnor U15668 (N_15668,N_12791,N_13472);
and U15669 (N_15669,N_12780,N_13938);
and U15670 (N_15670,N_14367,N_14358);
nand U15671 (N_15671,N_14754,N_12840);
nor U15672 (N_15672,N_14731,N_13596);
xnor U15673 (N_15673,N_12580,N_14448);
xnor U15674 (N_15674,N_12687,N_14462);
xnor U15675 (N_15675,N_13315,N_13950);
nor U15676 (N_15676,N_14564,N_14092);
and U15677 (N_15677,N_13215,N_14841);
and U15678 (N_15678,N_12974,N_12991);
nor U15679 (N_15679,N_14572,N_12704);
and U15680 (N_15680,N_13344,N_14413);
nand U15681 (N_15681,N_14211,N_14843);
or U15682 (N_15682,N_14547,N_14238);
nand U15683 (N_15683,N_14674,N_14403);
xnor U15684 (N_15684,N_12924,N_12824);
and U15685 (N_15685,N_14706,N_14457);
xor U15686 (N_15686,N_13733,N_13265);
or U15687 (N_15687,N_14217,N_13363);
xor U15688 (N_15688,N_14506,N_13844);
xor U15689 (N_15689,N_14799,N_13476);
or U15690 (N_15690,N_13529,N_12976);
and U15691 (N_15691,N_13790,N_13110);
xor U15692 (N_15692,N_14128,N_12723);
xor U15693 (N_15693,N_14508,N_14949);
nand U15694 (N_15694,N_12736,N_14819);
nand U15695 (N_15695,N_14113,N_12603);
or U15696 (N_15696,N_12554,N_12737);
and U15697 (N_15697,N_12785,N_14963);
xor U15698 (N_15698,N_12763,N_13896);
nor U15699 (N_15699,N_13901,N_13987);
or U15700 (N_15700,N_13289,N_12653);
nand U15701 (N_15701,N_13422,N_13904);
and U15702 (N_15702,N_14967,N_13047);
xnor U15703 (N_15703,N_13045,N_14772);
or U15704 (N_15704,N_13684,N_13670);
nand U15705 (N_15705,N_13003,N_14511);
or U15706 (N_15706,N_12674,N_12607);
xor U15707 (N_15707,N_14291,N_14284);
nand U15708 (N_15708,N_13100,N_14381);
nor U15709 (N_15709,N_12799,N_12895);
nand U15710 (N_15710,N_12709,N_13630);
nand U15711 (N_15711,N_14921,N_12813);
nand U15712 (N_15712,N_12869,N_13545);
nand U15713 (N_15713,N_14104,N_12776);
or U15714 (N_15714,N_14937,N_13179);
or U15715 (N_15715,N_14337,N_12797);
xor U15716 (N_15716,N_13404,N_12717);
nor U15717 (N_15717,N_13114,N_13856);
or U15718 (N_15718,N_14444,N_14278);
nor U15719 (N_15719,N_14515,N_14673);
xnor U15720 (N_15720,N_14688,N_13038);
nand U15721 (N_15721,N_13104,N_14456);
and U15722 (N_15722,N_14964,N_13958);
and U15723 (N_15723,N_13092,N_12689);
and U15724 (N_15724,N_12925,N_13444);
nor U15725 (N_15725,N_13148,N_14651);
or U15726 (N_15726,N_13663,N_14249);
and U15727 (N_15727,N_13998,N_14281);
nand U15728 (N_15728,N_13695,N_13966);
or U15729 (N_15729,N_13207,N_14165);
xnor U15730 (N_15730,N_14895,N_14620);
nand U15731 (N_15731,N_12781,N_14626);
nor U15732 (N_15732,N_13455,N_13099);
nor U15733 (N_15733,N_13532,N_13875);
nand U15734 (N_15734,N_12812,N_14459);
and U15735 (N_15735,N_14898,N_14742);
or U15736 (N_15736,N_12897,N_14105);
and U15737 (N_15737,N_14539,N_12530);
nor U15738 (N_15738,N_14720,N_13878);
or U15739 (N_15739,N_14894,N_13748);
xor U15740 (N_15740,N_13646,N_13248);
or U15741 (N_15741,N_12998,N_13071);
nand U15742 (N_15742,N_12842,N_13921);
and U15743 (N_15743,N_13204,N_12863);
nor U15744 (N_15744,N_13525,N_13926);
or U15745 (N_15745,N_14910,N_13046);
and U15746 (N_15746,N_13543,N_12921);
or U15747 (N_15747,N_14614,N_14704);
and U15748 (N_15748,N_13881,N_14184);
nor U15749 (N_15749,N_14866,N_14466);
or U15750 (N_15750,N_13414,N_14615);
or U15751 (N_15751,N_13750,N_12850);
nor U15752 (N_15752,N_14266,N_14201);
or U15753 (N_15753,N_13788,N_12832);
or U15754 (N_15754,N_13193,N_14000);
nor U15755 (N_15755,N_14770,N_13907);
or U15756 (N_15756,N_13868,N_13843);
xnor U15757 (N_15757,N_14134,N_13876);
or U15758 (N_15758,N_12675,N_14026);
nor U15759 (N_15759,N_13539,N_14172);
nor U15760 (N_15760,N_14766,N_13911);
nand U15761 (N_15761,N_14486,N_14083);
and U15762 (N_15762,N_13996,N_14733);
nand U15763 (N_15763,N_14613,N_14913);
xnor U15764 (N_15764,N_13836,N_13257);
and U15765 (N_15765,N_13258,N_13796);
xor U15766 (N_15766,N_13112,N_12977);
or U15767 (N_15767,N_12511,N_14599);
nand U15768 (N_15768,N_13572,N_12979);
nand U15769 (N_15769,N_13064,N_12679);
nor U15770 (N_15770,N_13634,N_13101);
nor U15771 (N_15771,N_12935,N_12815);
or U15772 (N_15772,N_12874,N_14907);
or U15773 (N_15773,N_12612,N_13887);
nand U15774 (N_15774,N_14555,N_14722);
nor U15775 (N_15775,N_13288,N_14062);
and U15776 (N_15776,N_13271,N_12556);
or U15777 (N_15777,N_13484,N_12680);
xnor U15778 (N_15778,N_13147,N_14237);
and U15779 (N_15779,N_13930,N_13552);
and U15780 (N_15780,N_13381,N_13255);
or U15781 (N_15781,N_13660,N_14476);
xor U15782 (N_15782,N_14196,N_14854);
nand U15783 (N_15783,N_14219,N_12846);
or U15784 (N_15784,N_13604,N_12505);
nor U15785 (N_15785,N_14845,N_13776);
nand U15786 (N_15786,N_13209,N_13145);
xor U15787 (N_15787,N_14227,N_12578);
nand U15788 (N_15788,N_12600,N_14980);
xor U15789 (N_15789,N_13347,N_12525);
nand U15790 (N_15790,N_12957,N_13609);
nand U15791 (N_15791,N_14192,N_13631);
or U15792 (N_15792,N_13228,N_13356);
and U15793 (N_15793,N_13501,N_14361);
nor U15794 (N_15794,N_12588,N_13927);
nor U15795 (N_15795,N_14132,N_13812);
or U15796 (N_15796,N_12823,N_13870);
nand U15797 (N_15797,N_13925,N_14077);
nand U15798 (N_15798,N_14997,N_13299);
and U15799 (N_15799,N_13626,N_13296);
and U15800 (N_15800,N_14147,N_13584);
nand U15801 (N_15801,N_14214,N_12975);
or U15802 (N_15802,N_12845,N_14676);
or U15803 (N_15803,N_13467,N_12699);
nor U15804 (N_15804,N_13821,N_14943);
or U15805 (N_15805,N_13074,N_13948);
nand U15806 (N_15806,N_13932,N_13366);
and U15807 (N_15807,N_13873,N_12646);
nor U15808 (N_15808,N_14072,N_14174);
or U15809 (N_15809,N_13139,N_14304);
nand U15810 (N_15810,N_12596,N_14906);
or U15811 (N_15811,N_13205,N_12972);
nand U15812 (N_15812,N_13738,N_13284);
or U15813 (N_15813,N_13375,N_13673);
or U15814 (N_15814,N_13089,N_14787);
xnor U15815 (N_15815,N_13473,N_12885);
and U15816 (N_15816,N_14471,N_13027);
nand U15817 (N_15817,N_14589,N_14376);
xnor U15818 (N_15818,N_14730,N_14848);
nor U15819 (N_15819,N_12817,N_13373);
nand U15820 (N_15820,N_14789,N_13920);
nand U15821 (N_15821,N_13886,N_13313);
nand U15822 (N_15822,N_13326,N_12543);
nand U15823 (N_15823,N_14517,N_12728);
nand U15824 (N_15824,N_14768,N_13558);
or U15825 (N_15825,N_14296,N_12542);
and U15826 (N_15826,N_13056,N_13222);
or U15827 (N_15827,N_14015,N_14178);
nor U15828 (N_15828,N_13741,N_13441);
nand U15829 (N_15829,N_14947,N_12512);
or U15830 (N_15830,N_14327,N_14022);
nor U15831 (N_15831,N_13322,N_13063);
xor U15832 (N_15832,N_13803,N_14566);
nand U15833 (N_15833,N_13934,N_13753);
or U15834 (N_15834,N_13354,N_14355);
xnor U15835 (N_15835,N_13170,N_14247);
nor U15836 (N_15836,N_13657,N_14612);
nand U15837 (N_15837,N_12537,N_13491);
nand U15838 (N_15838,N_14018,N_13721);
nor U15839 (N_15839,N_14133,N_13550);
or U15840 (N_15840,N_14223,N_14007);
xor U15841 (N_15841,N_13668,N_13661);
or U15842 (N_15842,N_13202,N_12540);
xnor U15843 (N_15843,N_13212,N_13617);
nor U15844 (N_15844,N_13048,N_14886);
and U15845 (N_15845,N_14529,N_14771);
and U15846 (N_15846,N_14586,N_14066);
nor U15847 (N_15847,N_14840,N_14293);
nand U15848 (N_15848,N_14909,N_14309);
xor U15849 (N_15849,N_14334,N_12820);
nor U15850 (N_15850,N_12576,N_13253);
and U15851 (N_15851,N_14885,N_13619);
nor U15852 (N_15852,N_14417,N_14677);
or U15853 (N_15853,N_14100,N_14911);
xnor U15854 (N_15854,N_14837,N_14320);
and U15855 (N_15855,N_13069,N_14627);
nand U15856 (N_15856,N_12923,N_13524);
and U15857 (N_15857,N_13132,N_14137);
and U15858 (N_15858,N_14051,N_14142);
or U15859 (N_15859,N_14725,N_13955);
xor U15860 (N_15860,N_13813,N_13127);
nand U15861 (N_15861,N_14694,N_13200);
nand U15862 (N_15862,N_12725,N_14230);
or U15863 (N_15863,N_13740,N_13013);
nor U15864 (N_15864,N_14047,N_14915);
nand U15865 (N_15865,N_13514,N_13316);
xnor U15866 (N_15866,N_14592,N_14094);
and U15867 (N_15867,N_12501,N_14155);
nor U15868 (N_15868,N_13078,N_14773);
and U15869 (N_15869,N_14087,N_14257);
nor U15870 (N_15870,N_14019,N_13500);
nand U15871 (N_15871,N_14621,N_14308);
xor U15872 (N_15872,N_13638,N_14726);
or U15873 (N_15873,N_13109,N_14098);
nand U15874 (N_15874,N_13480,N_14816);
nand U15875 (N_15875,N_12524,N_14931);
and U15876 (N_15876,N_14686,N_13361);
and U15877 (N_15877,N_14248,N_14347);
xnor U15878 (N_15878,N_13206,N_13869);
xnor U15879 (N_15879,N_12989,N_14563);
nor U15880 (N_15880,N_13188,N_14502);
nor U15881 (N_15881,N_13830,N_14561);
and U15882 (N_15882,N_13655,N_13429);
xor U15883 (N_15883,N_14877,N_14596);
and U15884 (N_15884,N_14027,N_14118);
or U15885 (N_15885,N_13153,N_14401);
nand U15886 (N_15886,N_13456,N_14460);
xnor U15887 (N_15887,N_12936,N_13131);
nand U15888 (N_15888,N_12749,N_12809);
and U15889 (N_15889,N_13989,N_14162);
nor U15890 (N_15890,N_13757,N_12821);
or U15891 (N_15891,N_13512,N_13307);
nand U15892 (N_15892,N_13909,N_12833);
nand U15893 (N_15893,N_12965,N_13040);
or U15894 (N_15894,N_13827,N_14958);
nor U15895 (N_15895,N_14585,N_14183);
nor U15896 (N_15896,N_14942,N_14778);
nor U15897 (N_15897,N_13535,N_12762);
xor U15898 (N_15898,N_12826,N_14380);
nor U15899 (N_15899,N_13900,N_13311);
xnor U15900 (N_15900,N_13437,N_12696);
and U15901 (N_15901,N_13022,N_13158);
or U15902 (N_15902,N_12796,N_12697);
nor U15903 (N_15903,N_14784,N_13849);
xnor U15904 (N_15904,N_14863,N_14431);
or U15905 (N_15905,N_14465,N_13409);
and U15906 (N_15906,N_14719,N_14666);
nor U15907 (N_15907,N_13314,N_13388);
or U15908 (N_15908,N_13055,N_13768);
nand U15909 (N_15909,N_14124,N_14655);
xor U15910 (N_15910,N_13587,N_13714);
nor U15911 (N_15911,N_14551,N_14263);
and U15912 (N_15912,N_13334,N_14405);
and U15913 (N_15913,N_14177,N_14043);
nor U15914 (N_15914,N_14473,N_13386);
nor U15915 (N_15915,N_14003,N_12771);
nand U15916 (N_15916,N_14383,N_13037);
nor U15917 (N_15917,N_12551,N_12705);
xnor U15918 (N_15918,N_13399,N_12549);
nor U15919 (N_15919,N_13124,N_12918);
xnor U15920 (N_15920,N_14681,N_12589);
or U15921 (N_15921,N_12614,N_14685);
xnor U15922 (N_15922,N_13234,N_14889);
nand U15923 (N_15923,N_14496,N_13567);
nor U15924 (N_15924,N_14794,N_13597);
nor U15925 (N_15925,N_12597,N_14995);
xnor U15926 (N_15926,N_14984,N_13277);
or U15927 (N_15927,N_12995,N_14781);
nor U15928 (N_15928,N_13614,N_12519);
nand U15929 (N_15929,N_14930,N_12983);
or U15930 (N_15930,N_13249,N_14813);
nor U15931 (N_15931,N_12562,N_12592);
nor U15932 (N_15932,N_14042,N_12730);
nor U15933 (N_15933,N_12841,N_13082);
xnor U15934 (N_15934,N_13105,N_13840);
and U15935 (N_15935,N_14783,N_13978);
xor U15936 (N_15936,N_13676,N_13635);
and U15937 (N_15937,N_13155,N_13023);
xor U15938 (N_15938,N_14808,N_14206);
and U15939 (N_15939,N_14233,N_14815);
nand U15940 (N_15940,N_12642,N_12541);
nand U15941 (N_15941,N_12814,N_13778);
xnor U15942 (N_15942,N_13459,N_12638);
nor U15943 (N_15943,N_12884,N_14501);
and U15944 (N_15944,N_14637,N_14807);
and U15945 (N_15945,N_14505,N_13563);
or U15946 (N_15946,N_14052,N_13688);
xor U15947 (N_15947,N_13086,N_12899);
or U15948 (N_15948,N_14146,N_14864);
and U15949 (N_15949,N_14810,N_12900);
nor U15950 (N_15950,N_12671,N_13144);
nand U15951 (N_15951,N_13465,N_13620);
xnor U15952 (N_15952,N_13895,N_14663);
nor U15953 (N_15953,N_13035,N_12758);
nor U15954 (N_15954,N_13530,N_13546);
xnor U15955 (N_15955,N_14976,N_13324);
and U15956 (N_15956,N_14185,N_12560);
nand U15957 (N_15957,N_14166,N_14795);
xnor U15958 (N_15958,N_14158,N_14786);
xor U15959 (N_15959,N_12594,N_13612);
or U15960 (N_15960,N_12875,N_13196);
or U15961 (N_15961,N_13861,N_13963);
nor U15962 (N_15962,N_14199,N_14101);
nor U15963 (N_15963,N_12940,N_14171);
xnor U15964 (N_15964,N_14695,N_14286);
or U15965 (N_15965,N_14440,N_14579);
or U15966 (N_15966,N_12641,N_14169);
nand U15967 (N_15967,N_14067,N_13421);
or U15968 (N_15968,N_14050,N_14892);
and U15969 (N_15969,N_13014,N_12630);
nor U15970 (N_15970,N_12822,N_14525);
or U15971 (N_15971,N_13935,N_14588);
xor U15972 (N_15972,N_12767,N_14528);
and U15973 (N_15973,N_13417,N_12720);
and U15974 (N_15974,N_12520,N_12857);
nand U15975 (N_15975,N_13403,N_14765);
nor U15976 (N_15976,N_12553,N_14687);
nand U15977 (N_15977,N_13995,N_13658);
or U15978 (N_15978,N_14479,N_14776);
and U15979 (N_15979,N_13972,N_13152);
and U15980 (N_15980,N_13418,N_14831);
nand U15981 (N_15981,N_13522,N_13918);
and U15982 (N_15982,N_14658,N_12564);
and U15983 (N_15983,N_14868,N_13262);
or U15984 (N_15984,N_14584,N_12650);
or U15985 (N_15985,N_14297,N_14775);
xor U15986 (N_15986,N_14929,N_12969);
xnor U15987 (N_15987,N_13916,N_13140);
nor U15988 (N_15988,N_14447,N_14253);
nand U15989 (N_15989,N_14922,N_12631);
xnor U15990 (N_15990,N_13059,N_13954);
or U15991 (N_15991,N_12539,N_12962);
or U15992 (N_15992,N_13679,N_12611);
xor U15993 (N_15993,N_13766,N_12803);
nand U15994 (N_15994,N_14546,N_14833);
nand U15995 (N_15995,N_12782,N_12973);
or U15996 (N_15996,N_14552,N_13555);
xor U15997 (N_15997,N_14438,N_13382);
and U15998 (N_15998,N_14699,N_13076);
xor U15999 (N_15999,N_14715,N_14544);
xor U16000 (N_16000,N_13968,N_13085);
nor U16001 (N_16001,N_13177,N_14872);
or U16002 (N_16002,N_13592,N_14828);
nor U16003 (N_16003,N_13675,N_12941);
and U16004 (N_16004,N_14250,N_14875);
nand U16005 (N_16005,N_13504,N_12575);
or U16006 (N_16006,N_14994,N_14664);
and U16007 (N_16007,N_12808,N_14241);
xnor U16008 (N_16008,N_13083,N_14635);
nand U16009 (N_16009,N_14106,N_14595);
and U16010 (N_16010,N_14756,N_12677);
xnor U16011 (N_16011,N_14095,N_13749);
nand U16012 (N_16012,N_13246,N_12877);
nor U16013 (N_16013,N_13066,N_14559);
nor U16014 (N_16014,N_14623,N_13126);
nor U16015 (N_16015,N_14650,N_13605);
nor U16016 (N_16016,N_12579,N_13122);
or U16017 (N_16017,N_13636,N_12685);
and U16018 (N_16018,N_14641,N_14269);
nand U16019 (N_16019,N_13773,N_14917);
and U16020 (N_16020,N_14955,N_12765);
nor U16021 (N_16021,N_14545,N_13641);
nand U16022 (N_16022,N_14670,N_14032);
and U16023 (N_16023,N_13582,N_13791);
or U16024 (N_16024,N_14103,N_13412);
nand U16025 (N_16025,N_14570,N_14558);
xnor U16026 (N_16026,N_14691,N_12827);
xnor U16027 (N_16027,N_14574,N_12660);
nor U16028 (N_16028,N_14439,N_12506);
xor U16029 (N_16029,N_14744,N_14180);
nand U16030 (N_16030,N_12847,N_14861);
nor U16031 (N_16031,N_12624,N_13330);
nor U16032 (N_16032,N_13727,N_13160);
xor U16033 (N_16033,N_14490,N_14130);
or U16034 (N_16034,N_13012,N_14136);
nand U16035 (N_16035,N_13378,N_14482);
or U16036 (N_16036,N_12945,N_14972);
nand U16037 (N_16037,N_13754,N_14896);
xor U16038 (N_16038,N_14484,N_13362);
or U16039 (N_16039,N_14316,N_14636);
or U16040 (N_16040,N_12860,N_14175);
or U16041 (N_16041,N_13117,N_13979);
xor U16042 (N_16042,N_12929,N_13171);
xnor U16043 (N_16043,N_14790,N_14239);
or U16044 (N_16044,N_13142,N_13216);
or U16045 (N_16045,N_12747,N_13164);
xor U16046 (N_16046,N_12768,N_12927);
nand U16047 (N_16047,N_14478,N_13922);
nand U16048 (N_16048,N_14179,N_13239);
xor U16049 (N_16049,N_12946,N_14901);
and U16050 (N_16050,N_14053,N_13329);
xnor U16051 (N_16051,N_14167,N_13396);
xnor U16052 (N_16052,N_14341,N_13643);
and U16053 (N_16053,N_14139,N_12652);
xnor U16054 (N_16054,N_14758,N_14683);
nor U16055 (N_16055,N_14307,N_13183);
nor U16056 (N_16056,N_14882,N_12544);
xor U16057 (N_16057,N_12779,N_14323);
and U16058 (N_16058,N_14567,N_12988);
nor U16059 (N_16059,N_13291,N_12643);
or U16060 (N_16060,N_13342,N_13775);
and U16061 (N_16061,N_14258,N_13372);
and U16062 (N_16062,N_13648,N_14011);
nor U16063 (N_16063,N_14045,N_13471);
or U16064 (N_16064,N_13270,N_14352);
or U16065 (N_16065,N_14990,N_12598);
xnor U16066 (N_16066,N_14254,N_13254);
and U16067 (N_16067,N_12609,N_13434);
xor U16068 (N_16068,N_14222,N_12843);
and U16069 (N_16069,N_13011,N_14313);
nand U16070 (N_16070,N_13338,N_14469);
xnor U16071 (N_16071,N_14803,N_12855);
nand U16072 (N_16072,N_14746,N_13479);
nor U16073 (N_16073,N_13716,N_12557);
nor U16074 (N_16074,N_13906,N_13846);
nor U16075 (N_16075,N_14855,N_13994);
and U16076 (N_16076,N_14497,N_12663);
xor U16077 (N_16077,N_13831,N_12909);
or U16078 (N_16078,N_14668,N_12623);
xnor U16079 (N_16079,N_14728,N_12835);
nor U16080 (N_16080,N_14853,N_14421);
nor U16081 (N_16081,N_14076,N_14300);
nor U16082 (N_16082,N_13415,N_14556);
and U16083 (N_16083,N_13601,N_12690);
nand U16084 (N_16084,N_12761,N_13487);
and U16085 (N_16085,N_13939,N_14667);
nor U16086 (N_16086,N_14126,N_12635);
nand U16087 (N_16087,N_13002,N_13460);
or U16088 (N_16088,N_14817,N_13097);
nor U16089 (N_16089,N_14424,N_13857);
and U16090 (N_16090,N_14419,N_13541);
and U16091 (N_16091,N_13944,N_12950);
xnor U16092 (N_16092,N_12968,N_13493);
xor U16093 (N_16093,N_14143,N_12938);
nor U16094 (N_16094,N_13295,N_13268);
and U16095 (N_16095,N_14303,N_14339);
nand U16096 (N_16096,N_12901,N_13138);
nand U16097 (N_16097,N_13488,N_13333);
xor U16098 (N_16098,N_12798,N_12548);
nand U16099 (N_16099,N_12754,N_13683);
nand U16100 (N_16100,N_14809,N_12893);
nand U16101 (N_16101,N_13393,N_13575);
and U16102 (N_16102,N_14212,N_12818);
nor U16103 (N_16103,N_12913,N_14074);
and U16104 (N_16104,N_12994,N_13221);
nand U16105 (N_16105,N_12732,N_13189);
and U16106 (N_16106,N_12966,N_12789);
xor U16107 (N_16107,N_12503,N_13961);
nor U16108 (N_16108,N_13752,N_14224);
or U16109 (N_16109,N_13115,N_14093);
xnor U16110 (N_16110,N_12517,N_13722);
xnor U16111 (N_16111,N_13822,N_14035);
nor U16112 (N_16112,N_14312,N_14252);
nand U16113 (N_16113,N_14780,N_12922);
nand U16114 (N_16114,N_14220,N_13693);
or U16115 (N_16115,N_14870,N_12751);
and U16116 (N_16116,N_13997,N_12866);
and U16117 (N_16117,N_13589,N_14879);
and U16118 (N_16118,N_14182,N_14880);
or U16119 (N_16119,N_14246,N_14532);
xor U16120 (N_16120,N_14499,N_13685);
xnor U16121 (N_16121,N_14371,N_14091);
or U16122 (N_16122,N_14436,N_14153);
nor U16123 (N_16123,N_12788,N_14767);
or U16124 (N_16124,N_14959,N_13842);
xnor U16125 (N_16125,N_12666,N_14952);
and U16126 (N_16126,N_14542,N_12746);
nor U16127 (N_16127,N_14033,N_14311);
nor U16128 (N_16128,N_14319,N_12632);
and U16129 (N_16129,N_14745,N_13298);
nor U16130 (N_16130,N_13423,N_14404);
nand U16131 (N_16131,N_14876,N_14121);
and U16132 (N_16132,N_13883,N_13406);
xor U16133 (N_16133,N_13021,N_12892);
or U16134 (N_16134,N_14640,N_14463);
nand U16135 (N_16135,N_12837,N_14708);
xnor U16136 (N_16136,N_14797,N_13513);
nand U16137 (N_16137,N_13804,N_14194);
xnor U16138 (N_16138,N_14261,N_14983);
nor U16139 (N_16139,N_12620,N_13838);
nand U16140 (N_16140,N_13302,N_13211);
nor U16141 (N_16141,N_13833,N_14714);
nand U16142 (N_16142,N_14427,N_14844);
or U16143 (N_16143,N_13419,N_13285);
and U16144 (N_16144,N_13411,N_14979);
and U16145 (N_16145,N_14344,N_12932);
or U16146 (N_16146,N_13367,N_14838);
xnor U16147 (N_16147,N_14449,N_14849);
nor U16148 (N_16148,N_14384,N_14245);
or U16149 (N_16149,N_13718,N_13862);
and U16150 (N_16150,N_13095,N_14630);
nor U16151 (N_16151,N_14836,N_14333);
xor U16152 (N_16152,N_13769,N_14330);
nor U16153 (N_16153,N_13556,N_13854);
nor U16154 (N_16154,N_14988,N_14859);
or U16155 (N_16155,N_13561,N_12854);
xor U16156 (N_16156,N_13391,N_13528);
nor U16157 (N_16157,N_14968,N_12647);
and U16158 (N_16158,N_14874,N_14624);
xor U16159 (N_16159,N_13426,N_12911);
or U16160 (N_16160,N_12558,N_14590);
or U16161 (N_16161,N_14234,N_12896);
nand U16162 (N_16162,N_14089,N_13300);
or U16163 (N_16163,N_13293,N_13402);
xnor U16164 (N_16164,N_13783,N_14593);
or U16165 (N_16165,N_14649,N_14749);
nand U16166 (N_16166,N_14186,N_13390);
or U16167 (N_16167,N_13885,N_13845);
and U16168 (N_16168,N_13533,N_13962);
nor U16169 (N_16169,N_14519,N_13229);
nand U16170 (N_16170,N_14543,N_13579);
xor U16171 (N_16171,N_13172,N_13725);
nand U16172 (N_16172,N_14305,N_12889);
xnor U16173 (N_16173,N_14777,N_12734);
nor U16174 (N_16174,N_14096,N_13051);
nand U16175 (N_16175,N_13573,N_13475);
and U16176 (N_16176,N_13659,N_13303);
nor U16177 (N_16177,N_13765,N_12831);
xor U16178 (N_16178,N_13489,N_13192);
nor U16179 (N_16179,N_14792,N_12879);
xnor U16180 (N_16180,N_12739,N_13369);
nor U16181 (N_16181,N_14443,N_14159);
xor U16182 (N_16182,N_12862,N_13502);
and U16183 (N_16183,N_12816,N_14396);
xor U16184 (N_16184,N_13637,N_14645);
xor U16185 (N_16185,N_14820,N_14982);
or U16186 (N_16186,N_14275,N_14873);
nand U16187 (N_16187,N_14374,N_12996);
nand U16188 (N_16188,N_14129,N_13755);
nor U16189 (N_16189,N_14205,N_14504);
nor U16190 (N_16190,N_14634,N_14657);
nor U16191 (N_16191,N_13705,N_13871);
and U16192 (N_16192,N_14491,N_14336);
nor U16193 (N_16193,N_13072,N_13724);
xor U16194 (N_16194,N_13050,N_14603);
or U16195 (N_16195,N_13442,N_13252);
nor U16196 (N_16196,N_13454,N_14289);
and U16197 (N_16197,N_13478,N_12522);
or U16198 (N_16198,N_13852,N_13433);
nand U16199 (N_16199,N_14372,N_13624);
nand U16200 (N_16200,N_13154,N_13061);
nand U16201 (N_16201,N_13506,N_14762);
nand U16202 (N_16202,N_14461,N_14839);
and U16203 (N_16203,N_14619,N_13195);
nand U16204 (N_16204,N_12617,N_14024);
or U16205 (N_16205,N_14422,N_12527);
nand U16206 (N_16206,N_13577,N_13713);
nand U16207 (N_16207,N_13815,N_14698);
or U16208 (N_16208,N_14321,N_13464);
nor U16209 (N_16209,N_14429,N_13208);
nor U16210 (N_16210,N_14867,N_14514);
or U16211 (N_16211,N_14985,N_13999);
or U16212 (N_16212,N_12914,N_14016);
nand U16213 (N_16213,N_13187,N_12876);
and U16214 (N_16214,N_13903,N_14878);
or U16215 (N_16215,N_14395,N_13068);
and U16216 (N_16216,N_13355,N_13031);
nand U16217 (N_16217,N_13190,N_12906);
or U16218 (N_16218,N_12555,N_13763);
nand U16219 (N_16219,N_14751,N_12920);
nor U16220 (N_16220,N_13353,N_13305);
or U16221 (N_16221,N_14392,N_14818);
nor U16222 (N_16222,N_14200,N_14534);
nand U16223 (N_16223,N_13667,N_14002);
and U16224 (N_16224,N_12574,N_14079);
or U16225 (N_16225,N_14315,N_14387);
nand U16226 (N_16226,N_14729,N_13823);
or U16227 (N_16227,N_14672,N_13440);
nand U16228 (N_16228,N_14306,N_14115);
nor U16229 (N_16229,N_12759,N_14604);
nor U16230 (N_16230,N_12662,N_13081);
and U16231 (N_16231,N_13899,N_14805);
nand U16232 (N_16232,N_14829,N_14717);
or U16233 (N_16233,N_13457,N_14225);
xor U16234 (N_16234,N_13320,N_12673);
and U16235 (N_16235,N_12608,N_12626);
or U16236 (N_16236,N_13853,N_12848);
or U16237 (N_16237,N_14609,N_14467);
nor U16238 (N_16238,N_13583,N_13509);
nor U16239 (N_16239,N_13549,N_12649);
or U16240 (N_16240,N_13235,N_14445);
xor U16241 (N_16241,N_14782,N_12707);
nor U16242 (N_16242,N_13696,N_14272);
or U16243 (N_16243,N_14059,N_13091);
or U16244 (N_16244,N_13820,N_14149);
and U16245 (N_16245,N_14522,N_13503);
xor U16246 (N_16246,N_13728,N_12851);
or U16247 (N_16247,N_14652,N_14852);
nor U16248 (N_16248,N_13498,N_14350);
or U16249 (N_16249,N_14712,N_14458);
nor U16250 (N_16250,N_13091,N_13568);
nand U16251 (N_16251,N_14442,N_14166);
xor U16252 (N_16252,N_14996,N_13005);
nor U16253 (N_16253,N_13843,N_14128);
xor U16254 (N_16254,N_13237,N_14844);
or U16255 (N_16255,N_12688,N_14783);
xnor U16256 (N_16256,N_13396,N_12569);
xnor U16257 (N_16257,N_14327,N_14750);
and U16258 (N_16258,N_13964,N_13168);
nor U16259 (N_16259,N_13562,N_13725);
or U16260 (N_16260,N_13670,N_12982);
or U16261 (N_16261,N_14443,N_13244);
nor U16262 (N_16262,N_14311,N_13540);
xnor U16263 (N_16263,N_14993,N_12553);
or U16264 (N_16264,N_14038,N_14519);
and U16265 (N_16265,N_14131,N_14386);
or U16266 (N_16266,N_14687,N_14880);
or U16267 (N_16267,N_13142,N_14195);
or U16268 (N_16268,N_13578,N_12876);
nor U16269 (N_16269,N_13674,N_13198);
xor U16270 (N_16270,N_14937,N_13268);
nand U16271 (N_16271,N_13147,N_13018);
nor U16272 (N_16272,N_12776,N_14757);
or U16273 (N_16273,N_14514,N_14120);
xor U16274 (N_16274,N_14512,N_14609);
nor U16275 (N_16275,N_14531,N_14907);
nand U16276 (N_16276,N_13532,N_13200);
and U16277 (N_16277,N_13148,N_13347);
and U16278 (N_16278,N_13767,N_12828);
nand U16279 (N_16279,N_14289,N_12806);
nand U16280 (N_16280,N_13990,N_12566);
and U16281 (N_16281,N_12901,N_14125);
nor U16282 (N_16282,N_14446,N_12996);
xnor U16283 (N_16283,N_13865,N_13217);
xnor U16284 (N_16284,N_13137,N_12904);
or U16285 (N_16285,N_13990,N_12929);
xor U16286 (N_16286,N_14173,N_14998);
nor U16287 (N_16287,N_14037,N_12564);
and U16288 (N_16288,N_13282,N_14262);
or U16289 (N_16289,N_13195,N_12683);
or U16290 (N_16290,N_14223,N_14320);
and U16291 (N_16291,N_14920,N_13758);
xnor U16292 (N_16292,N_14009,N_14904);
xnor U16293 (N_16293,N_13002,N_14847);
nor U16294 (N_16294,N_13449,N_13536);
or U16295 (N_16295,N_12531,N_13929);
and U16296 (N_16296,N_14529,N_14891);
nor U16297 (N_16297,N_13661,N_13778);
nor U16298 (N_16298,N_12573,N_14266);
and U16299 (N_16299,N_12959,N_12703);
nand U16300 (N_16300,N_14347,N_12766);
or U16301 (N_16301,N_13385,N_12641);
nor U16302 (N_16302,N_14359,N_14451);
nor U16303 (N_16303,N_12961,N_13682);
and U16304 (N_16304,N_13031,N_13486);
or U16305 (N_16305,N_14162,N_14546);
xor U16306 (N_16306,N_14819,N_13377);
or U16307 (N_16307,N_13863,N_14422);
and U16308 (N_16308,N_14242,N_13643);
xor U16309 (N_16309,N_13206,N_13858);
nor U16310 (N_16310,N_13150,N_13937);
and U16311 (N_16311,N_12583,N_12762);
nor U16312 (N_16312,N_14760,N_12574);
nand U16313 (N_16313,N_13232,N_14064);
xnor U16314 (N_16314,N_13306,N_13586);
and U16315 (N_16315,N_13168,N_13342);
nand U16316 (N_16316,N_13718,N_14386);
nand U16317 (N_16317,N_14361,N_14773);
or U16318 (N_16318,N_14113,N_13122);
nand U16319 (N_16319,N_13041,N_12668);
xor U16320 (N_16320,N_14974,N_14876);
xnor U16321 (N_16321,N_14167,N_13436);
nor U16322 (N_16322,N_13647,N_14650);
nor U16323 (N_16323,N_12766,N_13421);
nand U16324 (N_16324,N_13025,N_13584);
xnor U16325 (N_16325,N_13639,N_12561);
and U16326 (N_16326,N_13809,N_14117);
and U16327 (N_16327,N_14151,N_14900);
nor U16328 (N_16328,N_12630,N_14746);
and U16329 (N_16329,N_13028,N_12910);
and U16330 (N_16330,N_12841,N_13705);
nor U16331 (N_16331,N_14806,N_13941);
nand U16332 (N_16332,N_13687,N_12769);
or U16333 (N_16333,N_14641,N_14800);
xnor U16334 (N_16334,N_13275,N_14332);
nand U16335 (N_16335,N_13644,N_13642);
nand U16336 (N_16336,N_12692,N_14240);
nor U16337 (N_16337,N_13570,N_14577);
nand U16338 (N_16338,N_13454,N_14315);
nand U16339 (N_16339,N_14260,N_13602);
nand U16340 (N_16340,N_13353,N_12844);
nand U16341 (N_16341,N_14907,N_12635);
and U16342 (N_16342,N_14668,N_13650);
and U16343 (N_16343,N_14359,N_14733);
nand U16344 (N_16344,N_12739,N_12972);
nor U16345 (N_16345,N_14173,N_14838);
and U16346 (N_16346,N_12810,N_14266);
nor U16347 (N_16347,N_12501,N_12575);
xor U16348 (N_16348,N_13994,N_14907);
and U16349 (N_16349,N_14820,N_14707);
nand U16350 (N_16350,N_14422,N_13085);
and U16351 (N_16351,N_12649,N_14538);
nand U16352 (N_16352,N_14986,N_14319);
and U16353 (N_16353,N_12647,N_13330);
and U16354 (N_16354,N_13676,N_14979);
nor U16355 (N_16355,N_14294,N_14300);
or U16356 (N_16356,N_13139,N_13706);
and U16357 (N_16357,N_12898,N_12772);
nand U16358 (N_16358,N_14368,N_14401);
xnor U16359 (N_16359,N_14847,N_13970);
nand U16360 (N_16360,N_14517,N_12798);
and U16361 (N_16361,N_14031,N_12809);
and U16362 (N_16362,N_14042,N_12692);
xor U16363 (N_16363,N_14277,N_14261);
nand U16364 (N_16364,N_14104,N_14936);
nor U16365 (N_16365,N_14035,N_14690);
nor U16366 (N_16366,N_13660,N_13632);
nor U16367 (N_16367,N_14182,N_14871);
or U16368 (N_16368,N_13353,N_14524);
nand U16369 (N_16369,N_14617,N_14797);
nor U16370 (N_16370,N_14915,N_13941);
and U16371 (N_16371,N_12878,N_13581);
xor U16372 (N_16372,N_14298,N_14747);
nand U16373 (N_16373,N_12968,N_14535);
nand U16374 (N_16374,N_12797,N_14110);
nand U16375 (N_16375,N_13717,N_13098);
and U16376 (N_16376,N_13453,N_12731);
nand U16377 (N_16377,N_12977,N_14478);
nor U16378 (N_16378,N_14697,N_13976);
nand U16379 (N_16379,N_14020,N_14360);
nor U16380 (N_16380,N_13598,N_13836);
and U16381 (N_16381,N_14335,N_14546);
nand U16382 (N_16382,N_13054,N_13659);
or U16383 (N_16383,N_14895,N_13292);
nor U16384 (N_16384,N_13302,N_14751);
and U16385 (N_16385,N_14305,N_13902);
nand U16386 (N_16386,N_13422,N_13714);
nand U16387 (N_16387,N_12894,N_13840);
or U16388 (N_16388,N_14891,N_14241);
or U16389 (N_16389,N_14069,N_12767);
nand U16390 (N_16390,N_13882,N_13552);
nor U16391 (N_16391,N_14561,N_14605);
nor U16392 (N_16392,N_13811,N_13660);
xnor U16393 (N_16393,N_13051,N_13455);
xor U16394 (N_16394,N_13758,N_14962);
nand U16395 (N_16395,N_14256,N_13092);
or U16396 (N_16396,N_12817,N_12544);
xor U16397 (N_16397,N_13244,N_13340);
or U16398 (N_16398,N_12670,N_13186);
xor U16399 (N_16399,N_13790,N_13737);
nor U16400 (N_16400,N_13088,N_12822);
nand U16401 (N_16401,N_14682,N_14848);
nor U16402 (N_16402,N_13037,N_13725);
and U16403 (N_16403,N_12914,N_14443);
or U16404 (N_16404,N_13304,N_14007);
nor U16405 (N_16405,N_12808,N_13220);
and U16406 (N_16406,N_13246,N_13602);
and U16407 (N_16407,N_14119,N_14597);
nand U16408 (N_16408,N_14071,N_13418);
nor U16409 (N_16409,N_14433,N_14778);
or U16410 (N_16410,N_14266,N_14977);
nor U16411 (N_16411,N_14525,N_13534);
xnor U16412 (N_16412,N_14529,N_14985);
nand U16413 (N_16413,N_12742,N_13272);
xor U16414 (N_16414,N_13767,N_12692);
nor U16415 (N_16415,N_14270,N_13235);
or U16416 (N_16416,N_14036,N_14223);
or U16417 (N_16417,N_14893,N_14456);
and U16418 (N_16418,N_12646,N_13371);
nand U16419 (N_16419,N_12806,N_14612);
nand U16420 (N_16420,N_12939,N_14009);
xor U16421 (N_16421,N_13781,N_13170);
nor U16422 (N_16422,N_13843,N_13277);
or U16423 (N_16423,N_14169,N_14974);
nor U16424 (N_16424,N_14444,N_12998);
nand U16425 (N_16425,N_12801,N_13954);
nor U16426 (N_16426,N_12811,N_13906);
and U16427 (N_16427,N_12807,N_14765);
xor U16428 (N_16428,N_13098,N_13038);
xor U16429 (N_16429,N_12773,N_13394);
and U16430 (N_16430,N_13371,N_13773);
nand U16431 (N_16431,N_14247,N_14883);
nand U16432 (N_16432,N_14903,N_13098);
nand U16433 (N_16433,N_13811,N_14546);
nor U16434 (N_16434,N_13954,N_14792);
xor U16435 (N_16435,N_13993,N_13130);
xnor U16436 (N_16436,N_13761,N_12616);
nor U16437 (N_16437,N_13104,N_13002);
nor U16438 (N_16438,N_12781,N_14893);
and U16439 (N_16439,N_14150,N_14021);
or U16440 (N_16440,N_13432,N_13998);
nor U16441 (N_16441,N_12714,N_12904);
or U16442 (N_16442,N_13427,N_13972);
nor U16443 (N_16443,N_14477,N_13488);
or U16444 (N_16444,N_14184,N_14883);
xor U16445 (N_16445,N_14868,N_13751);
nor U16446 (N_16446,N_12621,N_14222);
or U16447 (N_16447,N_14465,N_13398);
nand U16448 (N_16448,N_13282,N_14813);
or U16449 (N_16449,N_14954,N_12629);
and U16450 (N_16450,N_13479,N_14083);
or U16451 (N_16451,N_14439,N_12918);
nor U16452 (N_16452,N_12655,N_13768);
or U16453 (N_16453,N_13126,N_14572);
or U16454 (N_16454,N_13901,N_14981);
nand U16455 (N_16455,N_14190,N_13613);
xnor U16456 (N_16456,N_14930,N_14872);
nor U16457 (N_16457,N_12787,N_13427);
or U16458 (N_16458,N_14815,N_14768);
xnor U16459 (N_16459,N_12641,N_14682);
or U16460 (N_16460,N_13375,N_14239);
xnor U16461 (N_16461,N_13485,N_13448);
and U16462 (N_16462,N_14508,N_13626);
or U16463 (N_16463,N_12617,N_14600);
and U16464 (N_16464,N_13713,N_14315);
nor U16465 (N_16465,N_13037,N_13738);
xor U16466 (N_16466,N_12884,N_13232);
nand U16467 (N_16467,N_13634,N_14620);
or U16468 (N_16468,N_13567,N_14953);
and U16469 (N_16469,N_14677,N_13417);
nor U16470 (N_16470,N_13029,N_12790);
nor U16471 (N_16471,N_14930,N_14678);
xor U16472 (N_16472,N_14932,N_13362);
xor U16473 (N_16473,N_14520,N_14340);
and U16474 (N_16474,N_12798,N_12910);
and U16475 (N_16475,N_13264,N_13825);
nor U16476 (N_16476,N_14724,N_13559);
nor U16477 (N_16477,N_14112,N_14578);
and U16478 (N_16478,N_14161,N_13132);
and U16479 (N_16479,N_12917,N_12918);
and U16480 (N_16480,N_13537,N_14206);
xor U16481 (N_16481,N_13805,N_13470);
xnor U16482 (N_16482,N_13848,N_14176);
xnor U16483 (N_16483,N_13300,N_14471);
and U16484 (N_16484,N_12785,N_13667);
xor U16485 (N_16485,N_13364,N_13062);
or U16486 (N_16486,N_12730,N_12680);
nand U16487 (N_16487,N_13221,N_14525);
or U16488 (N_16488,N_14003,N_14377);
xnor U16489 (N_16489,N_13125,N_14941);
nand U16490 (N_16490,N_14203,N_14957);
nand U16491 (N_16491,N_14919,N_14459);
nor U16492 (N_16492,N_14127,N_14935);
nand U16493 (N_16493,N_14250,N_12807);
and U16494 (N_16494,N_13867,N_14739);
nor U16495 (N_16495,N_14334,N_14103);
nand U16496 (N_16496,N_13032,N_13594);
nor U16497 (N_16497,N_13715,N_12571);
nand U16498 (N_16498,N_13261,N_14637);
nand U16499 (N_16499,N_14215,N_14743);
xor U16500 (N_16500,N_13092,N_12818);
or U16501 (N_16501,N_14295,N_13229);
nand U16502 (N_16502,N_12559,N_13888);
xor U16503 (N_16503,N_12740,N_13518);
nand U16504 (N_16504,N_13458,N_14586);
or U16505 (N_16505,N_14830,N_13739);
nor U16506 (N_16506,N_13725,N_12532);
or U16507 (N_16507,N_14224,N_14876);
or U16508 (N_16508,N_14369,N_12866);
nand U16509 (N_16509,N_14686,N_13127);
nand U16510 (N_16510,N_13118,N_12510);
and U16511 (N_16511,N_13411,N_14002);
and U16512 (N_16512,N_14625,N_12969);
nand U16513 (N_16513,N_13567,N_12852);
nor U16514 (N_16514,N_13462,N_13854);
and U16515 (N_16515,N_12874,N_14347);
nand U16516 (N_16516,N_13809,N_12929);
xnor U16517 (N_16517,N_14918,N_12520);
nor U16518 (N_16518,N_14720,N_12569);
nand U16519 (N_16519,N_13839,N_13981);
and U16520 (N_16520,N_13232,N_13686);
nand U16521 (N_16521,N_14229,N_13733);
xnor U16522 (N_16522,N_14939,N_14634);
and U16523 (N_16523,N_13712,N_13436);
and U16524 (N_16524,N_14118,N_13786);
and U16525 (N_16525,N_13740,N_13157);
xnor U16526 (N_16526,N_14583,N_13049);
xor U16527 (N_16527,N_13557,N_14346);
nand U16528 (N_16528,N_13205,N_12787);
and U16529 (N_16529,N_14988,N_12685);
nor U16530 (N_16530,N_13008,N_12656);
nand U16531 (N_16531,N_14379,N_13268);
nor U16532 (N_16532,N_13249,N_13515);
xor U16533 (N_16533,N_13861,N_14470);
nor U16534 (N_16534,N_13949,N_14805);
nor U16535 (N_16535,N_14940,N_13179);
or U16536 (N_16536,N_14748,N_12962);
or U16537 (N_16537,N_13502,N_12513);
xor U16538 (N_16538,N_14239,N_14558);
nand U16539 (N_16539,N_14363,N_14003);
nor U16540 (N_16540,N_13767,N_13802);
nor U16541 (N_16541,N_13710,N_13947);
nor U16542 (N_16542,N_13887,N_13448);
xor U16543 (N_16543,N_14368,N_12999);
xor U16544 (N_16544,N_12534,N_14865);
nand U16545 (N_16545,N_12923,N_12917);
xor U16546 (N_16546,N_14728,N_14398);
xnor U16547 (N_16547,N_12514,N_14184);
xor U16548 (N_16548,N_14356,N_14757);
xnor U16549 (N_16549,N_14077,N_14307);
and U16550 (N_16550,N_14765,N_14280);
or U16551 (N_16551,N_14731,N_14873);
or U16552 (N_16552,N_12799,N_14805);
and U16553 (N_16553,N_12914,N_14741);
xnor U16554 (N_16554,N_14489,N_14107);
nor U16555 (N_16555,N_14651,N_13500);
and U16556 (N_16556,N_13615,N_13026);
or U16557 (N_16557,N_12798,N_14392);
and U16558 (N_16558,N_13842,N_12514);
xor U16559 (N_16559,N_13153,N_13520);
or U16560 (N_16560,N_13938,N_14250);
xnor U16561 (N_16561,N_14106,N_14144);
nand U16562 (N_16562,N_14950,N_13397);
xor U16563 (N_16563,N_14505,N_14250);
and U16564 (N_16564,N_12809,N_12826);
nor U16565 (N_16565,N_13620,N_14051);
and U16566 (N_16566,N_14288,N_13749);
and U16567 (N_16567,N_12651,N_12959);
nor U16568 (N_16568,N_13064,N_13276);
xnor U16569 (N_16569,N_14494,N_13489);
nand U16570 (N_16570,N_12514,N_14632);
xnor U16571 (N_16571,N_13673,N_12834);
xor U16572 (N_16572,N_14712,N_14260);
nand U16573 (N_16573,N_14706,N_13091);
or U16574 (N_16574,N_13372,N_13718);
nand U16575 (N_16575,N_12714,N_12779);
or U16576 (N_16576,N_12906,N_13565);
and U16577 (N_16577,N_14401,N_13366);
xor U16578 (N_16578,N_14245,N_14666);
nor U16579 (N_16579,N_13591,N_12524);
or U16580 (N_16580,N_13689,N_14746);
xnor U16581 (N_16581,N_12817,N_14837);
xor U16582 (N_16582,N_14828,N_13659);
nor U16583 (N_16583,N_13354,N_14064);
or U16584 (N_16584,N_12832,N_14419);
and U16585 (N_16585,N_14078,N_13904);
and U16586 (N_16586,N_14746,N_13343);
nor U16587 (N_16587,N_13718,N_13594);
nand U16588 (N_16588,N_13897,N_12825);
nand U16589 (N_16589,N_12800,N_14525);
nand U16590 (N_16590,N_12748,N_13321);
xnor U16591 (N_16591,N_14646,N_14639);
or U16592 (N_16592,N_13179,N_14713);
nand U16593 (N_16593,N_14870,N_12679);
and U16594 (N_16594,N_14110,N_14958);
xnor U16595 (N_16595,N_14282,N_13927);
or U16596 (N_16596,N_13678,N_12943);
nor U16597 (N_16597,N_12624,N_12609);
or U16598 (N_16598,N_14078,N_13680);
nor U16599 (N_16599,N_14374,N_13837);
or U16600 (N_16600,N_14492,N_13951);
and U16601 (N_16601,N_13160,N_13573);
or U16602 (N_16602,N_14473,N_14983);
nor U16603 (N_16603,N_14560,N_14344);
nor U16604 (N_16604,N_12800,N_14206);
nor U16605 (N_16605,N_14505,N_13283);
nor U16606 (N_16606,N_14964,N_13021);
nor U16607 (N_16607,N_13384,N_13953);
nand U16608 (N_16608,N_14915,N_13176);
or U16609 (N_16609,N_14791,N_13321);
xnor U16610 (N_16610,N_14730,N_12931);
or U16611 (N_16611,N_14648,N_13410);
xnor U16612 (N_16612,N_12577,N_13322);
and U16613 (N_16613,N_14617,N_14049);
xnor U16614 (N_16614,N_13093,N_13483);
xor U16615 (N_16615,N_13776,N_14786);
nand U16616 (N_16616,N_13067,N_12800);
nor U16617 (N_16617,N_14760,N_14746);
and U16618 (N_16618,N_14131,N_13749);
or U16619 (N_16619,N_12555,N_12884);
or U16620 (N_16620,N_14672,N_12817);
nand U16621 (N_16621,N_13864,N_13615);
nor U16622 (N_16622,N_13444,N_14656);
nand U16623 (N_16623,N_14706,N_14292);
nor U16624 (N_16624,N_14113,N_13688);
nor U16625 (N_16625,N_13857,N_13334);
nor U16626 (N_16626,N_12938,N_12702);
or U16627 (N_16627,N_12838,N_12966);
or U16628 (N_16628,N_13152,N_14642);
or U16629 (N_16629,N_14350,N_13188);
and U16630 (N_16630,N_12845,N_14240);
and U16631 (N_16631,N_14220,N_14743);
nand U16632 (N_16632,N_13777,N_13417);
nor U16633 (N_16633,N_14989,N_14289);
nor U16634 (N_16634,N_14113,N_12894);
nor U16635 (N_16635,N_13996,N_13024);
nor U16636 (N_16636,N_13511,N_14750);
xnor U16637 (N_16637,N_14788,N_14263);
nand U16638 (N_16638,N_12646,N_14276);
nand U16639 (N_16639,N_12551,N_14956);
and U16640 (N_16640,N_14855,N_13107);
or U16641 (N_16641,N_12856,N_13016);
xnor U16642 (N_16642,N_12546,N_13616);
xor U16643 (N_16643,N_13574,N_12672);
or U16644 (N_16644,N_13699,N_12925);
and U16645 (N_16645,N_13908,N_14420);
nand U16646 (N_16646,N_13624,N_13470);
nand U16647 (N_16647,N_14200,N_13595);
nand U16648 (N_16648,N_13078,N_14485);
or U16649 (N_16649,N_12609,N_13373);
nand U16650 (N_16650,N_14076,N_12902);
and U16651 (N_16651,N_13428,N_14782);
or U16652 (N_16652,N_14495,N_12723);
and U16653 (N_16653,N_14217,N_13486);
nand U16654 (N_16654,N_13782,N_14089);
nor U16655 (N_16655,N_14086,N_13848);
nor U16656 (N_16656,N_13283,N_14698);
or U16657 (N_16657,N_14512,N_14518);
or U16658 (N_16658,N_14888,N_12713);
nand U16659 (N_16659,N_13173,N_14423);
or U16660 (N_16660,N_13744,N_12610);
and U16661 (N_16661,N_13836,N_14867);
or U16662 (N_16662,N_13400,N_14562);
nor U16663 (N_16663,N_14965,N_13697);
or U16664 (N_16664,N_13242,N_14454);
xor U16665 (N_16665,N_14325,N_13052);
xnor U16666 (N_16666,N_12928,N_12649);
nand U16667 (N_16667,N_13321,N_12684);
nor U16668 (N_16668,N_13424,N_14118);
and U16669 (N_16669,N_13090,N_13857);
xor U16670 (N_16670,N_14512,N_14921);
and U16671 (N_16671,N_13820,N_14961);
or U16672 (N_16672,N_14050,N_14479);
or U16673 (N_16673,N_14051,N_14330);
nand U16674 (N_16674,N_13455,N_14106);
nor U16675 (N_16675,N_14738,N_13834);
xnor U16676 (N_16676,N_14510,N_14707);
nand U16677 (N_16677,N_14546,N_13254);
nand U16678 (N_16678,N_12905,N_13701);
or U16679 (N_16679,N_13907,N_14738);
and U16680 (N_16680,N_13786,N_12673);
xor U16681 (N_16681,N_14672,N_13760);
xnor U16682 (N_16682,N_14386,N_13519);
xor U16683 (N_16683,N_13805,N_13036);
nand U16684 (N_16684,N_13797,N_13402);
and U16685 (N_16685,N_13940,N_14982);
nor U16686 (N_16686,N_14981,N_13065);
or U16687 (N_16687,N_13196,N_13580);
or U16688 (N_16688,N_12874,N_14392);
nand U16689 (N_16689,N_12869,N_14662);
and U16690 (N_16690,N_13198,N_13891);
nor U16691 (N_16691,N_13537,N_12804);
nor U16692 (N_16692,N_13997,N_13348);
and U16693 (N_16693,N_14293,N_13731);
and U16694 (N_16694,N_14902,N_14968);
and U16695 (N_16695,N_13628,N_14710);
xnor U16696 (N_16696,N_12919,N_14207);
and U16697 (N_16697,N_14746,N_13833);
and U16698 (N_16698,N_12937,N_13491);
and U16699 (N_16699,N_13613,N_14624);
xor U16700 (N_16700,N_12803,N_14184);
nand U16701 (N_16701,N_14581,N_14727);
and U16702 (N_16702,N_13764,N_12993);
xnor U16703 (N_16703,N_14142,N_13733);
or U16704 (N_16704,N_14622,N_12819);
or U16705 (N_16705,N_13495,N_13494);
or U16706 (N_16706,N_14354,N_14336);
and U16707 (N_16707,N_14820,N_13593);
and U16708 (N_16708,N_14190,N_12535);
or U16709 (N_16709,N_12751,N_14989);
xor U16710 (N_16710,N_14284,N_14503);
xnor U16711 (N_16711,N_13020,N_12838);
nand U16712 (N_16712,N_14790,N_14789);
xnor U16713 (N_16713,N_13054,N_13930);
and U16714 (N_16714,N_14299,N_13467);
nand U16715 (N_16715,N_14747,N_13642);
nor U16716 (N_16716,N_12675,N_13204);
nor U16717 (N_16717,N_13031,N_14643);
nand U16718 (N_16718,N_12691,N_14620);
and U16719 (N_16719,N_14471,N_14396);
xnor U16720 (N_16720,N_14986,N_14619);
nor U16721 (N_16721,N_13610,N_14054);
nor U16722 (N_16722,N_14007,N_13721);
nor U16723 (N_16723,N_14792,N_14671);
xnor U16724 (N_16724,N_13043,N_13638);
or U16725 (N_16725,N_14679,N_12921);
or U16726 (N_16726,N_13707,N_14748);
and U16727 (N_16727,N_13683,N_12628);
or U16728 (N_16728,N_13872,N_14891);
nand U16729 (N_16729,N_13940,N_13773);
xnor U16730 (N_16730,N_12826,N_13784);
nand U16731 (N_16731,N_12843,N_12900);
xnor U16732 (N_16732,N_14428,N_14271);
nor U16733 (N_16733,N_14651,N_13123);
or U16734 (N_16734,N_13699,N_14432);
nor U16735 (N_16735,N_13104,N_13496);
and U16736 (N_16736,N_13903,N_14294);
nor U16737 (N_16737,N_12856,N_13961);
nand U16738 (N_16738,N_14617,N_13166);
nor U16739 (N_16739,N_14032,N_12907);
nand U16740 (N_16740,N_13564,N_13583);
or U16741 (N_16741,N_14228,N_13348);
xor U16742 (N_16742,N_14508,N_12541);
nand U16743 (N_16743,N_14040,N_14132);
or U16744 (N_16744,N_13164,N_12504);
and U16745 (N_16745,N_14781,N_12661);
or U16746 (N_16746,N_13864,N_14686);
nor U16747 (N_16747,N_12600,N_13577);
nor U16748 (N_16748,N_12701,N_12616);
xor U16749 (N_16749,N_12819,N_13068);
nand U16750 (N_16750,N_14082,N_13924);
nor U16751 (N_16751,N_12629,N_12787);
nor U16752 (N_16752,N_13051,N_12808);
or U16753 (N_16753,N_14671,N_13285);
xor U16754 (N_16754,N_13173,N_12908);
or U16755 (N_16755,N_14555,N_14300);
nand U16756 (N_16756,N_13106,N_14859);
nor U16757 (N_16757,N_14934,N_14861);
nand U16758 (N_16758,N_13708,N_13058);
xnor U16759 (N_16759,N_14991,N_13946);
nor U16760 (N_16760,N_14064,N_14909);
or U16761 (N_16761,N_13757,N_14452);
nor U16762 (N_16762,N_14472,N_12561);
nor U16763 (N_16763,N_14112,N_13530);
nor U16764 (N_16764,N_14537,N_14884);
nor U16765 (N_16765,N_13178,N_13904);
nor U16766 (N_16766,N_14531,N_13137);
xnor U16767 (N_16767,N_14015,N_14351);
nor U16768 (N_16768,N_12506,N_13927);
xor U16769 (N_16769,N_14016,N_12679);
xnor U16770 (N_16770,N_14394,N_14969);
or U16771 (N_16771,N_12816,N_13459);
and U16772 (N_16772,N_14025,N_13802);
nand U16773 (N_16773,N_14775,N_12731);
and U16774 (N_16774,N_14430,N_14209);
and U16775 (N_16775,N_13670,N_14812);
nor U16776 (N_16776,N_13984,N_14384);
or U16777 (N_16777,N_12806,N_13297);
nand U16778 (N_16778,N_13539,N_14486);
xnor U16779 (N_16779,N_13822,N_12658);
xor U16780 (N_16780,N_13377,N_14787);
nor U16781 (N_16781,N_13339,N_14650);
or U16782 (N_16782,N_13946,N_13699);
xor U16783 (N_16783,N_13903,N_13058);
xnor U16784 (N_16784,N_13888,N_14995);
nor U16785 (N_16785,N_13943,N_14637);
or U16786 (N_16786,N_14744,N_13221);
and U16787 (N_16787,N_13335,N_14374);
nor U16788 (N_16788,N_13990,N_12737);
or U16789 (N_16789,N_13611,N_14671);
xnor U16790 (N_16790,N_14732,N_13556);
xor U16791 (N_16791,N_14115,N_13827);
and U16792 (N_16792,N_13687,N_13627);
or U16793 (N_16793,N_12517,N_14882);
nor U16794 (N_16794,N_14410,N_13295);
and U16795 (N_16795,N_13147,N_12603);
xor U16796 (N_16796,N_13733,N_14413);
nor U16797 (N_16797,N_14787,N_14526);
and U16798 (N_16798,N_13674,N_14353);
xor U16799 (N_16799,N_13303,N_13373);
xor U16800 (N_16800,N_12597,N_14856);
nand U16801 (N_16801,N_14032,N_13124);
nor U16802 (N_16802,N_14591,N_14399);
or U16803 (N_16803,N_14691,N_12860);
or U16804 (N_16804,N_13292,N_13182);
nand U16805 (N_16805,N_12784,N_13808);
nand U16806 (N_16806,N_14111,N_12804);
and U16807 (N_16807,N_14825,N_14270);
and U16808 (N_16808,N_13436,N_12546);
nand U16809 (N_16809,N_13775,N_14379);
or U16810 (N_16810,N_14297,N_14777);
nor U16811 (N_16811,N_12797,N_12895);
and U16812 (N_16812,N_14432,N_14306);
or U16813 (N_16813,N_13596,N_14664);
xnor U16814 (N_16814,N_14175,N_13978);
nand U16815 (N_16815,N_13915,N_12560);
or U16816 (N_16816,N_14399,N_13764);
nand U16817 (N_16817,N_14126,N_13406);
and U16818 (N_16818,N_12600,N_14155);
xnor U16819 (N_16819,N_14031,N_14095);
and U16820 (N_16820,N_14572,N_12671);
and U16821 (N_16821,N_12912,N_12817);
xor U16822 (N_16822,N_13848,N_13895);
nor U16823 (N_16823,N_13426,N_14757);
nand U16824 (N_16824,N_13831,N_14655);
xor U16825 (N_16825,N_14125,N_12850);
nor U16826 (N_16826,N_14462,N_12699);
or U16827 (N_16827,N_14414,N_13140);
and U16828 (N_16828,N_13521,N_14012);
and U16829 (N_16829,N_13408,N_12786);
xor U16830 (N_16830,N_12891,N_13707);
nand U16831 (N_16831,N_14270,N_13926);
and U16832 (N_16832,N_14522,N_13933);
nand U16833 (N_16833,N_13251,N_14584);
and U16834 (N_16834,N_12732,N_13086);
nand U16835 (N_16835,N_12691,N_12857);
nor U16836 (N_16836,N_14287,N_14893);
nand U16837 (N_16837,N_12948,N_14855);
nand U16838 (N_16838,N_13465,N_14058);
and U16839 (N_16839,N_13691,N_14319);
and U16840 (N_16840,N_14152,N_14527);
or U16841 (N_16841,N_13391,N_14387);
nor U16842 (N_16842,N_13784,N_12870);
nand U16843 (N_16843,N_13019,N_14747);
nor U16844 (N_16844,N_13175,N_14154);
and U16845 (N_16845,N_13159,N_12599);
and U16846 (N_16846,N_13993,N_14119);
nand U16847 (N_16847,N_14549,N_14731);
or U16848 (N_16848,N_13553,N_13629);
or U16849 (N_16849,N_14827,N_13749);
and U16850 (N_16850,N_12554,N_13601);
and U16851 (N_16851,N_12646,N_14017);
and U16852 (N_16852,N_12955,N_12740);
nand U16853 (N_16853,N_14772,N_13278);
or U16854 (N_16854,N_13251,N_14388);
or U16855 (N_16855,N_12944,N_14854);
and U16856 (N_16856,N_14204,N_13843);
and U16857 (N_16857,N_13446,N_12852);
nor U16858 (N_16858,N_14991,N_14786);
and U16859 (N_16859,N_14892,N_13882);
or U16860 (N_16860,N_13508,N_13421);
xor U16861 (N_16861,N_12985,N_14360);
nand U16862 (N_16862,N_13107,N_14132);
or U16863 (N_16863,N_14281,N_13233);
xnor U16864 (N_16864,N_14786,N_14874);
or U16865 (N_16865,N_12944,N_13879);
xnor U16866 (N_16866,N_13185,N_14408);
or U16867 (N_16867,N_14616,N_14088);
nand U16868 (N_16868,N_14266,N_13829);
and U16869 (N_16869,N_14504,N_14154);
nor U16870 (N_16870,N_12749,N_13205);
nor U16871 (N_16871,N_12814,N_13857);
or U16872 (N_16872,N_14485,N_13581);
or U16873 (N_16873,N_13504,N_14987);
or U16874 (N_16874,N_12617,N_14267);
or U16875 (N_16875,N_13978,N_13431);
xnor U16876 (N_16876,N_14413,N_12825);
or U16877 (N_16877,N_13815,N_13307);
xnor U16878 (N_16878,N_13842,N_12574);
xnor U16879 (N_16879,N_13977,N_12945);
or U16880 (N_16880,N_13605,N_12615);
nand U16881 (N_16881,N_14154,N_12661);
nand U16882 (N_16882,N_13369,N_12613);
nand U16883 (N_16883,N_14674,N_13057);
nand U16884 (N_16884,N_14390,N_13017);
nand U16885 (N_16885,N_14635,N_14158);
nor U16886 (N_16886,N_13301,N_14070);
and U16887 (N_16887,N_14510,N_14999);
or U16888 (N_16888,N_12807,N_12880);
or U16889 (N_16889,N_12931,N_14999);
xnor U16890 (N_16890,N_14950,N_13913);
nor U16891 (N_16891,N_13130,N_13707);
or U16892 (N_16892,N_12864,N_12512);
or U16893 (N_16893,N_14338,N_14543);
and U16894 (N_16894,N_14178,N_13984);
xor U16895 (N_16895,N_14616,N_13285);
and U16896 (N_16896,N_14658,N_13440);
or U16897 (N_16897,N_14352,N_13547);
xnor U16898 (N_16898,N_14204,N_13964);
or U16899 (N_16899,N_14709,N_12943);
nor U16900 (N_16900,N_14895,N_14102);
xnor U16901 (N_16901,N_12780,N_13949);
xnor U16902 (N_16902,N_13901,N_13223);
xnor U16903 (N_16903,N_12505,N_14793);
and U16904 (N_16904,N_12710,N_13731);
nand U16905 (N_16905,N_13478,N_12699);
nand U16906 (N_16906,N_13155,N_14177);
nor U16907 (N_16907,N_14806,N_14152);
and U16908 (N_16908,N_12887,N_14526);
nor U16909 (N_16909,N_13027,N_14367);
xnor U16910 (N_16910,N_13627,N_14996);
xor U16911 (N_16911,N_14691,N_12790);
or U16912 (N_16912,N_13351,N_14780);
and U16913 (N_16913,N_13107,N_13891);
and U16914 (N_16914,N_12509,N_13812);
or U16915 (N_16915,N_13189,N_14690);
or U16916 (N_16916,N_14888,N_13501);
and U16917 (N_16917,N_14139,N_13577);
nor U16918 (N_16918,N_13421,N_13867);
nand U16919 (N_16919,N_13734,N_13655);
or U16920 (N_16920,N_14213,N_13758);
and U16921 (N_16921,N_13565,N_12702);
and U16922 (N_16922,N_14942,N_13031);
nor U16923 (N_16923,N_13099,N_12996);
nand U16924 (N_16924,N_12503,N_12729);
or U16925 (N_16925,N_13114,N_13157);
or U16926 (N_16926,N_13845,N_13846);
and U16927 (N_16927,N_14745,N_14225);
and U16928 (N_16928,N_14589,N_13621);
xnor U16929 (N_16929,N_14713,N_14917);
xor U16930 (N_16930,N_13651,N_13114);
nand U16931 (N_16931,N_13537,N_12565);
nand U16932 (N_16932,N_12784,N_14619);
xor U16933 (N_16933,N_12616,N_14510);
xnor U16934 (N_16934,N_13687,N_13187);
and U16935 (N_16935,N_14706,N_14323);
nand U16936 (N_16936,N_13221,N_14298);
xor U16937 (N_16937,N_14446,N_13166);
nor U16938 (N_16938,N_14229,N_12646);
xnor U16939 (N_16939,N_14782,N_13303);
or U16940 (N_16940,N_14568,N_13870);
nand U16941 (N_16941,N_14765,N_13429);
xor U16942 (N_16942,N_14307,N_14862);
nand U16943 (N_16943,N_12811,N_14531);
xnor U16944 (N_16944,N_14828,N_12840);
or U16945 (N_16945,N_13319,N_13598);
nand U16946 (N_16946,N_13023,N_12579);
or U16947 (N_16947,N_12560,N_13832);
xor U16948 (N_16948,N_12606,N_13213);
or U16949 (N_16949,N_14366,N_12958);
and U16950 (N_16950,N_13896,N_13943);
or U16951 (N_16951,N_14388,N_13848);
and U16952 (N_16952,N_13809,N_12603);
or U16953 (N_16953,N_13990,N_14679);
nor U16954 (N_16954,N_13040,N_14551);
and U16955 (N_16955,N_12593,N_14329);
and U16956 (N_16956,N_13172,N_12608);
nand U16957 (N_16957,N_13614,N_13397);
nor U16958 (N_16958,N_13047,N_14521);
xnor U16959 (N_16959,N_12760,N_13124);
and U16960 (N_16960,N_13942,N_13700);
and U16961 (N_16961,N_13531,N_14620);
nand U16962 (N_16962,N_13876,N_13145);
nand U16963 (N_16963,N_12921,N_12926);
xor U16964 (N_16964,N_13836,N_13695);
nor U16965 (N_16965,N_14204,N_14881);
nor U16966 (N_16966,N_13595,N_14970);
nor U16967 (N_16967,N_14917,N_13259);
xor U16968 (N_16968,N_12633,N_14474);
or U16969 (N_16969,N_13140,N_14981);
nor U16970 (N_16970,N_14039,N_14478);
or U16971 (N_16971,N_14326,N_13866);
or U16972 (N_16972,N_12755,N_14665);
or U16973 (N_16973,N_14685,N_13053);
and U16974 (N_16974,N_13849,N_14290);
xor U16975 (N_16975,N_13133,N_14390);
xnor U16976 (N_16976,N_14595,N_13657);
or U16977 (N_16977,N_14152,N_14217);
nor U16978 (N_16978,N_14725,N_14395);
nand U16979 (N_16979,N_12543,N_14813);
or U16980 (N_16980,N_14192,N_14024);
nand U16981 (N_16981,N_13288,N_14641);
nand U16982 (N_16982,N_13097,N_12695);
xor U16983 (N_16983,N_14934,N_13204);
nor U16984 (N_16984,N_12731,N_13661);
and U16985 (N_16985,N_14793,N_13102);
or U16986 (N_16986,N_14764,N_13473);
or U16987 (N_16987,N_13150,N_12574);
nand U16988 (N_16988,N_14333,N_13242);
nand U16989 (N_16989,N_13502,N_13961);
and U16990 (N_16990,N_13000,N_13941);
xnor U16991 (N_16991,N_14086,N_14061);
and U16992 (N_16992,N_12596,N_14926);
and U16993 (N_16993,N_12582,N_12805);
nor U16994 (N_16994,N_14711,N_14910);
or U16995 (N_16995,N_12574,N_13096);
xor U16996 (N_16996,N_14328,N_12767);
nor U16997 (N_16997,N_14037,N_14863);
nand U16998 (N_16998,N_12986,N_14728);
xor U16999 (N_16999,N_14075,N_13270);
and U17000 (N_17000,N_12814,N_12830);
nor U17001 (N_17001,N_14292,N_14087);
xor U17002 (N_17002,N_14372,N_13304);
or U17003 (N_17003,N_13988,N_13499);
or U17004 (N_17004,N_13847,N_13896);
and U17005 (N_17005,N_13312,N_14222);
nor U17006 (N_17006,N_14911,N_13308);
nand U17007 (N_17007,N_13526,N_14910);
nand U17008 (N_17008,N_13934,N_13516);
or U17009 (N_17009,N_13145,N_13821);
or U17010 (N_17010,N_13688,N_14100);
and U17011 (N_17011,N_12616,N_13809);
and U17012 (N_17012,N_13556,N_12652);
nand U17013 (N_17013,N_13867,N_13856);
nand U17014 (N_17014,N_14887,N_14245);
and U17015 (N_17015,N_14745,N_12901);
nor U17016 (N_17016,N_14489,N_14611);
nand U17017 (N_17017,N_14236,N_14250);
nand U17018 (N_17018,N_12838,N_14159);
and U17019 (N_17019,N_14146,N_14548);
xnor U17020 (N_17020,N_14853,N_13471);
xor U17021 (N_17021,N_14072,N_13457);
nand U17022 (N_17022,N_12969,N_13366);
and U17023 (N_17023,N_12837,N_13609);
nor U17024 (N_17024,N_13525,N_13959);
or U17025 (N_17025,N_13200,N_12856);
nor U17026 (N_17026,N_14915,N_14034);
and U17027 (N_17027,N_14959,N_12957);
or U17028 (N_17028,N_13283,N_12978);
or U17029 (N_17029,N_13818,N_14124);
and U17030 (N_17030,N_14883,N_14144);
or U17031 (N_17031,N_12897,N_13262);
xnor U17032 (N_17032,N_14364,N_13587);
or U17033 (N_17033,N_13246,N_13021);
nor U17034 (N_17034,N_14105,N_12747);
nand U17035 (N_17035,N_12856,N_14766);
or U17036 (N_17036,N_14228,N_13384);
xor U17037 (N_17037,N_13853,N_13683);
and U17038 (N_17038,N_14514,N_13632);
nor U17039 (N_17039,N_12744,N_13987);
or U17040 (N_17040,N_13442,N_13974);
and U17041 (N_17041,N_13747,N_13651);
xor U17042 (N_17042,N_13593,N_14818);
xor U17043 (N_17043,N_14370,N_14853);
and U17044 (N_17044,N_14938,N_12511);
and U17045 (N_17045,N_13881,N_14545);
nor U17046 (N_17046,N_13851,N_12700);
and U17047 (N_17047,N_14063,N_13286);
and U17048 (N_17048,N_14118,N_13453);
or U17049 (N_17049,N_14397,N_13301);
nor U17050 (N_17050,N_14595,N_13689);
or U17051 (N_17051,N_14938,N_14967);
or U17052 (N_17052,N_12629,N_13462);
nor U17053 (N_17053,N_14905,N_14393);
or U17054 (N_17054,N_14845,N_13749);
nand U17055 (N_17055,N_13049,N_13968);
or U17056 (N_17056,N_13883,N_13551);
and U17057 (N_17057,N_12880,N_14502);
nor U17058 (N_17058,N_13478,N_14789);
or U17059 (N_17059,N_12726,N_13980);
xnor U17060 (N_17060,N_13846,N_14689);
nand U17061 (N_17061,N_14219,N_13615);
nor U17062 (N_17062,N_13847,N_12609);
xnor U17063 (N_17063,N_12637,N_13619);
xor U17064 (N_17064,N_14274,N_14672);
or U17065 (N_17065,N_14756,N_13485);
or U17066 (N_17066,N_14439,N_12720);
and U17067 (N_17067,N_13238,N_13353);
nand U17068 (N_17068,N_14785,N_12726);
nor U17069 (N_17069,N_14515,N_12630);
xor U17070 (N_17070,N_12561,N_14207);
or U17071 (N_17071,N_14820,N_14436);
nand U17072 (N_17072,N_13730,N_13165);
and U17073 (N_17073,N_14336,N_14417);
or U17074 (N_17074,N_13056,N_14574);
and U17075 (N_17075,N_14296,N_14269);
nand U17076 (N_17076,N_12784,N_14666);
nor U17077 (N_17077,N_14194,N_13897);
xnor U17078 (N_17078,N_14143,N_12751);
xor U17079 (N_17079,N_12718,N_13970);
and U17080 (N_17080,N_13647,N_12603);
nand U17081 (N_17081,N_13310,N_13126);
nor U17082 (N_17082,N_14147,N_14740);
and U17083 (N_17083,N_13310,N_12748);
and U17084 (N_17084,N_12918,N_14213);
nand U17085 (N_17085,N_14737,N_14387);
or U17086 (N_17086,N_13174,N_14870);
and U17087 (N_17087,N_14256,N_13293);
nor U17088 (N_17088,N_14439,N_13379);
or U17089 (N_17089,N_14394,N_13007);
xnor U17090 (N_17090,N_14874,N_13606);
xor U17091 (N_17091,N_14231,N_13903);
and U17092 (N_17092,N_12721,N_12869);
xnor U17093 (N_17093,N_13848,N_14261);
xor U17094 (N_17094,N_14442,N_13571);
and U17095 (N_17095,N_14645,N_14549);
nor U17096 (N_17096,N_14280,N_13262);
and U17097 (N_17097,N_12966,N_13977);
xnor U17098 (N_17098,N_13980,N_14188);
and U17099 (N_17099,N_13070,N_13025);
nand U17100 (N_17100,N_14082,N_13227);
nand U17101 (N_17101,N_13659,N_14404);
or U17102 (N_17102,N_14033,N_14397);
xnor U17103 (N_17103,N_13613,N_13410);
xor U17104 (N_17104,N_13082,N_12749);
xnor U17105 (N_17105,N_13846,N_14840);
nand U17106 (N_17106,N_13421,N_12517);
nand U17107 (N_17107,N_14573,N_12700);
nor U17108 (N_17108,N_13476,N_14944);
nand U17109 (N_17109,N_13603,N_14009);
or U17110 (N_17110,N_14894,N_14109);
xor U17111 (N_17111,N_13417,N_13696);
nor U17112 (N_17112,N_14936,N_14347);
nand U17113 (N_17113,N_13581,N_13881);
nand U17114 (N_17114,N_13910,N_14626);
and U17115 (N_17115,N_13183,N_14740);
xor U17116 (N_17116,N_14710,N_13923);
xor U17117 (N_17117,N_14848,N_13786);
and U17118 (N_17118,N_13571,N_14127);
nor U17119 (N_17119,N_13307,N_14020);
nor U17120 (N_17120,N_13393,N_13626);
or U17121 (N_17121,N_14465,N_13133);
xor U17122 (N_17122,N_12727,N_14795);
xor U17123 (N_17123,N_13781,N_14917);
and U17124 (N_17124,N_14916,N_13581);
or U17125 (N_17125,N_12618,N_13559);
nand U17126 (N_17126,N_13762,N_12712);
or U17127 (N_17127,N_14117,N_14232);
nor U17128 (N_17128,N_13650,N_13947);
or U17129 (N_17129,N_13623,N_12556);
and U17130 (N_17130,N_13875,N_13336);
or U17131 (N_17131,N_14325,N_13549);
or U17132 (N_17132,N_13394,N_12989);
xnor U17133 (N_17133,N_13497,N_12973);
or U17134 (N_17134,N_13072,N_13156);
and U17135 (N_17135,N_12700,N_13635);
nand U17136 (N_17136,N_12946,N_12767);
or U17137 (N_17137,N_13330,N_14552);
nor U17138 (N_17138,N_12753,N_13506);
nor U17139 (N_17139,N_13887,N_14344);
nor U17140 (N_17140,N_13092,N_14915);
xor U17141 (N_17141,N_14143,N_14978);
or U17142 (N_17142,N_12653,N_13598);
or U17143 (N_17143,N_14208,N_12742);
and U17144 (N_17144,N_13052,N_14426);
nand U17145 (N_17145,N_12713,N_13539);
nand U17146 (N_17146,N_13916,N_13926);
nor U17147 (N_17147,N_13119,N_14589);
xor U17148 (N_17148,N_14620,N_14774);
xor U17149 (N_17149,N_13694,N_13502);
nor U17150 (N_17150,N_14204,N_12501);
and U17151 (N_17151,N_12519,N_13800);
nand U17152 (N_17152,N_14042,N_13642);
or U17153 (N_17153,N_14830,N_13487);
and U17154 (N_17154,N_13551,N_13993);
nor U17155 (N_17155,N_13306,N_13078);
nand U17156 (N_17156,N_14489,N_13981);
and U17157 (N_17157,N_14218,N_13533);
nand U17158 (N_17158,N_13838,N_13762);
xnor U17159 (N_17159,N_13298,N_14625);
and U17160 (N_17160,N_14767,N_14134);
nor U17161 (N_17161,N_13635,N_14988);
and U17162 (N_17162,N_12956,N_14924);
or U17163 (N_17163,N_13811,N_14074);
nor U17164 (N_17164,N_14653,N_14631);
nor U17165 (N_17165,N_13927,N_14470);
xor U17166 (N_17166,N_12648,N_13624);
or U17167 (N_17167,N_14454,N_13013);
nand U17168 (N_17168,N_14795,N_14178);
and U17169 (N_17169,N_14710,N_12730);
xor U17170 (N_17170,N_14938,N_13066);
and U17171 (N_17171,N_13017,N_12743);
xor U17172 (N_17172,N_14203,N_12851);
nand U17173 (N_17173,N_13312,N_12933);
or U17174 (N_17174,N_12561,N_14113);
and U17175 (N_17175,N_14671,N_12650);
nor U17176 (N_17176,N_13070,N_14940);
or U17177 (N_17177,N_12689,N_13994);
nand U17178 (N_17178,N_14537,N_12821);
nor U17179 (N_17179,N_13656,N_13189);
or U17180 (N_17180,N_13987,N_13103);
xor U17181 (N_17181,N_13133,N_13330);
xor U17182 (N_17182,N_13522,N_14575);
nor U17183 (N_17183,N_13994,N_13488);
or U17184 (N_17184,N_14341,N_14722);
xnor U17185 (N_17185,N_14683,N_14810);
nand U17186 (N_17186,N_14808,N_12659);
and U17187 (N_17187,N_13777,N_12559);
or U17188 (N_17188,N_13935,N_12591);
or U17189 (N_17189,N_14205,N_14708);
xnor U17190 (N_17190,N_13231,N_13090);
nor U17191 (N_17191,N_14150,N_13222);
and U17192 (N_17192,N_12714,N_12889);
nor U17193 (N_17193,N_13045,N_13826);
or U17194 (N_17194,N_12726,N_13570);
or U17195 (N_17195,N_13362,N_14240);
xor U17196 (N_17196,N_14396,N_14695);
and U17197 (N_17197,N_14192,N_13339);
xnor U17198 (N_17198,N_14751,N_13150);
nor U17199 (N_17199,N_14136,N_13333);
or U17200 (N_17200,N_13319,N_14774);
and U17201 (N_17201,N_13119,N_13429);
nor U17202 (N_17202,N_14130,N_12821);
nand U17203 (N_17203,N_13923,N_14999);
and U17204 (N_17204,N_14905,N_12738);
xor U17205 (N_17205,N_13127,N_12675);
and U17206 (N_17206,N_14485,N_13474);
and U17207 (N_17207,N_12947,N_12962);
xnor U17208 (N_17208,N_12560,N_13654);
nor U17209 (N_17209,N_14441,N_14842);
nor U17210 (N_17210,N_13062,N_13997);
nand U17211 (N_17211,N_13322,N_14694);
nand U17212 (N_17212,N_13599,N_13959);
nor U17213 (N_17213,N_13204,N_14403);
and U17214 (N_17214,N_14717,N_14834);
xor U17215 (N_17215,N_12853,N_14946);
or U17216 (N_17216,N_14523,N_13674);
and U17217 (N_17217,N_14615,N_12524);
nor U17218 (N_17218,N_13506,N_13391);
or U17219 (N_17219,N_14306,N_13539);
nand U17220 (N_17220,N_14044,N_14707);
xnor U17221 (N_17221,N_13673,N_13726);
or U17222 (N_17222,N_14119,N_14670);
or U17223 (N_17223,N_14011,N_14251);
and U17224 (N_17224,N_12505,N_13556);
xnor U17225 (N_17225,N_13020,N_14893);
or U17226 (N_17226,N_14788,N_13201);
and U17227 (N_17227,N_14977,N_14276);
and U17228 (N_17228,N_14679,N_13453);
or U17229 (N_17229,N_13934,N_14164);
xor U17230 (N_17230,N_13431,N_13401);
and U17231 (N_17231,N_14136,N_13079);
or U17232 (N_17232,N_14498,N_12558);
nor U17233 (N_17233,N_14787,N_12586);
nor U17234 (N_17234,N_14800,N_14734);
nor U17235 (N_17235,N_12512,N_14035);
xnor U17236 (N_17236,N_12608,N_13675);
nand U17237 (N_17237,N_13550,N_13705);
nand U17238 (N_17238,N_14266,N_14826);
and U17239 (N_17239,N_12736,N_14521);
nand U17240 (N_17240,N_14016,N_13344);
or U17241 (N_17241,N_14494,N_14637);
nand U17242 (N_17242,N_14644,N_14059);
or U17243 (N_17243,N_14884,N_14577);
or U17244 (N_17244,N_13119,N_14318);
xor U17245 (N_17245,N_13015,N_14086);
or U17246 (N_17246,N_13284,N_13576);
xnor U17247 (N_17247,N_12889,N_13525);
nand U17248 (N_17248,N_14798,N_14416);
and U17249 (N_17249,N_13352,N_13495);
xnor U17250 (N_17250,N_13943,N_12926);
nor U17251 (N_17251,N_13089,N_13956);
and U17252 (N_17252,N_13488,N_13634);
nor U17253 (N_17253,N_13901,N_14730);
nand U17254 (N_17254,N_14023,N_13177);
xor U17255 (N_17255,N_13561,N_12616);
or U17256 (N_17256,N_13841,N_14075);
nand U17257 (N_17257,N_13911,N_12593);
nor U17258 (N_17258,N_13967,N_14976);
nor U17259 (N_17259,N_12921,N_13619);
nor U17260 (N_17260,N_12681,N_13120);
nor U17261 (N_17261,N_14878,N_14799);
xor U17262 (N_17262,N_12910,N_14911);
or U17263 (N_17263,N_14258,N_13145);
and U17264 (N_17264,N_12890,N_13427);
and U17265 (N_17265,N_14310,N_14904);
xnor U17266 (N_17266,N_12702,N_12879);
nand U17267 (N_17267,N_13914,N_12909);
nor U17268 (N_17268,N_13411,N_14916);
or U17269 (N_17269,N_13571,N_14265);
or U17270 (N_17270,N_13180,N_14455);
xnor U17271 (N_17271,N_14089,N_13735);
or U17272 (N_17272,N_14203,N_12972);
or U17273 (N_17273,N_13260,N_12859);
nor U17274 (N_17274,N_13817,N_14677);
and U17275 (N_17275,N_12888,N_12533);
and U17276 (N_17276,N_12798,N_13307);
nand U17277 (N_17277,N_14688,N_12719);
nor U17278 (N_17278,N_13224,N_14512);
nand U17279 (N_17279,N_12803,N_14857);
nand U17280 (N_17280,N_13542,N_13308);
xnor U17281 (N_17281,N_14835,N_12813);
nand U17282 (N_17282,N_14304,N_14277);
or U17283 (N_17283,N_12933,N_14513);
nor U17284 (N_17284,N_13553,N_13442);
or U17285 (N_17285,N_13844,N_13742);
xor U17286 (N_17286,N_13811,N_14554);
or U17287 (N_17287,N_12847,N_12905);
nor U17288 (N_17288,N_13641,N_14357);
nor U17289 (N_17289,N_14032,N_14066);
nor U17290 (N_17290,N_13517,N_14913);
xor U17291 (N_17291,N_14762,N_13387);
nand U17292 (N_17292,N_13561,N_14413);
or U17293 (N_17293,N_14931,N_13303);
nor U17294 (N_17294,N_13791,N_14279);
xor U17295 (N_17295,N_13261,N_14693);
nor U17296 (N_17296,N_12885,N_14807);
nor U17297 (N_17297,N_13211,N_13317);
and U17298 (N_17298,N_14756,N_14432);
and U17299 (N_17299,N_14842,N_14955);
or U17300 (N_17300,N_14850,N_14071);
or U17301 (N_17301,N_14491,N_14529);
nand U17302 (N_17302,N_14149,N_12802);
and U17303 (N_17303,N_14515,N_13953);
and U17304 (N_17304,N_13452,N_13178);
nand U17305 (N_17305,N_14397,N_13660);
and U17306 (N_17306,N_13104,N_13760);
and U17307 (N_17307,N_14620,N_13843);
xnor U17308 (N_17308,N_13184,N_14371);
nor U17309 (N_17309,N_14358,N_14816);
or U17310 (N_17310,N_14218,N_14396);
nor U17311 (N_17311,N_13831,N_14728);
or U17312 (N_17312,N_13517,N_13061);
nand U17313 (N_17313,N_14503,N_14895);
xor U17314 (N_17314,N_13214,N_12763);
nor U17315 (N_17315,N_13871,N_14617);
nor U17316 (N_17316,N_14626,N_14722);
nor U17317 (N_17317,N_14314,N_13243);
nand U17318 (N_17318,N_13102,N_12525);
and U17319 (N_17319,N_12568,N_13244);
nor U17320 (N_17320,N_12990,N_13695);
xor U17321 (N_17321,N_14950,N_13516);
or U17322 (N_17322,N_14900,N_14354);
and U17323 (N_17323,N_13371,N_13621);
nand U17324 (N_17324,N_14874,N_14878);
or U17325 (N_17325,N_13919,N_13160);
and U17326 (N_17326,N_13134,N_13649);
and U17327 (N_17327,N_14913,N_12595);
nor U17328 (N_17328,N_13745,N_14823);
and U17329 (N_17329,N_12682,N_13954);
nand U17330 (N_17330,N_13800,N_13398);
xor U17331 (N_17331,N_14960,N_13074);
nand U17332 (N_17332,N_12587,N_14001);
and U17333 (N_17333,N_13972,N_13175);
or U17334 (N_17334,N_13609,N_14235);
nand U17335 (N_17335,N_13673,N_13499);
or U17336 (N_17336,N_14458,N_14606);
nor U17337 (N_17337,N_12762,N_12549);
nor U17338 (N_17338,N_13437,N_12943);
or U17339 (N_17339,N_14933,N_12939);
nand U17340 (N_17340,N_13444,N_12702);
nand U17341 (N_17341,N_14294,N_13451);
nand U17342 (N_17342,N_13363,N_12874);
nor U17343 (N_17343,N_14858,N_14521);
xor U17344 (N_17344,N_13724,N_13888);
nor U17345 (N_17345,N_12599,N_12750);
nand U17346 (N_17346,N_12678,N_14843);
nor U17347 (N_17347,N_13302,N_13041);
nand U17348 (N_17348,N_14725,N_13157);
nand U17349 (N_17349,N_13389,N_13878);
and U17350 (N_17350,N_13144,N_13244);
nor U17351 (N_17351,N_13886,N_14999);
or U17352 (N_17352,N_12844,N_13226);
nand U17353 (N_17353,N_14429,N_14570);
nand U17354 (N_17354,N_14513,N_14766);
and U17355 (N_17355,N_14549,N_12542);
or U17356 (N_17356,N_13955,N_13454);
or U17357 (N_17357,N_14800,N_14211);
nand U17358 (N_17358,N_13672,N_13926);
nor U17359 (N_17359,N_14651,N_13670);
nor U17360 (N_17360,N_14763,N_14003);
and U17361 (N_17361,N_14399,N_13400);
nor U17362 (N_17362,N_14394,N_14301);
nand U17363 (N_17363,N_12736,N_14517);
or U17364 (N_17364,N_13442,N_13111);
or U17365 (N_17365,N_13372,N_14623);
and U17366 (N_17366,N_13919,N_13242);
nand U17367 (N_17367,N_14316,N_14280);
or U17368 (N_17368,N_12853,N_12567);
or U17369 (N_17369,N_13578,N_14416);
and U17370 (N_17370,N_13174,N_14775);
nor U17371 (N_17371,N_12978,N_13988);
xor U17372 (N_17372,N_14513,N_13261);
or U17373 (N_17373,N_14932,N_14723);
nand U17374 (N_17374,N_13231,N_12929);
nor U17375 (N_17375,N_12812,N_13878);
nor U17376 (N_17376,N_12658,N_12819);
nor U17377 (N_17377,N_13233,N_14969);
xor U17378 (N_17378,N_14958,N_13895);
or U17379 (N_17379,N_14806,N_12649);
xor U17380 (N_17380,N_14198,N_14605);
xnor U17381 (N_17381,N_14081,N_13849);
xnor U17382 (N_17382,N_13620,N_12526);
xnor U17383 (N_17383,N_13621,N_14397);
xor U17384 (N_17384,N_13558,N_13221);
or U17385 (N_17385,N_13769,N_14381);
xnor U17386 (N_17386,N_12905,N_14975);
nand U17387 (N_17387,N_13426,N_14003);
or U17388 (N_17388,N_14611,N_13884);
or U17389 (N_17389,N_14967,N_14046);
xor U17390 (N_17390,N_14539,N_13009);
and U17391 (N_17391,N_12724,N_13397);
nor U17392 (N_17392,N_14342,N_13928);
or U17393 (N_17393,N_13721,N_12568);
or U17394 (N_17394,N_14613,N_13175);
nand U17395 (N_17395,N_12711,N_12631);
xor U17396 (N_17396,N_13613,N_12728);
or U17397 (N_17397,N_13607,N_12603);
and U17398 (N_17398,N_14634,N_14071);
xor U17399 (N_17399,N_14378,N_12628);
and U17400 (N_17400,N_13783,N_14048);
and U17401 (N_17401,N_13665,N_12798);
nand U17402 (N_17402,N_14419,N_13747);
xnor U17403 (N_17403,N_14345,N_14256);
or U17404 (N_17404,N_14197,N_14113);
or U17405 (N_17405,N_14319,N_13502);
and U17406 (N_17406,N_14970,N_12785);
nor U17407 (N_17407,N_13800,N_14550);
xor U17408 (N_17408,N_14319,N_14364);
nand U17409 (N_17409,N_14933,N_14592);
nor U17410 (N_17410,N_14816,N_12532);
nor U17411 (N_17411,N_14709,N_12564);
xor U17412 (N_17412,N_14994,N_14286);
nor U17413 (N_17413,N_12827,N_13231);
nand U17414 (N_17414,N_13232,N_14833);
xor U17415 (N_17415,N_14058,N_13748);
xnor U17416 (N_17416,N_12793,N_14780);
nor U17417 (N_17417,N_13802,N_12981);
or U17418 (N_17418,N_13759,N_13600);
or U17419 (N_17419,N_13344,N_12860);
or U17420 (N_17420,N_14002,N_13507);
nor U17421 (N_17421,N_13019,N_12815);
xor U17422 (N_17422,N_13951,N_12900);
or U17423 (N_17423,N_13484,N_13870);
xor U17424 (N_17424,N_13533,N_12650);
nand U17425 (N_17425,N_13474,N_14333);
nor U17426 (N_17426,N_13973,N_13818);
xor U17427 (N_17427,N_13442,N_13751);
and U17428 (N_17428,N_12832,N_12885);
nand U17429 (N_17429,N_13671,N_14876);
xor U17430 (N_17430,N_13393,N_13852);
nor U17431 (N_17431,N_13901,N_14214);
xor U17432 (N_17432,N_13347,N_14759);
xnor U17433 (N_17433,N_14717,N_13010);
and U17434 (N_17434,N_14723,N_14003);
and U17435 (N_17435,N_14777,N_14042);
or U17436 (N_17436,N_14589,N_14488);
nor U17437 (N_17437,N_12767,N_13168);
or U17438 (N_17438,N_14531,N_13232);
nand U17439 (N_17439,N_13507,N_13404);
and U17440 (N_17440,N_12892,N_14562);
nor U17441 (N_17441,N_13344,N_14107);
nand U17442 (N_17442,N_12791,N_13927);
nand U17443 (N_17443,N_14937,N_13400);
or U17444 (N_17444,N_13593,N_14638);
nor U17445 (N_17445,N_13228,N_13309);
nor U17446 (N_17446,N_14843,N_13666);
or U17447 (N_17447,N_14082,N_14667);
xnor U17448 (N_17448,N_13049,N_14992);
and U17449 (N_17449,N_14149,N_12990);
or U17450 (N_17450,N_14541,N_13605);
xor U17451 (N_17451,N_14720,N_14138);
nand U17452 (N_17452,N_14370,N_12937);
or U17453 (N_17453,N_14773,N_14843);
nor U17454 (N_17454,N_14593,N_14565);
and U17455 (N_17455,N_14992,N_13934);
nand U17456 (N_17456,N_14649,N_13560);
xor U17457 (N_17457,N_14851,N_13093);
xor U17458 (N_17458,N_12590,N_12641);
and U17459 (N_17459,N_14970,N_13969);
nor U17460 (N_17460,N_12778,N_13407);
nor U17461 (N_17461,N_14231,N_13669);
nand U17462 (N_17462,N_13811,N_13158);
nand U17463 (N_17463,N_13495,N_14266);
or U17464 (N_17464,N_13265,N_13540);
or U17465 (N_17465,N_14770,N_12982);
nor U17466 (N_17466,N_14644,N_14027);
or U17467 (N_17467,N_13157,N_12631);
nand U17468 (N_17468,N_13157,N_12768);
and U17469 (N_17469,N_14055,N_13539);
nor U17470 (N_17470,N_13561,N_14460);
nor U17471 (N_17471,N_14854,N_13569);
nor U17472 (N_17472,N_13354,N_13423);
and U17473 (N_17473,N_12936,N_12776);
xnor U17474 (N_17474,N_14798,N_12888);
nand U17475 (N_17475,N_13595,N_12842);
nand U17476 (N_17476,N_12652,N_13470);
or U17477 (N_17477,N_12650,N_14728);
nand U17478 (N_17478,N_14280,N_12544);
or U17479 (N_17479,N_13508,N_12759);
xnor U17480 (N_17480,N_13818,N_12553);
or U17481 (N_17481,N_13756,N_14995);
xnor U17482 (N_17482,N_12954,N_14047);
nand U17483 (N_17483,N_13617,N_12897);
or U17484 (N_17484,N_13389,N_14335);
xnor U17485 (N_17485,N_14818,N_12843);
or U17486 (N_17486,N_13287,N_13705);
or U17487 (N_17487,N_13251,N_14960);
nand U17488 (N_17488,N_13467,N_14416);
nor U17489 (N_17489,N_14826,N_13662);
nand U17490 (N_17490,N_13155,N_12815);
and U17491 (N_17491,N_14703,N_13725);
or U17492 (N_17492,N_13136,N_13316);
nand U17493 (N_17493,N_13765,N_14542);
nor U17494 (N_17494,N_13934,N_14017);
nand U17495 (N_17495,N_12962,N_13381);
xnor U17496 (N_17496,N_13909,N_13314);
and U17497 (N_17497,N_12665,N_14108);
xnor U17498 (N_17498,N_13922,N_12775);
nand U17499 (N_17499,N_13711,N_14550);
and U17500 (N_17500,N_16699,N_16892);
or U17501 (N_17501,N_17457,N_17261);
and U17502 (N_17502,N_15509,N_17110);
or U17503 (N_17503,N_15828,N_15212);
nand U17504 (N_17504,N_15081,N_16840);
nand U17505 (N_17505,N_16603,N_16314);
or U17506 (N_17506,N_17438,N_15405);
or U17507 (N_17507,N_15132,N_17371);
xor U17508 (N_17508,N_15201,N_15978);
nor U17509 (N_17509,N_16083,N_16062);
and U17510 (N_17510,N_15693,N_15925);
or U17511 (N_17511,N_17471,N_15959);
nand U17512 (N_17512,N_16782,N_16248);
nand U17513 (N_17513,N_16673,N_15465);
or U17514 (N_17514,N_16135,N_15391);
nor U17515 (N_17515,N_16470,N_16285);
nor U17516 (N_17516,N_15311,N_16258);
and U17517 (N_17517,N_16515,N_16312);
xor U17518 (N_17518,N_16316,N_16236);
xor U17519 (N_17519,N_16755,N_17269);
or U17520 (N_17520,N_17421,N_16296);
or U17521 (N_17521,N_17419,N_16191);
xnor U17522 (N_17522,N_16768,N_16455);
xor U17523 (N_17523,N_15038,N_17299);
and U17524 (N_17524,N_15142,N_15744);
or U17525 (N_17525,N_15616,N_16299);
nor U17526 (N_17526,N_16981,N_15543);
xnor U17527 (N_17527,N_16852,N_16099);
xor U17528 (N_17528,N_15286,N_15253);
nand U17529 (N_17529,N_15900,N_17120);
or U17530 (N_17530,N_15618,N_17322);
nand U17531 (N_17531,N_16338,N_17332);
nor U17532 (N_17532,N_15528,N_15290);
xor U17533 (N_17533,N_15600,N_15851);
nand U17534 (N_17534,N_15944,N_16706);
and U17535 (N_17535,N_16129,N_15617);
xnor U17536 (N_17536,N_15283,N_15531);
nand U17537 (N_17537,N_15302,N_15957);
or U17538 (N_17538,N_16354,N_15464);
and U17539 (N_17539,N_16807,N_17343);
and U17540 (N_17540,N_16491,N_16272);
nor U17541 (N_17541,N_16082,N_17455);
nor U17542 (N_17542,N_16397,N_17445);
and U17543 (N_17543,N_15368,N_16737);
and U17544 (N_17544,N_15926,N_17070);
xnor U17545 (N_17545,N_15322,N_15039);
and U17546 (N_17546,N_16210,N_17287);
and U17547 (N_17547,N_15447,N_16731);
or U17548 (N_17548,N_16380,N_16475);
nor U17549 (N_17549,N_15104,N_15389);
and U17550 (N_17550,N_15517,N_17373);
or U17551 (N_17551,N_17138,N_15146);
nand U17552 (N_17552,N_16345,N_17391);
xor U17553 (N_17553,N_15143,N_15161);
or U17554 (N_17554,N_15868,N_15939);
nor U17555 (N_17555,N_15857,N_17192);
or U17556 (N_17556,N_15656,N_15558);
or U17557 (N_17557,N_16851,N_16105);
and U17558 (N_17558,N_17405,N_16683);
and U17559 (N_17559,N_17169,N_16412);
or U17560 (N_17560,N_17459,N_16434);
or U17561 (N_17561,N_16436,N_17270);
and U17562 (N_17562,N_17293,N_17402);
nor U17563 (N_17563,N_16487,N_16536);
or U17564 (N_17564,N_16367,N_17243);
xnor U17565 (N_17565,N_15280,N_17485);
nor U17566 (N_17566,N_16457,N_17426);
nand U17567 (N_17567,N_16224,N_15689);
xor U17568 (N_17568,N_15083,N_17202);
xnor U17569 (N_17569,N_15396,N_16254);
or U17570 (N_17570,N_15029,N_17338);
nor U17571 (N_17571,N_15999,N_15576);
or U17572 (N_17572,N_17190,N_17075);
xnor U17573 (N_17573,N_16313,N_16670);
nand U17574 (N_17574,N_16907,N_15605);
nand U17575 (N_17575,N_16844,N_15331);
and U17576 (N_17576,N_17022,N_16485);
or U17577 (N_17577,N_16421,N_17420);
nand U17578 (N_17578,N_15166,N_15830);
xor U17579 (N_17579,N_15947,N_16070);
and U17580 (N_17580,N_16494,N_15373);
nand U17581 (N_17581,N_15610,N_16030);
nand U17582 (N_17582,N_16938,N_15333);
and U17583 (N_17583,N_16647,N_17408);
nand U17584 (N_17584,N_17285,N_16574);
nand U17585 (N_17585,N_15510,N_15971);
and U17586 (N_17586,N_16905,N_16912);
xor U17587 (N_17587,N_16045,N_15293);
nand U17588 (N_17588,N_16588,N_17250);
nor U17589 (N_17589,N_16608,N_15766);
nand U17590 (N_17590,N_16169,N_16654);
or U17591 (N_17591,N_15043,N_15014);
nand U17592 (N_17592,N_15227,N_16866);
nor U17593 (N_17593,N_15025,N_16593);
or U17594 (N_17594,N_15582,N_16902);
nand U17595 (N_17595,N_16249,N_15845);
nor U17596 (N_17596,N_17074,N_15028);
nand U17597 (N_17597,N_16900,N_15108);
or U17598 (N_17598,N_17222,N_16996);
xnor U17599 (N_17599,N_17308,N_15898);
nand U17600 (N_17600,N_16268,N_15714);
and U17601 (N_17601,N_16960,N_15958);
nor U17602 (N_17602,N_16220,N_16143);
or U17603 (N_17603,N_15544,N_15238);
xnor U17604 (N_17604,N_17301,N_17443);
nor U17605 (N_17605,N_16097,N_15094);
and U17606 (N_17606,N_17311,N_15599);
xnor U17607 (N_17607,N_16971,N_15606);
nand U17608 (N_17608,N_17153,N_15437);
xnor U17609 (N_17609,N_15979,N_17076);
nand U17610 (N_17610,N_15813,N_16655);
or U17611 (N_17611,N_15296,N_17246);
nor U17612 (N_17612,N_16047,N_16766);
or U17613 (N_17613,N_17067,N_16857);
xnor U17614 (N_17614,N_15839,N_15810);
nand U17615 (N_17615,N_15187,N_17025);
or U17616 (N_17616,N_16595,N_15015);
or U17617 (N_17617,N_15512,N_15165);
nand U17618 (N_17618,N_15407,N_15946);
or U17619 (N_17619,N_17378,N_16921);
or U17620 (N_17620,N_15241,N_16335);
nor U17621 (N_17621,N_17206,N_15365);
and U17622 (N_17622,N_15778,N_15346);
or U17623 (N_17623,N_17215,N_16711);
nor U17624 (N_17624,N_16009,N_16898);
nand U17625 (N_17625,N_17048,N_17043);
or U17626 (N_17626,N_16445,N_15414);
nor U17627 (N_17627,N_17477,N_15923);
xnor U17628 (N_17628,N_17052,N_15360);
and U17629 (N_17629,N_17262,N_16454);
xnor U17630 (N_17630,N_15002,N_16435);
and U17631 (N_17631,N_16687,N_15119);
nand U17632 (N_17632,N_16743,N_17105);
or U17633 (N_17633,N_15593,N_16562);
xor U17634 (N_17634,N_16552,N_15927);
or U17635 (N_17635,N_15800,N_17440);
nand U17636 (N_17636,N_15224,N_16941);
and U17637 (N_17637,N_15031,N_15085);
or U17638 (N_17638,N_16462,N_17026);
or U17639 (N_17639,N_15769,N_15795);
nor U17640 (N_17640,N_17348,N_17144);
or U17641 (N_17641,N_15673,N_15730);
and U17642 (N_17642,N_15246,N_16138);
or U17643 (N_17643,N_17160,N_15106);
nand U17644 (N_17644,N_16280,N_15870);
or U17645 (N_17645,N_17042,N_16399);
nand U17646 (N_17646,N_17382,N_16858);
and U17647 (N_17647,N_15886,N_15847);
and U17648 (N_17648,N_17251,N_15190);
nand U17649 (N_17649,N_16478,N_16497);
and U17650 (N_17650,N_17424,N_16948);
nand U17651 (N_17651,N_15913,N_15220);
and U17652 (N_17652,N_16928,N_17054);
nor U17653 (N_17653,N_16327,N_15676);
nor U17654 (N_17654,N_17413,N_16292);
nand U17655 (N_17655,N_16295,N_15826);
nand U17656 (N_17656,N_17499,N_15881);
and U17657 (N_17657,N_15261,N_17028);
nand U17658 (N_17658,N_17156,N_15217);
nor U17659 (N_17659,N_17004,N_17142);
xor U17660 (N_17660,N_15788,N_15804);
xnor U17661 (N_17661,N_15079,N_16833);
or U17662 (N_17662,N_16617,N_15638);
nand U17663 (N_17663,N_17289,N_15747);
or U17664 (N_17664,N_15872,N_17410);
or U17665 (N_17665,N_15499,N_15228);
nand U17666 (N_17666,N_16108,N_15336);
and U17667 (N_17667,N_17235,N_16976);
and U17668 (N_17668,N_15622,N_15579);
and U17669 (N_17669,N_16714,N_16621);
and U17670 (N_17670,N_15249,N_17211);
or U17671 (N_17671,N_15055,N_15716);
xor U17672 (N_17672,N_17217,N_17008);
or U17673 (N_17673,N_15095,N_17312);
nor U17674 (N_17674,N_17490,N_17115);
nor U17675 (N_17675,N_15682,N_15129);
and U17676 (N_17676,N_15601,N_16170);
nor U17677 (N_17677,N_16011,N_16742);
or U17678 (N_17678,N_17053,N_16809);
nand U17679 (N_17679,N_16036,N_16919);
and U17680 (N_17680,N_15948,N_15646);
xnor U17681 (N_17681,N_15974,N_16350);
and U17682 (N_17682,N_17155,N_16127);
and U17683 (N_17683,N_17309,N_17104);
nand U17684 (N_17684,N_17205,N_15885);
or U17685 (N_17685,N_16270,N_17330);
or U17686 (N_17686,N_17363,N_16816);
xor U17687 (N_17687,N_17290,N_16599);
or U17688 (N_17688,N_16791,N_16391);
nand U17689 (N_17689,N_15774,N_17288);
nor U17690 (N_17690,N_16159,N_15073);
nand U17691 (N_17691,N_16999,N_17082);
and U17692 (N_17692,N_15571,N_16756);
xnor U17693 (N_17693,N_17129,N_17321);
and U17694 (N_17694,N_16310,N_16931);
nor U17695 (N_17695,N_15023,N_15047);
nand U17696 (N_17696,N_17461,N_15764);
and U17697 (N_17697,N_17116,N_16966);
or U17698 (N_17698,N_17009,N_15863);
and U17699 (N_17699,N_15861,N_17300);
and U17700 (N_17700,N_16799,N_16728);
nand U17701 (N_17701,N_15449,N_16010);
and U17702 (N_17702,N_16954,N_15723);
or U17703 (N_17703,N_16982,N_16665);
nor U17704 (N_17704,N_16309,N_16474);
nand U17705 (N_17705,N_16212,N_17035);
and U17706 (N_17706,N_15790,N_15294);
xor U17707 (N_17707,N_15300,N_16074);
and U17708 (N_17708,N_15197,N_17324);
or U17709 (N_17709,N_16183,N_15848);
nand U17710 (N_17710,N_15631,N_17049);
nand U17711 (N_17711,N_16707,N_15889);
xnor U17712 (N_17712,N_15147,N_16842);
or U17713 (N_17713,N_15595,N_15451);
nand U17714 (N_17714,N_16078,N_15829);
and U17715 (N_17715,N_16464,N_16409);
nor U17716 (N_17716,N_16775,N_15385);
xnor U17717 (N_17717,N_16698,N_17236);
nor U17718 (N_17718,N_17170,N_16572);
xor U17719 (N_17719,N_16160,N_15068);
xnor U17720 (N_17720,N_15727,N_15623);
nor U17721 (N_17721,N_16987,N_16479);
or U17722 (N_17722,N_17333,N_16218);
and U17723 (N_17723,N_16227,N_16172);
and U17724 (N_17724,N_15503,N_15022);
nand U17725 (N_17725,N_17468,N_16887);
and U17726 (N_17726,N_15572,N_16100);
and U17727 (N_17727,N_15907,N_15340);
nand U17728 (N_17728,N_15757,N_16984);
or U17729 (N_17729,N_16261,N_16754);
xor U17730 (N_17730,N_15113,N_15334);
nand U17731 (N_17731,N_17232,N_16146);
nor U17732 (N_17732,N_16771,N_16586);
or U17733 (N_17733,N_16583,N_16029);
xnor U17734 (N_17734,N_15021,N_16815);
xnor U17735 (N_17735,N_17086,N_15981);
nand U17736 (N_17736,N_15789,N_17123);
and U17737 (N_17737,N_15101,N_15678);
nand U17738 (N_17738,N_16517,N_16717);
nand U17739 (N_17739,N_16974,N_17329);
nor U17740 (N_17740,N_17249,N_17273);
nor U17741 (N_17741,N_15854,N_15289);
nor U17742 (N_17742,N_16795,N_15621);
nor U17743 (N_17743,N_16582,N_15592);
xor U17744 (N_17744,N_17024,N_16034);
or U17745 (N_17745,N_15928,N_15668);
nor U17746 (N_17746,N_15372,N_16181);
or U17747 (N_17747,N_15102,N_17464);
and U17748 (N_17748,N_15608,N_15399);
nor U17749 (N_17749,N_15674,N_17397);
or U17750 (N_17750,N_15341,N_15090);
and U17751 (N_17751,N_17336,N_16814);
and U17752 (N_17752,N_15235,N_16035);
nor U17753 (N_17753,N_16895,N_15887);
xnor U17754 (N_17754,N_16349,N_15538);
nand U17755 (N_17755,N_16323,N_16880);
or U17756 (N_17756,N_16416,N_16672);
nand U17757 (N_17757,N_15743,N_16050);
nand U17758 (N_17758,N_16525,N_17213);
or U17759 (N_17759,N_15214,N_16472);
nor U17760 (N_17760,N_15052,N_16612);
xnor U17761 (N_17761,N_15805,N_15403);
or U17762 (N_17762,N_16969,N_15075);
nor U17763 (N_17763,N_17061,N_17425);
xor U17764 (N_17764,N_16013,N_16547);
and U17765 (N_17765,N_17446,N_15415);
nor U17766 (N_17766,N_15033,N_16914);
nor U17767 (N_17767,N_16242,N_15359);
or U17768 (N_17768,N_16513,N_16827);
nand U17769 (N_17769,N_16774,N_16635);
and U17770 (N_17770,N_15797,N_16111);
and U17771 (N_17771,N_16631,N_16308);
or U17772 (N_17772,N_17429,N_16511);
nand U17773 (N_17773,N_15835,N_16489);
xor U17774 (N_17774,N_15194,N_16561);
nand U17775 (N_17775,N_16760,N_16422);
xnor U17776 (N_17776,N_15091,N_15097);
xor U17777 (N_17777,N_15547,N_16745);
or U17778 (N_17778,N_15375,N_17168);
nand U17779 (N_17779,N_17254,N_17282);
or U17780 (N_17780,N_16625,N_16972);
or U17781 (N_17781,N_15087,N_16629);
nor U17782 (N_17782,N_16957,N_15174);
or U17783 (N_17783,N_16266,N_16610);
nor U17784 (N_17784,N_15355,N_16509);
xor U17785 (N_17785,N_17242,N_16970);
nand U17786 (N_17786,N_15591,N_15353);
nand U17787 (N_17787,N_15222,N_17248);
or U17788 (N_17788,N_15771,N_16725);
and U17789 (N_17789,N_16550,N_15849);
or U17790 (N_17790,N_16546,N_15866);
and U17791 (N_17791,N_15140,N_16413);
xor U17792 (N_17792,N_17291,N_17342);
nand U17793 (N_17793,N_15715,N_15581);
and U17794 (N_17794,N_15658,N_16044);
or U17795 (N_17795,N_15257,N_15546);
or U17796 (N_17796,N_17186,N_17196);
nor U17797 (N_17797,N_15251,N_16897);
and U17798 (N_17798,N_17195,N_16376);
nand U17799 (N_17799,N_17452,N_17031);
xor U17800 (N_17800,N_17307,N_16607);
or U17801 (N_17801,N_17122,N_16787);
nand U17802 (N_17802,N_16040,N_17209);
and U17803 (N_17803,N_15019,N_16428);
xor U17804 (N_17804,N_16694,N_15476);
and U17805 (N_17805,N_16952,N_17069);
xor U17806 (N_17806,N_15423,N_16293);
nand U17807 (N_17807,N_16441,N_16400);
xnor U17808 (N_17808,N_15876,N_15793);
and U17809 (N_17809,N_16046,N_17210);
nor U17810 (N_17810,N_15781,N_16688);
nor U17811 (N_17811,N_15660,N_16051);
or U17812 (N_17812,N_15207,N_16689);
nand U17813 (N_17813,N_15298,N_16466);
nor U17814 (N_17814,N_15018,N_15619);
nand U17815 (N_17815,N_15148,N_15768);
nand U17816 (N_17816,N_16681,N_16734);
and U17817 (N_17817,N_15305,N_15344);
and U17818 (N_17818,N_17238,N_15908);
xor U17819 (N_17819,N_16753,N_16845);
xor U17820 (N_17820,N_17315,N_16788);
and U17821 (N_17821,N_17346,N_15583);
nand U17822 (N_17822,N_16748,N_16379);
or U17823 (N_17823,N_16680,N_17487);
or U17824 (N_17824,N_16802,N_16913);
and U17825 (N_17825,N_17239,N_16442);
and U17826 (N_17826,N_16879,N_16205);
and U17827 (N_17827,N_15310,N_16204);
or U17828 (N_17828,N_15628,N_15103);
or U17829 (N_17829,N_15342,N_16317);
xor U17830 (N_17830,N_16347,N_16708);
nand U17831 (N_17831,N_16219,N_16622);
xnor U17832 (N_17832,N_15798,N_16716);
nand U17833 (N_17833,N_16085,N_15016);
nor U17834 (N_17834,N_16839,N_17476);
nand U17835 (N_17835,N_16095,N_15244);
or U17836 (N_17836,N_17040,N_16739);
xor U17837 (N_17837,N_16076,N_15896);
or U17838 (N_17838,N_15669,N_15136);
and U17839 (N_17839,N_16141,N_16520);
nand U17840 (N_17840,N_16544,N_16449);
or U17841 (N_17841,N_15844,N_15785);
and U17842 (N_17842,N_16602,N_15185);
xnor U17843 (N_17843,N_15463,N_15240);
xnor U17844 (N_17844,N_16087,N_15349);
and U17845 (N_17845,N_15961,N_15522);
xnor U17846 (N_17846,N_17214,N_15534);
or U17847 (N_17847,N_16894,N_15485);
or U17848 (N_17848,N_16630,N_17014);
nand U17849 (N_17849,N_15472,N_17275);
or U17850 (N_17850,N_16573,N_17032);
nand U17851 (N_17851,N_15209,N_16824);
nor U17852 (N_17852,N_16637,N_15114);
xor U17853 (N_17853,N_17462,N_17354);
xnor U17854 (N_17854,N_17392,N_17398);
and U17855 (N_17855,N_15416,N_15221);
nand U17856 (N_17856,N_15722,N_16943);
xor U17857 (N_17857,N_16072,N_15681);
nand U17858 (N_17858,N_16558,N_15580);
or U17859 (N_17859,N_17005,N_15394);
xor U17860 (N_17860,N_16514,N_17302);
or U17861 (N_17861,N_15408,N_16658);
nor U17862 (N_17862,N_15168,N_16500);
xnor U17863 (N_17863,N_16329,N_15951);
nor U17864 (N_17864,N_15304,N_15281);
and U17865 (N_17865,N_15664,N_16168);
nor U17866 (N_17866,N_15919,N_16330);
nand U17867 (N_17867,N_16002,N_15930);
nor U17868 (N_17868,N_17197,N_16611);
nand U17869 (N_17869,N_17172,N_17379);
and U17870 (N_17870,N_16342,N_16729);
xor U17871 (N_17871,N_15526,N_16163);
nor U17872 (N_17872,N_16066,N_15452);
and U17873 (N_17873,N_15883,N_16618);
or U17874 (N_17874,N_17084,N_15356);
and U17875 (N_17875,N_15180,N_15731);
nor U17876 (N_17876,N_15125,N_16382);
nand U17877 (N_17877,N_16811,N_16736);
nand U17878 (N_17878,N_17316,N_16420);
nor U17879 (N_17879,N_16164,N_16398);
nand U17880 (N_17880,N_17470,N_15299);
xor U17881 (N_17881,N_15245,N_16956);
or U17882 (N_17882,N_15986,N_16355);
and U17883 (N_17883,N_15917,N_15823);
nor U17884 (N_17884,N_16817,N_16761);
xnor U17885 (N_17885,N_16649,N_15745);
nor U17886 (N_17886,N_15741,N_15285);
and U17887 (N_17887,N_16908,N_15977);
xnor U17888 (N_17888,N_15752,N_17298);
xor U17889 (N_17889,N_15429,N_15145);
and U17890 (N_17890,N_15318,N_15252);
nand U17891 (N_17891,N_17436,N_15124);
or U17892 (N_17892,N_16732,N_15066);
xnor U17893 (N_17893,N_15840,N_16041);
or U17894 (N_17894,N_16028,N_16214);
or U17895 (N_17895,N_16107,N_15869);
nand U17896 (N_17896,N_17451,N_17101);
xnor U17897 (N_17897,N_16819,N_16861);
and U17898 (N_17898,N_16823,N_15425);
and U17899 (N_17899,N_16886,N_16899);
nor U17900 (N_17900,N_15697,N_16678);
nand U17901 (N_17901,N_15192,N_15568);
nand U17902 (N_17902,N_15077,N_16978);
xnor U17903 (N_17903,N_15409,N_15903);
and U17904 (N_17904,N_17400,N_16196);
xnor U17905 (N_17905,N_17107,N_16580);
or U17906 (N_17906,N_16120,N_15157);
and U17907 (N_17907,N_16794,N_15684);
nand U17908 (N_17908,N_16175,N_15338);
nor U17909 (N_17909,N_17034,N_16796);
nor U17910 (N_17910,N_15648,N_16937);
and U17911 (N_17911,N_16257,N_16951);
or U17912 (N_17912,N_16179,N_16378);
xor U17913 (N_17913,N_17409,N_16439);
nand U17914 (N_17914,N_16140,N_16267);
nor U17915 (N_17915,N_15279,N_15306);
and U17916 (N_17916,N_17015,N_15291);
nand U17917 (N_17917,N_17260,N_16125);
nand U17918 (N_17918,N_17435,N_17177);
or U17919 (N_17919,N_17411,N_16888);
xor U17920 (N_17920,N_15042,N_16721);
nor U17921 (N_17921,N_15474,N_15972);
nor U17922 (N_17922,N_15645,N_16916);
or U17923 (N_17923,N_15559,N_15607);
nor U17924 (N_17924,N_16667,N_15817);
nor U17925 (N_17925,N_15864,N_17090);
or U17926 (N_17926,N_15761,N_17233);
nand U17927 (N_17927,N_17050,N_15941);
xor U17928 (N_17928,N_17231,N_16783);
nor U17929 (N_17929,N_15832,N_16302);
and U17930 (N_17930,N_16426,N_16480);
xor U17931 (N_17931,N_15560,N_17314);
nor U17932 (N_17932,N_16848,N_16702);
nor U17933 (N_17933,N_16167,N_16147);
nor U17934 (N_17934,N_15633,N_15351);
or U17935 (N_17935,N_17304,N_17184);
and U17936 (N_17936,N_15659,N_17334);
xnor U17937 (N_17937,N_16444,N_16243);
xnor U17938 (N_17938,N_16305,N_16674);
and U17939 (N_17939,N_16206,N_16300);
xnor U17940 (N_17940,N_15994,N_16022);
or U17941 (N_17941,N_16503,N_15902);
nor U17942 (N_17942,N_15369,N_16373);
nand U17943 (N_17943,N_15871,N_15702);
xnor U17944 (N_17944,N_16498,N_17447);
and U17945 (N_17945,N_16831,N_17360);
and U17946 (N_17946,N_16451,N_16340);
xor U17947 (N_17947,N_15775,N_16767);
or U17948 (N_17948,N_15397,N_17127);
nor U17949 (N_17949,N_15915,N_16634);
xnor U17950 (N_17950,N_17079,N_16311);
or U17951 (N_17951,N_15846,N_15430);
nand U17952 (N_17952,N_15226,N_16339);
nand U17953 (N_17953,N_15604,N_15250);
xor U17954 (N_17954,N_17029,N_16463);
or U17955 (N_17955,N_17220,N_16822);
and U17956 (N_17956,N_16686,N_15196);
xnor U17957 (N_17957,N_15552,N_15625);
and U17958 (N_17958,N_16226,N_16512);
and U17959 (N_17959,N_15096,N_15667);
or U17960 (N_17960,N_15953,N_15542);
and U17961 (N_17961,N_16402,N_15495);
or U17962 (N_17962,N_17416,N_17126);
nand U17963 (N_17963,N_16705,N_16777);
and U17964 (N_17964,N_17087,N_16324);
and U17965 (N_17965,N_16166,N_15058);
nand U17966 (N_17966,N_15811,N_16048);
nand U17967 (N_17967,N_16038,N_15204);
nand U17968 (N_17968,N_16229,N_16377);
xnor U17969 (N_17969,N_15710,N_16344);
xor U17970 (N_17970,N_15107,N_15382);
or U17971 (N_17971,N_15443,N_15824);
xnor U17972 (N_17972,N_15357,N_15343);
or U17973 (N_17973,N_15815,N_15910);
or U17974 (N_17974,N_16601,N_16244);
and U17975 (N_17975,N_15905,N_15720);
nor U17976 (N_17976,N_17041,N_15234);
or U17977 (N_17977,N_15772,N_16119);
nand U17978 (N_17978,N_16995,N_16980);
nor U17979 (N_17979,N_17203,N_16265);
nor U17980 (N_17980,N_17037,N_17492);
xor U17981 (N_17981,N_15494,N_17484);
xnor U17982 (N_17982,N_15276,N_15822);
and U17983 (N_17983,N_15609,N_15966);
nand U17984 (N_17984,N_16131,N_16661);
nand U17985 (N_17985,N_16019,N_16073);
or U17986 (N_17986,N_15037,N_15178);
and U17987 (N_17987,N_16854,N_16651);
and U17988 (N_17988,N_15945,N_17109);
and U17989 (N_17989,N_15991,N_15109);
nand U17990 (N_17990,N_15551,N_17078);
nor U17991 (N_17991,N_16785,N_15313);
xor U17992 (N_17992,N_16004,N_15700);
nand U17993 (N_17993,N_16077,N_16086);
and U17994 (N_17994,N_17033,N_16225);
nand U17995 (N_17995,N_17450,N_16709);
nor U17996 (N_17996,N_15418,N_15200);
and U17997 (N_17997,N_15363,N_15615);
nand U17998 (N_17998,N_15696,N_15470);
xor U17999 (N_17999,N_15162,N_15916);
or U18000 (N_18000,N_15262,N_15466);
xor U18001 (N_18001,N_15647,N_15973);
nand U18002 (N_18002,N_16123,N_16231);
and U18003 (N_18003,N_16128,N_15699);
xor U18004 (N_18004,N_15998,N_15492);
or U18005 (N_18005,N_17320,N_15514);
nand U18006 (N_18006,N_16568,N_16137);
xnor U18007 (N_18007,N_15807,N_15330);
nor U18008 (N_18008,N_15573,N_16704);
nor U18009 (N_18009,N_15962,N_15188);
or U18010 (N_18010,N_16033,N_15548);
xor U18011 (N_18011,N_15453,N_15882);
xor U18012 (N_18012,N_16564,N_17071);
or U18013 (N_18013,N_16690,N_15639);
nand U18014 (N_18014,N_15620,N_17389);
or U18015 (N_18015,N_15709,N_16692);
and U18016 (N_18016,N_16114,N_16883);
or U18017 (N_18017,N_15176,N_16089);
xor U18018 (N_18018,N_15171,N_16915);
nand U18019 (N_18019,N_16712,N_17384);
or U18020 (N_18020,N_16977,N_16863);
or U18021 (N_18021,N_15237,N_15737);
and U18022 (N_18022,N_15654,N_16057);
xnor U18023 (N_18023,N_15850,N_15537);
and U18024 (N_18024,N_15371,N_16410);
and U18025 (N_18025,N_16075,N_15006);
nor U18026 (N_18026,N_17474,N_16955);
or U18027 (N_18027,N_16738,N_15013);
xnor U18028 (N_18028,N_16154,N_17427);
and U18029 (N_18029,N_15801,N_16187);
nor U18030 (N_18030,N_15718,N_15602);
nor U18031 (N_18031,N_17357,N_15191);
nor U18032 (N_18032,N_17085,N_17162);
or U18033 (N_18033,N_17441,N_16189);
nor U18034 (N_18034,N_15632,N_16333);
or U18035 (N_18035,N_15335,N_15044);
and U18036 (N_18036,N_15007,N_17136);
and U18037 (N_18037,N_16896,N_15748);
nor U18038 (N_18038,N_16636,N_16798);
and U18039 (N_18039,N_15478,N_15045);
or U18040 (N_18040,N_15906,N_16770);
xnor U18041 (N_18041,N_16465,N_16860);
or U18042 (N_18042,N_16501,N_15753);
nor U18043 (N_18043,N_15692,N_16545);
xnor U18044 (N_18044,N_16904,N_15320);
nor U18045 (N_18045,N_16273,N_16023);
xor U18046 (N_18046,N_16505,N_17317);
nand U18047 (N_18047,N_16947,N_16384);
nor U18048 (N_18048,N_16430,N_17473);
nor U18049 (N_18049,N_16701,N_15878);
nand U18050 (N_18050,N_16101,N_15345);
xnor U18051 (N_18051,N_16090,N_17131);
nor U18052 (N_18052,N_17463,N_15501);
and U18053 (N_18053,N_16032,N_15894);
or U18054 (N_18054,N_15404,N_15856);
and U18055 (N_18055,N_15867,N_16805);
and U18056 (N_18056,N_16190,N_15093);
nor U18057 (N_18057,N_15386,N_16246);
and U18058 (N_18058,N_16158,N_15457);
and U18059 (N_18059,N_15268,N_15454);
nor U18060 (N_18060,N_15732,N_15545);
nand U18061 (N_18061,N_16719,N_16458);
or U18062 (N_18062,N_17318,N_15487);
nor U18063 (N_18063,N_17226,N_17157);
nand U18064 (N_18064,N_16838,N_15248);
xor U18065 (N_18065,N_15729,N_15420);
xnor U18066 (N_18066,N_17376,N_15713);
or U18067 (N_18067,N_16438,N_17060);
and U18068 (N_18068,N_16781,N_16666);
or U18069 (N_18069,N_15942,N_17362);
xnor U18070 (N_18070,N_15653,N_17258);
and U18071 (N_18071,N_16935,N_15057);
and U18072 (N_18072,N_15444,N_16882);
xnor U18073 (N_18073,N_16016,N_16765);
xnor U18074 (N_18074,N_16306,N_15160);
xor U18075 (N_18075,N_15965,N_16371);
or U18076 (N_18076,N_17189,N_15516);
xor U18077 (N_18077,N_16944,N_15377);
xor U18078 (N_18078,N_16116,N_16985);
and U18079 (N_18079,N_15215,N_16859);
nor U18080 (N_18080,N_16362,N_17181);
nor U18081 (N_18081,N_15536,N_15989);
xor U18082 (N_18082,N_16609,N_17292);
xnor U18083 (N_18083,N_16942,N_16973);
xnor U18084 (N_18084,N_15141,N_16202);
or U18085 (N_18085,N_15462,N_16132);
and U18086 (N_18086,N_16488,N_15642);
nand U18087 (N_18087,N_15049,N_16808);
nand U18088 (N_18088,N_16930,N_15489);
nor U18089 (N_18089,N_16806,N_16803);
xnor U18090 (N_18090,N_15450,N_16909);
xnor U18091 (N_18091,N_16992,N_15938);
or U18092 (N_18092,N_16348,N_17345);
nand U18093 (N_18093,N_16875,N_15005);
xor U18094 (N_18094,N_15666,N_16216);
nand U18095 (N_18095,N_15009,N_15169);
nand U18096 (N_18096,N_15374,N_15976);
nor U18097 (N_18097,N_17134,N_17125);
or U18098 (N_18098,N_17182,N_16113);
nand U18099 (N_18099,N_15164,N_15891);
nand U18100 (N_18100,N_16659,N_15473);
nor U18101 (N_18101,N_16933,N_16790);
nor U18102 (N_18102,N_16468,N_15831);
or U18103 (N_18103,N_16821,N_15553);
and U18104 (N_18104,N_16642,N_15445);
or U18105 (N_18105,N_16566,N_16628);
xnor U18106 (N_18106,N_16576,N_15827);
nor U18107 (N_18107,N_15802,N_15393);
nand U18108 (N_18108,N_15267,N_15367);
or U18109 (N_18109,N_16171,N_15198);
nand U18110 (N_18110,N_15036,N_15122);
or U18111 (N_18111,N_15446,N_15968);
nor U18112 (N_18112,N_16037,N_16968);
nor U18113 (N_18113,N_17394,N_16052);
and U18114 (N_18114,N_17349,N_15287);
nand U18115 (N_18115,N_15264,N_15624);
or U18116 (N_18116,N_15821,N_16055);
xnor U18117 (N_18117,N_17038,N_16627);
xnor U18118 (N_18118,N_16069,N_15184);
nor U18119 (N_18119,N_16122,N_15834);
and U18120 (N_18120,N_17486,N_15379);
or U18121 (N_18121,N_16518,N_15577);
nand U18122 (N_18122,N_17370,N_15392);
xor U18123 (N_18123,N_17108,N_16217);
and U18124 (N_18124,N_16786,N_17449);
nor U18125 (N_18125,N_16215,N_16331);
or U18126 (N_18126,N_15179,N_16405);
xnor U18127 (N_18127,N_15787,N_17296);
and U18128 (N_18128,N_15460,N_15032);
nand U18129 (N_18129,N_16153,N_16726);
nand U18130 (N_18130,N_16188,N_16553);
and U18131 (N_18131,N_15970,N_15524);
and U18132 (N_18132,N_17467,N_15139);
nor U18133 (N_18133,N_17208,N_17481);
or U18134 (N_18134,N_16255,N_15080);
nand U18135 (N_18135,N_17145,N_15627);
or U18136 (N_18136,N_15949,N_15337);
nand U18137 (N_18137,N_15154,N_16619);
or U18138 (N_18138,N_15370,N_15278);
or U18139 (N_18139,N_16144,N_17271);
nand U18140 (N_18140,N_17241,N_17223);
and U18141 (N_18141,N_16297,N_15270);
and U18142 (N_18142,N_16275,N_16508);
nor U18143 (N_18143,N_15206,N_15312);
or U18144 (N_18144,N_16337,N_15183);
xnor U18145 (N_18145,N_15943,N_15705);
and U18146 (N_18146,N_17281,N_16008);
nor U18147 (N_18147,N_16260,N_16910);
nand U18148 (N_18148,N_17191,N_16735);
or U18149 (N_18149,N_17063,N_16080);
and U18150 (N_18150,N_15488,N_17176);
nand U18151 (N_18151,N_15630,N_17058);
or U18152 (N_18152,N_16836,N_16063);
and U18153 (N_18153,N_15231,N_15578);
or U18154 (N_18154,N_16161,N_16727);
nand U18155 (N_18155,N_17430,N_15364);
or U18156 (N_18156,N_15575,N_15507);
xnor U18157 (N_18157,N_16949,N_17001);
or U18158 (N_18158,N_16156,N_16997);
nand U18159 (N_18159,N_17094,N_15410);
and U18160 (N_18160,N_15017,N_15964);
and U18161 (N_18161,N_15557,N_15651);
xor U18162 (N_18162,N_16133,N_15208);
nor U18163 (N_18163,N_17404,N_15275);
and U18164 (N_18164,N_15233,N_16741);
nor U18165 (N_18165,N_15859,N_16533);
and U18166 (N_18166,N_17140,N_16358);
or U18167 (N_18167,N_16406,N_16211);
nand U18168 (N_18168,N_15911,N_15156);
and U18169 (N_18169,N_15680,N_17114);
nor U18170 (N_18170,N_15020,N_17163);
and U18171 (N_18171,N_16091,N_16878);
nor U18172 (N_18172,N_15975,N_15649);
nand U18173 (N_18173,N_15159,N_16645);
nor U18174 (N_18174,N_15806,N_15247);
or U18175 (N_18175,N_16025,N_16891);
nand U18176 (N_18176,N_15255,N_17319);
xnor U18177 (N_18177,N_16762,N_15671);
xnor U18178 (N_18178,N_15088,N_16369);
and U18179 (N_18179,N_16633,N_15307);
and U18180 (N_18180,N_16094,N_17077);
and U18181 (N_18181,N_15508,N_17478);
and U18182 (N_18182,N_16098,N_15995);
xnor U18183 (N_18183,N_16890,N_16024);
or U18184 (N_18184,N_15763,N_15738);
or U18185 (N_18185,N_15862,N_15493);
nor U18186 (N_18186,N_17113,N_16730);
nand U18187 (N_18187,N_16526,N_15918);
xor U18188 (N_18188,N_17230,N_15967);
nor U18189 (N_18189,N_17150,N_16989);
nand U18190 (N_18190,N_16551,N_17372);
or U18191 (N_18191,N_15421,N_17256);
nor U18192 (N_18192,N_16059,N_15390);
nand U18193 (N_18193,N_15131,N_17178);
xnor U18194 (N_18194,N_17188,N_17387);
or U18195 (N_18195,N_15663,N_15111);
or U18196 (N_18196,N_16020,N_16423);
xnor U18197 (N_18197,N_17059,N_15909);
xnor U18198 (N_18198,N_17180,N_17385);
nor U18199 (N_18199,N_16669,N_16855);
nor U18200 (N_18200,N_16495,N_17159);
or U18201 (N_18201,N_17019,N_15843);
nor U18202 (N_18202,N_16366,N_16604);
nand U18203 (N_18203,N_16979,N_15505);
nand U18204 (N_18204,N_16492,N_16961);
or U18205 (N_18205,N_16950,N_15527);
nand U18206 (N_18206,N_16271,N_16646);
xor U18207 (N_18207,N_15782,N_16393);
nor U18208 (N_18208,N_17255,N_15765);
xor U18209 (N_18209,N_17167,N_16322);
xor U18210 (N_18210,N_16003,N_15486);
and U18211 (N_18211,N_15048,N_15644);
xor U18212 (N_18212,N_16278,N_17418);
nor U18213 (N_18213,N_16764,N_15613);
or U18214 (N_18214,N_16407,N_16364);
nand U18215 (N_18215,N_17147,N_17200);
nand U18216 (N_18216,N_16039,N_16117);
nor U18217 (N_18217,N_17359,N_17135);
and U18218 (N_18218,N_17276,N_17488);
and U18219 (N_18219,N_16600,N_15436);
or U18220 (N_18220,N_16460,N_15984);
xor U18221 (N_18221,N_15115,N_16549);
nand U18222 (N_18222,N_15940,N_15170);
nor U18223 (N_18223,N_16663,N_17480);
nand U18224 (N_18224,N_15596,N_17412);
and U18225 (N_18225,N_15888,N_15326);
and U18226 (N_18226,N_16800,N_16828);
and U18227 (N_18227,N_15662,N_17036);
nand U18228 (N_18228,N_16792,N_15417);
nand U18229 (N_18229,N_15679,N_16502);
or U18230 (N_18230,N_16209,N_17431);
or U18231 (N_18231,N_17434,N_16818);
nor U18232 (N_18232,N_15034,N_17207);
xor U18233 (N_18233,N_15996,N_15152);
nand U18234 (N_18234,N_17268,N_16555);
xnor U18235 (N_18235,N_15074,N_16639);
and U18236 (N_18236,N_15589,N_15099);
or U18237 (N_18237,N_15001,N_16328);
xor U18238 (N_18238,N_15189,N_16605);
xnor U18239 (N_18239,N_17103,N_15259);
nand U18240 (N_18240,N_16963,N_16126);
xnor U18241 (N_18241,N_17263,N_16849);
xnor U18242 (N_18242,N_15422,N_16440);
and U18243 (N_18243,N_16014,N_15323);
or U18244 (N_18244,N_16864,N_17439);
and U18245 (N_18245,N_16326,N_15936);
nand U18246 (N_18246,N_16290,N_15956);
nor U18247 (N_18247,N_15569,N_17091);
nor U18248 (N_18248,N_16920,N_15100);
xnor U18249 (N_18249,N_16291,N_16283);
nor U18250 (N_18250,N_16486,N_15321);
nor U18251 (N_18251,N_17002,N_16724);
xnor U18252 (N_18252,N_15636,N_15175);
nor U18253 (N_18253,N_16945,N_17350);
xor U18254 (N_18254,N_16862,N_16015);
nor U18255 (N_18255,N_17415,N_15983);
and U18256 (N_18256,N_15210,N_16162);
xnor U18257 (N_18257,N_16856,N_15541);
nand U18258 (N_18258,N_16652,N_15354);
nand U18259 (N_18259,N_16865,N_15825);
nand U18260 (N_18260,N_17161,N_17422);
and U18261 (N_18261,N_15329,N_16784);
nor U18262 (N_18262,N_15836,N_16539);
nand U18263 (N_18263,N_15796,N_16527);
nor U18264 (N_18264,N_16543,N_15491);
xor U18265 (N_18265,N_15523,N_17198);
nand U18266 (N_18266,N_16835,N_16589);
and U18267 (N_18267,N_15480,N_17092);
or U18268 (N_18268,N_16746,N_15315);
nand U18269 (N_18269,N_16847,N_16155);
xnor U18270 (N_18270,N_17007,N_15912);
and U18271 (N_18271,N_15000,N_15736);
nand U18272 (N_18272,N_15426,N_16769);
or U18273 (N_18273,N_16352,N_17356);
and U18274 (N_18274,N_16256,N_16247);
or U18275 (N_18275,N_15092,N_15467);
xor U18276 (N_18276,N_16810,N_17369);
nor U18277 (N_18277,N_17498,N_15123);
xnor U18278 (N_18278,N_15643,N_15728);
nand U18279 (N_18279,N_16287,N_16235);
and U18280 (N_18280,N_17102,N_16264);
nor U18281 (N_18281,N_16870,N_17458);
nand U18282 (N_18282,N_17124,N_15182);
xor U18283 (N_18283,N_15672,N_17219);
or U18284 (N_18284,N_15629,N_15529);
or U18285 (N_18285,N_17278,N_16521);
xor U18286 (N_18286,N_17229,N_15118);
and U18287 (N_18287,N_16843,N_16307);
nor U18288 (N_18288,N_16643,N_16901);
xnor U18289 (N_18289,N_15565,N_16026);
nand U18290 (N_18290,N_15598,N_17284);
xor U18291 (N_18291,N_16641,N_15758);
and U18292 (N_18292,N_15626,N_15483);
xnor U18293 (N_18293,N_16962,N_16165);
xor U18294 (N_18294,N_15490,N_17380);
or U18295 (N_18295,N_16682,N_15733);
and U18296 (N_18296,N_16776,N_17118);
nor U18297 (N_18297,N_17096,N_15969);
nand U18298 (N_18298,N_16232,N_15117);
or U18299 (N_18299,N_17164,N_15482);
xor U18300 (N_18300,N_15521,N_15762);
nand U18301 (N_18301,N_17327,N_16695);
xnor U18302 (N_18302,N_15428,N_16528);
xor U18303 (N_18303,N_15920,N_15634);
nor U18304 (N_18304,N_17133,N_17252);
and U18305 (N_18305,N_16343,N_16198);
nand U18306 (N_18306,N_16049,N_15812);
or U18307 (N_18307,N_15661,N_15742);
xor U18308 (N_18308,N_17080,N_16173);
xnor U18309 (N_18309,N_16424,N_15691);
xnor U18310 (N_18310,N_16124,N_15072);
or U18311 (N_18311,N_16079,N_15381);
and U18312 (N_18312,N_15173,N_17117);
xor U18313 (N_18313,N_15980,N_17212);
or U18314 (N_18314,N_15431,N_15308);
and U18315 (N_18315,N_17386,N_15071);
nor U18316 (N_18316,N_15067,N_15024);
nor U18317 (N_18317,N_16241,N_15929);
or U18318 (N_18318,N_16615,N_16403);
and U18319 (N_18319,N_16448,N_15712);
nand U18320 (N_18320,N_17347,N_15076);
and U18321 (N_18321,N_15706,N_16042);
or U18322 (N_18322,N_15586,N_16199);
nand U18323 (N_18323,N_16001,N_16176);
xor U18324 (N_18324,N_15860,N_16387);
or U18325 (N_18325,N_15698,N_15144);
nor U18326 (N_18326,N_15773,N_15701);
nand U18327 (N_18327,N_16394,N_17093);
and U18328 (N_18328,N_16408,N_15277);
xnor U18329 (N_18329,N_15652,N_16195);
and U18330 (N_18330,N_16263,N_17479);
or U18331 (N_18331,N_16253,N_15506);
nand U18332 (N_18332,N_15314,N_16504);
or U18333 (N_18333,N_16245,N_17460);
nand U18334 (N_18334,N_16740,N_15708);
or U18335 (N_18335,N_15688,N_16797);
nand U18336 (N_18336,N_16620,N_16060);
or U18337 (N_18337,N_15690,N_15530);
nor U18338 (N_18338,N_16230,N_15133);
nand U18339 (N_18339,N_15084,N_15027);
nand U18340 (N_18340,N_16676,N_15062);
xor U18341 (N_18341,N_15406,N_15126);
or U18342 (N_18342,N_17403,N_16885);
nor U18343 (N_18343,N_15461,N_16917);
or U18344 (N_18344,N_15711,N_17234);
xor U18345 (N_18345,N_15791,N_16370);
nand U18346 (N_18346,N_16395,N_17062);
or U18347 (N_18347,N_15383,N_16102);
xnor U18348 (N_18348,N_15366,N_15555);
nor U18349 (N_18349,N_15833,N_15395);
or U18350 (N_18350,N_16675,N_17377);
and U18351 (N_18351,N_17065,N_16749);
nand U18352 (N_18352,N_17469,N_15127);
xnor U18353 (N_18353,N_15086,N_17390);
nor U18354 (N_18354,N_16447,N_16418);
or U18355 (N_18355,N_16820,N_16940);
or U18356 (N_18356,N_16134,N_15469);
nor U18357 (N_18357,N_16353,N_16201);
xnor U18358 (N_18358,N_15402,N_16262);
nand U18359 (N_18359,N_15987,N_16906);
xnor U18360 (N_18360,N_16065,N_15232);
xnor U18361 (N_18361,N_15439,N_15332);
or U18362 (N_18362,N_15726,N_16832);
nand U18363 (N_18363,N_15818,N_15750);
nand U18364 (N_18364,N_16632,N_15358);
or U18365 (N_18365,N_15721,N_16804);
nor U18366 (N_18366,N_15328,N_16240);
nor U18367 (N_18367,N_15135,N_15303);
nand U18368 (N_18368,N_15441,N_16653);
nand U18369 (N_18369,N_16375,N_16151);
nand U18370 (N_18370,N_15520,N_16043);
and U18371 (N_18371,N_15167,N_15567);
xor U18372 (N_18372,N_15163,N_16288);
or U18373 (N_18373,N_15539,N_16677);
nand U18374 (N_18374,N_16983,N_15922);
xnor U18375 (N_18375,N_17407,N_15060);
nand U18376 (N_18376,N_16250,N_16927);
and U18377 (N_18377,N_17297,N_16357);
nand U18378 (N_18378,N_16103,N_16648);
nand U18379 (N_18379,N_17000,N_16184);
and U18380 (N_18380,N_16722,N_15703);
nor U18381 (N_18381,N_16121,N_15611);
nor U18382 (N_18382,N_17247,N_15500);
and U18383 (N_18383,N_16437,N_16207);
or U18384 (N_18384,N_17497,N_16873);
or U18385 (N_18385,N_15657,N_17279);
and U18386 (N_18386,N_16303,N_16027);
or U18387 (N_18387,N_17151,N_17475);
nor U18388 (N_18388,N_16778,N_15637);
or U18389 (N_18389,N_15153,N_16388);
and U18390 (N_18390,N_17340,N_17444);
nand U18391 (N_18391,N_16519,N_15260);
and U18392 (N_18392,N_16834,N_16320);
xor U18393 (N_18393,N_16507,N_16396);
nand U18394 (N_18394,N_15325,N_16149);
xor U18395 (N_18395,N_17003,N_15837);
nor U18396 (N_18396,N_16477,N_15053);
and U18397 (N_18397,N_17437,N_15070);
and U18398 (N_18398,N_16613,N_16579);
nor U18399 (N_18399,N_16304,N_17265);
and U18400 (N_18400,N_17310,N_16548);
xnor U18401 (N_18401,N_16994,N_16889);
nor U18402 (N_18402,N_15035,N_15181);
xnor U18403 (N_18403,N_17057,N_15477);
xnor U18404 (N_18404,N_17201,N_16145);
xnor U18405 (N_18405,N_15256,N_16592);
nand U18406 (N_18406,N_16456,N_17187);
nor U18407 (N_18407,N_17016,N_16991);
nor U18408 (N_18408,N_16556,N_16221);
and U18409 (N_18409,N_16365,N_15412);
nor U18410 (N_18410,N_16067,N_16829);
xor U18411 (N_18411,N_16993,N_16484);
nand U18412 (N_18412,N_16715,N_16239);
nor U18413 (N_18413,N_16876,N_17185);
nand U18414 (N_18414,N_15955,N_16483);
nand U18415 (N_18415,N_17154,N_15921);
nor U18416 (N_18416,N_16534,N_17325);
or U18417 (N_18417,N_15065,N_16325);
nand U18418 (N_18418,N_16203,N_16594);
and U18419 (N_18419,N_17013,N_17225);
or U18420 (N_18420,N_15549,N_16476);
and U18421 (N_18421,N_16174,N_17266);
nand U18422 (N_18422,N_17493,N_16499);
or U18423 (N_18423,N_15739,N_15993);
nand U18424 (N_18424,N_15458,N_16152);
xor U18425 (N_18425,N_15225,N_16139);
or U18426 (N_18426,N_17494,N_15041);
nor U18427 (N_18427,N_17072,N_16559);
and U18428 (N_18428,N_17088,N_17399);
xor U18429 (N_18429,N_16012,N_16431);
xor U18430 (N_18430,N_17010,N_15760);
or U18431 (N_18431,N_17472,N_16157);
or U18432 (N_18432,N_16868,N_16877);
nor U18433 (N_18433,N_17245,N_17199);
and U18434 (N_18434,N_15554,N_16801);
xor U18435 (N_18435,N_16869,N_16148);
and U18436 (N_18436,N_16846,N_15435);
xnor U18437 (N_18437,N_15475,N_15563);
and U18438 (N_18438,N_16830,N_16415);
and U18439 (N_18439,N_15193,N_17482);
or U18440 (N_18440,N_17337,N_15271);
nand U18441 (N_18441,N_17381,N_16581);
nor U18442 (N_18442,N_17364,N_16585);
and U18443 (N_18443,N_15400,N_17143);
and U18444 (N_18444,N_15138,N_15584);
or U18445 (N_18445,N_17056,N_16031);
nor U18446 (N_18446,N_15990,N_15852);
or U18447 (N_18447,N_15561,N_15950);
nor U18448 (N_18448,N_17326,N_16351);
nand U18449 (N_18449,N_17218,N_15258);
or U18450 (N_18450,N_15266,N_15317);
or U18451 (N_18451,N_17204,N_15515);
nand U18452 (N_18452,N_16194,N_15893);
and U18453 (N_18453,N_17355,N_16959);
and U18454 (N_18454,N_16874,N_16758);
and U18455 (N_18455,N_15026,N_16021);
and U18456 (N_18456,N_15361,N_15265);
or U18457 (N_18457,N_16638,N_16450);
nor U18458 (N_18458,N_15498,N_16660);
nand U18459 (N_18459,N_16092,N_15985);
or U18460 (N_18460,N_15899,N_16853);
or U18461 (N_18461,N_16926,N_16662);
xor U18462 (N_18462,N_17448,N_15056);
xor U18463 (N_18463,N_16922,N_16096);
xor U18464 (N_18464,N_16524,N_16567);
and U18465 (N_18465,N_17351,N_15413);
nand U18466 (N_18466,N_16237,N_15427);
xor U18467 (N_18467,N_16614,N_16007);
and U18468 (N_18468,N_15952,N_16998);
xor U18469 (N_18469,N_17194,N_16386);
nand U18470 (N_18470,N_15603,N_16744);
and U18471 (N_18471,N_15327,N_15059);
or U18472 (N_18472,N_16425,N_15873);
and U18473 (N_18473,N_15040,N_17174);
nor U18474 (N_18474,N_15069,N_15814);
xnor U18475 (N_18475,N_17323,N_15010);
nand U18476 (N_18476,N_15640,N_15786);
or U18477 (N_18477,N_17216,N_16531);
nand U18478 (N_18478,N_17051,N_16563);
and U18479 (N_18479,N_15540,N_17395);
nor U18480 (N_18480,N_15177,N_17367);
and U18481 (N_18481,N_17020,N_16274);
or U18482 (N_18482,N_17130,N_17361);
xnor U18483 (N_18483,N_16006,N_16720);
nand U18484 (N_18484,N_17294,N_15350);
or U18485 (N_18485,N_16118,N_15819);
and U18486 (N_18486,N_16881,N_15218);
or U18487 (N_18487,N_15479,N_15511);
or U18488 (N_18488,N_16685,N_16390);
nor U18489 (N_18489,N_16005,N_16893);
nand U18490 (N_18490,N_15982,N_17456);
and U18491 (N_18491,N_15924,N_16668);
nand U18492 (N_18492,N_15612,N_16017);
nor U18493 (N_18493,N_16238,N_15205);
and U18494 (N_18494,N_17453,N_17224);
nor U18495 (N_18495,N_15229,N_16136);
xnor U18496 (N_18496,N_16640,N_15242);
and U18497 (N_18497,N_15004,N_16054);
nor U18498 (N_18498,N_17030,N_16061);
xnor U18499 (N_18499,N_17221,N_17442);
xnor U18500 (N_18500,N_16789,N_15130);
and U18501 (N_18501,N_15471,N_17491);
xnor U18502 (N_18502,N_15566,N_16471);
and U18503 (N_18503,N_17175,N_15895);
xor U18504 (N_18504,N_16404,N_16710);
xnor U18505 (N_18505,N_16939,N_16884);
nor U18506 (N_18506,N_15078,N_15816);
and U18507 (N_18507,N_15932,N_15282);
nor U18508 (N_18508,N_16417,N_16469);
and U18509 (N_18509,N_16577,N_16779);
or U18510 (N_18510,N_16482,N_17017);
nor U18511 (N_18511,N_16334,N_17083);
nor U18512 (N_18512,N_15842,N_16522);
nand U18513 (N_18513,N_15082,N_15694);
nor U18514 (N_18514,N_15564,N_17139);
or U18515 (N_18515,N_17148,N_15838);
nand U18516 (N_18516,N_16289,N_15570);
and U18517 (N_18517,N_15213,N_16542);
or U18518 (N_18518,N_17428,N_17119);
xor U18519 (N_18519,N_15755,N_16911);
or U18520 (N_18520,N_16213,N_16336);
nand U18521 (N_18521,N_15865,N_16259);
nor U18522 (N_18522,N_17393,N_15388);
xnor U18523 (N_18523,N_17012,N_15203);
nand U18524 (N_18524,N_16538,N_16532);
nand U18525 (N_18525,N_16490,N_15456);
nor U18526 (N_18526,N_15219,N_15767);
nand U18527 (N_18527,N_17240,N_16578);
nand U18528 (N_18528,N_16671,N_15419);
nor U18529 (N_18529,N_16718,N_15433);
nand U18530 (N_18530,N_15594,N_15934);
and U18531 (N_18531,N_15779,N_17179);
nand U18532 (N_18532,N_16703,N_15858);
and U18533 (N_18533,N_15754,N_16452);
and U18534 (N_18534,N_15751,N_15438);
nand U18535 (N_18535,N_17305,N_16713);
or U18536 (N_18536,N_16813,N_15442);
or U18537 (N_18537,N_17055,N_17366);
or U18538 (N_18538,N_15064,N_16197);
nand U18539 (N_18539,N_16529,N_15112);
and U18540 (N_18540,N_15914,N_16965);
and U18541 (N_18541,N_15892,N_17280);
and U18542 (N_18542,N_16540,N_16359);
nor U18543 (N_18543,N_17021,N_15121);
nand U18544 (N_18544,N_16757,N_17272);
nand U18545 (N_18545,N_16453,N_17295);
nand U18546 (N_18546,N_16443,N_16294);
and U18547 (N_18547,N_17417,N_16185);
nor U18548 (N_18548,N_16286,N_16650);
or U18549 (N_18549,N_17283,N_15808);
or U18550 (N_18550,N_16432,N_16923);
and U18551 (N_18551,N_17006,N_17306);
or U18552 (N_18552,N_16372,N_15424);
and U18553 (N_18553,N_16361,N_15481);
xor U18554 (N_18554,N_16751,N_16368);
and U18555 (N_18555,N_15362,N_15319);
or U18556 (N_18556,N_15574,N_15525);
nand U18557 (N_18557,N_17227,N_15931);
nand U18558 (N_18558,N_15297,N_15137);
xnor U18559 (N_18559,N_16446,N_17098);
and U18560 (N_18560,N_16389,N_15316);
nand U18561 (N_18561,N_17018,N_15677);
xnor U18562 (N_18562,N_15675,N_15746);
xnor U18563 (N_18563,N_17112,N_16234);
and U18564 (N_18564,N_17027,N_16988);
nand U18565 (N_18565,N_16953,N_15061);
xnor U18566 (N_18566,N_17158,N_16252);
or U18567 (N_18567,N_16752,N_16461);
or U18568 (N_18568,N_15269,N_16812);
xnor U18569 (N_18569,N_17228,N_15874);
and U18570 (N_18570,N_16793,N_16867);
or U18571 (N_18571,N_16433,N_16773);
or U18572 (N_18572,N_15384,N_15853);
xor U18573 (N_18573,N_15518,N_16772);
nor U18574 (N_18574,N_16575,N_17341);
nand U18575 (N_18575,N_15288,N_16383);
xnor U18576 (N_18576,N_17388,N_15759);
nand U18577 (N_18577,N_15376,N_15134);
and U18578 (N_18578,N_16664,N_15432);
nand U18579 (N_18579,N_17489,N_15434);
nor U18580 (N_18580,N_16591,N_15273);
and U18581 (N_18581,N_15120,N_16319);
or U18582 (N_18582,N_17121,N_15695);
nand U18583 (N_18583,N_17335,N_16571);
or U18584 (N_18584,N_16506,N_17141);
nand U18585 (N_18585,N_16590,N_17368);
nand U18586 (N_18586,N_17277,N_15484);
or U18587 (N_18587,N_17152,N_17383);
or U18588 (N_18588,N_16570,N_15556);
and U18589 (N_18589,N_16109,N_16918);
nor U18590 (N_18590,N_17183,N_16233);
nor U18591 (N_18591,N_16298,N_16697);
and U18592 (N_18592,N_16200,N_17401);
xnor U18593 (N_18593,N_15195,N_15519);
or U18594 (N_18594,N_15230,N_15777);
or U18595 (N_18595,N_15063,N_15054);
nor U18596 (N_18596,N_17374,N_15502);
nor U18597 (N_18597,N_15254,N_15590);
or U18598 (N_18598,N_15783,N_15105);
and U18599 (N_18599,N_17106,N_15448);
nand U18600 (N_18600,N_16301,N_17432);
nand U18601 (N_18601,N_15011,N_15880);
nand U18602 (N_18602,N_16560,N_16269);
or U18603 (N_18603,N_15301,N_15614);
and U18604 (N_18604,N_15670,N_16850);
nand U18605 (N_18605,N_15960,N_16750);
or U18606 (N_18606,N_17011,N_17286);
and U18607 (N_18607,N_16341,N_15216);
and U18608 (N_18608,N_17353,N_16276);
and U18609 (N_18609,N_16064,N_16315);
nor U18610 (N_18610,N_16759,N_15550);
xnor U18611 (N_18611,N_17375,N_16068);
nor U18612 (N_18612,N_16616,N_16872);
and U18613 (N_18613,N_16747,N_16279);
nand U18614 (N_18614,N_16903,N_15272);
xnor U18615 (N_18615,N_16106,N_17237);
and U18616 (N_18616,N_17146,N_16557);
or U18617 (N_18617,N_16093,N_15236);
and U18618 (N_18618,N_17483,N_16523);
and U18619 (N_18619,N_16385,N_16318);
xor U18620 (N_18620,N_15030,N_17171);
or U18621 (N_18621,N_17406,N_16228);
or U18622 (N_18622,N_17173,N_15309);
or U18623 (N_18623,N_17149,N_16934);
and U18624 (N_18624,N_15398,N_16837);
nor U18625 (N_18625,N_17064,N_15440);
nand U18626 (N_18626,N_16374,N_15172);
nor U18627 (N_18627,N_16401,N_15380);
nor U18628 (N_18628,N_16392,N_16081);
xor U18629 (N_18629,N_15725,N_17365);
xor U18630 (N_18630,N_16088,N_16584);
xor U18631 (N_18631,N_15535,N_15585);
nand U18632 (N_18632,N_15051,N_17257);
nor U18633 (N_18633,N_15003,N_16986);
and U18634 (N_18634,N_15890,N_15717);
xnor U18635 (N_18635,N_15794,N_16623);
and U18636 (N_18636,N_17137,N_17165);
or U18637 (N_18637,N_16964,N_16826);
nand U18638 (N_18638,N_15799,N_15749);
nor U18639 (N_18639,N_17166,N_15784);
or U18640 (N_18640,N_17423,N_15295);
nand U18641 (N_18641,N_17045,N_15735);
nand U18642 (N_18642,N_17128,N_15997);
and U18643 (N_18643,N_16180,N_15050);
or U18644 (N_18644,N_15740,N_15339);
nand U18645 (N_18645,N_17244,N_16516);
nand U18646 (N_18646,N_16419,N_16554);
or U18647 (N_18647,N_15459,N_17313);
nor U18648 (N_18648,N_15089,N_16222);
nand U18649 (N_18649,N_15879,N_16277);
or U18650 (N_18650,N_16053,N_16356);
and U18651 (N_18651,N_15992,N_16018);
xor U18652 (N_18652,N_15046,N_17352);
nand U18653 (N_18653,N_15292,N_15455);
and U18654 (N_18654,N_17433,N_16284);
nor U18655 (N_18655,N_15963,N_16656);
or U18656 (N_18656,N_16110,N_15841);
nand U18657 (N_18657,N_16058,N_16193);
nor U18658 (N_18658,N_16929,N_15158);
xor U18659 (N_18659,N_16363,N_15504);
nor U18660 (N_18660,N_17099,N_15150);
or U18661 (N_18661,N_15884,N_15496);
nor U18662 (N_18662,N_15655,N_15933);
and U18663 (N_18663,N_16684,N_16644);
and U18664 (N_18664,N_16841,N_15348);
nand U18665 (N_18665,N_15707,N_16925);
or U18666 (N_18666,N_15562,N_16975);
nor U18667 (N_18667,N_15588,N_15468);
nand U18668 (N_18668,N_15352,N_17495);
nor U18669 (N_18669,N_16657,N_16691);
xnor U18670 (N_18670,N_15988,N_17264);
nand U18671 (N_18671,N_16186,N_16958);
or U18672 (N_18672,N_16535,N_15411);
nor U18673 (N_18673,N_15128,N_15685);
nor U18674 (N_18674,N_17073,N_15008);
or U18675 (N_18675,N_16598,N_15497);
and U18676 (N_18676,N_16360,N_17081);
or U18677 (N_18677,N_16182,N_17097);
nor U18678 (N_18678,N_15734,N_16150);
xnor U18679 (N_18679,N_15897,N_15151);
nand U18680 (N_18680,N_16427,N_15186);
or U18681 (N_18681,N_15378,N_15387);
xor U18682 (N_18682,N_15770,N_16946);
or U18683 (N_18683,N_17466,N_16763);
and U18684 (N_18684,N_15324,N_16056);
nand U18685 (N_18685,N_16251,N_15901);
or U18686 (N_18686,N_16429,N_15780);
or U18687 (N_18687,N_16679,N_17331);
or U18688 (N_18688,N_16192,N_17044);
xor U18689 (N_18689,N_17193,N_16700);
xor U18690 (N_18690,N_15809,N_15635);
or U18691 (N_18691,N_16084,N_17095);
nand U18692 (N_18692,N_16208,N_15724);
or U18693 (N_18693,N_15877,N_15855);
and U18694 (N_18694,N_15223,N_16130);
nand U18695 (N_18695,N_15513,N_17274);
and U18696 (N_18696,N_17396,N_16723);
xnor U18697 (N_18697,N_16597,N_16332);
or U18698 (N_18698,N_16142,N_17066);
nor U18699 (N_18699,N_17047,N_17454);
and U18700 (N_18700,N_16321,N_16541);
and U18701 (N_18701,N_17328,N_16177);
xor U18702 (N_18702,N_16281,N_15532);
xnor U18703 (N_18703,N_16696,N_15641);
nor U18704 (N_18704,N_15202,N_16178);
nand U18705 (N_18705,N_16467,N_15587);
nand U18706 (N_18706,N_15012,N_16624);
or U18707 (N_18707,N_16104,N_15650);
nor U18708 (N_18708,N_16587,N_16780);
xnor U18709 (N_18709,N_15756,N_15533);
and U18710 (N_18710,N_16626,N_16693);
xor U18711 (N_18711,N_16414,N_17132);
nand U18712 (N_18712,N_15904,N_16071);
or U18713 (N_18713,N_15239,N_15347);
nand U18714 (N_18714,N_15803,N_17303);
nor U18715 (N_18715,N_15199,N_16000);
or U18716 (N_18716,N_16282,N_17046);
or U18717 (N_18717,N_16967,N_16596);
and U18718 (N_18718,N_16733,N_15597);
and U18719 (N_18719,N_16871,N_15686);
or U18720 (N_18720,N_17465,N_15683);
and U18721 (N_18721,N_15155,N_17111);
xnor U18722 (N_18722,N_16496,N_16473);
nand U18723 (N_18723,N_16924,N_15935);
xor U18724 (N_18724,N_15149,N_15284);
and U18725 (N_18725,N_16411,N_16493);
and U18726 (N_18726,N_17339,N_15704);
or U18727 (N_18727,N_16481,N_16606);
or U18728 (N_18728,N_16932,N_17253);
xnor U18729 (N_18729,N_17068,N_16936);
xor U18730 (N_18730,N_16346,N_15719);
nand U18731 (N_18731,N_16115,N_15875);
or U18732 (N_18732,N_16569,N_16510);
nor U18733 (N_18733,N_17358,N_15954);
and U18734 (N_18734,N_15792,N_15401);
nand U18735 (N_18735,N_15274,N_15243);
nand U18736 (N_18736,N_16990,N_16223);
or U18737 (N_18737,N_15687,N_15211);
xnor U18738 (N_18738,N_16530,N_16537);
and U18739 (N_18739,N_16459,N_15820);
xor U18740 (N_18740,N_17023,N_15937);
nand U18741 (N_18741,N_15776,N_17100);
and U18742 (N_18742,N_17089,N_16381);
or U18743 (N_18743,N_16112,N_17267);
nor U18744 (N_18744,N_15665,N_15098);
xor U18745 (N_18745,N_17496,N_15263);
nand U18746 (N_18746,N_16565,N_15116);
and U18747 (N_18747,N_15110,N_17039);
nand U18748 (N_18748,N_17344,N_17414);
xnor U18749 (N_18749,N_17259,N_16825);
nor U18750 (N_18750,N_16460,N_16172);
nor U18751 (N_18751,N_15094,N_16540);
nand U18752 (N_18752,N_16724,N_17102);
and U18753 (N_18753,N_15807,N_15753);
and U18754 (N_18754,N_15675,N_16313);
xor U18755 (N_18755,N_15237,N_15082);
nor U18756 (N_18756,N_15711,N_17460);
nor U18757 (N_18757,N_16648,N_16984);
or U18758 (N_18758,N_15744,N_15344);
xnor U18759 (N_18759,N_16132,N_15898);
xnor U18760 (N_18760,N_17416,N_15801);
xor U18761 (N_18761,N_17077,N_15097);
or U18762 (N_18762,N_15873,N_15297);
nand U18763 (N_18763,N_15721,N_16560);
nor U18764 (N_18764,N_15101,N_17130);
xor U18765 (N_18765,N_16155,N_16504);
xor U18766 (N_18766,N_16083,N_15111);
nand U18767 (N_18767,N_15985,N_16409);
xnor U18768 (N_18768,N_16229,N_15195);
and U18769 (N_18769,N_16887,N_15193);
and U18770 (N_18770,N_15613,N_15744);
xnor U18771 (N_18771,N_17030,N_17366);
xnor U18772 (N_18772,N_16391,N_16416);
xor U18773 (N_18773,N_17033,N_16143);
nor U18774 (N_18774,N_17096,N_16330);
nor U18775 (N_18775,N_16049,N_16862);
or U18776 (N_18776,N_16131,N_16880);
nor U18777 (N_18777,N_16213,N_17207);
nor U18778 (N_18778,N_17084,N_16594);
nand U18779 (N_18779,N_15413,N_16292);
nand U18780 (N_18780,N_15957,N_16511);
and U18781 (N_18781,N_17428,N_17134);
or U18782 (N_18782,N_16987,N_17157);
and U18783 (N_18783,N_15699,N_16272);
and U18784 (N_18784,N_15754,N_15732);
and U18785 (N_18785,N_15623,N_17315);
and U18786 (N_18786,N_15394,N_15639);
or U18787 (N_18787,N_16450,N_17276);
or U18788 (N_18788,N_16252,N_17143);
nand U18789 (N_18789,N_16436,N_16425);
xnor U18790 (N_18790,N_16763,N_16752);
nand U18791 (N_18791,N_17310,N_15958);
and U18792 (N_18792,N_16782,N_16911);
xnor U18793 (N_18793,N_16431,N_16100);
xnor U18794 (N_18794,N_17098,N_15702);
or U18795 (N_18795,N_15369,N_16014);
nand U18796 (N_18796,N_15951,N_16554);
and U18797 (N_18797,N_17173,N_17260);
nor U18798 (N_18798,N_15902,N_15189);
nand U18799 (N_18799,N_17491,N_16641);
xor U18800 (N_18800,N_16667,N_17403);
nor U18801 (N_18801,N_15301,N_16024);
or U18802 (N_18802,N_16881,N_15341);
and U18803 (N_18803,N_16856,N_15447);
nor U18804 (N_18804,N_15290,N_16630);
nand U18805 (N_18805,N_15902,N_17263);
xor U18806 (N_18806,N_17453,N_15229);
nor U18807 (N_18807,N_15972,N_15415);
xnor U18808 (N_18808,N_16287,N_17011);
nor U18809 (N_18809,N_15534,N_16970);
nand U18810 (N_18810,N_16748,N_16283);
and U18811 (N_18811,N_17354,N_16012);
nand U18812 (N_18812,N_16383,N_16001);
nor U18813 (N_18813,N_16963,N_17113);
and U18814 (N_18814,N_17100,N_16921);
or U18815 (N_18815,N_17216,N_17325);
and U18816 (N_18816,N_16439,N_17372);
or U18817 (N_18817,N_16067,N_15867);
nand U18818 (N_18818,N_15766,N_16565);
nor U18819 (N_18819,N_16681,N_15940);
or U18820 (N_18820,N_16622,N_15078);
and U18821 (N_18821,N_15386,N_16961);
nand U18822 (N_18822,N_16882,N_16038);
xor U18823 (N_18823,N_15307,N_16876);
xor U18824 (N_18824,N_17200,N_16160);
nor U18825 (N_18825,N_16777,N_15578);
xor U18826 (N_18826,N_17353,N_15223);
nand U18827 (N_18827,N_15158,N_17262);
or U18828 (N_18828,N_15797,N_15917);
or U18829 (N_18829,N_16954,N_16485);
and U18830 (N_18830,N_15660,N_16399);
xnor U18831 (N_18831,N_15833,N_16828);
xnor U18832 (N_18832,N_15756,N_15761);
and U18833 (N_18833,N_15249,N_15204);
and U18834 (N_18834,N_15906,N_15635);
nor U18835 (N_18835,N_15639,N_17362);
or U18836 (N_18836,N_16690,N_17146);
nor U18837 (N_18837,N_16584,N_16243);
and U18838 (N_18838,N_15913,N_16876);
xnor U18839 (N_18839,N_15311,N_16721);
nand U18840 (N_18840,N_15684,N_16153);
and U18841 (N_18841,N_17030,N_16730);
nand U18842 (N_18842,N_15206,N_15477);
xnor U18843 (N_18843,N_16764,N_15234);
or U18844 (N_18844,N_15655,N_17023);
and U18845 (N_18845,N_15202,N_16645);
or U18846 (N_18846,N_17423,N_16323);
nand U18847 (N_18847,N_16313,N_16549);
xor U18848 (N_18848,N_16088,N_17286);
nor U18849 (N_18849,N_16352,N_16342);
nor U18850 (N_18850,N_16946,N_16230);
or U18851 (N_18851,N_16619,N_17337);
and U18852 (N_18852,N_16813,N_15981);
xnor U18853 (N_18853,N_17457,N_15434);
nand U18854 (N_18854,N_15830,N_16770);
nand U18855 (N_18855,N_17121,N_17320);
xor U18856 (N_18856,N_16642,N_16547);
and U18857 (N_18857,N_17105,N_16772);
or U18858 (N_18858,N_16161,N_16496);
or U18859 (N_18859,N_15482,N_16222);
or U18860 (N_18860,N_17327,N_15387);
nor U18861 (N_18861,N_15928,N_16652);
xnor U18862 (N_18862,N_17030,N_15036);
xnor U18863 (N_18863,N_16379,N_15574);
nand U18864 (N_18864,N_16204,N_16968);
and U18865 (N_18865,N_17280,N_16576);
xor U18866 (N_18866,N_15043,N_17290);
xnor U18867 (N_18867,N_15281,N_16269);
nand U18868 (N_18868,N_17193,N_17360);
and U18869 (N_18869,N_15216,N_15870);
nand U18870 (N_18870,N_15720,N_16919);
and U18871 (N_18871,N_16454,N_15755);
and U18872 (N_18872,N_17300,N_15640);
or U18873 (N_18873,N_16335,N_15591);
nand U18874 (N_18874,N_16856,N_17481);
or U18875 (N_18875,N_15081,N_16928);
nand U18876 (N_18876,N_16758,N_15131);
or U18877 (N_18877,N_15415,N_16423);
nor U18878 (N_18878,N_17092,N_16192);
or U18879 (N_18879,N_16811,N_15597);
or U18880 (N_18880,N_15817,N_16267);
and U18881 (N_18881,N_15774,N_15819);
and U18882 (N_18882,N_16086,N_15962);
nand U18883 (N_18883,N_15254,N_16562);
nor U18884 (N_18884,N_16158,N_15520);
and U18885 (N_18885,N_16628,N_16106);
xnor U18886 (N_18886,N_17475,N_16020);
xnor U18887 (N_18887,N_16220,N_17360);
nor U18888 (N_18888,N_15762,N_17087);
and U18889 (N_18889,N_15286,N_15696);
nand U18890 (N_18890,N_16573,N_15178);
xor U18891 (N_18891,N_16431,N_16679);
nor U18892 (N_18892,N_16515,N_16512);
nor U18893 (N_18893,N_15211,N_15484);
or U18894 (N_18894,N_16071,N_16053);
nand U18895 (N_18895,N_15179,N_15906);
nand U18896 (N_18896,N_15521,N_16860);
and U18897 (N_18897,N_16333,N_15954);
nand U18898 (N_18898,N_16376,N_15634);
nor U18899 (N_18899,N_16213,N_17173);
xnor U18900 (N_18900,N_15625,N_16093);
nand U18901 (N_18901,N_16332,N_16523);
nand U18902 (N_18902,N_15422,N_16277);
xor U18903 (N_18903,N_16013,N_16294);
and U18904 (N_18904,N_15219,N_15110);
and U18905 (N_18905,N_15930,N_16527);
nor U18906 (N_18906,N_16131,N_15901);
nor U18907 (N_18907,N_15651,N_16042);
and U18908 (N_18908,N_15285,N_16684);
xnor U18909 (N_18909,N_15252,N_16428);
and U18910 (N_18910,N_17151,N_15576);
nand U18911 (N_18911,N_16055,N_15308);
or U18912 (N_18912,N_15160,N_15116);
nor U18913 (N_18913,N_15285,N_16543);
nor U18914 (N_18914,N_15524,N_16788);
nor U18915 (N_18915,N_15725,N_17462);
and U18916 (N_18916,N_15896,N_15478);
nand U18917 (N_18917,N_15959,N_15412);
xor U18918 (N_18918,N_16694,N_16434);
and U18919 (N_18919,N_16949,N_16286);
nand U18920 (N_18920,N_17180,N_17179);
and U18921 (N_18921,N_17338,N_15627);
or U18922 (N_18922,N_17370,N_16342);
xor U18923 (N_18923,N_15359,N_16051);
xnor U18924 (N_18924,N_15175,N_16211);
xnor U18925 (N_18925,N_15294,N_17214);
nand U18926 (N_18926,N_16325,N_15886);
nand U18927 (N_18927,N_16210,N_16223);
and U18928 (N_18928,N_16810,N_16355);
or U18929 (N_18929,N_16883,N_15358);
or U18930 (N_18930,N_15917,N_16302);
nand U18931 (N_18931,N_16922,N_16478);
and U18932 (N_18932,N_15151,N_17098);
and U18933 (N_18933,N_15256,N_15434);
nor U18934 (N_18934,N_15861,N_17354);
and U18935 (N_18935,N_16637,N_15810);
xor U18936 (N_18936,N_15348,N_17044);
xnor U18937 (N_18937,N_15899,N_15677);
nand U18938 (N_18938,N_15470,N_17285);
and U18939 (N_18939,N_15621,N_16090);
and U18940 (N_18940,N_16409,N_17252);
xnor U18941 (N_18941,N_17264,N_15739);
or U18942 (N_18942,N_15550,N_16065);
nand U18943 (N_18943,N_16064,N_15609);
nand U18944 (N_18944,N_16426,N_16209);
nand U18945 (N_18945,N_15120,N_16180);
or U18946 (N_18946,N_15116,N_15426);
nand U18947 (N_18947,N_17116,N_17350);
nand U18948 (N_18948,N_16203,N_16667);
and U18949 (N_18949,N_16831,N_16445);
or U18950 (N_18950,N_15251,N_15958);
or U18951 (N_18951,N_15097,N_15704);
nand U18952 (N_18952,N_16708,N_15524);
or U18953 (N_18953,N_15621,N_17149);
nand U18954 (N_18954,N_16685,N_15706);
nor U18955 (N_18955,N_16905,N_15474);
nor U18956 (N_18956,N_17203,N_16254);
or U18957 (N_18957,N_16156,N_17212);
or U18958 (N_18958,N_17056,N_16437);
and U18959 (N_18959,N_16248,N_16031);
or U18960 (N_18960,N_16511,N_16353);
and U18961 (N_18961,N_17221,N_16480);
nor U18962 (N_18962,N_16870,N_16138);
xor U18963 (N_18963,N_16766,N_17104);
nor U18964 (N_18964,N_15647,N_17427);
xnor U18965 (N_18965,N_16961,N_15328);
or U18966 (N_18966,N_16592,N_17204);
xnor U18967 (N_18967,N_15054,N_15201);
nand U18968 (N_18968,N_16669,N_16693);
and U18969 (N_18969,N_15225,N_16584);
xor U18970 (N_18970,N_15835,N_15940);
nand U18971 (N_18971,N_15313,N_15195);
xnor U18972 (N_18972,N_15998,N_16124);
xor U18973 (N_18973,N_16753,N_15538);
or U18974 (N_18974,N_15006,N_16227);
nand U18975 (N_18975,N_15144,N_15826);
xnor U18976 (N_18976,N_16304,N_15023);
and U18977 (N_18977,N_15301,N_15024);
and U18978 (N_18978,N_15596,N_16416);
xnor U18979 (N_18979,N_15550,N_17474);
xnor U18980 (N_18980,N_17001,N_16197);
nor U18981 (N_18981,N_15211,N_16725);
nor U18982 (N_18982,N_17444,N_16626);
nand U18983 (N_18983,N_16223,N_15176);
or U18984 (N_18984,N_17440,N_15034);
or U18985 (N_18985,N_17306,N_15900);
nor U18986 (N_18986,N_15605,N_15555);
nor U18987 (N_18987,N_15753,N_15363);
or U18988 (N_18988,N_15479,N_17284);
nand U18989 (N_18989,N_15999,N_17109);
or U18990 (N_18990,N_16272,N_15887);
and U18991 (N_18991,N_16982,N_16491);
nor U18992 (N_18992,N_16320,N_17452);
nand U18993 (N_18993,N_16459,N_15814);
xnor U18994 (N_18994,N_16091,N_16139);
and U18995 (N_18995,N_15269,N_16579);
or U18996 (N_18996,N_17382,N_15949);
nor U18997 (N_18997,N_16298,N_17065);
or U18998 (N_18998,N_16499,N_16755);
and U18999 (N_18999,N_15005,N_16916);
or U19000 (N_19000,N_16998,N_16900);
or U19001 (N_19001,N_15186,N_17466);
xnor U19002 (N_19002,N_17378,N_15759);
nand U19003 (N_19003,N_15757,N_16019);
nor U19004 (N_19004,N_15181,N_16893);
nand U19005 (N_19005,N_17247,N_16628);
or U19006 (N_19006,N_15602,N_15161);
or U19007 (N_19007,N_16523,N_17392);
or U19008 (N_19008,N_16930,N_17239);
or U19009 (N_19009,N_16366,N_15890);
nand U19010 (N_19010,N_16237,N_15378);
nand U19011 (N_19011,N_15070,N_16374);
nand U19012 (N_19012,N_16075,N_15080);
or U19013 (N_19013,N_15343,N_15231);
nand U19014 (N_19014,N_15495,N_15210);
xor U19015 (N_19015,N_16612,N_16472);
or U19016 (N_19016,N_16532,N_16535);
nand U19017 (N_19017,N_15990,N_15671);
and U19018 (N_19018,N_15755,N_15416);
xor U19019 (N_19019,N_16983,N_15649);
xnor U19020 (N_19020,N_15567,N_16118);
xnor U19021 (N_19021,N_15912,N_16036);
or U19022 (N_19022,N_17119,N_15502);
xnor U19023 (N_19023,N_15633,N_15967);
or U19024 (N_19024,N_16956,N_15254);
nand U19025 (N_19025,N_16050,N_16744);
nand U19026 (N_19026,N_15432,N_16069);
xor U19027 (N_19027,N_15565,N_16646);
xor U19028 (N_19028,N_17229,N_15451);
and U19029 (N_19029,N_15412,N_15506);
xnor U19030 (N_19030,N_15778,N_16791);
nor U19031 (N_19031,N_15050,N_15992);
nand U19032 (N_19032,N_15426,N_15333);
nor U19033 (N_19033,N_15996,N_15771);
nand U19034 (N_19034,N_16000,N_16419);
xnor U19035 (N_19035,N_15577,N_15336);
and U19036 (N_19036,N_17065,N_15464);
and U19037 (N_19037,N_15378,N_15298);
xor U19038 (N_19038,N_16336,N_15891);
and U19039 (N_19039,N_15017,N_15565);
or U19040 (N_19040,N_15984,N_16917);
and U19041 (N_19041,N_16569,N_16208);
xor U19042 (N_19042,N_16291,N_16094);
nor U19043 (N_19043,N_17133,N_17411);
nor U19044 (N_19044,N_17211,N_16263);
nor U19045 (N_19045,N_17083,N_16110);
or U19046 (N_19046,N_16384,N_16310);
xor U19047 (N_19047,N_15753,N_17044);
and U19048 (N_19048,N_15764,N_16080);
nor U19049 (N_19049,N_17317,N_16269);
or U19050 (N_19050,N_15042,N_16505);
xor U19051 (N_19051,N_16020,N_15419);
nor U19052 (N_19052,N_16818,N_15228);
nor U19053 (N_19053,N_15268,N_15870);
or U19054 (N_19054,N_16369,N_16670);
nand U19055 (N_19055,N_15914,N_16176);
nand U19056 (N_19056,N_16641,N_17189);
or U19057 (N_19057,N_16664,N_16807);
nor U19058 (N_19058,N_16476,N_16408);
nand U19059 (N_19059,N_16953,N_16368);
nand U19060 (N_19060,N_16036,N_17299);
or U19061 (N_19061,N_16084,N_17186);
nand U19062 (N_19062,N_15741,N_15584);
xnor U19063 (N_19063,N_16707,N_15097);
nand U19064 (N_19064,N_16190,N_15694);
nor U19065 (N_19065,N_15318,N_16443);
xor U19066 (N_19066,N_16846,N_15238);
and U19067 (N_19067,N_15661,N_16523);
nor U19068 (N_19068,N_16168,N_16157);
nand U19069 (N_19069,N_16807,N_15254);
nor U19070 (N_19070,N_16023,N_15815);
nand U19071 (N_19071,N_16343,N_17202);
and U19072 (N_19072,N_16071,N_17332);
or U19073 (N_19073,N_15434,N_15785);
nor U19074 (N_19074,N_16136,N_17002);
or U19075 (N_19075,N_16660,N_15397);
or U19076 (N_19076,N_17450,N_16362);
and U19077 (N_19077,N_15090,N_16396);
nor U19078 (N_19078,N_15283,N_15511);
or U19079 (N_19079,N_15134,N_16370);
and U19080 (N_19080,N_15557,N_17086);
xor U19081 (N_19081,N_15732,N_16112);
xor U19082 (N_19082,N_16775,N_17310);
and U19083 (N_19083,N_17149,N_15510);
or U19084 (N_19084,N_17494,N_16485);
nor U19085 (N_19085,N_16725,N_16806);
or U19086 (N_19086,N_16633,N_15749);
nor U19087 (N_19087,N_15042,N_15251);
xor U19088 (N_19088,N_17094,N_15214);
and U19089 (N_19089,N_15769,N_16434);
nor U19090 (N_19090,N_16627,N_15485);
xor U19091 (N_19091,N_15686,N_17196);
and U19092 (N_19092,N_15574,N_15230);
nand U19093 (N_19093,N_16837,N_15092);
and U19094 (N_19094,N_15673,N_17488);
xnor U19095 (N_19095,N_17374,N_16449);
or U19096 (N_19096,N_16533,N_15702);
nor U19097 (N_19097,N_15455,N_16660);
and U19098 (N_19098,N_17237,N_16865);
nor U19099 (N_19099,N_15096,N_17008);
xor U19100 (N_19100,N_15743,N_15741);
nor U19101 (N_19101,N_15330,N_16176);
or U19102 (N_19102,N_15643,N_16579);
or U19103 (N_19103,N_15601,N_16255);
and U19104 (N_19104,N_15277,N_15648);
xnor U19105 (N_19105,N_17289,N_16190);
nand U19106 (N_19106,N_16889,N_15437);
xor U19107 (N_19107,N_15343,N_15925);
xnor U19108 (N_19108,N_15108,N_16904);
nor U19109 (N_19109,N_16507,N_16094);
and U19110 (N_19110,N_15519,N_17356);
xor U19111 (N_19111,N_16793,N_15923);
nor U19112 (N_19112,N_16522,N_15079);
nor U19113 (N_19113,N_16076,N_16691);
and U19114 (N_19114,N_17259,N_15295);
nor U19115 (N_19115,N_15140,N_16948);
xor U19116 (N_19116,N_16098,N_16610);
nor U19117 (N_19117,N_17391,N_16882);
and U19118 (N_19118,N_17311,N_16750);
nor U19119 (N_19119,N_16631,N_15816);
and U19120 (N_19120,N_16903,N_15259);
nor U19121 (N_19121,N_16896,N_15493);
nand U19122 (N_19122,N_15532,N_16141);
nand U19123 (N_19123,N_16950,N_15146);
and U19124 (N_19124,N_16440,N_15089);
or U19125 (N_19125,N_15202,N_17257);
xor U19126 (N_19126,N_16177,N_15736);
nor U19127 (N_19127,N_15604,N_15813);
nand U19128 (N_19128,N_15673,N_15794);
xor U19129 (N_19129,N_15695,N_15465);
nor U19130 (N_19130,N_15961,N_15216);
or U19131 (N_19131,N_16442,N_16834);
xnor U19132 (N_19132,N_15380,N_16445);
xor U19133 (N_19133,N_16403,N_17045);
and U19134 (N_19134,N_15345,N_16614);
and U19135 (N_19135,N_16094,N_16530);
nand U19136 (N_19136,N_17176,N_16476);
nand U19137 (N_19137,N_17251,N_17387);
xor U19138 (N_19138,N_16877,N_15558);
nand U19139 (N_19139,N_16764,N_15343);
or U19140 (N_19140,N_16688,N_16724);
and U19141 (N_19141,N_17213,N_16420);
nor U19142 (N_19142,N_15517,N_15144);
and U19143 (N_19143,N_15179,N_16425);
nor U19144 (N_19144,N_17383,N_16382);
or U19145 (N_19145,N_16266,N_16677);
nor U19146 (N_19146,N_16293,N_15775);
or U19147 (N_19147,N_15409,N_17145);
nand U19148 (N_19148,N_15328,N_16466);
nand U19149 (N_19149,N_15634,N_16142);
nand U19150 (N_19150,N_15426,N_16239);
and U19151 (N_19151,N_15502,N_16306);
and U19152 (N_19152,N_16892,N_15820);
or U19153 (N_19153,N_15611,N_16762);
or U19154 (N_19154,N_15399,N_15075);
nand U19155 (N_19155,N_15809,N_16520);
nand U19156 (N_19156,N_17311,N_15772);
or U19157 (N_19157,N_16519,N_16019);
nand U19158 (N_19158,N_15190,N_17400);
and U19159 (N_19159,N_16352,N_17000);
nand U19160 (N_19160,N_16063,N_15578);
and U19161 (N_19161,N_16403,N_17158);
and U19162 (N_19162,N_16187,N_15735);
and U19163 (N_19163,N_15638,N_15536);
and U19164 (N_19164,N_16312,N_17365);
nor U19165 (N_19165,N_16232,N_16754);
nor U19166 (N_19166,N_15097,N_15620);
nand U19167 (N_19167,N_17068,N_16885);
xor U19168 (N_19168,N_16345,N_17154);
and U19169 (N_19169,N_17175,N_15709);
xor U19170 (N_19170,N_15098,N_16795);
nand U19171 (N_19171,N_15519,N_15257);
xnor U19172 (N_19172,N_17044,N_17016);
xor U19173 (N_19173,N_15207,N_16390);
xnor U19174 (N_19174,N_16429,N_16294);
nor U19175 (N_19175,N_16219,N_16237);
nor U19176 (N_19176,N_16895,N_16757);
nand U19177 (N_19177,N_15003,N_16202);
xnor U19178 (N_19178,N_16836,N_17360);
or U19179 (N_19179,N_15024,N_15032);
nor U19180 (N_19180,N_16917,N_15185);
xnor U19181 (N_19181,N_15501,N_16626);
xor U19182 (N_19182,N_15415,N_15666);
and U19183 (N_19183,N_16299,N_17462);
nand U19184 (N_19184,N_15215,N_17065);
or U19185 (N_19185,N_16145,N_15496);
and U19186 (N_19186,N_16004,N_17219);
xnor U19187 (N_19187,N_15370,N_16343);
or U19188 (N_19188,N_16227,N_15209);
nand U19189 (N_19189,N_16151,N_15653);
and U19190 (N_19190,N_17248,N_17121);
or U19191 (N_19191,N_17340,N_15400);
xnor U19192 (N_19192,N_15663,N_16251);
nand U19193 (N_19193,N_16531,N_16251);
xnor U19194 (N_19194,N_15067,N_16715);
xor U19195 (N_19195,N_16968,N_15200);
and U19196 (N_19196,N_16942,N_16043);
nand U19197 (N_19197,N_16722,N_16776);
and U19198 (N_19198,N_15023,N_15450);
nor U19199 (N_19199,N_15348,N_15634);
nand U19200 (N_19200,N_15165,N_17110);
xnor U19201 (N_19201,N_15280,N_16776);
xor U19202 (N_19202,N_17097,N_17075);
and U19203 (N_19203,N_17196,N_16345);
or U19204 (N_19204,N_15508,N_16840);
or U19205 (N_19205,N_17474,N_16385);
xor U19206 (N_19206,N_15765,N_17487);
xnor U19207 (N_19207,N_16615,N_15342);
xnor U19208 (N_19208,N_15029,N_16381);
nand U19209 (N_19209,N_15475,N_16296);
xor U19210 (N_19210,N_16644,N_17260);
nor U19211 (N_19211,N_16846,N_15415);
and U19212 (N_19212,N_17452,N_15284);
xor U19213 (N_19213,N_16927,N_17307);
xnor U19214 (N_19214,N_16652,N_15762);
xnor U19215 (N_19215,N_15578,N_16243);
xnor U19216 (N_19216,N_16518,N_15557);
nand U19217 (N_19217,N_16281,N_15673);
nor U19218 (N_19218,N_15962,N_16899);
and U19219 (N_19219,N_17161,N_15956);
nand U19220 (N_19220,N_15283,N_15181);
nand U19221 (N_19221,N_15929,N_15612);
or U19222 (N_19222,N_16185,N_16243);
nand U19223 (N_19223,N_16388,N_16556);
nand U19224 (N_19224,N_17302,N_16506);
nor U19225 (N_19225,N_15136,N_16957);
nor U19226 (N_19226,N_15837,N_15451);
xnor U19227 (N_19227,N_15776,N_17363);
nor U19228 (N_19228,N_16701,N_16382);
nand U19229 (N_19229,N_16296,N_16992);
and U19230 (N_19230,N_16631,N_16281);
nor U19231 (N_19231,N_16606,N_17472);
or U19232 (N_19232,N_17379,N_16487);
nor U19233 (N_19233,N_16522,N_16417);
nand U19234 (N_19234,N_16627,N_15753);
xor U19235 (N_19235,N_17386,N_15855);
and U19236 (N_19236,N_16240,N_16925);
xor U19237 (N_19237,N_15284,N_16730);
and U19238 (N_19238,N_17236,N_16052);
and U19239 (N_19239,N_16805,N_17001);
nor U19240 (N_19240,N_15890,N_15899);
nor U19241 (N_19241,N_16587,N_16086);
and U19242 (N_19242,N_15690,N_15872);
or U19243 (N_19243,N_16362,N_17298);
nand U19244 (N_19244,N_16007,N_15654);
and U19245 (N_19245,N_15093,N_15932);
and U19246 (N_19246,N_17128,N_17121);
and U19247 (N_19247,N_16928,N_16584);
nor U19248 (N_19248,N_17241,N_15386);
or U19249 (N_19249,N_15005,N_16015);
xor U19250 (N_19250,N_16998,N_15773);
and U19251 (N_19251,N_15467,N_17365);
nand U19252 (N_19252,N_17224,N_16786);
nor U19253 (N_19253,N_15745,N_17474);
nor U19254 (N_19254,N_15061,N_15069);
nand U19255 (N_19255,N_17101,N_17430);
nand U19256 (N_19256,N_15128,N_15558);
and U19257 (N_19257,N_16597,N_16460);
nor U19258 (N_19258,N_16457,N_15018);
nor U19259 (N_19259,N_15916,N_15663);
nor U19260 (N_19260,N_16155,N_15517);
nand U19261 (N_19261,N_17337,N_15353);
xnor U19262 (N_19262,N_15804,N_17283);
and U19263 (N_19263,N_15149,N_16084);
xor U19264 (N_19264,N_17081,N_15561);
nand U19265 (N_19265,N_16400,N_16226);
and U19266 (N_19266,N_17410,N_17339);
nor U19267 (N_19267,N_17190,N_15533);
and U19268 (N_19268,N_15997,N_17315);
or U19269 (N_19269,N_16069,N_16929);
xnor U19270 (N_19270,N_16981,N_15728);
and U19271 (N_19271,N_15538,N_17047);
xnor U19272 (N_19272,N_16140,N_16991);
nor U19273 (N_19273,N_16322,N_15981);
and U19274 (N_19274,N_16883,N_16304);
and U19275 (N_19275,N_15719,N_15533);
and U19276 (N_19276,N_15945,N_15145);
nor U19277 (N_19277,N_15410,N_16497);
or U19278 (N_19278,N_16846,N_15879);
and U19279 (N_19279,N_15453,N_16242);
nor U19280 (N_19280,N_16535,N_15225);
xnor U19281 (N_19281,N_17195,N_15903);
nand U19282 (N_19282,N_16769,N_16490);
nor U19283 (N_19283,N_17285,N_16599);
nor U19284 (N_19284,N_16720,N_17205);
xor U19285 (N_19285,N_16035,N_15661);
nor U19286 (N_19286,N_15967,N_17270);
nor U19287 (N_19287,N_16582,N_15180);
and U19288 (N_19288,N_16562,N_16698);
or U19289 (N_19289,N_16428,N_16538);
or U19290 (N_19290,N_15879,N_17345);
nor U19291 (N_19291,N_15033,N_17161);
and U19292 (N_19292,N_17059,N_16657);
nor U19293 (N_19293,N_15186,N_15332);
or U19294 (N_19294,N_16846,N_15077);
nor U19295 (N_19295,N_15720,N_17078);
xor U19296 (N_19296,N_16852,N_15251);
or U19297 (N_19297,N_15822,N_15135);
or U19298 (N_19298,N_16002,N_16098);
xor U19299 (N_19299,N_16973,N_16301);
xnor U19300 (N_19300,N_15383,N_15332);
and U19301 (N_19301,N_16972,N_16472);
nand U19302 (N_19302,N_16340,N_15478);
nor U19303 (N_19303,N_15674,N_16016);
or U19304 (N_19304,N_15209,N_15726);
or U19305 (N_19305,N_15163,N_16077);
nand U19306 (N_19306,N_15327,N_16239);
and U19307 (N_19307,N_16755,N_17148);
or U19308 (N_19308,N_16460,N_15870);
or U19309 (N_19309,N_15312,N_17355);
nand U19310 (N_19310,N_16324,N_16891);
or U19311 (N_19311,N_16506,N_17148);
xnor U19312 (N_19312,N_17179,N_15209);
nand U19313 (N_19313,N_15661,N_15093);
nand U19314 (N_19314,N_15402,N_16426);
or U19315 (N_19315,N_16261,N_15160);
xnor U19316 (N_19316,N_16025,N_15033);
nand U19317 (N_19317,N_15340,N_17139);
nand U19318 (N_19318,N_16039,N_15562);
xnor U19319 (N_19319,N_15446,N_16362);
nand U19320 (N_19320,N_16945,N_17283);
nor U19321 (N_19321,N_15887,N_17040);
xnor U19322 (N_19322,N_15202,N_15777);
xor U19323 (N_19323,N_15948,N_17412);
and U19324 (N_19324,N_16614,N_15185);
nor U19325 (N_19325,N_15932,N_17205);
nand U19326 (N_19326,N_15040,N_15119);
nand U19327 (N_19327,N_16353,N_16697);
and U19328 (N_19328,N_17379,N_16929);
or U19329 (N_19329,N_16882,N_15645);
nor U19330 (N_19330,N_16434,N_15717);
xnor U19331 (N_19331,N_16827,N_15237);
nor U19332 (N_19332,N_15573,N_16715);
and U19333 (N_19333,N_15748,N_15553);
xnor U19334 (N_19334,N_15403,N_17088);
nand U19335 (N_19335,N_15333,N_16960);
or U19336 (N_19336,N_17136,N_15106);
and U19337 (N_19337,N_15090,N_16157);
nand U19338 (N_19338,N_16491,N_16010);
nand U19339 (N_19339,N_16554,N_15041);
or U19340 (N_19340,N_16991,N_15613);
nor U19341 (N_19341,N_17480,N_16154);
or U19342 (N_19342,N_15724,N_15544);
xor U19343 (N_19343,N_17142,N_17115);
or U19344 (N_19344,N_16199,N_17464);
nand U19345 (N_19345,N_15195,N_15185);
and U19346 (N_19346,N_16178,N_16108);
nand U19347 (N_19347,N_15363,N_15911);
xor U19348 (N_19348,N_16600,N_16195);
nand U19349 (N_19349,N_16992,N_16673);
nor U19350 (N_19350,N_17472,N_15384);
and U19351 (N_19351,N_17127,N_16619);
nand U19352 (N_19352,N_17131,N_17474);
xor U19353 (N_19353,N_16628,N_16133);
nor U19354 (N_19354,N_15666,N_16466);
xor U19355 (N_19355,N_15913,N_16045);
xnor U19356 (N_19356,N_16231,N_16117);
xor U19357 (N_19357,N_16448,N_15072);
and U19358 (N_19358,N_17005,N_15011);
nand U19359 (N_19359,N_16619,N_16394);
or U19360 (N_19360,N_17480,N_15140);
nand U19361 (N_19361,N_15105,N_16987);
nand U19362 (N_19362,N_15722,N_15493);
or U19363 (N_19363,N_15798,N_15175);
and U19364 (N_19364,N_15382,N_16721);
and U19365 (N_19365,N_16595,N_15576);
or U19366 (N_19366,N_17419,N_17059);
or U19367 (N_19367,N_17000,N_17022);
nor U19368 (N_19368,N_15207,N_16268);
or U19369 (N_19369,N_17110,N_16798);
or U19370 (N_19370,N_17261,N_16986);
nand U19371 (N_19371,N_15660,N_17060);
or U19372 (N_19372,N_16028,N_15661);
nor U19373 (N_19373,N_17026,N_17335);
and U19374 (N_19374,N_17076,N_15855);
and U19375 (N_19375,N_15341,N_15985);
and U19376 (N_19376,N_15161,N_17001);
xor U19377 (N_19377,N_15893,N_16749);
or U19378 (N_19378,N_16542,N_16084);
nand U19379 (N_19379,N_16011,N_16765);
nand U19380 (N_19380,N_16547,N_16353);
xnor U19381 (N_19381,N_16470,N_16474);
xor U19382 (N_19382,N_16506,N_16572);
xor U19383 (N_19383,N_16023,N_15031);
nor U19384 (N_19384,N_16242,N_15691);
nor U19385 (N_19385,N_16698,N_15643);
and U19386 (N_19386,N_17405,N_16436);
and U19387 (N_19387,N_15189,N_17073);
and U19388 (N_19388,N_17217,N_15840);
and U19389 (N_19389,N_16353,N_17039);
or U19390 (N_19390,N_16724,N_16781);
xor U19391 (N_19391,N_15081,N_17319);
and U19392 (N_19392,N_16779,N_16544);
or U19393 (N_19393,N_17232,N_16985);
nand U19394 (N_19394,N_15686,N_17242);
or U19395 (N_19395,N_15368,N_15557);
xor U19396 (N_19396,N_17496,N_16969);
or U19397 (N_19397,N_15342,N_15501);
or U19398 (N_19398,N_16478,N_16723);
nor U19399 (N_19399,N_16378,N_15890);
or U19400 (N_19400,N_17262,N_16660);
and U19401 (N_19401,N_16007,N_15295);
nor U19402 (N_19402,N_15666,N_17396);
nor U19403 (N_19403,N_16662,N_15724);
nor U19404 (N_19404,N_16244,N_15349);
nor U19405 (N_19405,N_17052,N_16134);
xnor U19406 (N_19406,N_15808,N_16365);
nor U19407 (N_19407,N_15161,N_17147);
and U19408 (N_19408,N_15856,N_16211);
or U19409 (N_19409,N_16809,N_17155);
or U19410 (N_19410,N_15313,N_15837);
nor U19411 (N_19411,N_16655,N_15181);
nand U19412 (N_19412,N_16542,N_16345);
xor U19413 (N_19413,N_15760,N_15426);
nand U19414 (N_19414,N_17454,N_15059);
nand U19415 (N_19415,N_16467,N_15479);
xor U19416 (N_19416,N_16920,N_15916);
or U19417 (N_19417,N_16665,N_15526);
nand U19418 (N_19418,N_16971,N_17357);
xor U19419 (N_19419,N_16724,N_16999);
nor U19420 (N_19420,N_16083,N_15698);
or U19421 (N_19421,N_15083,N_17075);
nor U19422 (N_19422,N_15365,N_16784);
and U19423 (N_19423,N_17288,N_16021);
nand U19424 (N_19424,N_15355,N_15114);
nand U19425 (N_19425,N_15912,N_16757);
xor U19426 (N_19426,N_15633,N_16235);
nand U19427 (N_19427,N_17424,N_15378);
and U19428 (N_19428,N_16095,N_17017);
or U19429 (N_19429,N_16019,N_15780);
nand U19430 (N_19430,N_16357,N_15042);
or U19431 (N_19431,N_16899,N_15904);
nand U19432 (N_19432,N_15305,N_16034);
nor U19433 (N_19433,N_17181,N_16179);
or U19434 (N_19434,N_16092,N_16041);
or U19435 (N_19435,N_16928,N_16548);
and U19436 (N_19436,N_15446,N_16613);
and U19437 (N_19437,N_16024,N_15055);
or U19438 (N_19438,N_15338,N_15624);
nor U19439 (N_19439,N_15705,N_15179);
nand U19440 (N_19440,N_16126,N_16513);
nor U19441 (N_19441,N_15759,N_16654);
nor U19442 (N_19442,N_15371,N_15399);
and U19443 (N_19443,N_15440,N_17305);
nand U19444 (N_19444,N_15895,N_15000);
xnor U19445 (N_19445,N_17208,N_16734);
nor U19446 (N_19446,N_15671,N_17014);
nor U19447 (N_19447,N_15157,N_17088);
and U19448 (N_19448,N_16163,N_17029);
nand U19449 (N_19449,N_16837,N_15364);
nand U19450 (N_19450,N_15317,N_17048);
xor U19451 (N_19451,N_15116,N_16237);
nand U19452 (N_19452,N_15804,N_15080);
and U19453 (N_19453,N_15203,N_16322);
xor U19454 (N_19454,N_15268,N_15592);
nand U19455 (N_19455,N_17294,N_17141);
nand U19456 (N_19456,N_16318,N_15713);
nor U19457 (N_19457,N_15959,N_16941);
or U19458 (N_19458,N_15025,N_16469);
nand U19459 (N_19459,N_16539,N_16032);
xor U19460 (N_19460,N_15065,N_17161);
xnor U19461 (N_19461,N_16400,N_15802);
and U19462 (N_19462,N_15677,N_16016);
or U19463 (N_19463,N_15368,N_16227);
nand U19464 (N_19464,N_15634,N_17262);
or U19465 (N_19465,N_17107,N_16569);
and U19466 (N_19466,N_15227,N_16282);
xor U19467 (N_19467,N_16015,N_17123);
nand U19468 (N_19468,N_17207,N_16728);
or U19469 (N_19469,N_15834,N_15800);
and U19470 (N_19470,N_15502,N_15339);
and U19471 (N_19471,N_15567,N_15714);
nand U19472 (N_19472,N_16635,N_15376);
nand U19473 (N_19473,N_16785,N_17328);
or U19474 (N_19474,N_16402,N_15451);
and U19475 (N_19475,N_17440,N_16663);
xor U19476 (N_19476,N_16670,N_17118);
nand U19477 (N_19477,N_16842,N_16653);
nand U19478 (N_19478,N_16363,N_16825);
nand U19479 (N_19479,N_15337,N_15738);
nand U19480 (N_19480,N_16743,N_15943);
nor U19481 (N_19481,N_16095,N_15373);
and U19482 (N_19482,N_15767,N_17417);
and U19483 (N_19483,N_15344,N_15395);
or U19484 (N_19484,N_15980,N_16525);
xnor U19485 (N_19485,N_17354,N_16742);
nand U19486 (N_19486,N_17387,N_15408);
nand U19487 (N_19487,N_17183,N_17226);
or U19488 (N_19488,N_16861,N_16888);
and U19489 (N_19489,N_16568,N_16157);
xor U19490 (N_19490,N_16054,N_16849);
nand U19491 (N_19491,N_16750,N_17244);
or U19492 (N_19492,N_15145,N_15019);
and U19493 (N_19493,N_16864,N_16195);
nor U19494 (N_19494,N_15985,N_15131);
or U19495 (N_19495,N_15586,N_17020);
and U19496 (N_19496,N_15356,N_15234);
nor U19497 (N_19497,N_16652,N_15453);
and U19498 (N_19498,N_16822,N_15438);
and U19499 (N_19499,N_17474,N_15126);
nor U19500 (N_19500,N_17046,N_16346);
and U19501 (N_19501,N_15362,N_15529);
and U19502 (N_19502,N_17019,N_16086);
xor U19503 (N_19503,N_15109,N_16752);
or U19504 (N_19504,N_15064,N_17057);
nor U19505 (N_19505,N_15128,N_16805);
and U19506 (N_19506,N_17062,N_15367);
nand U19507 (N_19507,N_15357,N_17423);
nor U19508 (N_19508,N_15785,N_15126);
and U19509 (N_19509,N_16970,N_17060);
nand U19510 (N_19510,N_16112,N_17425);
nand U19511 (N_19511,N_15050,N_15958);
nand U19512 (N_19512,N_16368,N_15859);
nor U19513 (N_19513,N_16457,N_16431);
nor U19514 (N_19514,N_15740,N_15685);
nand U19515 (N_19515,N_16248,N_17039);
nand U19516 (N_19516,N_17055,N_15850);
xor U19517 (N_19517,N_16098,N_16209);
xnor U19518 (N_19518,N_17371,N_16601);
or U19519 (N_19519,N_17122,N_15322);
nand U19520 (N_19520,N_15025,N_16691);
or U19521 (N_19521,N_16626,N_16791);
nand U19522 (N_19522,N_16250,N_15543);
nor U19523 (N_19523,N_15689,N_16520);
or U19524 (N_19524,N_15119,N_15580);
nor U19525 (N_19525,N_15183,N_15817);
and U19526 (N_19526,N_17230,N_16114);
or U19527 (N_19527,N_17108,N_15763);
xor U19528 (N_19528,N_17433,N_15297);
nor U19529 (N_19529,N_17014,N_16410);
nor U19530 (N_19530,N_16087,N_15291);
or U19531 (N_19531,N_17328,N_17212);
nand U19532 (N_19532,N_17304,N_15196);
or U19533 (N_19533,N_15158,N_16883);
xnor U19534 (N_19534,N_17014,N_15204);
and U19535 (N_19535,N_16055,N_16065);
nor U19536 (N_19536,N_16942,N_16209);
or U19537 (N_19537,N_15672,N_16911);
or U19538 (N_19538,N_16641,N_15607);
xnor U19539 (N_19539,N_15783,N_15364);
xnor U19540 (N_19540,N_16476,N_15750);
xnor U19541 (N_19541,N_16404,N_16831);
nand U19542 (N_19542,N_15339,N_17193);
xor U19543 (N_19543,N_15166,N_17472);
or U19544 (N_19544,N_16172,N_16020);
and U19545 (N_19545,N_15792,N_16459);
nor U19546 (N_19546,N_16988,N_15660);
xor U19547 (N_19547,N_17489,N_17259);
and U19548 (N_19548,N_17396,N_16786);
xor U19549 (N_19549,N_15992,N_16689);
nand U19550 (N_19550,N_15118,N_17130);
nor U19551 (N_19551,N_16082,N_16534);
and U19552 (N_19552,N_17494,N_17278);
xnor U19553 (N_19553,N_17274,N_16407);
nand U19554 (N_19554,N_16709,N_17031);
or U19555 (N_19555,N_16030,N_16399);
and U19556 (N_19556,N_16245,N_16861);
nand U19557 (N_19557,N_15582,N_16774);
nand U19558 (N_19558,N_15618,N_16343);
nor U19559 (N_19559,N_17139,N_16095);
xor U19560 (N_19560,N_15267,N_15247);
nor U19561 (N_19561,N_15857,N_16400);
nand U19562 (N_19562,N_16718,N_16431);
nand U19563 (N_19563,N_15191,N_16484);
nand U19564 (N_19564,N_16977,N_15618);
or U19565 (N_19565,N_17308,N_15257);
xnor U19566 (N_19566,N_15835,N_17094);
or U19567 (N_19567,N_16219,N_15734);
xor U19568 (N_19568,N_15731,N_16907);
or U19569 (N_19569,N_16335,N_16993);
or U19570 (N_19570,N_16658,N_16118);
xnor U19571 (N_19571,N_16586,N_17190);
nand U19572 (N_19572,N_15641,N_17074);
xor U19573 (N_19573,N_15127,N_15028);
xnor U19574 (N_19574,N_17434,N_15289);
nor U19575 (N_19575,N_15804,N_15747);
or U19576 (N_19576,N_15450,N_17220);
or U19577 (N_19577,N_15580,N_15469);
xnor U19578 (N_19578,N_16335,N_16688);
nand U19579 (N_19579,N_16797,N_16552);
and U19580 (N_19580,N_15717,N_15777);
or U19581 (N_19581,N_16408,N_15316);
xnor U19582 (N_19582,N_15448,N_16856);
or U19583 (N_19583,N_15743,N_17040);
xnor U19584 (N_19584,N_15860,N_15335);
or U19585 (N_19585,N_15820,N_15199);
xnor U19586 (N_19586,N_15376,N_17086);
and U19587 (N_19587,N_17425,N_15618);
and U19588 (N_19588,N_17298,N_16323);
xor U19589 (N_19589,N_15312,N_16095);
nand U19590 (N_19590,N_16051,N_15199);
nor U19591 (N_19591,N_17228,N_16023);
or U19592 (N_19592,N_17133,N_16389);
and U19593 (N_19593,N_15963,N_16239);
nor U19594 (N_19594,N_15447,N_15602);
and U19595 (N_19595,N_16357,N_16105);
xor U19596 (N_19596,N_16359,N_16124);
or U19597 (N_19597,N_15824,N_16239);
nand U19598 (N_19598,N_16805,N_16026);
nor U19599 (N_19599,N_16475,N_16602);
nor U19600 (N_19600,N_16851,N_16684);
xor U19601 (N_19601,N_17267,N_15754);
nand U19602 (N_19602,N_17363,N_15781);
or U19603 (N_19603,N_16554,N_17367);
and U19604 (N_19604,N_15984,N_16311);
nor U19605 (N_19605,N_15776,N_16449);
xor U19606 (N_19606,N_15084,N_15730);
and U19607 (N_19607,N_16108,N_16812);
and U19608 (N_19608,N_16599,N_17214);
or U19609 (N_19609,N_16324,N_17150);
xnor U19610 (N_19610,N_15222,N_15514);
or U19611 (N_19611,N_15494,N_17244);
and U19612 (N_19612,N_16811,N_15818);
xor U19613 (N_19613,N_15143,N_15892);
xor U19614 (N_19614,N_16521,N_16598);
nand U19615 (N_19615,N_15025,N_15324);
or U19616 (N_19616,N_16080,N_15228);
xor U19617 (N_19617,N_17052,N_16791);
and U19618 (N_19618,N_16399,N_16692);
nand U19619 (N_19619,N_17102,N_17198);
nor U19620 (N_19620,N_16856,N_16250);
xnor U19621 (N_19621,N_16013,N_16388);
nor U19622 (N_19622,N_17329,N_15414);
nand U19623 (N_19623,N_15010,N_15304);
nand U19624 (N_19624,N_16720,N_15599);
nor U19625 (N_19625,N_17380,N_16049);
xor U19626 (N_19626,N_15014,N_16884);
nand U19627 (N_19627,N_16078,N_16571);
and U19628 (N_19628,N_16439,N_15402);
or U19629 (N_19629,N_16274,N_15516);
and U19630 (N_19630,N_17354,N_17319);
or U19631 (N_19631,N_17470,N_15094);
nor U19632 (N_19632,N_16588,N_15497);
nor U19633 (N_19633,N_15872,N_15076);
and U19634 (N_19634,N_17155,N_17447);
xnor U19635 (N_19635,N_16791,N_15818);
xnor U19636 (N_19636,N_15252,N_16013);
and U19637 (N_19637,N_15611,N_16808);
xnor U19638 (N_19638,N_15549,N_16107);
or U19639 (N_19639,N_15565,N_16021);
or U19640 (N_19640,N_17471,N_15312);
xnor U19641 (N_19641,N_15192,N_15375);
xor U19642 (N_19642,N_17406,N_15440);
xnor U19643 (N_19643,N_17363,N_16777);
and U19644 (N_19644,N_16900,N_15905);
xor U19645 (N_19645,N_15418,N_15324);
nand U19646 (N_19646,N_16565,N_17228);
nor U19647 (N_19647,N_16340,N_15489);
or U19648 (N_19648,N_15927,N_16087);
nor U19649 (N_19649,N_16439,N_15462);
or U19650 (N_19650,N_15700,N_15346);
xor U19651 (N_19651,N_15200,N_16698);
nor U19652 (N_19652,N_15548,N_15899);
and U19653 (N_19653,N_16385,N_17102);
or U19654 (N_19654,N_15057,N_16442);
xnor U19655 (N_19655,N_16252,N_15041);
nand U19656 (N_19656,N_16539,N_17017);
or U19657 (N_19657,N_16929,N_17237);
nand U19658 (N_19658,N_15914,N_15721);
xor U19659 (N_19659,N_15805,N_17316);
and U19660 (N_19660,N_17467,N_16930);
or U19661 (N_19661,N_16334,N_16778);
nand U19662 (N_19662,N_15192,N_17007);
or U19663 (N_19663,N_16745,N_16833);
or U19664 (N_19664,N_15711,N_16226);
xnor U19665 (N_19665,N_16640,N_15209);
and U19666 (N_19666,N_17308,N_17488);
and U19667 (N_19667,N_17246,N_15952);
xor U19668 (N_19668,N_17074,N_15472);
nor U19669 (N_19669,N_15452,N_16270);
or U19670 (N_19670,N_15747,N_15772);
nand U19671 (N_19671,N_16620,N_16272);
nor U19672 (N_19672,N_16218,N_15942);
and U19673 (N_19673,N_16384,N_15255);
or U19674 (N_19674,N_15051,N_17294);
or U19675 (N_19675,N_17317,N_15824);
nor U19676 (N_19676,N_15355,N_17078);
nor U19677 (N_19677,N_15152,N_15878);
xnor U19678 (N_19678,N_15512,N_17227);
nand U19679 (N_19679,N_16418,N_15248);
xnor U19680 (N_19680,N_16180,N_17071);
xor U19681 (N_19681,N_15347,N_16840);
or U19682 (N_19682,N_16469,N_17405);
nor U19683 (N_19683,N_15948,N_16028);
nand U19684 (N_19684,N_15783,N_15412);
nor U19685 (N_19685,N_17439,N_17306);
and U19686 (N_19686,N_15666,N_16820);
xnor U19687 (N_19687,N_17071,N_15168);
and U19688 (N_19688,N_17125,N_16808);
xnor U19689 (N_19689,N_16247,N_17175);
xnor U19690 (N_19690,N_16844,N_17346);
and U19691 (N_19691,N_15288,N_17040);
xnor U19692 (N_19692,N_16784,N_17457);
nand U19693 (N_19693,N_15260,N_15994);
and U19694 (N_19694,N_16259,N_15441);
nor U19695 (N_19695,N_17368,N_16207);
or U19696 (N_19696,N_17377,N_16133);
xor U19697 (N_19697,N_17323,N_17047);
xnor U19698 (N_19698,N_16424,N_15325);
xor U19699 (N_19699,N_15229,N_16101);
nand U19700 (N_19700,N_15006,N_17482);
and U19701 (N_19701,N_15731,N_16568);
nor U19702 (N_19702,N_17463,N_16168);
or U19703 (N_19703,N_16708,N_15627);
nor U19704 (N_19704,N_15193,N_16474);
nor U19705 (N_19705,N_16110,N_17241);
nor U19706 (N_19706,N_16164,N_16090);
xor U19707 (N_19707,N_15990,N_16680);
xor U19708 (N_19708,N_16862,N_15699);
xor U19709 (N_19709,N_16270,N_16800);
or U19710 (N_19710,N_16641,N_16215);
nand U19711 (N_19711,N_15130,N_15446);
nand U19712 (N_19712,N_16914,N_17055);
and U19713 (N_19713,N_15431,N_15141);
or U19714 (N_19714,N_16692,N_17218);
xnor U19715 (N_19715,N_15339,N_15269);
and U19716 (N_19716,N_15737,N_15058);
or U19717 (N_19717,N_16842,N_15755);
xnor U19718 (N_19718,N_17417,N_15372);
nand U19719 (N_19719,N_15399,N_15789);
or U19720 (N_19720,N_15392,N_17260);
nor U19721 (N_19721,N_17388,N_16901);
or U19722 (N_19722,N_15984,N_16435);
nand U19723 (N_19723,N_15888,N_16650);
and U19724 (N_19724,N_15661,N_15226);
or U19725 (N_19725,N_17213,N_15078);
xnor U19726 (N_19726,N_16677,N_15859);
nor U19727 (N_19727,N_16941,N_16555);
or U19728 (N_19728,N_15693,N_17446);
nand U19729 (N_19729,N_16483,N_15641);
nand U19730 (N_19730,N_15008,N_15139);
nor U19731 (N_19731,N_17496,N_16387);
nand U19732 (N_19732,N_15079,N_16006);
nand U19733 (N_19733,N_15308,N_15361);
nand U19734 (N_19734,N_16299,N_16263);
and U19735 (N_19735,N_16092,N_16064);
nand U19736 (N_19736,N_15605,N_15480);
xor U19737 (N_19737,N_15966,N_15126);
nor U19738 (N_19738,N_15797,N_16917);
or U19739 (N_19739,N_15141,N_15136);
nor U19740 (N_19740,N_15917,N_16322);
or U19741 (N_19741,N_15620,N_17380);
nor U19742 (N_19742,N_16739,N_16950);
nand U19743 (N_19743,N_16338,N_16644);
or U19744 (N_19744,N_17007,N_16654);
nand U19745 (N_19745,N_15148,N_15161);
and U19746 (N_19746,N_17228,N_16196);
nand U19747 (N_19747,N_17447,N_16960);
and U19748 (N_19748,N_15607,N_17424);
xnor U19749 (N_19749,N_17130,N_17233);
nand U19750 (N_19750,N_15340,N_16669);
xor U19751 (N_19751,N_16664,N_16113);
or U19752 (N_19752,N_17338,N_15304);
nand U19753 (N_19753,N_16145,N_17237);
or U19754 (N_19754,N_16504,N_15149);
or U19755 (N_19755,N_16303,N_15373);
nor U19756 (N_19756,N_17348,N_15620);
xor U19757 (N_19757,N_15638,N_15122);
nor U19758 (N_19758,N_16966,N_17454);
xnor U19759 (N_19759,N_15738,N_15788);
or U19760 (N_19760,N_15890,N_16581);
nor U19761 (N_19761,N_16019,N_17012);
and U19762 (N_19762,N_15610,N_16944);
nor U19763 (N_19763,N_15391,N_16868);
nor U19764 (N_19764,N_15000,N_16184);
nor U19765 (N_19765,N_15811,N_16364);
nand U19766 (N_19766,N_17448,N_16034);
nor U19767 (N_19767,N_17368,N_17179);
xnor U19768 (N_19768,N_16591,N_16041);
or U19769 (N_19769,N_17145,N_16955);
nor U19770 (N_19770,N_16518,N_15274);
xor U19771 (N_19771,N_16031,N_17041);
nor U19772 (N_19772,N_17086,N_15198);
xor U19773 (N_19773,N_16740,N_16348);
nor U19774 (N_19774,N_16975,N_16526);
nor U19775 (N_19775,N_16841,N_15308);
or U19776 (N_19776,N_17173,N_15598);
nor U19777 (N_19777,N_17345,N_17232);
or U19778 (N_19778,N_15872,N_15237);
nand U19779 (N_19779,N_16946,N_15472);
and U19780 (N_19780,N_17106,N_16397);
and U19781 (N_19781,N_16316,N_15611);
or U19782 (N_19782,N_16547,N_15897);
xnor U19783 (N_19783,N_15584,N_15395);
nand U19784 (N_19784,N_17241,N_15941);
or U19785 (N_19785,N_17444,N_15564);
and U19786 (N_19786,N_15937,N_16879);
or U19787 (N_19787,N_16543,N_17057);
nor U19788 (N_19788,N_15289,N_17145);
nand U19789 (N_19789,N_15908,N_15815);
and U19790 (N_19790,N_16907,N_17214);
xnor U19791 (N_19791,N_15016,N_16026);
and U19792 (N_19792,N_16740,N_17408);
nand U19793 (N_19793,N_15717,N_15222);
nor U19794 (N_19794,N_16487,N_15427);
xnor U19795 (N_19795,N_17133,N_16721);
nand U19796 (N_19796,N_17051,N_15662);
and U19797 (N_19797,N_15719,N_16835);
or U19798 (N_19798,N_16578,N_15988);
nor U19799 (N_19799,N_15435,N_15378);
xnor U19800 (N_19800,N_17327,N_16928);
or U19801 (N_19801,N_15295,N_15688);
xor U19802 (N_19802,N_16749,N_15506);
nor U19803 (N_19803,N_17347,N_15030);
and U19804 (N_19804,N_16170,N_16676);
and U19805 (N_19805,N_16147,N_15192);
and U19806 (N_19806,N_15972,N_15975);
and U19807 (N_19807,N_17290,N_15838);
or U19808 (N_19808,N_15198,N_15389);
nor U19809 (N_19809,N_16232,N_16955);
nand U19810 (N_19810,N_15334,N_17225);
nand U19811 (N_19811,N_16119,N_16556);
xnor U19812 (N_19812,N_15504,N_15169);
or U19813 (N_19813,N_16214,N_15048);
nand U19814 (N_19814,N_15627,N_16241);
xnor U19815 (N_19815,N_16705,N_15527);
xnor U19816 (N_19816,N_16665,N_15255);
nand U19817 (N_19817,N_16957,N_15016);
nor U19818 (N_19818,N_15805,N_15743);
nand U19819 (N_19819,N_15529,N_15292);
nand U19820 (N_19820,N_16680,N_17443);
nand U19821 (N_19821,N_15039,N_17148);
or U19822 (N_19822,N_17438,N_15483);
nand U19823 (N_19823,N_16029,N_16936);
or U19824 (N_19824,N_15268,N_16894);
nand U19825 (N_19825,N_17160,N_17222);
and U19826 (N_19826,N_16584,N_16955);
or U19827 (N_19827,N_16556,N_17345);
or U19828 (N_19828,N_15238,N_15683);
nand U19829 (N_19829,N_15959,N_16400);
nor U19830 (N_19830,N_16328,N_15548);
nor U19831 (N_19831,N_17111,N_17394);
and U19832 (N_19832,N_16164,N_15960);
nor U19833 (N_19833,N_17255,N_16689);
and U19834 (N_19834,N_15997,N_15208);
and U19835 (N_19835,N_17018,N_15694);
and U19836 (N_19836,N_15648,N_17301);
and U19837 (N_19837,N_15999,N_16306);
and U19838 (N_19838,N_15532,N_15127);
xnor U19839 (N_19839,N_15174,N_16722);
nand U19840 (N_19840,N_16157,N_17095);
nand U19841 (N_19841,N_17291,N_16097);
nor U19842 (N_19842,N_15314,N_17236);
or U19843 (N_19843,N_15692,N_16507);
and U19844 (N_19844,N_15480,N_16842);
or U19845 (N_19845,N_15879,N_15130);
xnor U19846 (N_19846,N_17302,N_15128);
nor U19847 (N_19847,N_15489,N_17413);
xnor U19848 (N_19848,N_15614,N_15248);
nand U19849 (N_19849,N_16070,N_15279);
and U19850 (N_19850,N_16202,N_17071);
and U19851 (N_19851,N_15514,N_15964);
nor U19852 (N_19852,N_16864,N_17362);
nand U19853 (N_19853,N_16812,N_16942);
or U19854 (N_19854,N_17013,N_15246);
xor U19855 (N_19855,N_16930,N_16549);
nor U19856 (N_19856,N_16192,N_16900);
xnor U19857 (N_19857,N_15847,N_17196);
nor U19858 (N_19858,N_15292,N_17127);
or U19859 (N_19859,N_15059,N_16439);
or U19860 (N_19860,N_15473,N_16332);
nor U19861 (N_19861,N_15883,N_15843);
and U19862 (N_19862,N_16002,N_17085);
xor U19863 (N_19863,N_15662,N_16674);
xnor U19864 (N_19864,N_16287,N_15951);
nor U19865 (N_19865,N_16226,N_15558);
and U19866 (N_19866,N_15934,N_16381);
xor U19867 (N_19867,N_16598,N_15993);
nand U19868 (N_19868,N_16518,N_16644);
and U19869 (N_19869,N_16584,N_17282);
xor U19870 (N_19870,N_16811,N_15075);
nor U19871 (N_19871,N_15527,N_15602);
or U19872 (N_19872,N_16540,N_15195);
xor U19873 (N_19873,N_16225,N_17303);
nor U19874 (N_19874,N_17115,N_16818);
nor U19875 (N_19875,N_15873,N_15142);
xor U19876 (N_19876,N_16592,N_16892);
nor U19877 (N_19877,N_15113,N_15713);
and U19878 (N_19878,N_15371,N_16314);
and U19879 (N_19879,N_16353,N_17096);
nand U19880 (N_19880,N_16433,N_16765);
nand U19881 (N_19881,N_16572,N_15115);
nand U19882 (N_19882,N_16972,N_15653);
or U19883 (N_19883,N_17227,N_16803);
nand U19884 (N_19884,N_15582,N_17141);
or U19885 (N_19885,N_17189,N_17239);
nand U19886 (N_19886,N_15756,N_16626);
nand U19887 (N_19887,N_17441,N_17149);
nand U19888 (N_19888,N_15516,N_17490);
nor U19889 (N_19889,N_16721,N_16691);
or U19890 (N_19890,N_17296,N_17423);
or U19891 (N_19891,N_15010,N_17168);
nor U19892 (N_19892,N_17158,N_15973);
and U19893 (N_19893,N_16604,N_15419);
nand U19894 (N_19894,N_17323,N_15474);
nand U19895 (N_19895,N_16442,N_16994);
or U19896 (N_19896,N_15011,N_16317);
nand U19897 (N_19897,N_17486,N_16737);
or U19898 (N_19898,N_15441,N_15435);
nand U19899 (N_19899,N_15362,N_15340);
and U19900 (N_19900,N_17077,N_16070);
xor U19901 (N_19901,N_15968,N_15331);
nor U19902 (N_19902,N_16379,N_16657);
or U19903 (N_19903,N_16656,N_17436);
xor U19904 (N_19904,N_15077,N_15251);
nor U19905 (N_19905,N_15356,N_17214);
xor U19906 (N_19906,N_15528,N_16349);
or U19907 (N_19907,N_17034,N_16945);
nor U19908 (N_19908,N_16748,N_16001);
xnor U19909 (N_19909,N_16636,N_15455);
and U19910 (N_19910,N_16348,N_17000);
or U19911 (N_19911,N_16660,N_16155);
xnor U19912 (N_19912,N_15436,N_16340);
and U19913 (N_19913,N_17334,N_16201);
nand U19914 (N_19914,N_17355,N_17078);
or U19915 (N_19915,N_16848,N_15361);
and U19916 (N_19916,N_17242,N_17105);
or U19917 (N_19917,N_16658,N_16374);
nand U19918 (N_19918,N_17305,N_17074);
or U19919 (N_19919,N_15112,N_16983);
nand U19920 (N_19920,N_16477,N_17008);
nand U19921 (N_19921,N_17028,N_15183);
nor U19922 (N_19922,N_16268,N_15069);
and U19923 (N_19923,N_15677,N_16932);
or U19924 (N_19924,N_15751,N_15185);
and U19925 (N_19925,N_15647,N_16163);
or U19926 (N_19926,N_15035,N_15860);
or U19927 (N_19927,N_16022,N_15780);
or U19928 (N_19928,N_17468,N_15998);
xor U19929 (N_19929,N_15524,N_16183);
or U19930 (N_19930,N_15340,N_17128);
or U19931 (N_19931,N_17244,N_15573);
nor U19932 (N_19932,N_16761,N_15920);
or U19933 (N_19933,N_17140,N_17099);
and U19934 (N_19934,N_16249,N_15952);
or U19935 (N_19935,N_16840,N_16849);
nand U19936 (N_19936,N_16641,N_15686);
nand U19937 (N_19937,N_17213,N_16379);
or U19938 (N_19938,N_15503,N_16777);
nand U19939 (N_19939,N_15248,N_15467);
nor U19940 (N_19940,N_15996,N_15144);
xnor U19941 (N_19941,N_16357,N_15852);
and U19942 (N_19942,N_16388,N_15640);
xor U19943 (N_19943,N_17092,N_16574);
or U19944 (N_19944,N_15874,N_16198);
and U19945 (N_19945,N_16232,N_16330);
or U19946 (N_19946,N_15834,N_15557);
xnor U19947 (N_19947,N_16347,N_17179);
nand U19948 (N_19948,N_16401,N_16229);
and U19949 (N_19949,N_16418,N_16186);
nand U19950 (N_19950,N_16107,N_15919);
nor U19951 (N_19951,N_15148,N_16130);
xor U19952 (N_19952,N_16867,N_15970);
nor U19953 (N_19953,N_17279,N_17253);
nor U19954 (N_19954,N_15995,N_17300);
nor U19955 (N_19955,N_16964,N_15071);
nand U19956 (N_19956,N_17474,N_15383);
and U19957 (N_19957,N_15008,N_15404);
and U19958 (N_19958,N_17319,N_16354);
and U19959 (N_19959,N_15563,N_16152);
or U19960 (N_19960,N_17281,N_15555);
and U19961 (N_19961,N_17182,N_15150);
or U19962 (N_19962,N_15463,N_16747);
or U19963 (N_19963,N_16953,N_16058);
or U19964 (N_19964,N_16791,N_16981);
and U19965 (N_19965,N_16661,N_16227);
or U19966 (N_19966,N_16416,N_16555);
and U19967 (N_19967,N_16992,N_16272);
nor U19968 (N_19968,N_17058,N_16630);
nand U19969 (N_19969,N_16388,N_17085);
xor U19970 (N_19970,N_17249,N_16948);
and U19971 (N_19971,N_17153,N_15425);
and U19972 (N_19972,N_16121,N_17024);
or U19973 (N_19973,N_17341,N_16071);
xor U19974 (N_19974,N_16710,N_17157);
or U19975 (N_19975,N_15776,N_16236);
nor U19976 (N_19976,N_15811,N_15781);
nand U19977 (N_19977,N_16816,N_15207);
nor U19978 (N_19978,N_17043,N_17402);
nor U19979 (N_19979,N_16336,N_17372);
nor U19980 (N_19980,N_16558,N_16877);
nor U19981 (N_19981,N_17337,N_15334);
nor U19982 (N_19982,N_15045,N_15831);
and U19983 (N_19983,N_17273,N_15182);
xor U19984 (N_19984,N_17005,N_16567);
or U19985 (N_19985,N_16010,N_16080);
and U19986 (N_19986,N_15038,N_16034);
or U19987 (N_19987,N_15487,N_15697);
and U19988 (N_19988,N_17492,N_15386);
nor U19989 (N_19989,N_17266,N_16147);
nand U19990 (N_19990,N_16641,N_17227);
nand U19991 (N_19991,N_16978,N_15182);
or U19992 (N_19992,N_15020,N_17138);
nand U19993 (N_19993,N_15856,N_15599);
or U19994 (N_19994,N_15562,N_15215);
xnor U19995 (N_19995,N_16544,N_15251);
nand U19996 (N_19996,N_17190,N_16034);
or U19997 (N_19997,N_15037,N_16579);
nor U19998 (N_19998,N_15203,N_17141);
or U19999 (N_19999,N_16457,N_17435);
or U20000 (N_20000,N_18365,N_18256);
or U20001 (N_20001,N_19109,N_17807);
xnor U20002 (N_20002,N_17681,N_17861);
nor U20003 (N_20003,N_19447,N_19485);
and U20004 (N_20004,N_17565,N_19985);
nor U20005 (N_20005,N_18509,N_18890);
nor U20006 (N_20006,N_18571,N_18054);
xnor U20007 (N_20007,N_18168,N_18134);
and U20008 (N_20008,N_19092,N_18645);
nor U20009 (N_20009,N_19004,N_18133);
xor U20010 (N_20010,N_19384,N_17976);
and U20011 (N_20011,N_19978,N_19334);
or U20012 (N_20012,N_19193,N_18640);
nor U20013 (N_20013,N_19101,N_19127);
nand U20014 (N_20014,N_18292,N_17599);
nor U20015 (N_20015,N_19573,N_19096);
and U20016 (N_20016,N_18630,N_19887);
xor U20017 (N_20017,N_19215,N_17970);
or U20018 (N_20018,N_18723,N_19824);
and U20019 (N_20019,N_19584,N_19613);
nand U20020 (N_20020,N_19874,N_18677);
nor U20021 (N_20021,N_19498,N_19748);
nor U20022 (N_20022,N_19247,N_19585);
xor U20023 (N_20023,N_18759,N_19347);
nor U20024 (N_20024,N_18880,N_18388);
or U20025 (N_20025,N_19944,N_17820);
xor U20026 (N_20026,N_17783,N_18730);
xor U20027 (N_20027,N_18982,N_17730);
or U20028 (N_20028,N_19697,N_19021);
and U20029 (N_20029,N_17602,N_18592);
xor U20030 (N_20030,N_19465,N_19449);
nor U20031 (N_20031,N_19346,N_19624);
and U20032 (N_20032,N_19828,N_19512);
or U20033 (N_20033,N_17985,N_19185);
or U20034 (N_20034,N_19150,N_19927);
xnor U20035 (N_20035,N_19020,N_19408);
and U20036 (N_20036,N_18091,N_18065);
nor U20037 (N_20037,N_19280,N_19983);
nor U20038 (N_20038,N_18310,N_17764);
or U20039 (N_20039,N_18455,N_18503);
nand U20040 (N_20040,N_18359,N_17962);
nand U20041 (N_20041,N_17611,N_19474);
nand U20042 (N_20042,N_19800,N_18439);
and U20043 (N_20043,N_18076,N_19926);
xnor U20044 (N_20044,N_18385,N_19745);
xor U20045 (N_20045,N_17541,N_18375);
or U20046 (N_20046,N_18196,N_19501);
nor U20047 (N_20047,N_19161,N_19626);
xor U20048 (N_20048,N_19296,N_18353);
xor U20049 (N_20049,N_18719,N_18979);
or U20050 (N_20050,N_19289,N_18458);
nand U20051 (N_20051,N_19272,N_19151);
nor U20052 (N_20052,N_18729,N_18824);
nor U20053 (N_20053,N_19012,N_18098);
nand U20054 (N_20054,N_19237,N_17750);
nand U20055 (N_20055,N_19362,N_18915);
nand U20056 (N_20056,N_19736,N_17514);
and U20057 (N_20057,N_18403,N_19484);
and U20058 (N_20058,N_19596,N_19071);
nor U20059 (N_20059,N_17589,N_19231);
xor U20060 (N_20060,N_18247,N_18610);
nor U20061 (N_20061,N_18790,N_19300);
or U20062 (N_20062,N_19470,N_18056);
and U20063 (N_20063,N_18984,N_17718);
nor U20064 (N_20064,N_18620,N_19067);
nand U20065 (N_20065,N_18823,N_19803);
or U20066 (N_20066,N_18899,N_18290);
nor U20067 (N_20067,N_18794,N_18102);
and U20068 (N_20068,N_19661,N_19743);
nor U20069 (N_20069,N_17708,N_18024);
nand U20070 (N_20070,N_17935,N_19212);
nor U20071 (N_20071,N_18844,N_18502);
or U20072 (N_20072,N_19271,N_18976);
nor U20073 (N_20073,N_18431,N_18371);
xnor U20074 (N_20074,N_19541,N_17663);
nand U20075 (N_20075,N_17926,N_17548);
and U20076 (N_20076,N_18528,N_18298);
xnor U20077 (N_20077,N_19112,N_19250);
xnor U20078 (N_20078,N_19899,N_18514);
and U20079 (N_20079,N_18676,N_17886);
and U20080 (N_20080,N_18483,N_19788);
xnor U20081 (N_20081,N_19201,N_17812);
or U20082 (N_20082,N_19122,N_17907);
or U20083 (N_20083,N_18021,N_17826);
xor U20084 (N_20084,N_19062,N_17527);
or U20085 (N_20085,N_18272,N_18917);
or U20086 (N_20086,N_19494,N_17638);
nor U20087 (N_20087,N_19049,N_18243);
xor U20088 (N_20088,N_18861,N_18116);
xnor U20089 (N_20089,N_18025,N_18320);
nand U20090 (N_20090,N_17978,N_19763);
nor U20091 (N_20091,N_18323,N_17662);
and U20092 (N_20092,N_17659,N_18888);
nor U20093 (N_20093,N_18387,N_19889);
or U20094 (N_20094,N_18548,N_19960);
nor U20095 (N_20095,N_19908,N_19931);
nand U20096 (N_20096,N_17518,N_17752);
or U20097 (N_20097,N_19973,N_19235);
or U20098 (N_20098,N_19715,N_17869);
xor U20099 (N_20099,N_19380,N_18672);
nor U20100 (N_20100,N_17661,N_18713);
xnor U20101 (N_20101,N_18921,N_19050);
nand U20102 (N_20102,N_18002,N_18209);
nand U20103 (N_20103,N_19790,N_18588);
nor U20104 (N_20104,N_17914,N_19665);
nor U20105 (N_20105,N_17794,N_18760);
nor U20106 (N_20106,N_18094,N_17846);
nor U20107 (N_20107,N_18027,N_17637);
nor U20108 (N_20108,N_19907,N_18328);
xor U20109 (N_20109,N_18873,N_18662);
xor U20110 (N_20110,N_18705,N_17797);
nor U20111 (N_20111,N_17606,N_19947);
or U20112 (N_20112,N_17557,N_19292);
xnor U20113 (N_20113,N_18579,N_18496);
and U20114 (N_20114,N_19495,N_18546);
xor U20115 (N_20115,N_18977,N_18161);
or U20116 (N_20116,N_18832,N_17691);
nand U20117 (N_20117,N_19844,N_17529);
nor U20118 (N_20118,N_19104,N_18657);
or U20119 (N_20119,N_19725,N_19354);
nand U20120 (N_20120,N_18518,N_19328);
or U20121 (N_20121,N_19367,N_19262);
nand U20122 (N_20122,N_18220,N_18433);
xnor U20123 (N_20123,N_17946,N_19135);
nor U20124 (N_20124,N_19809,N_19701);
or U20125 (N_20125,N_18810,N_17617);
xor U20126 (N_20126,N_18520,N_18034);
or U20127 (N_20127,N_19849,N_17871);
nor U20128 (N_20128,N_18124,N_18679);
and U20129 (N_20129,N_18975,N_19586);
or U20130 (N_20130,N_19473,N_19276);
and U20131 (N_20131,N_19270,N_18476);
or U20132 (N_20132,N_18249,N_17645);
nor U20133 (N_20133,N_19464,N_18831);
and U20134 (N_20134,N_17819,N_19941);
xnor U20135 (N_20135,N_17977,N_19209);
xor U20136 (N_20136,N_19079,N_19623);
xor U20137 (N_20137,N_17688,N_18892);
xor U20138 (N_20138,N_19674,N_18229);
xor U20139 (N_20139,N_18391,N_17535);
and U20140 (N_20140,N_19784,N_18750);
nor U20141 (N_20141,N_18270,N_18636);
or U20142 (N_20142,N_17593,N_18318);
or U20143 (N_20143,N_17753,N_18495);
and U20144 (N_20144,N_18752,N_17536);
nand U20145 (N_20145,N_19398,N_18346);
or U20146 (N_20146,N_17702,N_18408);
nor U20147 (N_20147,N_19649,N_19432);
nor U20148 (N_20148,N_18327,N_18966);
and U20149 (N_20149,N_18113,N_18908);
xnor U20150 (N_20150,N_19675,N_18747);
or U20151 (N_20151,N_19144,N_18036);
nand U20152 (N_20152,N_18783,N_18374);
nand U20153 (N_20153,N_18464,N_19469);
or U20154 (N_20154,N_18281,N_19366);
and U20155 (N_20155,N_19006,N_19597);
xor U20156 (N_20156,N_18813,N_17858);
nor U20157 (N_20157,N_18505,N_17626);
xnor U20158 (N_20158,N_18972,N_18178);
and U20159 (N_20159,N_19571,N_18597);
xnor U20160 (N_20160,N_19815,N_17740);
nor U20161 (N_20161,N_17903,N_19344);
or U20162 (N_20162,N_19162,N_19595);
or U20163 (N_20163,N_18405,N_19190);
nand U20164 (N_20164,N_19910,N_17845);
xnor U20165 (N_20165,N_19836,N_18781);
nor U20166 (N_20166,N_17988,N_18448);
and U20167 (N_20167,N_18923,N_18423);
xnor U20168 (N_20168,N_17705,N_18289);
and U20169 (N_20169,N_19037,N_19919);
xor U20170 (N_20170,N_18066,N_17574);
and U20171 (N_20171,N_18087,N_18266);
xor U20172 (N_20172,N_19379,N_19695);
nor U20173 (N_20173,N_19940,N_18830);
or U20174 (N_20174,N_19489,N_18782);
nand U20175 (N_20175,N_18119,N_18086);
or U20176 (N_20176,N_17749,N_19967);
and U20177 (N_20177,N_19094,N_19313);
xnor U20178 (N_20178,N_19901,N_17631);
and U20179 (N_20179,N_18635,N_18363);
and U20180 (N_20180,N_18842,N_19738);
and U20181 (N_20181,N_18803,N_17580);
or U20182 (N_20182,N_19574,N_18085);
or U20183 (N_20183,N_18165,N_18399);
nand U20184 (N_20184,N_19604,N_17891);
nand U20185 (N_20185,N_18093,N_18775);
or U20186 (N_20186,N_19991,N_18356);
or U20187 (N_20187,N_17568,N_18659);
or U20188 (N_20188,N_18061,N_17668);
xnor U20189 (N_20189,N_17774,N_18724);
xnor U20190 (N_20190,N_18334,N_18572);
or U20191 (N_20191,N_18602,N_18500);
xnor U20192 (N_20192,N_18965,N_18732);
xnor U20193 (N_20193,N_19838,N_18501);
and U20194 (N_20194,N_18567,N_18083);
or U20195 (N_20195,N_17605,N_17919);
nor U20196 (N_20196,N_19284,N_18988);
and U20197 (N_20197,N_19582,N_18802);
nand U20198 (N_20198,N_17870,N_17844);
xor U20199 (N_20199,N_18115,N_19389);
xor U20200 (N_20200,N_19396,N_19837);
nand U20201 (N_20201,N_19822,N_19418);
and U20202 (N_20202,N_19205,N_18598);
xor U20203 (N_20203,N_18302,N_19923);
xor U20204 (N_20204,N_18473,N_17513);
xnor U20205 (N_20205,N_18584,N_19554);
nand U20206 (N_20206,N_18383,N_19723);
and U20207 (N_20207,N_19047,N_18358);
nand U20208 (N_20208,N_18507,N_18955);
xor U20209 (N_20209,N_19275,N_19671);
and U20210 (N_20210,N_19444,N_19427);
and U20211 (N_20211,N_18032,N_18916);
xnor U20212 (N_20212,N_18770,N_19456);
or U20213 (N_20213,N_17725,N_19939);
or U20214 (N_20214,N_19064,N_17887);
and U20215 (N_20215,N_19206,N_17581);
nand U20216 (N_20216,N_18226,N_18935);
xor U20217 (N_20217,N_18845,N_18421);
or U20218 (N_20218,N_18671,N_18943);
or U20219 (N_20219,N_19035,N_18394);
or U20220 (N_20220,N_18190,N_17639);
and U20221 (N_20221,N_19873,N_18513);
and U20222 (N_20222,N_18118,N_19841);
and U20223 (N_20223,N_19664,N_18714);
xnor U20224 (N_20224,N_18217,N_17939);
and U20225 (N_20225,N_19070,N_19607);
and U20226 (N_20226,N_17649,N_17893);
or U20227 (N_20227,N_18666,N_19142);
or U20228 (N_20228,N_19424,N_19269);
or U20229 (N_20229,N_18044,N_19188);
nor U20230 (N_20230,N_19816,N_17963);
nor U20231 (N_20231,N_19945,N_19369);
xnor U20232 (N_20232,N_19785,N_19986);
xor U20233 (N_20233,N_19957,N_17524);
xnor U20234 (N_20234,N_19351,N_18583);
nor U20235 (N_20235,N_17851,N_18905);
and U20236 (N_20236,N_18453,N_19093);
and U20237 (N_20237,N_18774,N_18527);
xnor U20238 (N_20238,N_17614,N_17900);
or U20239 (N_20239,N_17704,N_18199);
or U20240 (N_20240,N_19783,N_17890);
or U20241 (N_20241,N_18684,N_19042);
xnor U20242 (N_20242,N_19297,N_19400);
xor U20243 (N_20243,N_17627,N_19542);
or U20244 (N_20244,N_19528,N_17863);
xnor U20245 (N_20245,N_18858,N_19360);
xor U20246 (N_20246,N_17501,N_19214);
or U20247 (N_20247,N_19324,N_18967);
nand U20248 (N_20248,N_18817,N_18751);
and U20249 (N_20249,N_19529,N_19365);
xnor U20250 (N_20250,N_18038,N_19103);
nand U20251 (N_20251,N_19544,N_18735);
nor U20252 (N_20252,N_17947,N_18710);
nor U20253 (N_20253,N_18681,N_17759);
nor U20254 (N_20254,N_18784,N_17735);
and U20255 (N_20255,N_18067,N_18838);
xor U20256 (N_20256,N_19443,N_19057);
nand U20257 (N_20257,N_17966,N_19204);
nand U20258 (N_20258,N_19515,N_17839);
or U20259 (N_20259,N_18361,N_19606);
nor U20260 (N_20260,N_19306,N_18516);
or U20261 (N_20261,N_17687,N_18039);
xnor U20262 (N_20262,N_18929,N_19490);
nor U20263 (N_20263,N_19123,N_18996);
nor U20264 (N_20264,N_19618,N_19920);
and U20265 (N_20265,N_19130,N_18764);
nand U20266 (N_20266,N_17621,N_18139);
xnor U20267 (N_20267,N_17507,N_18575);
xor U20268 (N_20268,N_19031,N_18234);
nor U20269 (N_20269,N_19390,N_19787);
and U20270 (N_20270,N_19199,N_19587);
nand U20271 (N_20271,N_19955,N_19508);
nand U20272 (N_20272,N_19349,N_17902);
nor U20273 (N_20273,N_18733,N_19716);
nand U20274 (N_20274,N_18853,N_18815);
or U20275 (N_20275,N_18211,N_17762);
nor U20276 (N_20276,N_19871,N_17642);
xor U20277 (N_20277,N_19662,N_19976);
xnor U20278 (N_20278,N_17833,N_19381);
or U20279 (N_20279,N_19029,N_18779);
xnor U20280 (N_20280,N_17953,N_18690);
xnor U20281 (N_20281,N_19909,N_19108);
and U20282 (N_20282,N_19930,N_19722);
xor U20283 (N_20283,N_18763,N_19705);
xor U20284 (N_20284,N_19090,N_19720);
nand U20285 (N_20285,N_19011,N_19264);
xnor U20286 (N_20286,N_19823,N_17697);
nand U20287 (N_20287,N_17531,N_19255);
nor U20288 (N_20288,N_19463,N_18885);
nor U20289 (N_20289,N_19061,N_18325);
xnor U20290 (N_20290,N_18801,N_19224);
xor U20291 (N_20291,N_19014,N_18904);
and U20292 (N_20292,N_18664,N_18321);
and U20293 (N_20293,N_19412,N_18898);
or U20294 (N_20294,N_19861,N_18278);
and U20295 (N_20295,N_17784,N_18212);
xnor U20296 (N_20296,N_19640,N_19886);
xor U20297 (N_20297,N_19737,N_19752);
or U20298 (N_20298,N_18656,N_19038);
or U20299 (N_20299,N_19538,N_19942);
and U20300 (N_20300,N_18000,N_18541);
xnor U20301 (N_20301,N_18601,N_19892);
xnor U20302 (N_20302,N_19533,N_19343);
and U20303 (N_20303,N_19796,N_17873);
or U20304 (N_20304,N_18128,N_17545);
nor U20305 (N_20305,N_17622,N_18538);
or U20306 (N_20306,N_18275,N_19537);
nor U20307 (N_20307,N_17944,N_19726);
nor U20308 (N_20308,N_18887,N_17525);
and U20309 (N_20309,N_18668,N_18953);
xnor U20310 (N_20310,N_17629,N_18562);
xnor U20311 (N_20311,N_18412,N_17558);
nor U20312 (N_20312,N_18990,N_18218);
or U20313 (N_20313,N_18169,N_17633);
or U20314 (N_20314,N_19027,N_18262);
nor U20315 (N_20315,N_18046,N_17619);
nor U20316 (N_20316,N_18581,N_18855);
and U20317 (N_20317,N_19073,N_19797);
or U20318 (N_20318,N_18075,N_18092);
xnor U20319 (N_20319,N_19691,N_19876);
nor U20320 (N_20320,N_19018,N_19277);
or U20321 (N_20321,N_18633,N_19700);
and U20322 (N_20322,N_17930,N_18340);
xor U20323 (N_20323,N_19374,N_18867);
and U20324 (N_20324,N_19416,N_18060);
nor U20325 (N_20325,N_18693,N_19307);
nand U20326 (N_20326,N_18931,N_19592);
or U20327 (N_20327,N_17726,N_17595);
nor U20328 (N_20328,N_17672,N_18089);
and U20329 (N_20329,N_17984,N_18658);
nor U20330 (N_20330,N_19041,N_19023);
or U20331 (N_20331,N_19000,N_18293);
or U20332 (N_20332,N_18132,N_18191);
nand U20333 (N_20333,N_19616,N_18015);
or U20334 (N_20334,N_18629,N_19835);
and U20335 (N_20335,N_18158,N_19091);
nand U20336 (N_20336,N_17651,N_19747);
and U20337 (N_20337,N_18969,N_19866);
xnor U20338 (N_20338,N_17888,N_18879);
nor U20339 (N_20339,N_18902,N_18761);
or U20340 (N_20340,N_18376,N_17745);
nor U20341 (N_20341,N_19245,N_17882);
nand U20342 (N_20342,N_19753,N_18531);
nor U20343 (N_20343,N_19352,N_18700);
xnor U20344 (N_20344,N_18947,N_19656);
xnor U20345 (N_20345,N_18612,N_19966);
nor U20346 (N_20346,N_19546,N_17588);
and U20347 (N_20347,N_19677,N_18740);
nand U20348 (N_20348,N_18985,N_19928);
or U20349 (N_20349,N_18603,N_18703);
or U20350 (N_20350,N_19750,N_17905);
or U20351 (N_20351,N_19197,N_19744);
nand U20352 (N_20352,N_19405,N_18426);
nand U20353 (N_20353,N_18582,N_19786);
nand U20354 (N_20354,N_18755,N_18626);
and U20355 (N_20355,N_19709,N_19184);
nand U20356 (N_20356,N_18793,N_19633);
or U20357 (N_20357,N_17895,N_17610);
or U20358 (N_20358,N_17789,N_19713);
nand U20359 (N_20359,N_19363,N_18995);
or U20360 (N_20360,N_19252,N_19046);
and U20361 (N_20361,N_18295,N_18846);
or U20362 (N_20362,N_19682,N_18787);
and U20363 (N_20363,N_18160,N_19581);
nor U20364 (N_20364,N_19100,N_18674);
nor U20365 (N_20365,N_18205,N_17575);
and U20366 (N_20366,N_18063,N_17554);
xor U20367 (N_20367,N_17742,N_17958);
nand U20368 (N_20368,N_18030,N_17987);
nand U20369 (N_20369,N_19666,N_17813);
xor U20370 (N_20370,N_17578,N_18045);
or U20371 (N_20371,N_19195,N_18026);
nand U20372 (N_20372,N_18607,N_19403);
and U20373 (N_20373,N_18143,N_19323);
xor U20374 (N_20374,N_17562,N_19283);
nand U20375 (N_20375,N_19336,N_17785);
nand U20376 (N_20376,N_19082,N_18324);
xor U20377 (N_20377,N_19234,N_19806);
xnor U20378 (N_20378,N_19840,N_18973);
nand U20379 (N_20379,N_18654,N_17528);
nor U20380 (N_20380,N_18717,N_19478);
nand U20381 (N_20381,N_18042,N_19520);
and U20382 (N_20382,N_19680,N_17802);
and U20383 (N_20383,N_18534,N_17832);
nand U20384 (N_20384,N_17679,N_19793);
xnor U20385 (N_20385,N_17694,N_17921);
or U20386 (N_20386,N_18216,N_19539);
or U20387 (N_20387,N_18699,N_19243);
nor U20388 (N_20388,N_17954,N_19053);
or U20389 (N_20389,N_19111,N_18682);
or U20390 (N_20390,N_17915,N_19414);
or U20391 (N_20391,N_19918,N_18155);
nor U20392 (N_20392,N_19801,N_18484);
xor U20393 (N_20393,N_19285,N_18568);
or U20394 (N_20394,N_19702,N_19022);
nor U20395 (N_20395,N_18930,N_19411);
xor U20396 (N_20396,N_17855,N_17847);
xnor U20397 (N_20397,N_19043,N_18702);
xnor U20398 (N_20398,N_19954,N_19001);
and U20399 (N_20399,N_18315,N_18429);
nand U20400 (N_20400,N_19331,N_19648);
nor U20401 (N_20401,N_19159,N_18849);
or U20402 (N_20402,N_18378,N_19423);
and U20403 (N_20403,N_19036,N_19293);
and U20404 (N_20404,N_18494,N_18377);
nor U20405 (N_20405,N_19105,N_19211);
or U20406 (N_20406,N_18616,N_18778);
nand U20407 (N_20407,N_18914,N_19653);
or U20408 (N_20408,N_17940,N_19827);
and U20409 (N_20409,N_18925,N_19461);
and U20410 (N_20410,N_18559,N_19847);
xor U20411 (N_20411,N_19877,N_18043);
xor U20412 (N_20412,N_18558,N_18456);
or U20413 (N_20413,N_19830,N_19536);
nor U20414 (N_20414,N_18753,N_18422);
nor U20415 (N_20415,N_18069,N_19239);
xnor U20416 (N_20416,N_19173,N_18767);
or U20417 (N_20417,N_17597,N_19359);
nand U20418 (N_20418,N_19905,N_17771);
xnor U20419 (N_20419,N_18937,N_17692);
nand U20420 (N_20420,N_19817,N_19168);
xor U20421 (N_20421,N_18194,N_19076);
and U20422 (N_20422,N_19436,N_19672);
or U20423 (N_20423,N_19413,N_18362);
and U20424 (N_20424,N_19754,N_18077);
nor U20425 (N_20425,N_18569,N_17773);
nor U20426 (N_20426,N_18669,N_18949);
or U20427 (N_20427,N_18712,N_19060);
or U20428 (N_20428,N_19575,N_18286);
nor U20429 (N_20429,N_17751,N_17722);
xor U20430 (N_20430,N_18058,N_19005);
or U20431 (N_20431,N_19263,N_18663);
or U20432 (N_20432,N_17996,N_18847);
and U20433 (N_20433,N_18487,N_18285);
nor U20434 (N_20434,N_18167,N_18406);
xnor U20435 (N_20435,N_19959,N_18192);
nand U20436 (N_20436,N_19274,N_19730);
and U20437 (N_20437,N_19453,N_19467);
nand U20438 (N_20438,N_19812,N_18333);
or U20439 (N_20439,N_19792,N_19932);
xnor U20440 (N_20440,N_19566,N_19459);
nand U20441 (N_20441,N_19769,N_18020);
nor U20442 (N_20442,N_19415,N_18430);
nand U20443 (N_20443,N_18573,N_19721);
and U20444 (N_20444,N_19632,N_19862);
nand U20445 (N_20445,N_19688,N_17505);
nor U20446 (N_20446,N_19951,N_19580);
and U20447 (N_20447,N_18418,N_19439);
xnor U20448 (N_20448,N_17721,N_19593);
and U20449 (N_20449,N_18314,N_18150);
nor U20450 (N_20450,N_19392,N_19570);
nor U20451 (N_20451,N_19179,N_17618);
nor U20452 (N_20452,N_19825,N_19768);
and U20453 (N_20453,N_18267,N_18644);
or U20454 (N_20454,N_18263,N_18329);
or U20455 (N_20455,N_17965,N_17714);
and U20456 (N_20456,N_18010,N_19371);
nand U20457 (N_20457,N_19420,N_19232);
or U20458 (N_20458,N_18499,N_18401);
and U20459 (N_20459,N_19388,N_17768);
nor U20460 (N_20460,N_19821,N_19226);
and U20461 (N_20461,N_18586,N_19492);
xnor U20462 (N_20462,N_19914,N_18820);
nand U20463 (N_20463,N_18909,N_17728);
xor U20464 (N_20464,N_19098,N_19856);
and U20465 (N_20465,N_19791,N_19106);
and U20466 (N_20466,N_18860,N_19475);
xor U20467 (N_20467,N_19971,N_17916);
nor U20468 (N_20468,N_18806,N_18313);
and U20469 (N_20469,N_19394,N_17711);
or U20470 (N_20470,N_19891,N_19683);
and U20471 (N_20471,N_17526,N_19650);
xor U20472 (N_20472,N_18563,N_19798);
nand U20473 (N_20473,N_18303,N_18198);
or U20474 (N_20474,N_18550,N_18184);
nor U20475 (N_20475,N_19335,N_18952);
nand U20476 (N_20476,N_18008,N_19807);
or U20477 (N_20477,N_18291,N_17678);
or U20478 (N_20478,N_18479,N_19045);
nand U20479 (N_20479,N_19658,N_18454);
xor U20480 (N_20480,N_18622,N_18153);
or U20481 (N_20481,N_19503,N_18738);
nor U20482 (N_20482,N_18366,N_18736);
or U20483 (N_20483,N_19916,N_17511);
nand U20484 (N_20484,N_19767,N_19222);
xor U20485 (N_20485,N_19227,N_17701);
nor U20486 (N_20486,N_19998,N_19969);
xnor U20487 (N_20487,N_17555,N_19353);
or U20488 (N_20488,N_19997,N_19114);
nor U20489 (N_20489,N_17624,N_17650);
nand U20490 (N_20490,N_19514,N_18555);
xnor U20491 (N_20491,N_18591,N_18523);
and U20492 (N_20492,N_18337,N_19339);
xnor U20493 (N_20493,N_17543,N_18900);
nand U20494 (N_20494,N_18731,N_18825);
or U20495 (N_20495,N_19545,N_18031);
nor U20496 (N_20496,N_17937,N_18543);
or U20497 (N_20497,N_18389,N_18163);
nand U20498 (N_20498,N_18342,N_19448);
or U20499 (N_20499,N_18590,N_17594);
xnor U20500 (N_20500,N_19729,N_19875);
xnor U20501 (N_20501,N_18308,N_18339);
and U20502 (N_20502,N_18344,N_18331);
xor U20503 (N_20503,N_19898,N_18593);
xnor U20504 (N_20504,N_19724,N_17959);
and U20505 (N_20505,N_18227,N_17550);
nor U20506 (N_20506,N_17816,N_17778);
and U20507 (N_20507,N_19808,N_18741);
nand U20508 (N_20508,N_19513,N_18386);
and U20509 (N_20509,N_18224,N_17696);
and U20510 (N_20510,N_18874,N_18404);
xnor U20511 (N_20511,N_19175,N_19140);
xor U20512 (N_20512,N_17998,N_19938);
nor U20513 (N_20513,N_17883,N_19718);
or U20514 (N_20514,N_19719,N_18517);
xnor U20515 (N_20515,N_17537,N_19314);
and U20516 (N_20516,N_18457,N_18012);
xnor U20517 (N_20517,N_18106,N_18193);
nor U20518 (N_20518,N_18718,N_19869);
nor U20519 (N_20519,N_17885,N_19177);
nand U20520 (N_20520,N_17840,N_17500);
and U20521 (N_20521,N_19572,N_18539);
nor U20522 (N_20522,N_17941,N_19975);
nand U20523 (N_20523,N_17655,N_18745);
and U20524 (N_20524,N_19192,N_17837);
nor U20525 (N_20525,N_18754,N_19348);
nand U20526 (N_20526,N_18114,N_18987);
or U20527 (N_20527,N_19483,N_18230);
and U20528 (N_20528,N_17549,N_19794);
or U20529 (N_20529,N_18246,N_18241);
and U20530 (N_20530,N_19259,N_18960);
nor U20531 (N_20531,N_19107,N_18283);
nand U20532 (N_20532,N_17931,N_17918);
or U20533 (N_20533,N_18631,N_19281);
xnor U20534 (N_20534,N_18452,N_17635);
or U20535 (N_20535,N_18251,N_19131);
and U20536 (N_20536,N_18839,N_18660);
and U20537 (N_20537,N_17779,N_18814);
nand U20538 (N_20538,N_19660,N_19854);
xnor U20539 (N_20539,N_19727,N_18604);
nand U20540 (N_20540,N_19804,N_18400);
or U20541 (N_20541,N_18609,N_18138);
or U20542 (N_20542,N_17652,N_17573);
and U20543 (N_20543,N_17607,N_19652);
or U20544 (N_20544,N_19576,N_18309);
and U20545 (N_20545,N_18126,N_18107);
and U20546 (N_20546,N_17828,N_18271);
xor U20547 (N_20547,N_19864,N_19069);
nand U20548 (N_20548,N_18554,N_18792);
or U20549 (N_20549,N_18561,N_18511);
xor U20550 (N_20550,N_19717,N_19422);
or U20551 (N_20551,N_17741,N_17553);
and U20552 (N_20552,N_18670,N_19774);
and U20553 (N_20553,N_17664,N_18013);
or U20554 (N_20554,N_19126,N_18442);
nand U20555 (N_20555,N_19312,N_19863);
and U20556 (N_20556,N_18615,N_19814);
nor U20557 (N_20557,N_18749,N_19684);
or U20558 (N_20558,N_19407,N_19634);
nand U20559 (N_20559,N_17856,N_18424);
and U20560 (N_20560,N_17862,N_18637);
and U20561 (N_20561,N_18033,N_19317);
or U20562 (N_20562,N_17600,N_19052);
xor U20563 (N_20563,N_19834,N_18438);
xor U20564 (N_20564,N_18854,N_17734);
xnor U20565 (N_20565,N_18619,N_18260);
nor U20566 (N_20566,N_18282,N_18022);
nand U20567 (N_20567,N_19589,N_18840);
and U20568 (N_20568,N_18074,N_18207);
and U20569 (N_20569,N_18201,N_19765);
and U20570 (N_20570,N_17590,N_18533);
xor U20571 (N_20571,N_19054,N_19426);
xor U20572 (N_20572,N_18242,N_17712);
nand U20573 (N_20573,N_17677,N_18050);
and U20574 (N_20574,N_17927,N_18866);
xnor U20575 (N_20575,N_18341,N_19385);
nand U20576 (N_20576,N_19337,N_18183);
and U20577 (N_20577,N_17506,N_19419);
xor U20578 (N_20578,N_18997,N_18147);
or U20579 (N_20579,N_18130,N_18653);
or U20580 (N_20580,N_19133,N_19885);
nor U20581 (N_20581,N_17604,N_17803);
or U20582 (N_20582,N_17512,N_19387);
or U20583 (N_20583,N_19288,N_19523);
or U20584 (N_20584,N_19246,N_17654);
nor U20585 (N_20585,N_19166,N_19316);
xor U20586 (N_20586,N_18665,N_18940);
or U20587 (N_20587,N_17991,N_19831);
and U20588 (N_20588,N_19615,N_18962);
or U20589 (N_20589,N_19525,N_18739);
or U20590 (N_20590,N_18112,N_19181);
and U20591 (N_20591,N_17698,N_17719);
nand U20592 (N_20592,N_18372,N_19707);
nor U20593 (N_20593,N_18379,N_19696);
or U20594 (N_20594,N_19320,N_19386);
nor U20595 (N_20595,N_17955,N_18912);
xor U20596 (N_20596,N_17867,N_18156);
nor U20597 (N_20597,N_18070,N_19013);
xor U20598 (N_20598,N_19878,N_19601);
xnor U20599 (N_20599,N_17733,N_19621);
xor U20600 (N_20600,N_17936,N_18449);
or U20601 (N_20601,N_19116,N_19240);
nand U20602 (N_20602,N_19989,N_17969);
nand U20603 (N_20603,N_19377,N_18848);
nand U20604 (N_20604,N_18557,N_18079);
and U20605 (N_20605,N_18233,N_19619);
or U20606 (N_20606,N_18189,N_18088);
and U20607 (N_20607,N_19147,N_18639);
nor U20608 (N_20608,N_17786,N_17875);
nand U20609 (N_20609,N_19242,N_19668);
nand U20610 (N_20610,N_19198,N_17564);
nor U20611 (N_20611,N_18944,N_18773);
xor U20612 (N_20612,N_18478,N_18142);
nor U20613 (N_20613,N_19120,N_18151);
nand U20614 (N_20614,N_17715,N_19692);
xor U20615 (N_20615,N_19438,N_19309);
nor U20616 (N_20616,N_18445,N_18011);
nor U20617 (N_20617,N_17674,N_18299);
xor U20618 (N_20618,N_19870,N_17676);
nand U20619 (N_20619,N_19605,N_18675);
nand U20620 (N_20620,N_18109,N_18715);
xnor U20621 (N_20621,N_18390,N_17710);
or U20622 (N_20622,N_19517,N_18882);
xnor U20623 (N_20623,N_17841,N_17612);
xnor U20624 (N_20624,N_18617,N_19879);
and U20625 (N_20625,N_19251,N_17818);
or U20626 (N_20626,N_17615,N_19301);
nor U20627 (N_20627,N_18440,N_19534);
nand U20628 (N_20628,N_19450,N_19654);
xnor U20629 (N_20629,N_18304,N_19933);
nor U20630 (N_20630,N_18051,N_18566);
xnor U20631 (N_20631,N_18822,N_17878);
xor U20632 (N_20632,N_19099,N_18686);
nand U20633 (N_20633,N_19897,N_19775);
nand U20634 (N_20634,N_18721,N_19678);
or U20635 (N_20635,N_18059,N_18173);
or U20636 (N_20636,N_19376,N_19180);
nand U20637 (N_20637,N_18488,N_18529);
nor U20638 (N_20638,N_18336,N_19258);
and U20639 (N_20639,N_18255,N_17656);
and U20640 (N_20640,N_19636,N_19210);
nand U20641 (N_20641,N_19458,N_19476);
nor U20642 (N_20642,N_18231,N_17673);
or U20643 (N_20643,N_19155,N_17630);
nand U20644 (N_20644,N_18906,N_18667);
and U20645 (N_20645,N_19773,N_19055);
nand U20646 (N_20646,N_18223,N_19462);
or U20647 (N_20647,N_18851,N_18652);
or U20648 (N_20648,N_18073,N_18796);
nor U20649 (N_20649,N_19097,N_17508);
and U20650 (N_20650,N_17964,N_18709);
xnor U20651 (N_20651,N_18918,N_18037);
nor U20652 (N_20652,N_18970,N_18127);
nand U20653 (N_20653,N_18470,N_19551);
xor U20654 (N_20654,N_18095,N_18235);
xor U20655 (N_20655,N_19992,N_18041);
and U20656 (N_20656,N_18785,N_18498);
and U20657 (N_20657,N_17758,N_19081);
nand U20658 (N_20658,N_18948,N_19903);
nor U20659 (N_20659,N_17925,N_19228);
or U20660 (N_20660,N_18510,N_19780);
nand U20661 (N_20661,N_19267,N_18980);
or U20662 (N_20662,N_18884,N_19552);
nand U20663 (N_20663,N_19762,N_19095);
xor U20664 (N_20664,N_17906,N_18347);
nand U20665 (N_20665,N_18570,N_19433);
xor U20666 (N_20666,N_18552,N_19890);
and U20667 (N_20667,N_18435,N_19033);
nand U20668 (N_20668,N_19756,N_17866);
or U20669 (N_20669,N_18203,N_18903);
xnor U20670 (N_20670,N_18893,N_19466);
or U20671 (N_20671,N_19364,N_19757);
nand U20672 (N_20672,N_18701,N_17857);
or U20673 (N_20673,N_18553,N_19802);
nor U20674 (N_20674,N_19977,N_17972);
nand U20675 (N_20675,N_19260,N_19084);
xnor U20676 (N_20676,N_18023,N_19010);
nand U20677 (N_20677,N_19635,N_19040);
nor U20678 (N_20678,N_19163,N_19764);
or U20679 (N_20679,N_18722,N_18176);
xnor U20680 (N_20680,N_17653,N_19826);
and U20681 (N_20681,N_18472,N_18945);
nand U20682 (N_20682,N_18549,N_18742);
or U20683 (N_20683,N_18485,N_19026);
xnor U20684 (N_20684,N_18141,N_19888);
or U20685 (N_20685,N_19017,N_18895);
or U20686 (N_20686,N_19617,N_18522);
nor U20687 (N_20687,N_19357,N_18919);
nor U20688 (N_20688,N_19074,N_18963);
and U20689 (N_20689,N_17572,N_19404);
nand U20690 (N_20690,N_19961,N_19282);
or U20691 (N_20691,N_18068,N_17584);
or U20692 (N_20692,N_19089,N_17761);
or U20693 (N_20693,N_19016,N_17788);
nor U20694 (N_20694,N_19442,N_19007);
and U20695 (N_20695,N_19409,N_18933);
or U20696 (N_20696,N_17569,N_18277);
and U20697 (N_20697,N_19818,N_19614);
nand U20698 (N_20698,N_18974,N_19025);
or U20699 (N_20699,N_17707,N_18121);
nor U20700 (N_20700,N_17960,N_18475);
nor U20701 (N_20701,N_19236,N_18661);
xor U20702 (N_20702,N_18288,N_17909);
or U20703 (N_20703,N_18148,N_18350);
nor U20704 (N_20704,N_18427,N_19667);
xnor U20705 (N_20705,N_19531,N_19686);
xor U20706 (N_20706,N_19507,N_19002);
xor U20707 (N_20707,N_18691,N_19777);
nor U20708 (N_20708,N_19518,N_18795);
and U20709 (N_20709,N_19999,N_17806);
and U20710 (N_20710,N_19921,N_17776);
nor U20711 (N_20711,N_18232,N_18197);
nor U20712 (N_20712,N_19118,N_17994);
nor U20713 (N_20713,N_17566,N_18367);
or U20714 (N_20714,N_18447,N_19303);
xnor U20715 (N_20715,N_18186,N_19431);
and U20716 (N_20716,N_19711,N_19567);
and U20717 (N_20717,N_19279,N_18618);
nand U20718 (N_20718,N_19319,N_19833);
or U20719 (N_20719,N_17823,N_18870);
or U20720 (N_20720,N_18480,N_19710);
nor U20721 (N_20721,N_17860,N_19839);
and U20722 (N_20722,N_19169,N_19851);
and U20723 (N_20723,N_19034,N_17747);
nor U20724 (N_20724,N_17798,N_18828);
xor U20725 (N_20725,N_18131,N_18504);
or U20726 (N_20726,N_17879,N_19225);
nand U20727 (N_20727,N_19970,N_18380);
or U20728 (N_20728,N_18250,N_17760);
nand U20729 (N_20729,N_18411,N_18055);
nand U20730 (N_20730,N_18646,N_17829);
nor U20731 (N_20731,N_19603,N_18624);
or U20732 (N_20732,N_18248,N_17700);
or U20733 (N_20733,N_17517,N_17709);
or U20734 (N_20734,N_19468,N_19981);
nand U20735 (N_20735,N_19481,N_19860);
nor U20736 (N_20736,N_17834,N_19852);
nor U20737 (N_20737,N_19772,N_17968);
or U20738 (N_20738,N_19657,N_17644);
and U20739 (N_20739,N_17929,N_19521);
xnor U20740 (N_20740,N_18704,N_17684);
nand U20741 (N_20741,N_18294,N_18875);
nor U20742 (N_20742,N_19524,N_18938);
nand U20743 (N_20743,N_19454,N_19644);
and U20744 (N_20744,N_17997,N_18574);
nand U20745 (N_20745,N_17608,N_18181);
xnor U20746 (N_20746,N_18961,N_19445);
xor U20747 (N_20747,N_19556,N_17825);
nand U20748 (N_20748,N_17587,N_18461);
and U20749 (N_20749,N_18613,N_17804);
nand U20750 (N_20750,N_19086,N_19216);
or U20751 (N_20751,N_17838,N_19217);
nor U20752 (N_20752,N_19712,N_18525);
nand U20753 (N_20753,N_19156,N_17620);
nor U20754 (N_20754,N_19083,N_18382);
and U20755 (N_20755,N_17552,N_18869);
nor U20756 (N_20756,N_18606,N_18913);
xnor U20757 (N_20757,N_19311,N_19642);
and U20758 (N_20758,N_19813,N_19558);
and U20759 (N_20759,N_19375,N_19315);
nor U20760 (N_20760,N_17713,N_19322);
nor U20761 (N_20761,N_18687,N_18765);
nor U20762 (N_20762,N_17975,N_19766);
nor U20763 (N_20763,N_19213,N_17868);
nand U20764 (N_20764,N_19598,N_18986);
and U20765 (N_20765,N_17579,N_19059);
or U20766 (N_20766,N_19491,N_19333);
nand U20767 (N_20767,N_18019,N_19148);
xor U20768 (N_20768,N_19555,N_18345);
nand U20769 (N_20769,N_17522,N_17756);
nand U20770 (N_20770,N_19611,N_19638);
xnor U20771 (N_20771,N_17854,N_18300);
or U20772 (N_20772,N_18180,N_19799);
nor U20773 (N_20773,N_17884,N_19340);
or U20774 (N_20774,N_19670,N_18519);
nand U20775 (N_20775,N_18542,N_17669);
and U20776 (N_20776,N_19220,N_18185);
and U20777 (N_20777,N_18650,N_17942);
or U20778 (N_20778,N_19516,N_18252);
and U20779 (N_20779,N_18210,N_18343);
nand U20780 (N_20780,N_17519,N_18145);
xnor U20781 (N_20781,N_17534,N_19295);
and U20782 (N_20782,N_18208,N_19631);
xnor U20783 (N_20783,N_18253,N_18491);
nor U20784 (N_20784,N_19134,N_17791);
or U20785 (N_20785,N_17769,N_19048);
nor U20786 (N_20786,N_19115,N_19742);
xor U20787 (N_20787,N_19924,N_18415);
nand U20788 (N_20788,N_17796,N_18829);
nand U20789 (N_20789,N_19395,N_18090);
or U20790 (N_20790,N_18711,N_18117);
and U20791 (N_20791,N_19609,N_19187);
xor U20792 (N_20792,N_19855,N_18727);
or U20793 (N_20793,N_19987,N_17737);
nor U20794 (N_20794,N_18307,N_18437);
nor U20795 (N_20795,N_18863,N_19810);
and U20796 (N_20796,N_18240,N_18605);
nand U20797 (N_20797,N_17641,N_18195);
or U20798 (N_20798,N_19170,N_19894);
xnor U20799 (N_20799,N_19435,N_19627);
nand U20800 (N_20800,N_19859,N_18228);
xnor U20801 (N_20801,N_19950,N_18744);
nand U20802 (N_20802,N_17961,N_18540);
nand U20803 (N_20803,N_17973,N_18469);
and U20804 (N_20804,N_18460,N_17724);
nand U20805 (N_20805,N_17945,N_18941);
xnor U20806 (N_20806,N_19132,N_19789);
xnor U20807 (N_20807,N_18071,N_18072);
or U20808 (N_20808,N_18788,N_18896);
or U20809 (N_20809,N_18360,N_18099);
and U20810 (N_20810,N_17904,N_19771);
xor U20811 (N_20811,N_18311,N_17646);
xor U20812 (N_20812,N_19532,N_18120);
or U20813 (N_20813,N_17989,N_17666);
xnor U20814 (N_20814,N_18018,N_19962);
nor U20815 (N_20815,N_17908,N_17736);
xor U20816 (N_20816,N_18819,N_18971);
nand U20817 (N_20817,N_19327,N_18110);
or U20818 (N_20818,N_18152,N_19401);
xor U20819 (N_20819,N_19157,N_19778);
xnor U20820 (N_20820,N_19540,N_18301);
nand U20821 (N_20821,N_18436,N_19437);
and U20822 (N_20822,N_18035,N_19610);
nor U20823 (N_20823,N_18535,N_18780);
xnor U20824 (N_20824,N_17532,N_19172);
and U20825 (N_20825,N_18578,N_19153);
and U20826 (N_20826,N_17755,N_19294);
and U20827 (N_20827,N_18100,N_17981);
nand U20828 (N_20828,N_18547,N_17986);
nor U20829 (N_20829,N_19171,N_18798);
nor U20830 (N_20830,N_18381,N_17993);
xor U20831 (N_20831,N_17658,N_18576);
and U20832 (N_20832,N_19178,N_18524);
nand U20833 (N_20833,N_19562,N_18384);
xnor U20834 (N_20834,N_17729,N_17949);
and U20835 (N_20835,N_18287,N_18136);
xor U20836 (N_20836,N_19527,N_18244);
or U20837 (N_20837,N_18685,N_19072);
nor U20838 (N_20838,N_18868,N_18135);
or U20839 (N_20839,N_19857,N_18596);
and U20840 (N_20840,N_18428,N_17717);
or U20841 (N_20841,N_18544,N_19330);
nor U20842 (N_20842,N_18608,N_17800);
xor U20843 (N_20843,N_17842,N_19972);
xnor U20844 (N_20844,N_17623,N_19425);
xnor U20845 (N_20845,N_17790,N_19990);
or U20846 (N_20846,N_17952,N_18215);
and U20847 (N_20847,N_18466,N_19428);
xnor U20848 (N_20848,N_19673,N_19620);
or U20849 (N_20849,N_18734,N_17853);
xor U20850 (N_20850,N_19488,N_18694);
nor U20851 (N_20851,N_18857,N_18883);
nand U20852 (N_20852,N_19588,N_19843);
or U20853 (N_20853,N_18316,N_17699);
and U20854 (N_20854,N_19325,N_19268);
xnor U20855 (N_20855,N_19406,N_19039);
nand U20856 (N_20856,N_18978,N_18799);
xnor U20857 (N_20857,N_19510,N_18170);
nand U20858 (N_20858,N_17934,N_19867);
nor U20859 (N_20859,N_19749,N_18532);
xor U20860 (N_20860,N_18417,N_19679);
xor U20861 (N_20861,N_19882,N_19728);
nor U20862 (N_20862,N_19577,N_19497);
xor U20863 (N_20863,N_19948,N_19760);
and U20864 (N_20864,N_18297,N_18595);
or U20865 (N_20865,N_19689,N_17660);
xor U20866 (N_20866,N_18239,N_18911);
nand U20867 (N_20867,N_19548,N_18936);
xnor U20868 (N_20868,N_19965,N_18807);
nor U20869 (N_20869,N_17643,N_19912);
xnor U20870 (N_20870,N_19030,N_18843);
nor U20871 (N_20871,N_17766,N_18707);
nand U20872 (N_20872,N_19113,N_18482);
xor U20873 (N_20873,N_18332,N_18258);
nor U20874 (N_20874,N_19522,N_17703);
nand U20875 (N_20875,N_17894,N_18129);
nor U20876 (N_20876,N_18649,N_19068);
or U20877 (N_20877,N_18284,N_18515);
nor U20878 (N_20878,N_19058,N_18078);
nand U20879 (N_20879,N_18179,N_19740);
nand U20880 (N_20880,N_17515,N_19714);
xor U20881 (N_20881,N_19087,N_17913);
nand U20882 (N_20882,N_18164,N_17924);
nand U20883 (N_20883,N_19883,N_18040);
xor U20884 (N_20884,N_18768,N_18826);
or U20885 (N_20885,N_18108,N_17757);
and U20886 (N_20886,N_19669,N_19391);
nand U20887 (N_20887,N_18420,N_18958);
xnor U20888 (N_20888,N_19056,N_17932);
nand U20889 (N_20889,N_19291,N_18276);
xor U20890 (N_20890,N_18105,N_17881);
and U20891 (N_20891,N_18326,N_19964);
nor U20892 (N_20892,N_19564,N_17748);
nand U20893 (N_20893,N_19751,N_18621);
nand U20894 (N_20894,N_17503,N_17971);
xor U20895 (N_20895,N_19630,N_17690);
nor U20896 (N_20896,N_18808,N_19622);
xor U20897 (N_20897,N_18103,N_18236);
nand U20898 (N_20898,N_17547,N_17613);
nand U20899 (N_20899,N_17917,N_18413);
nand U20900 (N_20900,N_18123,N_19811);
xnor U20901 (N_20901,N_18084,N_18907);
xnor U20902 (N_20902,N_19203,N_18312);
xnor U20903 (N_20903,N_17585,N_18957);
nand U20904 (N_20904,N_18398,N_18279);
nand U20905 (N_20905,N_17583,N_17628);
nor U20906 (N_20906,N_17850,N_18521);
xnor U20907 (N_20907,N_19553,N_19846);
and U20908 (N_20908,N_19779,N_19044);
nand U20909 (N_20909,N_17792,N_19158);
nor U20910 (N_20910,N_18743,N_18004);
or U20911 (N_20911,N_18481,N_18052);
and U20912 (N_20912,N_17567,N_18206);
nand U20913 (N_20913,N_18697,N_19651);
or U20914 (N_20914,N_19119,N_17542);
xor U20915 (N_20915,N_18450,N_19065);
xor U20916 (N_20916,N_17636,N_17933);
and U20917 (N_20917,N_19608,N_18471);
nor U20918 (N_20918,N_17695,N_18708);
and U20919 (N_20919,N_19741,N_19591);
xnor U20920 (N_20920,N_17510,N_18202);
and U20921 (N_20921,N_19136,N_17546);
xnor U20922 (N_20922,N_19165,N_19451);
or U20923 (N_20923,N_17625,N_17551);
and U20924 (N_20924,N_18812,N_18894);
and U20925 (N_20925,N_18425,N_19003);
nand U20926 (N_20926,N_18009,N_19647);
nor U20927 (N_20927,N_19600,N_19261);
nand U20928 (N_20928,N_19832,N_18737);
xnor U20929 (N_20929,N_18082,N_18643);
xnor U20930 (N_20930,N_19829,N_18154);
nand U20931 (N_20931,N_19511,N_19191);
nor U20932 (N_20932,N_19578,N_18599);
or U20933 (N_20933,N_18409,N_17938);
or U20934 (N_20934,N_19308,N_19499);
xnor U20935 (N_20935,N_18393,N_19399);
nor U20936 (N_20936,N_19968,N_17723);
xnor U20937 (N_20937,N_19602,N_19287);
nand U20938 (N_20938,N_17706,N_19996);
and U20939 (N_20939,N_18140,N_17732);
xor U20940 (N_20940,N_17980,N_19141);
nand U20941 (N_20941,N_19565,N_18776);
nand U20942 (N_20942,N_17731,N_18756);
xnor U20943 (N_20943,N_19594,N_17727);
and U20944 (N_20944,N_17999,N_17504);
or U20945 (N_20945,N_17808,N_19229);
xor U20946 (N_20946,N_18881,N_18274);
nor U20947 (N_20947,N_17896,N_17538);
or U20948 (N_20948,N_18348,N_18410);
xor U20949 (N_20949,N_17632,N_18797);
or U20950 (N_20950,N_18444,N_19590);
or U20951 (N_20951,N_18769,N_19560);
xnor U20952 (N_20952,N_17634,N_18551);
xor U20953 (N_20953,N_18766,N_17570);
nand U20954 (N_20954,N_19984,N_18490);
nand U20955 (N_20955,N_18219,N_19486);
or U20956 (N_20956,N_18237,N_17667);
nand U20957 (N_20957,N_18414,N_19526);
xnor U20958 (N_20958,N_19900,N_19805);
nor U20959 (N_20959,N_18432,N_18594);
nand U20960 (N_20960,N_17880,N_18992);
nor U20961 (N_20961,N_19174,N_18122);
nand U20962 (N_20962,N_19350,N_18818);
or U20963 (N_20963,N_18872,N_17516);
xnor U20964 (N_20964,N_19373,N_19244);
and U20965 (N_20965,N_18688,N_19221);
nor U20966 (N_20966,N_17799,N_19066);
xor U20967 (N_20967,N_18852,N_18726);
or U20968 (N_20968,N_17686,N_18934);
or U20969 (N_20969,N_19699,N_18200);
xor U20970 (N_20970,N_19477,N_19472);
nor U20971 (N_20971,N_18991,N_18695);
and U20972 (N_20972,N_17831,N_19694);
nor U20973 (N_20973,N_18545,N_19505);
and U20974 (N_20974,N_19152,N_19761);
nor U20975 (N_20975,N_18564,N_18354);
and U20976 (N_20976,N_19645,N_19937);
or U20977 (N_20977,N_19963,N_17530);
nand U20978 (N_20978,N_18338,N_19176);
nor U20979 (N_20979,N_18623,N_18305);
and U20980 (N_20980,N_19509,N_19943);
and U20981 (N_20981,N_17693,N_17772);
nand U20982 (N_20982,N_17876,N_17591);
nand U20983 (N_20983,N_19341,N_18081);
nand U20984 (N_20984,N_18878,N_18182);
or U20985 (N_20985,N_17683,N_18589);
xor U20986 (N_20986,N_18330,N_19500);
and U20987 (N_20987,N_19378,N_18771);
and U20988 (N_20988,N_18910,N_17951);
xor U20989 (N_20989,N_19078,N_18451);
or U20990 (N_20990,N_17827,N_17811);
or U20991 (N_20991,N_18680,N_19421);
and U20992 (N_20992,N_19440,N_18474);
and U20993 (N_20993,N_17897,N_19819);
nand U20994 (N_20994,N_17586,N_19739);
nor U20995 (N_20995,N_18862,N_17821);
or U20996 (N_20996,N_19583,N_18804);
nand U20997 (N_20997,N_17502,N_18580);
and U20998 (N_20998,N_17912,N_18512);
and U20999 (N_20999,N_19299,N_18625);
nor U21000 (N_21000,N_18648,N_18368);
nand U21001 (N_21001,N_19075,N_17787);
and U21002 (N_21002,N_18392,N_18922);
or U21003 (N_21003,N_18402,N_17864);
or U21004 (N_21004,N_18942,N_19504);
xnor U21005 (N_21005,N_17922,N_19646);
nand U21006 (N_21006,N_17665,N_17577);
xnor U21007 (N_21007,N_17872,N_18146);
or U21008 (N_21008,N_18269,N_18407);
xnor U21009 (N_21009,N_18791,N_17874);
and U21010 (N_21010,N_19457,N_19629);
xor U21011 (N_21011,N_19139,N_18259);
nor U21012 (N_21012,N_18556,N_18889);
or U21013 (N_21013,N_19776,N_19286);
nand U21014 (N_21014,N_17814,N_19383);
nor U21015 (N_21015,N_18273,N_19257);
nand U21016 (N_21016,N_19547,N_17746);
nor U21017 (N_21017,N_17899,N_18611);
nor U21018 (N_21018,N_17822,N_17739);
nand U21019 (N_21019,N_18064,N_18062);
nand U21020 (N_21020,N_18628,N_17815);
and U21021 (N_21021,N_17848,N_19795);
or U21022 (N_21022,N_19273,N_18956);
nor U21023 (N_21023,N_18746,N_18526);
and U21024 (N_21024,N_18634,N_19988);
or U21025 (N_21025,N_17770,N_18213);
or U21026 (N_21026,N_18397,N_18716);
and U21027 (N_21027,N_19561,N_18317);
or U21028 (N_21028,N_19393,N_19361);
nand U21029 (N_21029,N_18280,N_17852);
or U21030 (N_21030,N_18172,N_18638);
or U21031 (N_21031,N_18355,N_19506);
nor U21032 (N_21032,N_18174,N_19290);
nand U21033 (N_21033,N_18254,N_19253);
nand U21034 (N_21034,N_18096,N_18261);
nor U21035 (N_21035,N_17979,N_18689);
or U21036 (N_21036,N_19117,N_19088);
nor U21037 (N_21037,N_19915,N_18101);
and U21038 (N_21038,N_17967,N_19189);
nand U21039 (N_21039,N_18536,N_17910);
nor U21040 (N_21040,N_18692,N_19952);
xor U21041 (N_21041,N_19880,N_19956);
nand U21042 (N_21042,N_19993,N_19628);
xor U21043 (N_21043,N_18465,N_18296);
nor U21044 (N_21044,N_19128,N_19356);
xor U21045 (N_21045,N_19872,N_19884);
nor U21046 (N_21046,N_19208,N_17520);
nor U21047 (N_21047,N_18125,N_18600);
xor U21048 (N_21048,N_18748,N_19196);
or U21049 (N_21049,N_19254,N_19865);
nor U21050 (N_21050,N_17716,N_19842);
nor U21051 (N_21051,N_17720,N_18777);
nand U21052 (N_21052,N_19685,N_18627);
nand U21053 (N_21053,N_18506,N_18459);
nand U21054 (N_21054,N_18683,N_18614);
or U21055 (N_21055,N_19329,N_19326);
or U21056 (N_21056,N_19278,N_18489);
or U21057 (N_21057,N_19051,N_17810);
and U21058 (N_21058,N_18370,N_19223);
nand U21059 (N_21059,N_18836,N_18642);
or U21060 (N_21060,N_17738,N_19429);
nor U21061 (N_21061,N_19681,N_19676);
and U21062 (N_21062,N_18585,N_19904);
and U21063 (N_21063,N_17920,N_18886);
and U21064 (N_21064,N_17974,N_18993);
xnor U21065 (N_21065,N_19434,N_19200);
xor U21066 (N_21066,N_17559,N_19452);
nand U21067 (N_21067,N_18306,N_19881);
nor U21068 (N_21068,N_19183,N_19164);
and U21069 (N_21069,N_19249,N_19238);
nand U21070 (N_21070,N_19559,N_17983);
or U21071 (N_21071,N_18335,N_19704);
or U21072 (N_21072,N_18641,N_19569);
or U21073 (N_21073,N_17777,N_19641);
nor U21074 (N_21074,N_19979,N_18222);
or U21075 (N_21075,N_19345,N_18137);
or U21076 (N_21076,N_19032,N_17923);
and U21077 (N_21077,N_18757,N_17877);
nand U21078 (N_21078,N_18950,N_18876);
and U21079 (N_21079,N_18007,N_18821);
or U21080 (N_21080,N_17763,N_19655);
and U21081 (N_21081,N_19735,N_19639);
or U21082 (N_21082,N_19557,N_18443);
or U21083 (N_21083,N_17582,N_18959);
xor U21084 (N_21084,N_19372,N_19758);
or U21085 (N_21085,N_19102,N_19746);
nor U21086 (N_21086,N_18678,N_17995);
nand U21087 (N_21087,N_17948,N_19202);
or U21088 (N_21088,N_18655,N_17601);
nor U21089 (N_21089,N_17892,N_18789);
xor U21090 (N_21090,N_19417,N_17943);
and U21091 (N_21091,N_17744,N_17754);
xnor U21092 (N_21092,N_19755,N_19687);
and U21093 (N_21093,N_17640,N_18351);
nand U21094 (N_21094,N_18419,N_18587);
nand U21095 (N_21095,N_18998,N_19706);
or U21096 (N_21096,N_18264,N_18850);
or U21097 (N_21097,N_18053,N_18014);
or U21098 (N_21098,N_18728,N_19302);
nand U21099 (N_21099,N_18188,N_19194);
nand U21100 (N_21100,N_19759,N_17849);
or U21101 (N_21101,N_18901,N_18891);
nand U21102 (N_21102,N_17596,N_19820);
or U21103 (N_21103,N_19936,N_18946);
xor U21104 (N_21104,N_18349,N_17603);
and U21105 (N_21105,N_19368,N_17648);
or U21106 (N_21106,N_19906,N_19893);
nor U21107 (N_21107,N_19219,N_18983);
nor U21108 (N_21108,N_19355,N_18016);
or U21109 (N_21109,N_19659,N_19024);
nand U21110 (N_21110,N_18238,N_18468);
xor U21111 (N_21111,N_17843,N_19935);
nand U21112 (N_21112,N_19549,N_17992);
nand U21113 (N_21113,N_19953,N_18416);
nor U21114 (N_21114,N_19858,N_17685);
or U21115 (N_21115,N_17560,N_18999);
and U21116 (N_21116,N_18268,N_17743);
nand U21117 (N_21117,N_19471,N_19690);
xor U21118 (N_21118,N_19782,N_17670);
xor U21119 (N_21119,N_19124,N_18492);
or U21120 (N_21120,N_18673,N_18373);
nor U21121 (N_21121,N_17859,N_18111);
xor U21122 (N_21122,N_19902,N_17865);
nand U21123 (N_21123,N_19781,N_18467);
or U21124 (N_21124,N_19063,N_18939);
and U21125 (N_21125,N_19974,N_18057);
nor U21126 (N_21126,N_19994,N_18434);
nor U21127 (N_21127,N_17539,N_17889);
and U21128 (N_21128,N_18049,N_18560);
and U21129 (N_21129,N_19009,N_18187);
and U21130 (N_21130,N_19637,N_19008);
nand U21131 (N_21131,N_18841,N_17775);
or U21132 (N_21132,N_19731,N_17540);
xor U21133 (N_21133,N_18396,N_19265);
xor U21134 (N_21134,N_19480,N_18725);
and U21135 (N_21135,N_19868,N_19358);
and U21136 (N_21136,N_19248,N_17782);
nor U21137 (N_21137,N_18029,N_19460);
xnor U21138 (N_21138,N_19625,N_18837);
and U21139 (N_21139,N_18462,N_19995);
xnor U21140 (N_21140,N_19332,N_18865);
or U21141 (N_21141,N_19693,N_19146);
xor U21142 (N_21142,N_18758,N_19310);
xor U21143 (N_21143,N_19543,N_19305);
or U21144 (N_21144,N_17616,N_19441);
or U21145 (N_21145,N_18877,N_19342);
or U21146 (N_21146,N_18497,N_18006);
xor U21147 (N_21147,N_19911,N_19663);
and U21148 (N_21148,N_17592,N_17795);
nand U21149 (N_21149,N_17563,N_18786);
and U21150 (N_21150,N_19946,N_19848);
xnor U21151 (N_21151,N_18871,N_18706);
or U21152 (N_21152,N_17657,N_17801);
and U21153 (N_21153,N_17765,N_19321);
nor U21154 (N_21154,N_17682,N_17609);
xnor U21155 (N_21155,N_18364,N_19929);
xor U21156 (N_21156,N_19733,N_17835);
nand U21157 (N_21157,N_19917,N_18159);
and U21158 (N_21158,N_18003,N_19125);
and U21159 (N_21159,N_19643,N_19934);
or U21160 (N_21160,N_19085,N_18698);
and U21161 (N_21161,N_18225,N_18856);
nand U21162 (N_21162,N_18834,N_19218);
xnor U21163 (N_21163,N_19304,N_19080);
xnor U21164 (N_21164,N_17824,N_19446);
and U21165 (N_21165,N_19770,N_19563);
xnor U21166 (N_21166,N_19980,N_17680);
nor U21167 (N_21167,N_19167,N_18859);
nand U21168 (N_21168,N_17523,N_19493);
nor U21169 (N_21169,N_19703,N_18835);
xor U21170 (N_21170,N_18097,N_18047);
nand U21171 (N_21171,N_18265,N_18319);
nor U21172 (N_21172,N_18864,N_18827);
nand U21173 (N_21173,N_17561,N_19121);
nor U21174 (N_21174,N_19028,N_17647);
xor U21175 (N_21175,N_17793,N_18647);
xor U21176 (N_21176,N_17671,N_17689);
xor U21177 (N_21177,N_19318,N_19455);
nand U21178 (N_21178,N_19487,N_19550);
nand U21179 (N_21179,N_18017,N_18162);
or U21180 (N_21180,N_18772,N_18245);
and U21181 (N_21181,N_19925,N_17805);
nand U21182 (N_21182,N_18149,N_17950);
or U21183 (N_21183,N_18651,N_19734);
nor U21184 (N_21184,N_19599,N_19853);
or U21185 (N_21185,N_19850,N_19922);
or U21186 (N_21186,N_17830,N_19496);
xnor U21187 (N_21187,N_17509,N_19145);
xor U21188 (N_21188,N_18446,N_18508);
nand U21189 (N_21189,N_17544,N_18928);
or U21190 (N_21190,N_19535,N_18805);
and U21191 (N_21191,N_18927,N_19382);
nand U21192 (N_21192,N_19207,N_18897);
nor U21193 (N_21193,N_17675,N_19397);
xnor U21194 (N_21194,N_17817,N_19241);
and U21195 (N_21195,N_19732,N_17521);
and U21196 (N_21196,N_18493,N_18214);
xor U21197 (N_21197,N_17780,N_19949);
and U21198 (N_21198,N_18221,N_18577);
xnor U21199 (N_21199,N_18048,N_18157);
nand U21200 (N_21200,N_18920,N_19530);
xor U21201 (N_21201,N_18811,N_18932);
and U21202 (N_21202,N_19182,N_18696);
xnor U21203 (N_21203,N_19149,N_17928);
xnor U21204 (N_21204,N_17571,N_19019);
nor U21205 (N_21205,N_17957,N_19230);
or U21206 (N_21206,N_18395,N_18954);
and U21207 (N_21207,N_18530,N_18357);
and U21208 (N_21208,N_19015,N_18171);
nand U21209 (N_21209,N_18166,N_18951);
and U21210 (N_21210,N_19579,N_18964);
nand U21211 (N_21211,N_19186,N_18028);
xnor U21212 (N_21212,N_18080,N_19845);
or U21213 (N_21213,N_19568,N_17767);
and U21214 (N_21214,N_19430,N_17898);
nor U21215 (N_21215,N_18989,N_18477);
or U21216 (N_21216,N_19256,N_17598);
nor U21217 (N_21217,N_17990,N_17533);
nand U21218 (N_21218,N_18809,N_18981);
nor U21219 (N_21219,N_19502,N_18632);
nor U21220 (N_21220,N_19370,N_18565);
and U21221 (N_21221,N_19143,N_18001);
nor U21222 (N_21222,N_18994,N_18924);
nor U21223 (N_21223,N_19266,N_19233);
nand U21224 (N_21224,N_18720,N_17982);
xor U21225 (N_21225,N_18144,N_18175);
nand U21226 (N_21226,N_18177,N_17911);
or U21227 (N_21227,N_18463,N_19479);
and U21228 (N_21228,N_18762,N_18322);
xnor U21229 (N_21229,N_17901,N_19110);
xor U21230 (N_21230,N_18486,N_19137);
nand U21231 (N_21231,N_19402,N_19612);
nand U21232 (N_21232,N_19154,N_17956);
nand U21233 (N_21233,N_17576,N_18005);
nor U21234 (N_21234,N_19129,N_17836);
xnor U21235 (N_21235,N_18537,N_18926);
xor U21236 (N_21236,N_18816,N_19708);
or U21237 (N_21237,N_19698,N_19982);
and U21238 (N_21238,N_18104,N_19298);
or U21239 (N_21239,N_19896,N_18441);
nand U21240 (N_21240,N_18204,N_17809);
and U21241 (N_21241,N_17781,N_18257);
or U21242 (N_21242,N_18352,N_19077);
xnor U21243 (N_21243,N_19958,N_19160);
and U21244 (N_21244,N_18369,N_19519);
nor U21245 (N_21245,N_17556,N_19138);
nor U21246 (N_21246,N_19482,N_18800);
nor U21247 (N_21247,N_19895,N_19410);
or U21248 (N_21248,N_18968,N_19338);
nor U21249 (N_21249,N_19913,N_18833);
nand U21250 (N_21250,N_19620,N_19982);
nand U21251 (N_21251,N_18158,N_18369);
xor U21252 (N_21252,N_19459,N_19724);
and U21253 (N_21253,N_17559,N_17699);
xnor U21254 (N_21254,N_18266,N_18748);
and U21255 (N_21255,N_19249,N_19074);
or U21256 (N_21256,N_18962,N_18195);
nor U21257 (N_21257,N_18237,N_19978);
and U21258 (N_21258,N_18668,N_19520);
nor U21259 (N_21259,N_18165,N_18367);
xor U21260 (N_21260,N_18047,N_19696);
nand U21261 (N_21261,N_18367,N_19512);
or U21262 (N_21262,N_19388,N_18247);
nand U21263 (N_21263,N_19737,N_19975);
and U21264 (N_21264,N_18690,N_18440);
or U21265 (N_21265,N_19320,N_19407);
nand U21266 (N_21266,N_17513,N_19818);
and U21267 (N_21267,N_18703,N_18011);
or U21268 (N_21268,N_19766,N_19050);
xor U21269 (N_21269,N_19434,N_18743);
and U21270 (N_21270,N_18902,N_19096);
and U21271 (N_21271,N_19919,N_18467);
xor U21272 (N_21272,N_17833,N_17887);
nor U21273 (N_21273,N_17647,N_19104);
xnor U21274 (N_21274,N_17805,N_19610);
nand U21275 (N_21275,N_17961,N_17764);
nor U21276 (N_21276,N_18925,N_18632);
xor U21277 (N_21277,N_18382,N_17691);
nand U21278 (N_21278,N_17528,N_18983);
and U21279 (N_21279,N_17632,N_19913);
nor U21280 (N_21280,N_17869,N_18469);
xor U21281 (N_21281,N_19122,N_17723);
or U21282 (N_21282,N_17910,N_19970);
xnor U21283 (N_21283,N_19569,N_18316);
nand U21284 (N_21284,N_19774,N_17690);
and U21285 (N_21285,N_18024,N_19202);
nor U21286 (N_21286,N_18029,N_19930);
and U21287 (N_21287,N_18095,N_19532);
and U21288 (N_21288,N_19319,N_18375);
xnor U21289 (N_21289,N_18181,N_19341);
nor U21290 (N_21290,N_18778,N_19478);
nand U21291 (N_21291,N_18245,N_18266);
nand U21292 (N_21292,N_18313,N_17817);
and U21293 (N_21293,N_18253,N_17703);
and U21294 (N_21294,N_19171,N_19333);
and U21295 (N_21295,N_19120,N_17883);
and U21296 (N_21296,N_18576,N_18196);
nor U21297 (N_21297,N_19500,N_18495);
xor U21298 (N_21298,N_19626,N_18286);
xor U21299 (N_21299,N_18715,N_18853);
xnor U21300 (N_21300,N_18722,N_19760);
nand U21301 (N_21301,N_19672,N_19651);
nor U21302 (N_21302,N_19142,N_19346);
nor U21303 (N_21303,N_19786,N_19346);
nor U21304 (N_21304,N_18391,N_18512);
xnor U21305 (N_21305,N_19407,N_17522);
xor U21306 (N_21306,N_17615,N_18132);
nand U21307 (N_21307,N_18244,N_19465);
nor U21308 (N_21308,N_18974,N_19734);
and U21309 (N_21309,N_19861,N_19717);
xnor U21310 (N_21310,N_17621,N_17655);
xnor U21311 (N_21311,N_19722,N_19619);
nor U21312 (N_21312,N_17506,N_18153);
nand U21313 (N_21313,N_18663,N_19069);
nand U21314 (N_21314,N_19487,N_18928);
nand U21315 (N_21315,N_19174,N_18354);
nand U21316 (N_21316,N_19867,N_17672);
nor U21317 (N_21317,N_18909,N_19021);
nor U21318 (N_21318,N_18136,N_19208);
and U21319 (N_21319,N_18678,N_17804);
and U21320 (N_21320,N_18475,N_17735);
and U21321 (N_21321,N_18831,N_19975);
or U21322 (N_21322,N_19661,N_18460);
or U21323 (N_21323,N_18443,N_19269);
nor U21324 (N_21324,N_18331,N_18963);
or U21325 (N_21325,N_19892,N_19462);
nand U21326 (N_21326,N_17918,N_19623);
and U21327 (N_21327,N_18814,N_18832);
or U21328 (N_21328,N_19670,N_19789);
nor U21329 (N_21329,N_19904,N_18646);
nor U21330 (N_21330,N_17626,N_18390);
xor U21331 (N_21331,N_18355,N_18149);
xor U21332 (N_21332,N_19354,N_19254);
or U21333 (N_21333,N_18441,N_18477);
nand U21334 (N_21334,N_17599,N_19542);
nand U21335 (N_21335,N_18266,N_18723);
and U21336 (N_21336,N_18589,N_17705);
nand U21337 (N_21337,N_19629,N_19000);
xnor U21338 (N_21338,N_18439,N_18545);
and U21339 (N_21339,N_19937,N_18579);
or U21340 (N_21340,N_17992,N_18817);
or U21341 (N_21341,N_19015,N_18497);
xor U21342 (N_21342,N_17789,N_17693);
or U21343 (N_21343,N_18451,N_19789);
xor U21344 (N_21344,N_17909,N_17689);
and U21345 (N_21345,N_18577,N_18321);
and U21346 (N_21346,N_19576,N_19942);
or U21347 (N_21347,N_19758,N_18352);
nand U21348 (N_21348,N_18294,N_18249);
nor U21349 (N_21349,N_18868,N_18193);
or U21350 (N_21350,N_18136,N_18605);
nand U21351 (N_21351,N_19133,N_19372);
and U21352 (N_21352,N_17555,N_19202);
nand U21353 (N_21353,N_18514,N_18825);
and U21354 (N_21354,N_19529,N_17926);
and U21355 (N_21355,N_19741,N_18149);
nor U21356 (N_21356,N_18037,N_17859);
and U21357 (N_21357,N_19462,N_19740);
nor U21358 (N_21358,N_19649,N_19176);
nand U21359 (N_21359,N_18983,N_19376);
nand U21360 (N_21360,N_17995,N_19818);
or U21361 (N_21361,N_18766,N_18354);
nor U21362 (N_21362,N_18693,N_19173);
nand U21363 (N_21363,N_17666,N_19936);
and U21364 (N_21364,N_19810,N_19539);
and U21365 (N_21365,N_19163,N_18030);
nor U21366 (N_21366,N_19990,N_19883);
or U21367 (N_21367,N_19697,N_17573);
and U21368 (N_21368,N_18466,N_18476);
nor U21369 (N_21369,N_18107,N_19943);
nor U21370 (N_21370,N_18666,N_19722);
nor U21371 (N_21371,N_19413,N_17760);
or U21372 (N_21372,N_17795,N_18416);
nor U21373 (N_21373,N_19997,N_17546);
and U21374 (N_21374,N_18763,N_19519);
nor U21375 (N_21375,N_17697,N_19748);
xnor U21376 (N_21376,N_19144,N_19400);
nand U21377 (N_21377,N_19278,N_18907);
and U21378 (N_21378,N_18452,N_18277);
or U21379 (N_21379,N_17863,N_18431);
nor U21380 (N_21380,N_17697,N_18332);
and U21381 (N_21381,N_19940,N_18625);
or U21382 (N_21382,N_17896,N_17730);
nand U21383 (N_21383,N_18879,N_17570);
nand U21384 (N_21384,N_18082,N_18446);
nand U21385 (N_21385,N_18509,N_19131);
xor U21386 (N_21386,N_19326,N_18237);
nand U21387 (N_21387,N_17514,N_19296);
nor U21388 (N_21388,N_17894,N_17672);
xnor U21389 (N_21389,N_19303,N_19429);
and U21390 (N_21390,N_18814,N_19007);
nand U21391 (N_21391,N_19623,N_17838);
or U21392 (N_21392,N_19914,N_17602);
nor U21393 (N_21393,N_19923,N_17660);
or U21394 (N_21394,N_19149,N_19073);
xnor U21395 (N_21395,N_18621,N_19898);
nor U21396 (N_21396,N_19228,N_19857);
xor U21397 (N_21397,N_19585,N_19595);
and U21398 (N_21398,N_19809,N_18547);
and U21399 (N_21399,N_19730,N_18548);
xnor U21400 (N_21400,N_18043,N_18118);
nand U21401 (N_21401,N_19524,N_19264);
xor U21402 (N_21402,N_18644,N_18838);
nand U21403 (N_21403,N_18024,N_18711);
nand U21404 (N_21404,N_18642,N_19425);
nor U21405 (N_21405,N_19507,N_18440);
nor U21406 (N_21406,N_18138,N_18930);
nand U21407 (N_21407,N_19449,N_18574);
xnor U21408 (N_21408,N_19078,N_19498);
xor U21409 (N_21409,N_18222,N_18950);
nand U21410 (N_21410,N_18299,N_18586);
nor U21411 (N_21411,N_19293,N_18589);
xor U21412 (N_21412,N_19180,N_19678);
nor U21413 (N_21413,N_18580,N_18870);
and U21414 (N_21414,N_18381,N_18309);
and U21415 (N_21415,N_18483,N_17795);
nand U21416 (N_21416,N_18158,N_18887);
nor U21417 (N_21417,N_18684,N_19532);
or U21418 (N_21418,N_18808,N_19816);
or U21419 (N_21419,N_18872,N_18486);
nor U21420 (N_21420,N_17810,N_19421);
or U21421 (N_21421,N_18309,N_18211);
xnor U21422 (N_21422,N_18006,N_19551);
and U21423 (N_21423,N_18506,N_19578);
nor U21424 (N_21424,N_18077,N_19574);
nand U21425 (N_21425,N_19575,N_19944);
or U21426 (N_21426,N_19752,N_18005);
nor U21427 (N_21427,N_18137,N_17968);
and U21428 (N_21428,N_18076,N_19326);
nand U21429 (N_21429,N_17983,N_18957);
or U21430 (N_21430,N_17808,N_19620);
nand U21431 (N_21431,N_17981,N_18918);
nand U21432 (N_21432,N_18449,N_19424);
nor U21433 (N_21433,N_18716,N_18956);
xor U21434 (N_21434,N_19965,N_19121);
and U21435 (N_21435,N_19898,N_19806);
nor U21436 (N_21436,N_18654,N_18955);
xor U21437 (N_21437,N_19192,N_17679);
or U21438 (N_21438,N_19334,N_18368);
and U21439 (N_21439,N_17906,N_18979);
or U21440 (N_21440,N_19148,N_19086);
and U21441 (N_21441,N_19803,N_18104);
or U21442 (N_21442,N_18851,N_17846);
nand U21443 (N_21443,N_19051,N_19178);
nand U21444 (N_21444,N_19271,N_18103);
or U21445 (N_21445,N_19849,N_19322);
xor U21446 (N_21446,N_18468,N_18848);
and U21447 (N_21447,N_19663,N_19673);
or U21448 (N_21448,N_19515,N_18915);
or U21449 (N_21449,N_17774,N_19195);
nor U21450 (N_21450,N_18849,N_19811);
nor U21451 (N_21451,N_17964,N_18826);
nor U21452 (N_21452,N_18313,N_17863);
or U21453 (N_21453,N_18911,N_19853);
and U21454 (N_21454,N_18606,N_19997);
xnor U21455 (N_21455,N_19452,N_18504);
or U21456 (N_21456,N_18459,N_17708);
xnor U21457 (N_21457,N_19862,N_17847);
and U21458 (N_21458,N_19621,N_18147);
xnor U21459 (N_21459,N_18067,N_19625);
or U21460 (N_21460,N_18039,N_18173);
nor U21461 (N_21461,N_17536,N_18760);
and U21462 (N_21462,N_19097,N_19738);
nor U21463 (N_21463,N_18353,N_18097);
or U21464 (N_21464,N_19981,N_17588);
or U21465 (N_21465,N_19673,N_19753);
nor U21466 (N_21466,N_19669,N_18704);
nor U21467 (N_21467,N_19825,N_18156);
xnor U21468 (N_21468,N_19004,N_19663);
or U21469 (N_21469,N_17603,N_19329);
or U21470 (N_21470,N_19832,N_19585);
xor U21471 (N_21471,N_17612,N_18839);
nand U21472 (N_21472,N_19546,N_17623);
nand U21473 (N_21473,N_17769,N_18511);
xnor U21474 (N_21474,N_17659,N_18904);
xnor U21475 (N_21475,N_18829,N_17810);
or U21476 (N_21476,N_19184,N_18444);
and U21477 (N_21477,N_19661,N_19295);
nor U21478 (N_21478,N_18434,N_19228);
nor U21479 (N_21479,N_17746,N_19440);
nor U21480 (N_21480,N_17915,N_19678);
and U21481 (N_21481,N_17754,N_17734);
or U21482 (N_21482,N_17828,N_19833);
and U21483 (N_21483,N_17933,N_19084);
and U21484 (N_21484,N_18852,N_18613);
and U21485 (N_21485,N_18905,N_18244);
nor U21486 (N_21486,N_17633,N_19592);
xnor U21487 (N_21487,N_18092,N_18659);
nand U21488 (N_21488,N_18000,N_19982);
or U21489 (N_21489,N_19676,N_19578);
nor U21490 (N_21490,N_18109,N_18852);
xor U21491 (N_21491,N_18936,N_18520);
xor U21492 (N_21492,N_19066,N_19582);
nand U21493 (N_21493,N_19568,N_19372);
nand U21494 (N_21494,N_18556,N_17775);
nand U21495 (N_21495,N_17616,N_17953);
nand U21496 (N_21496,N_18905,N_19814);
and U21497 (N_21497,N_18814,N_18117);
xor U21498 (N_21498,N_18587,N_18718);
xor U21499 (N_21499,N_17740,N_19195);
and U21500 (N_21500,N_18533,N_19516);
xor U21501 (N_21501,N_18407,N_17779);
and U21502 (N_21502,N_19504,N_19878);
xnor U21503 (N_21503,N_19403,N_17797);
or U21504 (N_21504,N_19128,N_18742);
xor U21505 (N_21505,N_18676,N_17912);
and U21506 (N_21506,N_17521,N_19566);
or U21507 (N_21507,N_18411,N_19361);
nand U21508 (N_21508,N_18329,N_17970);
and U21509 (N_21509,N_19529,N_19406);
and U21510 (N_21510,N_19467,N_18483);
xnor U21511 (N_21511,N_18688,N_19356);
and U21512 (N_21512,N_18950,N_19373);
and U21513 (N_21513,N_17738,N_19026);
nor U21514 (N_21514,N_18617,N_18093);
nand U21515 (N_21515,N_17756,N_19147);
xor U21516 (N_21516,N_19634,N_19926);
nand U21517 (N_21517,N_19762,N_19701);
nand U21518 (N_21518,N_18469,N_19331);
or U21519 (N_21519,N_18579,N_18299);
xor U21520 (N_21520,N_17595,N_19198);
or U21521 (N_21521,N_19687,N_17729);
nand U21522 (N_21522,N_19749,N_17871);
nor U21523 (N_21523,N_19167,N_19451);
or U21524 (N_21524,N_17685,N_19429);
or U21525 (N_21525,N_19683,N_17963);
nand U21526 (N_21526,N_18584,N_18259);
and U21527 (N_21527,N_18094,N_19159);
or U21528 (N_21528,N_19407,N_17753);
xor U21529 (N_21529,N_18325,N_17543);
nor U21530 (N_21530,N_19276,N_18570);
or U21531 (N_21531,N_18215,N_17518);
nand U21532 (N_21532,N_18382,N_19979);
nor U21533 (N_21533,N_18710,N_19314);
nand U21534 (N_21534,N_18214,N_19297);
or U21535 (N_21535,N_19477,N_18524);
or U21536 (N_21536,N_19510,N_19016);
nand U21537 (N_21537,N_17660,N_18077);
or U21538 (N_21538,N_18083,N_18591);
xor U21539 (N_21539,N_18937,N_19204);
and U21540 (N_21540,N_19635,N_17737);
xnor U21541 (N_21541,N_19905,N_19584);
or U21542 (N_21542,N_19556,N_18496);
xnor U21543 (N_21543,N_18444,N_19533);
nor U21544 (N_21544,N_19374,N_18637);
nor U21545 (N_21545,N_18909,N_17614);
or U21546 (N_21546,N_19980,N_19431);
or U21547 (N_21547,N_18481,N_19466);
xor U21548 (N_21548,N_18486,N_17748);
and U21549 (N_21549,N_17705,N_18246);
nand U21550 (N_21550,N_19177,N_18178);
nor U21551 (N_21551,N_19220,N_18551);
nand U21552 (N_21552,N_17566,N_18683);
nor U21553 (N_21553,N_18770,N_19228);
nor U21554 (N_21554,N_19742,N_17900);
and U21555 (N_21555,N_17560,N_19141);
and U21556 (N_21556,N_19056,N_19233);
nand U21557 (N_21557,N_19277,N_19623);
xnor U21558 (N_21558,N_17939,N_19585);
or U21559 (N_21559,N_18281,N_18104);
nor U21560 (N_21560,N_18163,N_18416);
nor U21561 (N_21561,N_19111,N_17931);
or U21562 (N_21562,N_18819,N_19713);
nor U21563 (N_21563,N_19677,N_18608);
and U21564 (N_21564,N_17559,N_17896);
nor U21565 (N_21565,N_18837,N_18781);
nand U21566 (N_21566,N_19053,N_19801);
xor U21567 (N_21567,N_18808,N_19867);
nor U21568 (N_21568,N_17800,N_19987);
xor U21569 (N_21569,N_19099,N_18050);
nor U21570 (N_21570,N_19099,N_18596);
nor U21571 (N_21571,N_18660,N_17693);
and U21572 (N_21572,N_19426,N_19239);
and U21573 (N_21573,N_18053,N_19070);
nor U21574 (N_21574,N_17703,N_18291);
or U21575 (N_21575,N_18902,N_18379);
xnor U21576 (N_21576,N_18786,N_18894);
xor U21577 (N_21577,N_18082,N_19977);
xnor U21578 (N_21578,N_18525,N_18631);
xnor U21579 (N_21579,N_19767,N_18825);
and U21580 (N_21580,N_19373,N_18904);
xnor U21581 (N_21581,N_18880,N_18663);
nand U21582 (N_21582,N_18918,N_19722);
and U21583 (N_21583,N_18785,N_19164);
and U21584 (N_21584,N_18649,N_17644);
and U21585 (N_21585,N_17687,N_18799);
or U21586 (N_21586,N_18630,N_19319);
and U21587 (N_21587,N_19725,N_19835);
and U21588 (N_21588,N_19399,N_19440);
nor U21589 (N_21589,N_18912,N_17741);
and U21590 (N_21590,N_19888,N_17822);
or U21591 (N_21591,N_19952,N_18711);
nor U21592 (N_21592,N_18008,N_19789);
nand U21593 (N_21593,N_18122,N_18501);
and U21594 (N_21594,N_18772,N_18453);
or U21595 (N_21595,N_17966,N_19409);
xnor U21596 (N_21596,N_19516,N_18975);
nor U21597 (N_21597,N_19629,N_18013);
nand U21598 (N_21598,N_19077,N_18373);
or U21599 (N_21599,N_19300,N_19168);
and U21600 (N_21600,N_18992,N_17798);
or U21601 (N_21601,N_19496,N_18665);
nor U21602 (N_21602,N_19608,N_19477);
or U21603 (N_21603,N_19601,N_18639);
nand U21604 (N_21604,N_19853,N_17631);
or U21605 (N_21605,N_18969,N_18454);
and U21606 (N_21606,N_18795,N_19137);
or U21607 (N_21607,N_18393,N_19953);
or U21608 (N_21608,N_17735,N_18355);
and U21609 (N_21609,N_19453,N_19251);
or U21610 (N_21610,N_18361,N_18402);
or U21611 (N_21611,N_17662,N_18925);
nor U21612 (N_21612,N_18900,N_19408);
or U21613 (N_21613,N_17554,N_18548);
and U21614 (N_21614,N_19285,N_19682);
and U21615 (N_21615,N_17763,N_19760);
and U21616 (N_21616,N_18752,N_19513);
xnor U21617 (N_21617,N_17761,N_19357);
nor U21618 (N_21618,N_19261,N_18376);
xor U21619 (N_21619,N_19823,N_18528);
nor U21620 (N_21620,N_19141,N_19059);
and U21621 (N_21621,N_19574,N_19270);
xor U21622 (N_21622,N_18851,N_18792);
or U21623 (N_21623,N_19898,N_17942);
or U21624 (N_21624,N_19307,N_18528);
or U21625 (N_21625,N_17547,N_19040);
and U21626 (N_21626,N_18567,N_18833);
or U21627 (N_21627,N_19332,N_19218);
nor U21628 (N_21628,N_19528,N_17876);
and U21629 (N_21629,N_19194,N_19652);
nor U21630 (N_21630,N_19283,N_18059);
or U21631 (N_21631,N_18597,N_17688);
nand U21632 (N_21632,N_17749,N_19381);
or U21633 (N_21633,N_19468,N_17833);
or U21634 (N_21634,N_18738,N_19809);
nand U21635 (N_21635,N_18336,N_17944);
or U21636 (N_21636,N_17756,N_18003);
or U21637 (N_21637,N_19622,N_17907);
nor U21638 (N_21638,N_19869,N_19664);
xor U21639 (N_21639,N_18122,N_18552);
and U21640 (N_21640,N_19324,N_18818);
xnor U21641 (N_21641,N_17783,N_18773);
xnor U21642 (N_21642,N_19835,N_18361);
and U21643 (N_21643,N_19008,N_19162);
or U21644 (N_21644,N_19890,N_17533);
nor U21645 (N_21645,N_19148,N_17839);
and U21646 (N_21646,N_19265,N_17895);
and U21647 (N_21647,N_18917,N_18771);
nand U21648 (N_21648,N_19656,N_19544);
and U21649 (N_21649,N_19959,N_18003);
xnor U21650 (N_21650,N_19108,N_19802);
or U21651 (N_21651,N_19463,N_18089);
and U21652 (N_21652,N_17758,N_18664);
nand U21653 (N_21653,N_18593,N_19425);
xor U21654 (N_21654,N_18706,N_17750);
and U21655 (N_21655,N_17885,N_18921);
xor U21656 (N_21656,N_17645,N_19987);
nand U21657 (N_21657,N_19276,N_18210);
nor U21658 (N_21658,N_19349,N_18230);
xnor U21659 (N_21659,N_18744,N_19219);
and U21660 (N_21660,N_18204,N_18331);
or U21661 (N_21661,N_18850,N_19827);
or U21662 (N_21662,N_18229,N_19951);
nand U21663 (N_21663,N_17977,N_19848);
or U21664 (N_21664,N_19984,N_18102);
xnor U21665 (N_21665,N_17938,N_18569);
and U21666 (N_21666,N_18384,N_19287);
and U21667 (N_21667,N_17963,N_18545);
nand U21668 (N_21668,N_19239,N_19616);
or U21669 (N_21669,N_19378,N_18827);
nor U21670 (N_21670,N_18691,N_18967);
or U21671 (N_21671,N_18584,N_19517);
xnor U21672 (N_21672,N_17915,N_18018);
nand U21673 (N_21673,N_18378,N_19793);
nor U21674 (N_21674,N_19982,N_18165);
xor U21675 (N_21675,N_18624,N_19815);
xnor U21676 (N_21676,N_18885,N_19633);
and U21677 (N_21677,N_17754,N_19210);
and U21678 (N_21678,N_18937,N_17900);
nand U21679 (N_21679,N_19826,N_17941);
and U21680 (N_21680,N_19007,N_19486);
and U21681 (N_21681,N_18912,N_19665);
xnor U21682 (N_21682,N_17869,N_19081);
or U21683 (N_21683,N_18116,N_18949);
nor U21684 (N_21684,N_17528,N_19336);
nand U21685 (N_21685,N_18890,N_18245);
and U21686 (N_21686,N_18216,N_18314);
and U21687 (N_21687,N_19592,N_17769);
and U21688 (N_21688,N_17654,N_19562);
nor U21689 (N_21689,N_18726,N_18724);
or U21690 (N_21690,N_19438,N_18821);
or U21691 (N_21691,N_17731,N_19873);
xor U21692 (N_21692,N_18830,N_18194);
or U21693 (N_21693,N_19002,N_18763);
nor U21694 (N_21694,N_17784,N_19906);
xnor U21695 (N_21695,N_18910,N_19152);
or U21696 (N_21696,N_19966,N_19416);
and U21697 (N_21697,N_18993,N_19233);
and U21698 (N_21698,N_18143,N_19234);
or U21699 (N_21699,N_19508,N_19931);
nor U21700 (N_21700,N_18036,N_17895);
xor U21701 (N_21701,N_18579,N_18407);
and U21702 (N_21702,N_18133,N_18898);
xor U21703 (N_21703,N_19470,N_19562);
nand U21704 (N_21704,N_17557,N_19675);
or U21705 (N_21705,N_19301,N_17705);
xor U21706 (N_21706,N_17663,N_18634);
and U21707 (N_21707,N_17673,N_18633);
or U21708 (N_21708,N_18174,N_18180);
and U21709 (N_21709,N_18480,N_18819);
or U21710 (N_21710,N_19216,N_17642);
nand U21711 (N_21711,N_17556,N_17824);
and U21712 (N_21712,N_18615,N_19145);
nor U21713 (N_21713,N_19042,N_18116);
or U21714 (N_21714,N_19237,N_18578);
and U21715 (N_21715,N_17500,N_18185);
nor U21716 (N_21716,N_18018,N_18472);
and U21717 (N_21717,N_18662,N_18279);
or U21718 (N_21718,N_18992,N_19269);
nor U21719 (N_21719,N_17601,N_19215);
nand U21720 (N_21720,N_18880,N_18600);
nand U21721 (N_21721,N_18203,N_18458);
and U21722 (N_21722,N_19117,N_19820);
nor U21723 (N_21723,N_18467,N_18155);
and U21724 (N_21724,N_19548,N_19428);
nand U21725 (N_21725,N_18316,N_18656);
or U21726 (N_21726,N_18638,N_19292);
nand U21727 (N_21727,N_17697,N_18688);
xor U21728 (N_21728,N_18734,N_17878);
nor U21729 (N_21729,N_18503,N_19294);
nand U21730 (N_21730,N_18606,N_18437);
xnor U21731 (N_21731,N_19647,N_18012);
and U21732 (N_21732,N_18951,N_18764);
and U21733 (N_21733,N_19550,N_17827);
xor U21734 (N_21734,N_18693,N_17687);
xor U21735 (N_21735,N_19134,N_19756);
nand U21736 (N_21736,N_18344,N_19106);
nand U21737 (N_21737,N_19051,N_17785);
nor U21738 (N_21738,N_18435,N_17504);
nand U21739 (N_21739,N_18998,N_19590);
and U21740 (N_21740,N_18789,N_17739);
nor U21741 (N_21741,N_19341,N_19840);
or U21742 (N_21742,N_18370,N_18146);
and U21743 (N_21743,N_17865,N_18744);
nand U21744 (N_21744,N_19794,N_19353);
xor U21745 (N_21745,N_19621,N_18174);
or U21746 (N_21746,N_18636,N_18834);
and U21747 (N_21747,N_19908,N_18370);
and U21748 (N_21748,N_18175,N_17822);
and U21749 (N_21749,N_18246,N_17647);
nor U21750 (N_21750,N_17679,N_19715);
or U21751 (N_21751,N_19874,N_19432);
nand U21752 (N_21752,N_19981,N_17561);
nor U21753 (N_21753,N_19781,N_17961);
nor U21754 (N_21754,N_19480,N_19849);
nand U21755 (N_21755,N_18557,N_19549);
nand U21756 (N_21756,N_19719,N_19811);
and U21757 (N_21757,N_18052,N_18530);
xnor U21758 (N_21758,N_19440,N_19401);
nand U21759 (N_21759,N_17848,N_19919);
xnor U21760 (N_21760,N_18294,N_19799);
nand U21761 (N_21761,N_19705,N_18319);
and U21762 (N_21762,N_19143,N_18972);
and U21763 (N_21763,N_17661,N_19432);
or U21764 (N_21764,N_17557,N_19992);
and U21765 (N_21765,N_19043,N_18805);
and U21766 (N_21766,N_19208,N_19348);
or U21767 (N_21767,N_17607,N_19504);
or U21768 (N_21768,N_18280,N_19491);
xor U21769 (N_21769,N_18616,N_19967);
nor U21770 (N_21770,N_18313,N_17667);
xor U21771 (N_21771,N_19544,N_19573);
nand U21772 (N_21772,N_18052,N_19288);
xnor U21773 (N_21773,N_19051,N_17643);
nor U21774 (N_21774,N_19916,N_19909);
xnor U21775 (N_21775,N_19094,N_19998);
and U21776 (N_21776,N_17844,N_17849);
and U21777 (N_21777,N_18161,N_18319);
or U21778 (N_21778,N_18031,N_17592);
nand U21779 (N_21779,N_19277,N_17884);
xor U21780 (N_21780,N_17714,N_18455);
xor U21781 (N_21781,N_19003,N_17792);
and U21782 (N_21782,N_18658,N_18182);
or U21783 (N_21783,N_17779,N_18836);
nand U21784 (N_21784,N_17633,N_17814);
and U21785 (N_21785,N_18683,N_18050);
and U21786 (N_21786,N_18084,N_19118);
nor U21787 (N_21787,N_19982,N_17599);
xnor U21788 (N_21788,N_19834,N_19052);
xnor U21789 (N_21789,N_19604,N_17912);
xnor U21790 (N_21790,N_19455,N_18894);
nand U21791 (N_21791,N_17604,N_18095);
and U21792 (N_21792,N_18470,N_19778);
nand U21793 (N_21793,N_17679,N_18218);
or U21794 (N_21794,N_19843,N_18042);
or U21795 (N_21795,N_19170,N_18054);
nand U21796 (N_21796,N_17656,N_17684);
and U21797 (N_21797,N_18854,N_18148);
nor U21798 (N_21798,N_17586,N_18630);
xnor U21799 (N_21799,N_17677,N_18049);
nand U21800 (N_21800,N_18761,N_18986);
and U21801 (N_21801,N_19075,N_18161);
nand U21802 (N_21802,N_18166,N_19923);
nor U21803 (N_21803,N_18438,N_19070);
or U21804 (N_21804,N_19809,N_17927);
nand U21805 (N_21805,N_19536,N_18791);
nor U21806 (N_21806,N_19898,N_19292);
nor U21807 (N_21807,N_18794,N_18847);
or U21808 (N_21808,N_19444,N_19799);
xor U21809 (N_21809,N_18553,N_19783);
and U21810 (N_21810,N_19081,N_19843);
xor U21811 (N_21811,N_19807,N_18217);
or U21812 (N_21812,N_19191,N_18272);
xnor U21813 (N_21813,N_18612,N_19105);
or U21814 (N_21814,N_18778,N_19895);
nor U21815 (N_21815,N_17937,N_17690);
and U21816 (N_21816,N_17546,N_19650);
and U21817 (N_21817,N_18336,N_19753);
xor U21818 (N_21818,N_17592,N_18437);
or U21819 (N_21819,N_18283,N_19200);
and U21820 (N_21820,N_18248,N_19725);
and U21821 (N_21821,N_19857,N_19336);
xor U21822 (N_21822,N_17859,N_19849);
nand U21823 (N_21823,N_18469,N_18473);
nand U21824 (N_21824,N_18125,N_18133);
xnor U21825 (N_21825,N_18297,N_19498);
nor U21826 (N_21826,N_18487,N_18154);
nor U21827 (N_21827,N_18002,N_18251);
nand U21828 (N_21828,N_18435,N_19930);
or U21829 (N_21829,N_18244,N_18953);
or U21830 (N_21830,N_18623,N_19600);
nor U21831 (N_21831,N_17624,N_19428);
nor U21832 (N_21832,N_17621,N_18148);
or U21833 (N_21833,N_17556,N_19529);
or U21834 (N_21834,N_17649,N_19061);
xnor U21835 (N_21835,N_18842,N_19072);
nand U21836 (N_21836,N_18096,N_17997);
nor U21837 (N_21837,N_19226,N_17592);
xnor U21838 (N_21838,N_17500,N_18930);
nor U21839 (N_21839,N_18890,N_19185);
nor U21840 (N_21840,N_18468,N_18128);
or U21841 (N_21841,N_18077,N_18564);
or U21842 (N_21842,N_18478,N_18912);
xnor U21843 (N_21843,N_17977,N_18601);
nand U21844 (N_21844,N_17649,N_17860);
and U21845 (N_21845,N_18761,N_19015);
nor U21846 (N_21846,N_18319,N_19741);
xnor U21847 (N_21847,N_18488,N_18806);
and U21848 (N_21848,N_19747,N_18635);
nand U21849 (N_21849,N_18156,N_18742);
xor U21850 (N_21850,N_18155,N_19926);
nand U21851 (N_21851,N_19149,N_18974);
xor U21852 (N_21852,N_18818,N_18261);
or U21853 (N_21853,N_17985,N_18717);
nor U21854 (N_21854,N_19025,N_19330);
nand U21855 (N_21855,N_19292,N_19154);
and U21856 (N_21856,N_19535,N_17675);
nand U21857 (N_21857,N_18035,N_18071);
and U21858 (N_21858,N_19554,N_19561);
nand U21859 (N_21859,N_19032,N_18817);
and U21860 (N_21860,N_19936,N_18809);
xor U21861 (N_21861,N_17937,N_18834);
and U21862 (N_21862,N_17979,N_17840);
nor U21863 (N_21863,N_18185,N_19304);
or U21864 (N_21864,N_18569,N_19636);
or U21865 (N_21865,N_17648,N_19562);
xor U21866 (N_21866,N_17743,N_17858);
or U21867 (N_21867,N_18966,N_19242);
xor U21868 (N_21868,N_18259,N_17845);
or U21869 (N_21869,N_19128,N_19460);
and U21870 (N_21870,N_19355,N_19375);
or U21871 (N_21871,N_19436,N_18371);
and U21872 (N_21872,N_18553,N_19265);
nor U21873 (N_21873,N_19981,N_17854);
or U21874 (N_21874,N_17585,N_18322);
xnor U21875 (N_21875,N_19068,N_18770);
and U21876 (N_21876,N_18395,N_18885);
nand U21877 (N_21877,N_18374,N_19377);
xor U21878 (N_21878,N_18429,N_18537);
xor U21879 (N_21879,N_18194,N_18746);
nor U21880 (N_21880,N_17935,N_18963);
and U21881 (N_21881,N_18042,N_18729);
xnor U21882 (N_21882,N_19427,N_19040);
and U21883 (N_21883,N_18786,N_19470);
and U21884 (N_21884,N_18710,N_18453);
and U21885 (N_21885,N_18689,N_17597);
nor U21886 (N_21886,N_18331,N_19434);
xor U21887 (N_21887,N_18232,N_19384);
nand U21888 (N_21888,N_17593,N_19651);
xnor U21889 (N_21889,N_18401,N_17836);
xor U21890 (N_21890,N_18009,N_19796);
and U21891 (N_21891,N_19766,N_19521);
nand U21892 (N_21892,N_17536,N_19393);
nor U21893 (N_21893,N_17630,N_18917);
and U21894 (N_21894,N_18167,N_18797);
or U21895 (N_21895,N_18474,N_18306);
and U21896 (N_21896,N_19054,N_18988);
xor U21897 (N_21897,N_19151,N_19902);
nor U21898 (N_21898,N_19133,N_17872);
nor U21899 (N_21899,N_18948,N_19880);
nand U21900 (N_21900,N_17504,N_18754);
and U21901 (N_21901,N_19673,N_17733);
xor U21902 (N_21902,N_19740,N_17527);
nor U21903 (N_21903,N_19320,N_18038);
nor U21904 (N_21904,N_19566,N_19199);
nand U21905 (N_21905,N_17614,N_19156);
nand U21906 (N_21906,N_18520,N_18621);
or U21907 (N_21907,N_17745,N_19898);
nand U21908 (N_21908,N_19128,N_19750);
nor U21909 (N_21909,N_19213,N_19900);
nand U21910 (N_21910,N_18524,N_17632);
nor U21911 (N_21911,N_18794,N_19976);
nor U21912 (N_21912,N_18042,N_19961);
or U21913 (N_21913,N_17919,N_18136);
xnor U21914 (N_21914,N_18479,N_19827);
xnor U21915 (N_21915,N_19124,N_19780);
nand U21916 (N_21916,N_19785,N_17734);
nand U21917 (N_21917,N_19241,N_19914);
nand U21918 (N_21918,N_17751,N_18192);
or U21919 (N_21919,N_18167,N_18192);
xnor U21920 (N_21920,N_17972,N_18301);
nand U21921 (N_21921,N_19789,N_18359);
xnor U21922 (N_21922,N_18595,N_19506);
xor U21923 (N_21923,N_18514,N_19524);
nand U21924 (N_21924,N_18081,N_19579);
nand U21925 (N_21925,N_19512,N_19793);
and U21926 (N_21926,N_17669,N_18566);
nor U21927 (N_21927,N_19516,N_19447);
and U21928 (N_21928,N_19635,N_19289);
or U21929 (N_21929,N_18580,N_19272);
xnor U21930 (N_21930,N_18741,N_18319);
xnor U21931 (N_21931,N_19897,N_17757);
nand U21932 (N_21932,N_19753,N_17739);
nor U21933 (N_21933,N_18070,N_19016);
nor U21934 (N_21934,N_19837,N_17766);
xor U21935 (N_21935,N_19632,N_17749);
or U21936 (N_21936,N_19236,N_19971);
or U21937 (N_21937,N_19973,N_19798);
or U21938 (N_21938,N_19629,N_18304);
nor U21939 (N_21939,N_19058,N_18164);
and U21940 (N_21940,N_19915,N_19925);
and U21941 (N_21941,N_17516,N_18796);
or U21942 (N_21942,N_19692,N_18288);
xnor U21943 (N_21943,N_17651,N_18401);
nor U21944 (N_21944,N_18137,N_18122);
or U21945 (N_21945,N_19836,N_19521);
nand U21946 (N_21946,N_18296,N_18641);
xnor U21947 (N_21947,N_19710,N_17867);
nor U21948 (N_21948,N_19144,N_19614);
xor U21949 (N_21949,N_18450,N_19674);
and U21950 (N_21950,N_17537,N_18521);
or U21951 (N_21951,N_17565,N_19978);
or U21952 (N_21952,N_17806,N_19263);
or U21953 (N_21953,N_19559,N_18360);
nor U21954 (N_21954,N_18245,N_19301);
nand U21955 (N_21955,N_19935,N_18096);
nor U21956 (N_21956,N_18627,N_18363);
nor U21957 (N_21957,N_19978,N_17530);
or U21958 (N_21958,N_18634,N_18455);
and U21959 (N_21959,N_18329,N_18984);
nand U21960 (N_21960,N_19733,N_18573);
nor U21961 (N_21961,N_18998,N_18087);
and U21962 (N_21962,N_18479,N_18440);
and U21963 (N_21963,N_19713,N_18744);
nand U21964 (N_21964,N_18014,N_17988);
xnor U21965 (N_21965,N_19875,N_17556);
nor U21966 (N_21966,N_18366,N_17801);
or U21967 (N_21967,N_18341,N_19164);
nand U21968 (N_21968,N_17666,N_19934);
or U21969 (N_21969,N_18008,N_17868);
and U21970 (N_21970,N_18694,N_19010);
nor U21971 (N_21971,N_17625,N_18544);
and U21972 (N_21972,N_18246,N_19413);
nand U21973 (N_21973,N_18348,N_18559);
xor U21974 (N_21974,N_17532,N_19158);
nor U21975 (N_21975,N_17815,N_19869);
nor U21976 (N_21976,N_19556,N_18767);
xor U21977 (N_21977,N_17623,N_19773);
nor U21978 (N_21978,N_18449,N_19004);
xor U21979 (N_21979,N_18638,N_19309);
nand U21980 (N_21980,N_19051,N_19771);
nand U21981 (N_21981,N_19681,N_17926);
nand U21982 (N_21982,N_18778,N_19067);
nand U21983 (N_21983,N_19140,N_18160);
nor U21984 (N_21984,N_17843,N_17603);
xor U21985 (N_21985,N_19743,N_18776);
or U21986 (N_21986,N_17778,N_17698);
nand U21987 (N_21987,N_19190,N_18495);
nor U21988 (N_21988,N_19924,N_17635);
and U21989 (N_21989,N_19692,N_19552);
nor U21990 (N_21990,N_17811,N_18030);
nand U21991 (N_21991,N_18938,N_18428);
nor U21992 (N_21992,N_19127,N_19860);
nor U21993 (N_21993,N_18586,N_17767);
and U21994 (N_21994,N_19018,N_19492);
and U21995 (N_21995,N_19939,N_18079);
nor U21996 (N_21996,N_17949,N_17669);
nand U21997 (N_21997,N_17704,N_19088);
nor U21998 (N_21998,N_19295,N_18897);
nor U21999 (N_21999,N_18521,N_19496);
nand U22000 (N_22000,N_18561,N_18509);
and U22001 (N_22001,N_19941,N_19632);
nor U22002 (N_22002,N_19602,N_19813);
and U22003 (N_22003,N_18883,N_18323);
nor U22004 (N_22004,N_18275,N_18100);
and U22005 (N_22005,N_18188,N_19759);
nand U22006 (N_22006,N_18030,N_17791);
and U22007 (N_22007,N_18095,N_18483);
and U22008 (N_22008,N_17861,N_18196);
xor U22009 (N_22009,N_19890,N_17586);
xnor U22010 (N_22010,N_19529,N_19460);
or U22011 (N_22011,N_19718,N_19499);
nand U22012 (N_22012,N_19265,N_19706);
and U22013 (N_22013,N_18436,N_19553);
nor U22014 (N_22014,N_18855,N_18391);
nor U22015 (N_22015,N_18255,N_19397);
or U22016 (N_22016,N_17559,N_19751);
and U22017 (N_22017,N_17772,N_17754);
xor U22018 (N_22018,N_17590,N_18421);
nor U22019 (N_22019,N_19492,N_18010);
and U22020 (N_22020,N_18396,N_17692);
and U22021 (N_22021,N_19057,N_18215);
nand U22022 (N_22022,N_19441,N_18327);
and U22023 (N_22023,N_17658,N_19059);
nand U22024 (N_22024,N_19148,N_19752);
nor U22025 (N_22025,N_18883,N_19777);
and U22026 (N_22026,N_18128,N_17614);
and U22027 (N_22027,N_18491,N_17847);
xnor U22028 (N_22028,N_18492,N_19660);
nand U22029 (N_22029,N_19684,N_19688);
and U22030 (N_22030,N_18093,N_17604);
and U22031 (N_22031,N_19956,N_18529);
nand U22032 (N_22032,N_19586,N_19031);
nor U22033 (N_22033,N_19467,N_19894);
nand U22034 (N_22034,N_17976,N_18365);
and U22035 (N_22035,N_19780,N_19214);
and U22036 (N_22036,N_18610,N_19315);
nor U22037 (N_22037,N_19788,N_18133);
xor U22038 (N_22038,N_18341,N_17842);
and U22039 (N_22039,N_19450,N_18040);
nor U22040 (N_22040,N_17737,N_19443);
nor U22041 (N_22041,N_19143,N_19098);
xor U22042 (N_22042,N_18874,N_17863);
nor U22043 (N_22043,N_18718,N_18923);
nand U22044 (N_22044,N_19056,N_17952);
nand U22045 (N_22045,N_19096,N_17793);
nand U22046 (N_22046,N_19465,N_18944);
and U22047 (N_22047,N_18022,N_19959);
xor U22048 (N_22048,N_18198,N_17973);
and U22049 (N_22049,N_19134,N_19346);
xor U22050 (N_22050,N_18111,N_18558);
nor U22051 (N_22051,N_18539,N_17945);
or U22052 (N_22052,N_19597,N_19852);
nand U22053 (N_22053,N_19767,N_17885);
and U22054 (N_22054,N_17612,N_18019);
nor U22055 (N_22055,N_17882,N_19892);
and U22056 (N_22056,N_19253,N_19841);
or U22057 (N_22057,N_17711,N_18535);
and U22058 (N_22058,N_18448,N_18853);
nand U22059 (N_22059,N_18559,N_19525);
and U22060 (N_22060,N_19544,N_19170);
nand U22061 (N_22061,N_17857,N_18141);
and U22062 (N_22062,N_19541,N_19809);
nor U22063 (N_22063,N_17622,N_17562);
nand U22064 (N_22064,N_18663,N_19773);
or U22065 (N_22065,N_17819,N_18219);
and U22066 (N_22066,N_18811,N_18240);
and U22067 (N_22067,N_18407,N_19370);
xor U22068 (N_22068,N_18843,N_18035);
xor U22069 (N_22069,N_17605,N_18683);
or U22070 (N_22070,N_19035,N_18004);
nand U22071 (N_22071,N_17806,N_18970);
xnor U22072 (N_22072,N_17861,N_19190);
nor U22073 (N_22073,N_17687,N_18118);
or U22074 (N_22074,N_19099,N_18210);
nand U22075 (N_22075,N_17528,N_19672);
nand U22076 (N_22076,N_19240,N_18535);
nor U22077 (N_22077,N_18136,N_19856);
nand U22078 (N_22078,N_17685,N_17960);
and U22079 (N_22079,N_19113,N_17955);
nand U22080 (N_22080,N_18840,N_18948);
or U22081 (N_22081,N_18742,N_19390);
and U22082 (N_22082,N_18660,N_19801);
and U22083 (N_22083,N_19036,N_19451);
nor U22084 (N_22084,N_17931,N_19089);
and U22085 (N_22085,N_18514,N_19762);
and U22086 (N_22086,N_19774,N_19797);
xor U22087 (N_22087,N_18748,N_19010);
and U22088 (N_22088,N_18993,N_17846);
xor U22089 (N_22089,N_18700,N_18055);
nand U22090 (N_22090,N_19237,N_18991);
nor U22091 (N_22091,N_18120,N_18630);
nor U22092 (N_22092,N_18111,N_19669);
and U22093 (N_22093,N_17590,N_19996);
nor U22094 (N_22094,N_19089,N_19078);
or U22095 (N_22095,N_19199,N_19218);
xor U22096 (N_22096,N_17975,N_17928);
or U22097 (N_22097,N_18248,N_19704);
xnor U22098 (N_22098,N_17732,N_19000);
nand U22099 (N_22099,N_19976,N_18009);
xor U22100 (N_22100,N_18652,N_19020);
nand U22101 (N_22101,N_18273,N_19536);
nor U22102 (N_22102,N_17917,N_19178);
xor U22103 (N_22103,N_19360,N_19112);
and U22104 (N_22104,N_17765,N_17592);
or U22105 (N_22105,N_17931,N_19153);
and U22106 (N_22106,N_19388,N_18189);
or U22107 (N_22107,N_18651,N_18385);
nor U22108 (N_22108,N_19107,N_19193);
xor U22109 (N_22109,N_19468,N_18142);
or U22110 (N_22110,N_18597,N_19098);
or U22111 (N_22111,N_19111,N_19806);
nand U22112 (N_22112,N_17578,N_17758);
and U22113 (N_22113,N_19104,N_17959);
or U22114 (N_22114,N_19230,N_18848);
and U22115 (N_22115,N_18326,N_19156);
or U22116 (N_22116,N_18652,N_18889);
or U22117 (N_22117,N_19314,N_19626);
xnor U22118 (N_22118,N_19277,N_18072);
nand U22119 (N_22119,N_18402,N_18203);
nand U22120 (N_22120,N_17505,N_19894);
or U22121 (N_22121,N_19264,N_18432);
nand U22122 (N_22122,N_17542,N_17560);
nor U22123 (N_22123,N_19629,N_18183);
xnor U22124 (N_22124,N_19377,N_19147);
nand U22125 (N_22125,N_19300,N_18718);
or U22126 (N_22126,N_18491,N_18874);
nand U22127 (N_22127,N_19492,N_19694);
xnor U22128 (N_22128,N_18860,N_18313);
and U22129 (N_22129,N_19270,N_19806);
or U22130 (N_22130,N_17927,N_18705);
and U22131 (N_22131,N_19392,N_19166);
xnor U22132 (N_22132,N_18164,N_19519);
xor U22133 (N_22133,N_19489,N_19662);
and U22134 (N_22134,N_18582,N_18894);
and U22135 (N_22135,N_19910,N_18781);
or U22136 (N_22136,N_19771,N_19907);
and U22137 (N_22137,N_19915,N_18093);
and U22138 (N_22138,N_18673,N_17693);
and U22139 (N_22139,N_17727,N_19657);
or U22140 (N_22140,N_19721,N_18688);
or U22141 (N_22141,N_19856,N_19281);
nor U22142 (N_22142,N_18595,N_18538);
or U22143 (N_22143,N_19828,N_19238);
and U22144 (N_22144,N_17823,N_19867);
or U22145 (N_22145,N_18636,N_19567);
or U22146 (N_22146,N_19143,N_19722);
or U22147 (N_22147,N_19682,N_18751);
and U22148 (N_22148,N_19727,N_19455);
and U22149 (N_22149,N_19631,N_18264);
nand U22150 (N_22150,N_19243,N_19776);
nand U22151 (N_22151,N_18294,N_19073);
nor U22152 (N_22152,N_19704,N_19046);
nand U22153 (N_22153,N_18591,N_17742);
xor U22154 (N_22154,N_19546,N_19703);
nand U22155 (N_22155,N_18109,N_18547);
and U22156 (N_22156,N_17699,N_19881);
nor U22157 (N_22157,N_18864,N_17690);
nor U22158 (N_22158,N_19559,N_19923);
nor U22159 (N_22159,N_18047,N_18322);
nor U22160 (N_22160,N_19046,N_19467);
nor U22161 (N_22161,N_19832,N_18907);
xor U22162 (N_22162,N_17947,N_17797);
or U22163 (N_22163,N_17668,N_19942);
nor U22164 (N_22164,N_18305,N_19161);
xnor U22165 (N_22165,N_18722,N_18880);
and U22166 (N_22166,N_18102,N_19433);
and U22167 (N_22167,N_19162,N_18108);
or U22168 (N_22168,N_19974,N_19381);
and U22169 (N_22169,N_18853,N_17574);
xnor U22170 (N_22170,N_18351,N_17826);
and U22171 (N_22171,N_18871,N_19048);
and U22172 (N_22172,N_19008,N_18666);
xnor U22173 (N_22173,N_18753,N_18757);
nor U22174 (N_22174,N_19323,N_18688);
or U22175 (N_22175,N_18055,N_18404);
and U22176 (N_22176,N_19088,N_19011);
or U22177 (N_22177,N_18748,N_17882);
nand U22178 (N_22178,N_19097,N_18726);
or U22179 (N_22179,N_17966,N_19176);
and U22180 (N_22180,N_17868,N_19820);
xor U22181 (N_22181,N_19667,N_18555);
xnor U22182 (N_22182,N_17996,N_19620);
nor U22183 (N_22183,N_17546,N_17514);
nor U22184 (N_22184,N_19460,N_19936);
nand U22185 (N_22185,N_19920,N_19064);
xnor U22186 (N_22186,N_17985,N_19816);
nor U22187 (N_22187,N_19072,N_19038);
xor U22188 (N_22188,N_18583,N_18799);
nand U22189 (N_22189,N_17629,N_18226);
and U22190 (N_22190,N_17557,N_18234);
nor U22191 (N_22191,N_18961,N_19062);
and U22192 (N_22192,N_19508,N_19055);
or U22193 (N_22193,N_18650,N_19039);
or U22194 (N_22194,N_19700,N_19748);
nor U22195 (N_22195,N_19402,N_17529);
and U22196 (N_22196,N_19926,N_18566);
nor U22197 (N_22197,N_19189,N_19787);
and U22198 (N_22198,N_17542,N_18820);
or U22199 (N_22199,N_17579,N_19412);
nand U22200 (N_22200,N_19523,N_18153);
xor U22201 (N_22201,N_19123,N_19267);
nand U22202 (N_22202,N_19549,N_18987);
nor U22203 (N_22203,N_17964,N_19201);
or U22204 (N_22204,N_19991,N_19273);
xnor U22205 (N_22205,N_19372,N_17893);
nand U22206 (N_22206,N_19742,N_18770);
nand U22207 (N_22207,N_19582,N_19294);
or U22208 (N_22208,N_19098,N_18797);
and U22209 (N_22209,N_17505,N_19765);
nor U22210 (N_22210,N_19980,N_19624);
nand U22211 (N_22211,N_18088,N_18953);
or U22212 (N_22212,N_18047,N_19042);
nor U22213 (N_22213,N_18511,N_19735);
and U22214 (N_22214,N_17803,N_18240);
or U22215 (N_22215,N_18144,N_19477);
nor U22216 (N_22216,N_19227,N_19482);
or U22217 (N_22217,N_18794,N_19312);
xor U22218 (N_22218,N_17699,N_17957);
xnor U22219 (N_22219,N_19516,N_18072);
nor U22220 (N_22220,N_18494,N_18047);
xor U22221 (N_22221,N_17506,N_19590);
nor U22222 (N_22222,N_19151,N_19834);
xnor U22223 (N_22223,N_17957,N_17960);
nor U22224 (N_22224,N_19675,N_19022);
nand U22225 (N_22225,N_18586,N_17850);
nor U22226 (N_22226,N_19827,N_19955);
nor U22227 (N_22227,N_18024,N_17904);
and U22228 (N_22228,N_18547,N_19531);
nand U22229 (N_22229,N_19599,N_17933);
xor U22230 (N_22230,N_19171,N_17671);
nor U22231 (N_22231,N_17806,N_19195);
xor U22232 (N_22232,N_19184,N_18174);
or U22233 (N_22233,N_17504,N_19288);
nand U22234 (N_22234,N_19352,N_19840);
xor U22235 (N_22235,N_18561,N_17524);
and U22236 (N_22236,N_18035,N_19790);
and U22237 (N_22237,N_17675,N_18598);
nand U22238 (N_22238,N_18602,N_19687);
or U22239 (N_22239,N_17861,N_19325);
and U22240 (N_22240,N_19532,N_19071);
xnor U22241 (N_22241,N_18505,N_18038);
nor U22242 (N_22242,N_19432,N_18678);
and U22243 (N_22243,N_17722,N_18037);
xor U22244 (N_22244,N_19333,N_19790);
nand U22245 (N_22245,N_18672,N_18939);
nor U22246 (N_22246,N_18961,N_19940);
xor U22247 (N_22247,N_17660,N_17936);
or U22248 (N_22248,N_19244,N_19821);
and U22249 (N_22249,N_19216,N_18779);
or U22250 (N_22250,N_17933,N_18037);
and U22251 (N_22251,N_19040,N_19660);
nor U22252 (N_22252,N_17915,N_17607);
xnor U22253 (N_22253,N_17822,N_18147);
nor U22254 (N_22254,N_19116,N_19511);
nor U22255 (N_22255,N_18343,N_19450);
nor U22256 (N_22256,N_19838,N_18238);
xnor U22257 (N_22257,N_19034,N_18581);
nand U22258 (N_22258,N_19652,N_19240);
or U22259 (N_22259,N_18562,N_19528);
or U22260 (N_22260,N_18961,N_19846);
nand U22261 (N_22261,N_19095,N_19836);
xnor U22262 (N_22262,N_18647,N_19633);
or U22263 (N_22263,N_17560,N_19161);
nand U22264 (N_22264,N_19088,N_17711);
nor U22265 (N_22265,N_18447,N_19952);
nand U22266 (N_22266,N_19817,N_18046);
nand U22267 (N_22267,N_19309,N_19091);
nand U22268 (N_22268,N_19793,N_17857);
nand U22269 (N_22269,N_18305,N_19822);
nand U22270 (N_22270,N_19746,N_19241);
nand U22271 (N_22271,N_17560,N_18550);
and U22272 (N_22272,N_19616,N_18433);
xor U22273 (N_22273,N_19295,N_19191);
nand U22274 (N_22274,N_18252,N_18677);
and U22275 (N_22275,N_19636,N_18361);
nor U22276 (N_22276,N_17924,N_18404);
nor U22277 (N_22277,N_19358,N_18662);
nor U22278 (N_22278,N_19063,N_19560);
nand U22279 (N_22279,N_19099,N_17980);
or U22280 (N_22280,N_19141,N_18739);
or U22281 (N_22281,N_18525,N_17855);
or U22282 (N_22282,N_18743,N_18544);
xnor U22283 (N_22283,N_17824,N_18767);
xor U22284 (N_22284,N_17858,N_18244);
and U22285 (N_22285,N_18249,N_19359);
nand U22286 (N_22286,N_19956,N_17946);
and U22287 (N_22287,N_18679,N_18387);
xor U22288 (N_22288,N_19014,N_19345);
or U22289 (N_22289,N_18743,N_18982);
or U22290 (N_22290,N_17718,N_19837);
and U22291 (N_22291,N_18039,N_18847);
nor U22292 (N_22292,N_17796,N_19824);
xnor U22293 (N_22293,N_17566,N_18326);
nor U22294 (N_22294,N_18595,N_17684);
or U22295 (N_22295,N_18319,N_19176);
and U22296 (N_22296,N_19236,N_19231);
or U22297 (N_22297,N_17898,N_17923);
xnor U22298 (N_22298,N_18481,N_18839);
nor U22299 (N_22299,N_17839,N_19409);
and U22300 (N_22300,N_19293,N_19326);
nor U22301 (N_22301,N_17806,N_17513);
xor U22302 (N_22302,N_18529,N_17746);
xor U22303 (N_22303,N_17505,N_18611);
or U22304 (N_22304,N_17688,N_18661);
nor U22305 (N_22305,N_19240,N_18938);
and U22306 (N_22306,N_18280,N_19543);
xnor U22307 (N_22307,N_18366,N_18389);
nand U22308 (N_22308,N_17759,N_18099);
xnor U22309 (N_22309,N_18961,N_17921);
or U22310 (N_22310,N_18839,N_17649);
or U22311 (N_22311,N_17857,N_17784);
and U22312 (N_22312,N_19392,N_19792);
and U22313 (N_22313,N_18800,N_19112);
xnor U22314 (N_22314,N_18981,N_19238);
or U22315 (N_22315,N_18011,N_19673);
nand U22316 (N_22316,N_18723,N_18148);
nand U22317 (N_22317,N_17821,N_19797);
and U22318 (N_22318,N_18744,N_18986);
and U22319 (N_22319,N_18770,N_19602);
or U22320 (N_22320,N_17549,N_19226);
nand U22321 (N_22321,N_18150,N_19224);
nor U22322 (N_22322,N_19220,N_19538);
nor U22323 (N_22323,N_18999,N_17840);
or U22324 (N_22324,N_19994,N_18575);
nand U22325 (N_22325,N_19301,N_18554);
and U22326 (N_22326,N_19773,N_19473);
or U22327 (N_22327,N_19818,N_19560);
nor U22328 (N_22328,N_18872,N_19597);
nor U22329 (N_22329,N_18342,N_18861);
xnor U22330 (N_22330,N_19320,N_18413);
or U22331 (N_22331,N_18781,N_18765);
xor U22332 (N_22332,N_19627,N_19699);
nor U22333 (N_22333,N_19945,N_19454);
nor U22334 (N_22334,N_19701,N_17721);
xor U22335 (N_22335,N_18048,N_19645);
and U22336 (N_22336,N_17590,N_17604);
nor U22337 (N_22337,N_18188,N_18367);
or U22338 (N_22338,N_18889,N_17914);
xnor U22339 (N_22339,N_18669,N_17921);
nor U22340 (N_22340,N_19190,N_18168);
nor U22341 (N_22341,N_18325,N_18949);
nor U22342 (N_22342,N_17796,N_19535);
xor U22343 (N_22343,N_17511,N_17864);
and U22344 (N_22344,N_17557,N_18069);
and U22345 (N_22345,N_17554,N_18307);
nor U22346 (N_22346,N_19682,N_18680);
nand U22347 (N_22347,N_19388,N_19769);
nor U22348 (N_22348,N_17779,N_17618);
nor U22349 (N_22349,N_19576,N_18351);
or U22350 (N_22350,N_18055,N_18185);
and U22351 (N_22351,N_19236,N_19021);
nor U22352 (N_22352,N_19571,N_18386);
xnor U22353 (N_22353,N_18110,N_19966);
or U22354 (N_22354,N_19474,N_18641);
nor U22355 (N_22355,N_18820,N_18014);
or U22356 (N_22356,N_18677,N_18337);
or U22357 (N_22357,N_18347,N_18718);
nor U22358 (N_22358,N_19883,N_19843);
nand U22359 (N_22359,N_19300,N_19946);
and U22360 (N_22360,N_17894,N_17658);
nand U22361 (N_22361,N_18398,N_19550);
and U22362 (N_22362,N_19447,N_19438);
xnor U22363 (N_22363,N_17636,N_18241);
nor U22364 (N_22364,N_17927,N_17766);
nor U22365 (N_22365,N_19053,N_19717);
nor U22366 (N_22366,N_18743,N_18268);
nor U22367 (N_22367,N_18986,N_19283);
nor U22368 (N_22368,N_18261,N_19098);
xnor U22369 (N_22369,N_17567,N_19699);
nor U22370 (N_22370,N_19828,N_19651);
and U22371 (N_22371,N_18143,N_18015);
nor U22372 (N_22372,N_18420,N_18604);
xor U22373 (N_22373,N_19560,N_18049);
nor U22374 (N_22374,N_18853,N_17834);
nand U22375 (N_22375,N_18708,N_19952);
xnor U22376 (N_22376,N_18453,N_18474);
xor U22377 (N_22377,N_19031,N_17631);
nor U22378 (N_22378,N_17919,N_19854);
xor U22379 (N_22379,N_18612,N_19135);
and U22380 (N_22380,N_19754,N_19679);
or U22381 (N_22381,N_19269,N_17857);
nand U22382 (N_22382,N_19830,N_19337);
nand U22383 (N_22383,N_19621,N_18237);
xnor U22384 (N_22384,N_19965,N_19574);
xor U22385 (N_22385,N_18657,N_18842);
xnor U22386 (N_22386,N_19333,N_19516);
xor U22387 (N_22387,N_19274,N_17765);
xor U22388 (N_22388,N_19285,N_19784);
or U22389 (N_22389,N_17546,N_18172);
nand U22390 (N_22390,N_18834,N_19014);
xnor U22391 (N_22391,N_18823,N_18920);
or U22392 (N_22392,N_18559,N_19095);
and U22393 (N_22393,N_19072,N_18147);
nand U22394 (N_22394,N_19085,N_18241);
and U22395 (N_22395,N_18809,N_19951);
xor U22396 (N_22396,N_19348,N_17645);
nand U22397 (N_22397,N_18080,N_17536);
nand U22398 (N_22398,N_19324,N_19254);
and U22399 (N_22399,N_17700,N_18027);
and U22400 (N_22400,N_19826,N_19364);
xnor U22401 (N_22401,N_19593,N_17668);
and U22402 (N_22402,N_18860,N_18068);
xnor U22403 (N_22403,N_19340,N_18735);
and U22404 (N_22404,N_17602,N_19445);
xnor U22405 (N_22405,N_17788,N_18029);
or U22406 (N_22406,N_19979,N_17653);
and U22407 (N_22407,N_19311,N_19035);
and U22408 (N_22408,N_18975,N_18267);
nor U22409 (N_22409,N_18692,N_19675);
nand U22410 (N_22410,N_19512,N_18614);
or U22411 (N_22411,N_18548,N_18895);
and U22412 (N_22412,N_18548,N_19788);
or U22413 (N_22413,N_18480,N_18652);
nand U22414 (N_22414,N_17588,N_18053);
or U22415 (N_22415,N_17813,N_17587);
and U22416 (N_22416,N_19101,N_18618);
nor U22417 (N_22417,N_18238,N_17928);
nor U22418 (N_22418,N_19262,N_18416);
and U22419 (N_22419,N_19335,N_18643);
or U22420 (N_22420,N_19857,N_19809);
or U22421 (N_22421,N_17643,N_18881);
nor U22422 (N_22422,N_19104,N_18829);
xnor U22423 (N_22423,N_18394,N_18032);
xor U22424 (N_22424,N_19190,N_17987);
and U22425 (N_22425,N_19121,N_19637);
nand U22426 (N_22426,N_19803,N_18805);
nand U22427 (N_22427,N_17759,N_17880);
or U22428 (N_22428,N_18993,N_18493);
xor U22429 (N_22429,N_19991,N_19738);
xor U22430 (N_22430,N_19140,N_18495);
or U22431 (N_22431,N_17538,N_19631);
or U22432 (N_22432,N_19593,N_17509);
xor U22433 (N_22433,N_17687,N_19153);
or U22434 (N_22434,N_18249,N_17963);
or U22435 (N_22435,N_19499,N_17916);
nor U22436 (N_22436,N_19019,N_18319);
xnor U22437 (N_22437,N_18316,N_18808);
nand U22438 (N_22438,N_18389,N_18106);
or U22439 (N_22439,N_18345,N_19796);
and U22440 (N_22440,N_19516,N_19886);
xnor U22441 (N_22441,N_17837,N_19387);
nand U22442 (N_22442,N_19914,N_17642);
or U22443 (N_22443,N_19870,N_17535);
xor U22444 (N_22444,N_18008,N_17527);
nor U22445 (N_22445,N_19884,N_18471);
or U22446 (N_22446,N_18919,N_19667);
and U22447 (N_22447,N_17612,N_18033);
nor U22448 (N_22448,N_17941,N_17601);
nand U22449 (N_22449,N_17937,N_19274);
and U22450 (N_22450,N_19458,N_18725);
and U22451 (N_22451,N_18781,N_18512);
xnor U22452 (N_22452,N_19803,N_19173);
and U22453 (N_22453,N_19686,N_18854);
nand U22454 (N_22454,N_19589,N_18968);
xor U22455 (N_22455,N_17949,N_18282);
nand U22456 (N_22456,N_19251,N_19896);
nand U22457 (N_22457,N_19654,N_18958);
nand U22458 (N_22458,N_18735,N_18363);
nor U22459 (N_22459,N_17641,N_18522);
and U22460 (N_22460,N_19741,N_18000);
or U22461 (N_22461,N_18565,N_19115);
xnor U22462 (N_22462,N_19797,N_17942);
nor U22463 (N_22463,N_18388,N_19346);
nor U22464 (N_22464,N_18116,N_19621);
nand U22465 (N_22465,N_17791,N_19008);
and U22466 (N_22466,N_17955,N_17639);
xnor U22467 (N_22467,N_19708,N_19459);
nand U22468 (N_22468,N_17511,N_17944);
and U22469 (N_22469,N_18594,N_19484);
or U22470 (N_22470,N_18126,N_17775);
or U22471 (N_22471,N_17650,N_18816);
or U22472 (N_22472,N_17689,N_19369);
and U22473 (N_22473,N_19927,N_18656);
and U22474 (N_22474,N_19116,N_19455);
nor U22475 (N_22475,N_19043,N_18766);
nor U22476 (N_22476,N_18398,N_18062);
or U22477 (N_22477,N_19639,N_19946);
xor U22478 (N_22478,N_18125,N_18559);
or U22479 (N_22479,N_17927,N_19897);
nor U22480 (N_22480,N_19105,N_19712);
nor U22481 (N_22481,N_19895,N_18308);
nor U22482 (N_22482,N_19913,N_19228);
xor U22483 (N_22483,N_19558,N_18692);
nor U22484 (N_22484,N_18339,N_19759);
xnor U22485 (N_22485,N_19798,N_18572);
nand U22486 (N_22486,N_18356,N_18435);
nand U22487 (N_22487,N_19309,N_18305);
xor U22488 (N_22488,N_19178,N_18689);
nor U22489 (N_22489,N_19032,N_18837);
nand U22490 (N_22490,N_18679,N_17928);
xnor U22491 (N_22491,N_19985,N_19924);
nor U22492 (N_22492,N_19794,N_18326);
nand U22493 (N_22493,N_18815,N_17914);
and U22494 (N_22494,N_18834,N_18797);
or U22495 (N_22495,N_18609,N_18732);
nor U22496 (N_22496,N_19681,N_18330);
nor U22497 (N_22497,N_19381,N_18556);
or U22498 (N_22498,N_18838,N_18808);
nor U22499 (N_22499,N_19033,N_19626);
nor U22500 (N_22500,N_21096,N_20740);
nor U22501 (N_22501,N_20893,N_20887);
and U22502 (N_22502,N_21013,N_21171);
nor U22503 (N_22503,N_20478,N_21558);
or U22504 (N_22504,N_21764,N_20675);
and U22505 (N_22505,N_20421,N_21742);
or U22506 (N_22506,N_20597,N_21791);
nor U22507 (N_22507,N_22332,N_20070);
xnor U22508 (N_22508,N_22055,N_21535);
nor U22509 (N_22509,N_21018,N_22366);
or U22510 (N_22510,N_21399,N_21426);
nand U22511 (N_22511,N_20767,N_21626);
nor U22512 (N_22512,N_21800,N_21323);
and U22513 (N_22513,N_22165,N_20814);
or U22514 (N_22514,N_21882,N_21395);
and U22515 (N_22515,N_22313,N_22365);
or U22516 (N_22516,N_21089,N_21133);
nand U22517 (N_22517,N_21037,N_20377);
xnor U22518 (N_22518,N_21246,N_21852);
and U22519 (N_22519,N_22259,N_21364);
nand U22520 (N_22520,N_21310,N_22018);
and U22521 (N_22521,N_20164,N_21505);
and U22522 (N_22522,N_21935,N_22217);
nor U22523 (N_22523,N_20585,N_20372);
xor U22524 (N_22524,N_20475,N_22150);
or U22525 (N_22525,N_20707,N_21795);
nor U22526 (N_22526,N_22193,N_21451);
nand U22527 (N_22527,N_20084,N_20205);
and U22528 (N_22528,N_20045,N_20752);
nor U22529 (N_22529,N_20474,N_22236);
xor U22530 (N_22530,N_21555,N_20050);
xor U22531 (N_22531,N_22022,N_20267);
and U22532 (N_22532,N_22068,N_20548);
nand U22533 (N_22533,N_20854,N_22435);
nand U22534 (N_22534,N_22324,N_21066);
nor U22535 (N_22535,N_21416,N_20677);
nand U22536 (N_22536,N_20510,N_20998);
nor U22537 (N_22537,N_20047,N_22104);
nor U22538 (N_22538,N_21633,N_22306);
xnor U22539 (N_22539,N_21636,N_21298);
or U22540 (N_22540,N_22132,N_20036);
nand U22541 (N_22541,N_22491,N_20097);
nor U22542 (N_22542,N_22134,N_22117);
or U22543 (N_22543,N_20590,N_20865);
nand U22544 (N_22544,N_20604,N_20052);
or U22545 (N_22545,N_21990,N_21065);
xnor U22546 (N_22546,N_21352,N_21726);
nor U22547 (N_22547,N_20243,N_20837);
and U22548 (N_22548,N_20336,N_21022);
xnor U22549 (N_22549,N_21290,N_21327);
and U22550 (N_22550,N_22384,N_20704);
nand U22551 (N_22551,N_21069,N_21942);
nand U22552 (N_22552,N_21039,N_20227);
or U22553 (N_22553,N_20215,N_20713);
or U22554 (N_22554,N_22394,N_22181);
nor U22555 (N_22555,N_20182,N_21024);
xnor U22556 (N_22556,N_22347,N_20549);
nand U22557 (N_22557,N_21015,N_20957);
or U22558 (N_22558,N_20757,N_21149);
and U22559 (N_22559,N_22005,N_21255);
nand U22560 (N_22560,N_21357,N_21927);
nand U22561 (N_22561,N_20016,N_20134);
and U22562 (N_22562,N_20771,N_21048);
nand U22563 (N_22563,N_21411,N_21932);
and U22564 (N_22564,N_20044,N_22326);
xnor U22565 (N_22565,N_20608,N_20090);
xnor U22566 (N_22566,N_21509,N_21554);
xnor U22567 (N_22567,N_20820,N_20127);
xnor U22568 (N_22568,N_21773,N_21602);
and U22569 (N_22569,N_22002,N_20932);
or U22570 (N_22570,N_20408,N_20672);
nor U22571 (N_22571,N_20412,N_20892);
nor U22572 (N_22572,N_20295,N_20742);
nor U22573 (N_22573,N_20329,N_21785);
nand U22574 (N_22574,N_21100,N_21944);
nor U22575 (N_22575,N_21432,N_21518);
nor U22576 (N_22576,N_20493,N_21784);
xor U22577 (N_22577,N_22454,N_20456);
nor U22578 (N_22578,N_21590,N_20866);
xnor U22579 (N_22579,N_20853,N_20149);
and U22580 (N_22580,N_20646,N_22270);
and U22581 (N_22581,N_21288,N_20225);
and U22582 (N_22582,N_21506,N_21651);
or U22583 (N_22583,N_21193,N_22076);
or U22584 (N_22584,N_20682,N_22239);
or U22585 (N_22585,N_22354,N_21036);
or U22586 (N_22586,N_20207,N_20003);
xnor U22587 (N_22587,N_20150,N_21946);
or U22588 (N_22588,N_20235,N_21978);
or U22589 (N_22589,N_21603,N_20944);
nand U22590 (N_22590,N_21094,N_22119);
xor U22591 (N_22591,N_22231,N_21152);
xnor U22592 (N_22592,N_22249,N_20147);
nand U22593 (N_22593,N_20739,N_21214);
xor U22594 (N_22594,N_21588,N_21861);
nand U22595 (N_22595,N_20249,N_20934);
nor U22596 (N_22596,N_21582,N_20844);
nand U22597 (N_22597,N_22393,N_21286);
xnor U22598 (N_22598,N_21786,N_22344);
nand U22599 (N_22599,N_21804,N_20253);
xnor U22600 (N_22600,N_22112,N_20762);
nor U22601 (N_22601,N_20393,N_20831);
nor U22602 (N_22602,N_21621,N_20744);
nor U22603 (N_22603,N_21869,N_20361);
nor U22604 (N_22604,N_20492,N_21315);
and U22605 (N_22605,N_21546,N_22311);
nor U22606 (N_22606,N_21049,N_20547);
nand U22607 (N_22607,N_22466,N_20068);
and U22608 (N_22608,N_21997,N_22097);
nand U22609 (N_22609,N_20032,N_21261);
or U22610 (N_22610,N_21106,N_20165);
xnor U22611 (N_22611,N_20530,N_21139);
nor U22612 (N_22612,N_20055,N_20064);
nand U22613 (N_22613,N_21428,N_20426);
or U22614 (N_22614,N_20335,N_20968);
nand U22615 (N_22615,N_22277,N_21635);
xnor U22616 (N_22616,N_22352,N_20157);
nor U22617 (N_22617,N_22314,N_22173);
nand U22618 (N_22618,N_20507,N_21318);
or U22619 (N_22619,N_20572,N_21964);
nor U22620 (N_22620,N_21335,N_21911);
nand U22621 (N_22621,N_20895,N_20786);
and U22622 (N_22622,N_20795,N_22014);
or U22623 (N_22623,N_22212,N_21445);
or U22624 (N_22624,N_21185,N_20722);
and U22625 (N_22625,N_20119,N_20277);
xnor U22626 (N_22626,N_22368,N_22362);
nand U22627 (N_22627,N_22448,N_22090);
nor U22628 (N_22628,N_20755,N_21977);
nor U22629 (N_22629,N_22310,N_21282);
or U22630 (N_22630,N_21908,N_21697);
nand U22631 (N_22631,N_20730,N_22462);
and U22632 (N_22632,N_20857,N_22082);
nand U22633 (N_22633,N_21652,N_22098);
or U22634 (N_22634,N_20930,N_20317);
xnor U22635 (N_22635,N_21517,N_21910);
or U22636 (N_22636,N_20297,N_21482);
or U22637 (N_22637,N_21731,N_20287);
nand U22638 (N_22638,N_20240,N_20031);
nand U22639 (N_22639,N_21166,N_20557);
or U22640 (N_22640,N_21741,N_20982);
or U22641 (N_22641,N_20327,N_22035);
xor U22642 (N_22642,N_21980,N_22091);
xor U22643 (N_22643,N_21688,N_20138);
xor U22644 (N_22644,N_20712,N_21712);
nand U22645 (N_22645,N_21141,N_20625);
and U22646 (N_22646,N_21940,N_20966);
or U22647 (N_22647,N_21394,N_21873);
xnor U22648 (N_22648,N_22229,N_20644);
or U22649 (N_22649,N_20439,N_20914);
nor U22650 (N_22650,N_21016,N_21306);
xnor U22651 (N_22651,N_20954,N_21706);
nor U22652 (N_22652,N_20735,N_21271);
nand U22653 (N_22653,N_21281,N_20034);
or U22654 (N_22654,N_22093,N_22070);
nor U22655 (N_22655,N_21787,N_22095);
nand U22656 (N_22656,N_22279,N_20635);
xor U22657 (N_22657,N_22413,N_21081);
nand U22658 (N_22658,N_22260,N_21299);
xnor U22659 (N_22659,N_20656,N_21272);
and U22660 (N_22660,N_21189,N_21027);
and U22661 (N_22661,N_21328,N_22139);
xor U22662 (N_22662,N_20542,N_21462);
nand U22663 (N_22663,N_22322,N_22382);
nor U22664 (N_22664,N_21711,N_21478);
xor U22665 (N_22665,N_22088,N_21347);
xor U22666 (N_22666,N_20875,N_21543);
nand U22667 (N_22667,N_21296,N_20759);
and U22668 (N_22668,N_22375,N_20734);
and U22669 (N_22669,N_20897,N_22419);
nor U22670 (N_22670,N_20621,N_20663);
or U22671 (N_22671,N_22490,N_20444);
and U22672 (N_22672,N_21629,N_20867);
xnor U22673 (N_22673,N_21115,N_21632);
or U22674 (N_22674,N_21471,N_22497);
and U22675 (N_22675,N_21441,N_22301);
or U22676 (N_22676,N_22201,N_21470);
nor U22677 (N_22677,N_21893,N_21040);
or U22678 (N_22678,N_20494,N_20670);
nand U22679 (N_22679,N_20271,N_21914);
nor U22680 (N_22680,N_21884,N_22308);
nand U22681 (N_22681,N_20738,N_21289);
or U22682 (N_22682,N_22111,N_21304);
or U22683 (N_22683,N_21937,N_22267);
and U22684 (N_22684,N_20912,N_20749);
xor U22685 (N_22685,N_21332,N_21538);
and U22686 (N_22686,N_20168,N_20180);
nand U22687 (N_22687,N_22226,N_21539);
nand U22688 (N_22688,N_20343,N_20501);
nor U22689 (N_22689,N_20567,N_21113);
nor U22690 (N_22690,N_21091,N_20030);
xor U22691 (N_22691,N_21684,N_20940);
nand U22692 (N_22692,N_20356,N_20679);
or U22693 (N_22693,N_22464,N_21803);
and U22694 (N_22694,N_20552,N_20888);
xor U22695 (N_22695,N_22333,N_21475);
nand U22696 (N_22696,N_22460,N_21301);
xnor U22697 (N_22697,N_21233,N_21544);
xor U22698 (N_22698,N_20623,N_21634);
xor U22699 (N_22699,N_20841,N_21278);
xnor U22700 (N_22700,N_20963,N_21370);
or U22701 (N_22701,N_21740,N_21936);
xnor U22702 (N_22702,N_21384,N_21906);
nor U22703 (N_22703,N_20580,N_22123);
xor U22704 (N_22704,N_21235,N_21553);
and U22705 (N_22705,N_21616,N_20109);
nand U22706 (N_22706,N_20595,N_22284);
xnor U22707 (N_22707,N_20194,N_20141);
nor U22708 (N_22708,N_21147,N_21524);
nor U22709 (N_22709,N_21270,N_22494);
and U22710 (N_22710,N_20654,N_20469);
nand U22711 (N_22711,N_20156,N_21656);
xnor U22712 (N_22712,N_20950,N_21584);
nand U22713 (N_22713,N_21051,N_21231);
nor U22714 (N_22714,N_20024,N_20487);
nor U22715 (N_22715,N_20276,N_22476);
or U22716 (N_22716,N_20201,N_20238);
nor U22717 (N_22717,N_22079,N_21236);
nor U22718 (N_22718,N_21960,N_21161);
nor U22719 (N_22719,N_20371,N_22012);
or U22720 (N_22720,N_22355,N_21947);
and U22721 (N_22721,N_20354,N_22264);
nand U22722 (N_22722,N_21685,N_20971);
nor U22723 (N_22723,N_22010,N_20220);
and U22724 (N_22724,N_20155,N_20203);
and U22725 (N_22725,N_20234,N_20079);
or U22726 (N_22726,N_21502,N_20946);
nand U22727 (N_22727,N_21026,N_21950);
or U22728 (N_22728,N_22161,N_20471);
nand U22729 (N_22729,N_20221,N_22475);
nand U22730 (N_22730,N_22081,N_21070);
xor U22731 (N_22731,N_21447,N_21552);
nor U22732 (N_22732,N_21537,N_21494);
nor U22733 (N_22733,N_22292,N_20925);
and U22734 (N_22734,N_22027,N_21153);
and U22735 (N_22735,N_21003,N_22183);
and U22736 (N_22736,N_21614,N_20299);
xnor U22737 (N_22737,N_22445,N_20233);
nand U22738 (N_22738,N_22361,N_21190);
nand U22739 (N_22739,N_20571,N_21720);
nand U22740 (N_22740,N_21611,N_20918);
or U22741 (N_22741,N_20649,N_22402);
nand U22742 (N_22742,N_20489,N_21401);
nor U22743 (N_22743,N_20922,N_20216);
and U22744 (N_22744,N_22468,N_22189);
or U22745 (N_22745,N_20063,N_22047);
nand U22746 (N_22746,N_22387,N_21234);
and U22747 (N_22747,N_21268,N_20651);
or U22748 (N_22748,N_20962,N_20929);
nand U22749 (N_22749,N_22015,N_20190);
and U22750 (N_22750,N_21188,N_21686);
nand U22751 (N_22751,N_21607,N_21930);
nand U22752 (N_22752,N_20696,N_22137);
nand U22753 (N_22753,N_21928,N_22498);
xor U22754 (N_22754,N_20890,N_21424);
xnor U22755 (N_22755,N_20796,N_22381);
or U22756 (N_22756,N_21446,N_20396);
nor U22757 (N_22757,N_20562,N_20442);
and U22758 (N_22758,N_21759,N_21510);
nand U22759 (N_22759,N_20671,N_22374);
nand U22760 (N_22760,N_20842,N_22458);
or U22761 (N_22761,N_21004,N_21929);
nor U22762 (N_22762,N_20222,N_20258);
nand U22763 (N_22763,N_20816,N_20037);
or U22764 (N_22764,N_20637,N_21067);
xor U22765 (N_22765,N_20010,N_22258);
nor U22766 (N_22766,N_21837,N_22084);
or U22767 (N_22767,N_20579,N_20454);
and U22768 (N_22768,N_20710,N_20839);
nand U22769 (N_22769,N_20450,N_22395);
nor U22770 (N_22770,N_21647,N_21644);
and U22771 (N_22771,N_22042,N_22272);
xor U22772 (N_22772,N_21182,N_20368);
nand U22773 (N_22773,N_22431,N_22009);
nor U22774 (N_22774,N_20272,N_21668);
nor U22775 (N_22775,N_21485,N_21209);
nor U22776 (N_22776,N_20486,N_21339);
nand U22777 (N_22777,N_20268,N_21995);
xor U22778 (N_22778,N_20942,N_21843);
or U22779 (N_22779,N_20163,N_20613);
or U22780 (N_22780,N_21245,N_20809);
or U22781 (N_22781,N_20583,N_20452);
xnor U22782 (N_22782,N_21736,N_21704);
xnor U22783 (N_22783,N_20414,N_21824);
and U22784 (N_22784,N_22020,N_21158);
or U22785 (N_22785,N_21413,N_21799);
nand U22786 (N_22786,N_20462,N_20695);
and U22787 (N_22787,N_21259,N_22116);
and U22788 (N_22788,N_20296,N_21904);
nor U22789 (N_22789,N_20514,N_21788);
or U22790 (N_22790,N_22167,N_20555);
and U22791 (N_22791,N_21131,N_22335);
and U22792 (N_22792,N_20959,N_22390);
nor U22793 (N_22793,N_22053,N_21643);
and U22794 (N_22794,N_21679,N_20758);
xor U22795 (N_22795,N_21576,N_20697);
and U22796 (N_22796,N_22210,N_22298);
nor U22797 (N_22797,N_20999,N_22321);
xnor U22798 (N_22798,N_20110,N_20324);
or U22799 (N_22799,N_20259,N_20404);
or U22800 (N_22800,N_20169,N_21253);
nor U22801 (N_22801,N_22232,N_21354);
and U22802 (N_22802,N_20525,N_22453);
or U22803 (N_22803,N_20995,N_21126);
nand U22804 (N_22804,N_20676,N_20433);
xnor U22805 (N_22805,N_21872,N_20325);
and U22806 (N_22806,N_20978,N_21257);
or U22807 (N_22807,N_20559,N_21962);
nor U22808 (N_22808,N_20199,N_20680);
xnor U22809 (N_22809,N_20383,N_20062);
and U22810 (N_22810,N_21609,N_20184);
or U22811 (N_22811,N_20148,N_22101);
nor U22812 (N_22812,N_22338,N_21194);
nor U22813 (N_22813,N_21695,N_20927);
xor U22814 (N_22814,N_21710,N_20049);
or U22815 (N_22815,N_22248,N_21279);
nand U22816 (N_22816,N_20691,N_22320);
and U22817 (N_22817,N_21284,N_20065);
and U22818 (N_22818,N_22031,N_21488);
xnor U22819 (N_22819,N_20975,N_21682);
nand U22820 (N_22820,N_20799,N_20241);
and U22821 (N_22821,N_20883,N_21312);
nand U22822 (N_22822,N_20774,N_21409);
nor U22823 (N_22823,N_20951,N_20939);
nor U22824 (N_22824,N_21489,N_20123);
nand U22825 (N_22825,N_20619,N_20901);
and U22826 (N_22826,N_21247,N_21833);
nand U22827 (N_22827,N_20424,N_21949);
and U22828 (N_22828,N_21056,N_21766);
xnor U22829 (N_22829,N_21573,N_21496);
nor U22830 (N_22830,N_21368,N_22000);
nor U22831 (N_22831,N_20535,N_21307);
nand U22832 (N_22832,N_21993,N_22273);
xor U22833 (N_22833,N_21693,N_22124);
and U22834 (N_22834,N_21892,N_22440);
or U22835 (N_22835,N_20896,N_20095);
or U22836 (N_22836,N_20881,N_21503);
or U22837 (N_22837,N_20202,N_20224);
xnor U22838 (N_22838,N_22108,N_21750);
or U22839 (N_22839,N_20262,N_20121);
nor U22840 (N_22840,N_21835,N_20385);
xor U22841 (N_22841,N_20230,N_20632);
nor U22842 (N_22842,N_20360,N_22001);
nor U22843 (N_22843,N_21516,N_20440);
nor U22844 (N_22844,N_21515,N_22144);
and U22845 (N_22845,N_21659,N_20290);
or U22846 (N_22846,N_20345,N_22004);
or U22847 (N_22847,N_20428,N_21177);
and U22848 (N_22848,N_21009,N_21522);
nand U22849 (N_22849,N_20705,N_21464);
or U22850 (N_22850,N_21373,N_22415);
nand U22851 (N_22851,N_21528,N_20878);
or U22852 (N_22852,N_21753,N_20791);
xor U22853 (N_22853,N_20591,N_20573);
and U22854 (N_22854,N_22160,N_21292);
nor U22855 (N_22855,N_20822,N_21640);
nor U22856 (N_22856,N_21976,N_22305);
nor U22857 (N_22857,N_21438,N_22323);
and U22858 (N_22858,N_21959,N_20790);
xor U22859 (N_22859,N_20394,N_21701);
xnor U22860 (N_22860,N_20298,N_22450);
nor U22861 (N_22861,N_20639,N_21330);
or U22862 (N_22862,N_20470,N_20025);
nor U22863 (N_22863,N_21549,N_22444);
and U22864 (N_22864,N_20674,N_21680);
and U22865 (N_22865,N_22472,N_20174);
nor U22866 (N_22866,N_20126,N_21252);
and U22867 (N_22867,N_20273,N_21690);
or U22868 (N_22868,N_22396,N_20524);
or U22869 (N_22869,N_21689,N_20466);
or U22870 (N_22870,N_22253,N_20872);
and U22871 (N_22871,N_21826,N_21638);
nand U22872 (N_22872,N_22030,N_21560);
nor U22873 (N_22873,N_21500,N_21010);
nor U22874 (N_22874,N_21823,N_20099);
nor U22875 (N_22875,N_21250,N_21989);
xnor U22876 (N_22876,N_21810,N_20815);
nor U22877 (N_22877,N_21902,N_21385);
and U22878 (N_22878,N_20005,N_20529);
xor U22879 (N_22879,N_21174,N_21479);
xnor U22880 (N_22880,N_20609,N_20533);
nor U22881 (N_22881,N_21698,N_20136);
xnor U22882 (N_22882,N_21992,N_20826);
nor U22883 (N_22883,N_20350,N_22023);
and U22884 (N_22884,N_20779,N_21317);
or U22885 (N_22885,N_22192,N_20443);
and U22886 (N_22886,N_21397,N_21021);
and U22887 (N_22887,N_20379,N_20133);
xor U22888 (N_22888,N_21703,N_22271);
and U22889 (N_22889,N_20192,N_21076);
nor U22890 (N_22890,N_21080,N_21455);
and U22891 (N_22891,N_21566,N_22100);
and U22892 (N_22892,N_20517,N_22078);
and U22893 (N_22893,N_20027,N_21206);
xnor U22894 (N_22894,N_20022,N_20989);
or U22895 (N_22895,N_22296,N_21822);
or U22896 (N_22896,N_22049,N_20485);
xor U22897 (N_22897,N_22222,N_21569);
and U22898 (N_22898,N_21311,N_21001);
xor U22899 (N_22899,N_20611,N_20231);
and U22900 (N_22900,N_21913,N_21111);
or U22901 (N_22901,N_22357,N_21264);
and U22902 (N_22902,N_22437,N_22159);
nor U22903 (N_22903,N_21877,N_21196);
nor U22904 (N_22904,N_21765,N_22265);
nor U22905 (N_22905,N_22479,N_21863);
nand U22906 (N_22906,N_22461,N_21867);
or U22907 (N_22907,N_21897,N_20871);
nor U22908 (N_22908,N_22441,N_22372);
nor U22909 (N_22909,N_21376,N_22044);
nor U22910 (N_22910,N_20536,N_21237);
xnor U22911 (N_22911,N_22037,N_21672);
or U22912 (N_22912,N_20515,N_21987);
or U22913 (N_22913,N_22213,N_20122);
and U22914 (N_22914,N_21073,N_21933);
nor U22915 (N_22915,N_22268,N_20128);
xor U22916 (N_22916,N_20178,N_21587);
nand U22917 (N_22917,N_21406,N_21329);
and U22918 (N_22918,N_21109,N_21466);
nand U22919 (N_22919,N_21776,N_20288);
xnor U22920 (N_22920,N_20622,N_20523);
or U22921 (N_22921,N_20596,N_21673);
or U22922 (N_22922,N_22032,N_20229);
nor U22923 (N_22923,N_21974,N_20745);
nor U22924 (N_22924,N_22171,N_21961);
xor U22925 (N_22925,N_20082,N_20505);
or U22926 (N_22926,N_20568,N_22094);
and U22927 (N_22927,N_22056,N_21477);
or U22928 (N_22928,N_20952,N_20112);
nand U22929 (N_22929,N_20907,N_20638);
or U22930 (N_22930,N_22285,N_22398);
xor U22931 (N_22931,N_20429,N_20006);
xor U22932 (N_22932,N_21727,N_21374);
nand U22933 (N_22933,N_20056,N_20316);
or U22934 (N_22934,N_21657,N_20223);
xor U22935 (N_22935,N_20076,N_20728);
or U22936 (N_22936,N_21570,N_20137);
nand U22937 (N_22937,N_21827,N_21782);
nand U22938 (N_22938,N_21028,N_22128);
nor U22939 (N_22939,N_22028,N_20172);
or U22940 (N_22940,N_20197,N_21601);
and U22941 (N_22941,N_21392,N_21865);
nor U22942 (N_22942,N_21223,N_21020);
nand U22943 (N_22943,N_20798,N_20577);
nor U22944 (N_22944,N_20096,N_21599);
xnor U22945 (N_22945,N_22289,N_21118);
nor U22946 (N_22946,N_20804,N_21350);
nor U22947 (N_22947,N_22457,N_21291);
xor U22948 (N_22948,N_20627,N_21232);
nand U22949 (N_22949,N_20666,N_21414);
and U22950 (N_22950,N_22169,N_20565);
nor U22951 (N_22951,N_21107,N_21430);
or U22952 (N_22952,N_20342,N_20092);
and U22953 (N_22953,N_22083,N_20448);
and U22954 (N_22954,N_20900,N_20924);
xor U22955 (N_22955,N_21501,N_21775);
and U22956 (N_22956,N_21275,N_21755);
and U22957 (N_22957,N_21982,N_22294);
or U22958 (N_22958,N_21000,N_22168);
nor U22959 (N_22959,N_21497,N_20793);
and U22960 (N_22960,N_20208,N_20630);
xnor U22961 (N_22961,N_20449,N_21079);
nor U22962 (N_22962,N_20313,N_21207);
nor U22963 (N_22963,N_21739,N_20000);
nor U22964 (N_22964,N_21641,N_20800);
xor U22965 (N_22965,N_22247,N_20323);
nand U22966 (N_22966,N_22484,N_20375);
and U22967 (N_22967,N_20094,N_20019);
and U22968 (N_22968,N_21269,N_22151);
nand U22969 (N_22969,N_22307,N_20617);
and U22970 (N_22970,N_21388,N_21305);
nor U22971 (N_22971,N_21487,N_21919);
xnor U22972 (N_22972,N_21658,N_22007);
nor U22973 (N_22973,N_21205,N_21924);
and U22974 (N_22974,N_20495,N_20560);
or U22975 (N_22975,N_21963,N_20303);
or U22976 (N_22976,N_21922,N_21103);
and U22977 (N_22977,N_21772,N_20960);
and U22978 (N_22978,N_20768,N_22051);
xor U22979 (N_22979,N_21894,N_22399);
xor U22980 (N_22980,N_22131,N_21619);
nor U22981 (N_22981,N_21322,N_21956);
nor U22982 (N_22982,N_20283,N_21197);
xor U22983 (N_22983,N_21366,N_21763);
or U22984 (N_22984,N_21481,N_21807);
xor U22985 (N_22985,N_20935,N_20703);
nand U22986 (N_22986,N_22029,N_21890);
and U22987 (N_22987,N_20154,N_21716);
xor U22988 (N_22988,N_20279,N_21415);
nor U22989 (N_22989,N_21238,N_20551);
nand U22990 (N_22990,N_20824,N_20188);
nor U22991 (N_22991,N_22152,N_20280);
or U22992 (N_22992,N_21217,N_22367);
nor U22993 (N_22993,N_21905,N_21805);
or U22994 (N_22994,N_20144,N_20021);
xnor U22995 (N_22995,N_22345,N_20491);
or U22996 (N_22996,N_21941,N_22489);
nand U22997 (N_22997,N_20254,N_21142);
or U22998 (N_22998,N_21075,N_22470);
and U22999 (N_22999,N_21586,N_21917);
and U23000 (N_23000,N_21043,N_21276);
nand U23001 (N_23001,N_21160,N_20806);
or U23002 (N_23002,N_22302,N_21457);
and U23003 (N_23003,N_21201,N_21938);
nand U23004 (N_23004,N_20943,N_22045);
nor U23005 (N_23005,N_21915,N_21101);
nor U23006 (N_23006,N_21592,N_20080);
or U23007 (N_23007,N_20100,N_20973);
nand U23008 (N_23008,N_20964,N_20801);
and U23009 (N_23009,N_20242,N_20576);
xor U23010 (N_23010,N_21155,N_22166);
nor U23011 (N_23011,N_21058,N_21386);
and U23012 (N_23012,N_22172,N_20789);
xnor U23013 (N_23013,N_21885,N_20472);
or U23014 (N_23014,N_21337,N_20906);
nand U23015 (N_23015,N_21801,N_22337);
or U23016 (N_23016,N_21631,N_21965);
nor U23017 (N_23017,N_20873,N_20833);
and U23018 (N_23018,N_21474,N_20863);
nand U23019 (N_23019,N_21886,N_22401);
nor U23020 (N_23020,N_21577,N_20318);
and U23021 (N_23021,N_20537,N_22219);
nand U23022 (N_23022,N_21719,N_21469);
nor U23023 (N_23023,N_20118,N_21796);
or U23024 (N_23024,N_21921,N_20415);
or U23025 (N_23025,N_21912,N_21624);
and U23026 (N_23026,N_20502,N_20282);
and U23027 (N_23027,N_21984,N_20664);
xnor U23028 (N_23028,N_20257,N_20382);
or U23029 (N_23029,N_20349,N_20775);
nand U23030 (N_23030,N_22436,N_21398);
nor U23031 (N_23031,N_21574,N_20843);
nand U23032 (N_23032,N_22425,N_20477);
nor U23033 (N_23033,N_21721,N_20782);
nor U23034 (N_23034,N_22471,N_20086);
nor U23035 (N_23035,N_21114,N_20248);
xnor U23036 (N_23036,N_21165,N_21148);
nor U23037 (N_23037,N_22325,N_20177);
nor U23038 (N_23038,N_20880,N_21467);
nand U23039 (N_23039,N_21319,N_20285);
xor U23040 (N_23040,N_20293,N_21723);
xor U23041 (N_23041,N_21983,N_21396);
nand U23042 (N_23042,N_21162,N_20176);
nor U23043 (N_23043,N_21340,N_20586);
xor U23044 (N_23044,N_21751,N_20965);
and U23045 (N_23045,N_21239,N_20001);
nor U23046 (N_23046,N_20526,N_22486);
nor U23047 (N_23047,N_21814,N_21654);
xor U23048 (N_23048,N_22426,N_21154);
nor U23049 (N_23049,N_21754,N_20756);
nand U23050 (N_23050,N_20167,N_20009);
nor U23051 (N_23051,N_21220,N_20765);
or U23052 (N_23052,N_21559,N_21622);
or U23053 (N_23053,N_20850,N_21175);
xnor U23054 (N_23054,N_20884,N_20648);
and U23055 (N_23055,N_21520,N_20026);
nand U23056 (N_23056,N_20512,N_21006);
xnor U23057 (N_23057,N_20628,N_22304);
xnor U23058 (N_23058,N_20642,N_21041);
xnor U23059 (N_23059,N_22250,N_20761);
and U23060 (N_23060,N_20633,N_20075);
nor U23061 (N_23061,N_21598,N_20459);
xnor U23062 (N_23062,N_21898,N_20818);
nor U23063 (N_23063,N_21699,N_21637);
and U23064 (N_23064,N_22140,N_21211);
nand U23065 (N_23065,N_20985,N_22184);
nor U23066 (N_23066,N_21901,N_21729);
nand U23067 (N_23067,N_21889,N_20300);
xor U23068 (N_23068,N_22343,N_20331);
or U23069 (N_23069,N_21314,N_21092);
and U23070 (N_23070,N_21864,N_21630);
nor U23071 (N_23071,N_22113,N_21846);
or U23072 (N_23072,N_21498,N_21743);
nor U23073 (N_23073,N_20690,N_20556);
or U23074 (N_23074,N_22269,N_22385);
or U23075 (N_23075,N_21427,N_21053);
nand U23076 (N_23076,N_22065,N_20920);
or U23077 (N_23077,N_20700,N_22295);
and U23078 (N_23078,N_21511,N_20020);
nor U23079 (N_23079,N_20849,N_21575);
nand U23080 (N_23080,N_22157,N_20463);
nand U23081 (N_23081,N_20969,N_21295);
nand U23082 (N_23082,N_21356,N_20714);
nor U23083 (N_23083,N_21361,N_21653);
nand U23084 (N_23084,N_21888,N_20131);
and U23085 (N_23085,N_21547,N_20480);
nor U23086 (N_23086,N_20228,N_20983);
or U23087 (N_23087,N_20784,N_21243);
or U23088 (N_23088,N_20956,N_21216);
and U23089 (N_23089,N_22371,N_20067);
nor U23090 (N_23090,N_20832,N_22349);
nor U23091 (N_23091,N_21140,N_20365);
and U23092 (N_23092,N_22225,N_21098);
xnor U23093 (N_23093,N_22228,N_20183);
nand U23094 (N_23094,N_21953,N_22242);
nand U23095 (N_23095,N_22334,N_21325);
and U23096 (N_23096,N_21124,N_21047);
xor U23097 (N_23097,N_20093,N_21019);
and U23098 (N_23098,N_20719,N_20330);
and U23099 (N_23099,N_20747,N_21733);
or U23100 (N_23100,N_21563,N_21858);
or U23101 (N_23101,N_21879,N_20936);
nand U23102 (N_23102,N_21596,N_21187);
xnor U23103 (N_23103,N_22359,N_20661);
nor U23104 (N_23104,N_22062,N_22218);
nand U23105 (N_23105,N_21844,N_20540);
xnor U23106 (N_23106,N_22455,N_21859);
xor U23107 (N_23107,N_21351,N_20447);
nand U23108 (N_23108,N_20432,N_20255);
or U23109 (N_23109,N_21513,N_20902);
or U23110 (N_23110,N_21419,N_20088);
nor U23111 (N_23111,N_22174,N_20933);
nor U23112 (N_23112,N_22016,N_22341);
xor U23113 (N_23113,N_21831,N_21338);
nor U23114 (N_23114,N_20823,N_20105);
or U23115 (N_23115,N_20506,N_21725);
xor U23116 (N_23116,N_22110,N_21988);
nor U23117 (N_23117,N_21724,N_21745);
and U23118 (N_23118,N_20980,N_20399);
or U23119 (N_23119,N_22059,N_20794);
xor U23120 (N_23120,N_21608,N_20659);
or U23121 (N_23121,N_22439,N_20384);
nand U23122 (N_23122,N_21709,N_20885);
nand U23123 (N_23123,N_20724,N_21875);
nand U23124 (N_23124,N_20864,N_20104);
nand U23125 (N_23125,N_20008,N_21343);
and U23126 (N_23126,N_21064,N_21903);
xnor U23127 (N_23127,N_21714,N_21229);
or U23128 (N_23128,N_21808,N_21121);
or U23129 (N_23129,N_21971,N_22388);
xor U23130 (N_23130,N_20304,N_22432);
xor U23131 (N_23131,N_21815,N_22328);
xor U23132 (N_23132,N_22223,N_22203);
or U23133 (N_23133,N_21757,N_22103);
nand U23134 (N_23134,N_21564,N_22077);
nand U23135 (N_23135,N_21594,N_21512);
and U23136 (N_23136,N_21032,N_20473);
and U23137 (N_23137,N_22149,N_22067);
and U23138 (N_23138,N_22099,N_22411);
nor U23139 (N_23139,N_20481,N_21551);
or U23140 (N_23140,N_21896,N_20620);
xor U23141 (N_23141,N_20718,N_22003);
nor U23142 (N_23142,N_20499,N_20923);
and U23143 (N_23143,N_20101,N_20270);
nand U23144 (N_23144,N_21344,N_21156);
nor U23145 (N_23145,N_21748,N_21849);
and U23146 (N_23146,N_20693,N_22118);
and U23147 (N_23147,N_21204,N_21561);
xor U23148 (N_23148,N_22224,N_20476);
xnor U23149 (N_23149,N_21151,N_21244);
and U23150 (N_23150,N_21143,N_20294);
nor U23151 (N_23151,N_21747,N_20601);
or U23152 (N_23152,N_22061,N_21277);
and U23153 (N_23153,N_21403,N_20400);
nand U23154 (N_23154,N_21737,N_22478);
and U23155 (N_23155,N_20405,N_21514);
xnor U23156 (N_23156,N_20836,N_20351);
and U23157 (N_23157,N_21097,N_21078);
xor U23158 (N_23158,N_22255,N_21666);
and U23159 (N_23159,N_21958,N_22106);
or U23160 (N_23160,N_20129,N_21135);
or U23161 (N_23161,N_21105,N_20825);
or U23162 (N_23162,N_22447,N_21665);
and U23163 (N_23163,N_21381,N_22069);
nand U23164 (N_23164,N_21007,N_21011);
xor U23165 (N_23165,N_20981,N_20792);
xnor U23166 (N_23166,N_22350,N_22196);
nand U23167 (N_23167,N_20852,N_20435);
or U23168 (N_23168,N_20143,N_22185);
nor U23169 (N_23169,N_21023,N_21033);
and U23170 (N_23170,N_20668,N_20389);
xor U23171 (N_23171,N_21429,N_21618);
and U23172 (N_23172,N_21210,N_20500);
nor U23173 (N_23173,N_20497,N_21074);
xor U23174 (N_23174,N_21838,N_21878);
and U23175 (N_23175,N_22046,N_21117);
or U23176 (N_23176,N_21781,N_22073);
xor U23177 (N_23177,N_20977,N_20403);
xor U23178 (N_23178,N_21540,N_20417);
or U23179 (N_23179,N_21851,N_20140);
nand U23180 (N_23180,N_20539,N_20731);
xnor U23181 (N_23181,N_20120,N_20306);
or U23182 (N_23182,N_20598,N_22237);
or U23183 (N_23183,N_20610,N_21192);
and U23184 (N_23184,N_22377,N_20308);
nand U23185 (N_23185,N_21042,N_20059);
nor U23186 (N_23186,N_20321,N_20015);
nor U23187 (N_23187,N_22380,N_20427);
and U23188 (N_23188,N_22405,N_20986);
or U23189 (N_23189,N_21985,N_20701);
xor U23190 (N_23190,N_20061,N_20315);
or U23191 (N_23191,N_22058,N_20014);
and U23192 (N_23192,N_21393,N_21600);
nor U23193 (N_23193,N_21157,N_21083);
xor U23194 (N_23194,N_20185,N_20310);
or U23195 (N_23195,N_22170,N_20013);
nor U23196 (N_23196,N_21044,N_21715);
nor U23197 (N_23197,N_20904,N_22017);
and U23198 (N_23198,N_20314,N_20416);
and U23199 (N_23199,N_20419,N_21050);
nand U23200 (N_23200,N_21678,N_20388);
or U23201 (N_23201,N_20819,N_22474);
or U23202 (N_23202,N_22329,N_20662);
nand U23203 (N_23203,N_20699,N_21655);
and U23204 (N_23204,N_20083,N_21945);
or U23205 (N_23205,N_22422,N_20732);
nand U23206 (N_23206,N_22026,N_22330);
nand U23207 (N_23207,N_20915,N_21931);
nand U23208 (N_23208,N_21055,N_21670);
and U23209 (N_23209,N_21533,N_22105);
nor U23210 (N_23210,N_20239,N_20132);
or U23211 (N_23211,N_20187,N_20496);
and U23212 (N_23212,N_21418,N_22481);
and U23213 (N_23213,N_20987,N_20990);
and U23214 (N_23214,N_22163,N_20363);
nand U23215 (N_23215,N_22075,N_20364);
nand U23216 (N_23216,N_21504,N_20054);
nor U23217 (N_23217,N_21830,N_22175);
nand U23218 (N_23218,N_22013,N_22200);
nor U23219 (N_23219,N_20594,N_21660);
nor U23220 (N_23220,N_20751,N_22358);
and U23221 (N_23221,N_20437,N_21874);
nand U23222 (N_23222,N_20217,N_20508);
and U23223 (N_23223,N_21274,N_20051);
xnor U23224 (N_23224,N_22488,N_20029);
nor U23225 (N_23225,N_21579,N_20717);
and U23226 (N_23226,N_20236,N_22048);
nand U23227 (N_23227,N_21183,N_21578);
nand U23228 (N_23228,N_21358,N_21422);
and U23229 (N_23229,N_21735,N_21379);
xor U23230 (N_23230,N_22403,N_22300);
xnor U23231 (N_23231,N_20289,N_21095);
nor U23232 (N_23232,N_20802,N_22465);
xor U23233 (N_23233,N_20721,N_22418);
xnor U23234 (N_23234,N_21536,N_21829);
and U23235 (N_23235,N_22467,N_21491);
and U23236 (N_23236,N_21060,N_20078);
xor U23237 (N_23237,N_21324,N_20750);
and U23238 (N_23238,N_21420,N_20286);
or U23239 (N_23239,N_21839,N_20592);
and U23240 (N_23240,N_20171,N_21567);
nand U23241 (N_23241,N_20991,N_22162);
nand U23242 (N_23242,N_21173,N_21597);
nand U23243 (N_23243,N_20012,N_22071);
nor U23244 (N_23244,N_22188,N_21265);
xnor U23245 (N_23245,N_21663,N_21480);
xor U23246 (N_23246,N_20048,N_22442);
nor U23247 (N_23247,N_21077,N_21181);
nand U23248 (N_23248,N_20113,N_20593);
or U23249 (N_23249,N_22317,N_21572);
nor U23250 (N_23250,N_20210,N_20307);
nor U23251 (N_23251,N_22254,N_21866);
nand U23252 (N_23252,N_22319,N_22011);
or U23253 (N_23253,N_20687,N_22208);
and U23254 (N_23254,N_20057,N_22257);
or U23255 (N_23255,N_20042,N_21473);
xor U23256 (N_23256,N_22266,N_21132);
and U23257 (N_23257,N_20773,N_20152);
and U23258 (N_23258,N_22276,N_20200);
nor U23259 (N_23259,N_21648,N_20769);
xor U23260 (N_23260,N_20938,N_21819);
and U23261 (N_23261,N_20195,N_20527);
nand U23262 (N_23262,N_20333,N_20334);
or U23263 (N_23263,N_20961,N_21955);
or U23264 (N_23264,N_21059,N_20069);
or U23265 (N_23265,N_21359,N_20587);
or U23266 (N_23266,N_22430,N_20753);
or U23267 (N_23267,N_21589,N_20214);
and U23268 (N_23268,N_20645,N_20028);
and U23269 (N_23269,N_21308,N_21203);
xnor U23270 (N_23270,N_22180,N_22233);
xor U23271 (N_23271,N_20777,N_20247);
and U23272 (N_23272,N_21082,N_20410);
nand U23273 (N_23273,N_22133,N_20589);
nor U23274 (N_23274,N_20851,N_21110);
nor U23275 (N_23275,N_21675,N_21671);
and U23276 (N_23276,N_20035,N_20953);
and U23277 (N_23277,N_21968,N_21186);
nor U23278 (N_23278,N_20618,N_20937);
and U23279 (N_23279,N_22186,N_21326);
and U23280 (N_23280,N_21891,N_21526);
nand U23281 (N_23281,N_20733,N_21375);
nor U23282 (N_23282,N_20746,N_21405);
and U23283 (N_23283,N_22283,N_21408);
nand U23284 (N_23284,N_22376,N_20362);
nor U23285 (N_23285,N_20503,N_21951);
nor U23286 (N_23286,N_21439,N_22198);
xnor U23287 (N_23287,N_21390,N_22179);
or U23288 (N_23288,N_20846,N_20278);
or U23289 (N_23289,N_20905,N_22316);
or U23290 (N_23290,N_21484,N_21421);
nor U23291 (N_23291,N_20401,N_20488);
or U23292 (N_23292,N_21200,N_20909);
xor U23293 (N_23293,N_22052,N_21565);
and U23294 (N_23294,N_22041,N_20252);
xnor U23295 (N_23295,N_20616,N_20889);
nand U23296 (N_23296,N_21119,N_20673);
xnor U23297 (N_23297,N_21542,N_22025);
xor U23298 (N_23298,N_22176,N_22370);
xor U23299 (N_23299,N_21248,N_21130);
and U23300 (N_23300,N_21939,N_21267);
and U23301 (N_23301,N_20958,N_21122);
nand U23302 (N_23302,N_20479,N_21163);
xnor U23303 (N_23303,N_22039,N_20624);
and U23304 (N_23304,N_20206,N_20458);
and U23305 (N_23305,N_20453,N_22299);
xnor U23306 (N_23306,N_22434,N_21966);
or U23307 (N_23307,N_21345,N_20570);
and U23308 (N_23308,N_22040,N_21845);
nand U23309 (N_23309,N_21499,N_20275);
xor U23310 (N_23310,N_22204,N_21531);
nor U23311 (N_23311,N_22339,N_21692);
nor U23312 (N_23312,N_20709,N_20669);
nor U23313 (N_23313,N_22054,N_21899);
nand U23314 (N_23314,N_20541,N_20160);
or U23315 (N_23315,N_21676,N_21090);
nor U23316 (N_23316,N_21262,N_20337);
nand U23317 (N_23317,N_21129,N_21732);
and U23318 (N_23318,N_21258,N_20359);
or U23319 (N_23319,N_20380,N_20921);
or U23320 (N_23320,N_20748,N_21818);
nand U23321 (N_23321,N_22096,N_20153);
nor U23322 (N_23322,N_21127,N_21694);
nand U23323 (N_23323,N_22281,N_20033);
and U23324 (N_23324,N_20422,N_20467);
nand U23325 (N_23325,N_21840,N_21998);
or U23326 (N_23326,N_21790,N_21456);
nand U23327 (N_23327,N_20776,N_22211);
and U23328 (N_23328,N_20139,N_21460);
xnor U23329 (N_23329,N_21730,N_21625);
nor U23330 (N_23330,N_21926,N_21783);
xnor U23331 (N_23331,N_22033,N_20151);
xnor U23332 (N_23332,N_21969,N_22187);
nor U23333 (N_23333,N_22477,N_20322);
and U23334 (N_23334,N_22364,N_20898);
and U23335 (N_23335,N_21468,N_20726);
nor U23336 (N_23336,N_22288,N_20647);
nor U23337 (N_23337,N_20561,N_20212);
xor U23338 (N_23338,N_21226,N_20600);
nor U23339 (N_23339,N_21834,N_20353);
nand U23340 (N_23340,N_20420,N_21778);
or U23341 (N_23341,N_20835,N_22282);
and U23342 (N_23342,N_21123,N_21880);
and U23343 (N_23343,N_20856,N_21465);
and U23344 (N_23344,N_20868,N_22407);
and U23345 (N_23345,N_22373,N_21030);
and U23346 (N_23346,N_20213,N_21014);
nand U23347 (N_23347,N_20347,N_21138);
and U23348 (N_23348,N_20107,N_21365);
xor U23349 (N_23349,N_21717,N_22057);
xnor U23350 (N_23350,N_21568,N_20615);
nor U23351 (N_23351,N_21794,N_21280);
nand U23352 (N_23352,N_20575,N_21198);
or U23353 (N_23353,N_20931,N_20513);
and U23354 (N_23354,N_20232,N_20626);
nand U23355 (N_23355,N_21854,N_20772);
nand U23356 (N_23356,N_20398,N_20711);
xor U23357 (N_23357,N_20715,N_20683);
xnor U23358 (N_23358,N_22206,N_20358);
nand U23359 (N_23359,N_20588,N_21832);
nand U23360 (N_23360,N_20332,N_20817);
or U23361 (N_23361,N_20812,N_21303);
and U23362 (N_23362,N_21591,N_20847);
or U23363 (N_23363,N_22391,N_20855);
nand U23364 (N_23364,N_22109,N_21495);
or U23365 (N_23365,N_21970,N_21948);
nand U23366 (N_23366,N_21313,N_21002);
nand U23367 (N_23367,N_20830,N_20102);
nand U23368 (N_23368,N_21125,N_20984);
nand U23369 (N_23369,N_20244,N_21809);
xor U23370 (N_23370,N_20518,N_21150);
or U23371 (N_23371,N_21628,N_21136);
xor U23372 (N_23372,N_20043,N_21057);
nor U23373 (N_23373,N_21400,N_20103);
and U23374 (N_23374,N_21793,N_22130);
and U23375 (N_23375,N_21134,N_21881);
and U23376 (N_23376,N_20098,N_20729);
nand U23377 (N_23377,N_20702,N_21256);
and U23378 (N_23378,N_21225,N_22410);
xor U23379 (N_23379,N_22456,N_22351);
nand U23380 (N_23380,N_20302,N_20861);
or U23381 (N_23381,N_22245,N_21486);
and U23382 (N_23382,N_21178,N_20698);
or U23383 (N_23383,N_22156,N_20411);
nand U23384 (N_23384,N_22404,N_20538);
nand U23385 (N_23385,N_22063,N_22499);
and U23386 (N_23386,N_22487,N_21797);
nor U23387 (N_23387,N_20108,N_20369);
or U23388 (N_23388,N_21452,N_21108);
nor U23389 (N_23389,N_20928,N_22417);
nand U23390 (N_23390,N_20522,N_21718);
nor U23391 (N_23391,N_22080,N_21771);
xnor U23392 (N_23392,N_21128,N_20189);
nand U23393 (N_23393,N_20941,N_21615);
nor U23394 (N_23394,N_20348,N_20446);
xor U23395 (N_23395,N_22278,N_20544);
nand U23396 (N_23396,N_20218,N_20269);
or U23397 (N_23397,N_22114,N_20166);
or U23398 (N_23398,N_20908,N_22019);
and U23399 (N_23399,N_20545,N_22064);
xnor U23400 (N_23400,N_20340,N_21164);
xnor U23401 (N_23401,N_20720,N_21585);
and U23402 (N_23402,N_21362,N_20409);
and U23403 (N_23403,N_22107,N_21179);
nor U23404 (N_23404,N_21012,N_21167);
xor U23405 (N_23405,N_20870,N_21556);
and U23406 (N_23406,N_21595,N_22446);
nor U23407 (N_23407,N_20423,N_22406);
nor U23408 (N_23408,N_20584,N_20451);
nand U23409 (N_23409,N_21159,N_21072);
or U23410 (N_23410,N_21333,N_21450);
xor U23411 (N_23411,N_20879,N_21664);
xnor U23412 (N_23412,N_20736,N_22414);
or U23413 (N_23413,N_20563,N_20948);
and U23414 (N_23414,N_20554,N_21035);
nand U23415 (N_23415,N_22409,N_21779);
nand U23416 (N_23416,N_21360,N_21461);
nor U23417 (N_23417,N_20550,N_21789);
xor U23418 (N_23418,N_20972,N_20209);
xnor U23419 (N_23419,N_22197,N_22331);
nor U23420 (N_23420,N_21378,N_21382);
xnor U23421 (N_23421,N_20264,N_21883);
nor U23422 (N_23422,N_21769,N_20261);
nor U23423 (N_23423,N_21062,N_21410);
and U23424 (N_23424,N_20498,N_20760);
nand U23425 (N_23425,N_20263,N_21492);
nor U23426 (N_23426,N_20785,N_20805);
or U23427 (N_23427,N_22315,N_21583);
nor U23428 (N_23428,N_22492,N_20081);
nand U23429 (N_23429,N_20810,N_20787);
or U23430 (N_23430,N_20418,N_21483);
xnor U23431 (N_23431,N_21213,N_20116);
nor U23432 (N_23432,N_21847,N_20516);
or U23433 (N_23433,N_21918,N_20468);
nand U23434 (N_23434,N_22369,N_20685);
nand U23435 (N_23435,N_20911,N_20041);
or U23436 (N_23436,N_21523,N_21909);
or U23437 (N_23437,N_21355,N_21802);
and U23438 (N_23438,N_21444,N_21853);
and U23439 (N_23439,N_20370,N_22340);
nor U23440 (N_23440,N_20366,N_20997);
or U23441 (N_23441,N_22389,N_22243);
or U23442 (N_23442,N_21623,N_20490);
nor U23443 (N_23443,N_22074,N_20519);
xor U23444 (N_23444,N_21336,N_22043);
nand U23445 (N_23445,N_20993,N_22146);
xor U23446 (N_23446,N_20460,N_20862);
or U23447 (N_23447,N_21377,N_21862);
nor U23448 (N_23448,N_20445,N_22138);
xnor U23449 (N_23449,N_21240,N_20274);
and U23450 (N_23450,N_21593,N_20284);
xnor U23451 (N_23451,N_21876,N_20341);
or U23452 (N_23452,N_21241,N_20091);
xor U23453 (N_23453,N_22148,N_21562);
nand U23454 (N_23454,N_20115,N_21667);
xnor U23455 (N_23455,N_22240,N_20326);
or U23456 (N_23456,N_20219,N_21169);
and U23457 (N_23457,N_20874,N_22164);
nor U23458 (N_23458,N_22275,N_21087);
xnor U23459 (N_23459,N_20011,N_21391);
nor U23460 (N_23460,N_22286,N_21871);
nand U23461 (N_23461,N_21266,N_21943);
and U23462 (N_23462,N_21525,N_21841);
or U23463 (N_23463,N_20546,N_22353);
and U23464 (N_23464,N_20813,N_21242);
and U23465 (N_23465,N_22092,N_22309);
nor U23466 (N_23466,N_22121,N_22209);
or U23467 (N_23467,N_21346,N_20643);
nor U23468 (N_23468,N_20574,N_20641);
and U23469 (N_23469,N_21722,N_20534);
nand U23470 (N_23470,N_20521,N_20581);
nand U23471 (N_23471,N_21979,N_21812);
and U23472 (N_23472,N_22261,N_20657);
xnor U23473 (N_23473,N_20599,N_21052);
and U23474 (N_23474,N_22087,N_22427);
xnor U23475 (N_23475,N_21677,N_20509);
and U23476 (N_23476,N_20319,N_20603);
nand U23477 (N_23477,N_22195,N_20175);
xnor U23478 (N_23478,N_21137,N_20464);
nand U23479 (N_23479,N_20250,N_20357);
xnor U23480 (N_23480,N_21981,N_22234);
and U23481 (N_23481,N_21855,N_22378);
and U23482 (N_23482,N_22202,N_20146);
nand U23483 (N_23483,N_21320,N_22473);
nand U23484 (N_23484,N_21008,N_22220);
xor U23485 (N_23485,N_20655,N_22400);
xor U23486 (N_23486,N_21068,N_21172);
nor U23487 (N_23487,N_20612,N_20882);
nand U23488 (N_23488,N_21813,N_21448);
and U23489 (N_23489,N_20374,N_21669);
nand U23490 (N_23490,N_21650,N_21642);
nand U23491 (N_23491,N_22493,N_21145);
nand U23492 (N_23492,N_20631,N_20338);
nor U23493 (N_23493,N_22482,N_20910);
and U23494 (N_23494,N_20483,N_20894);
or U23495 (N_23495,N_21530,N_22129);
or U23496 (N_23496,N_20511,N_21848);
nand U23497 (N_23497,N_20976,N_21507);
nor U23498 (N_23498,N_20260,N_21251);
xnor U23499 (N_23499,N_20191,N_21300);
nor U23500 (N_23500,N_21817,N_20992);
and U23501 (N_23501,N_21973,N_21613);
xor U23502 (N_23502,N_21437,N_21309);
xnor U23503 (N_23503,N_21571,N_21371);
or U23504 (N_23504,N_20004,N_21084);
and U23505 (N_23505,N_20226,N_21402);
xor U23506 (N_23506,N_20198,N_22423);
or U23507 (N_23507,N_20629,N_20754);
and U23508 (N_23508,N_21825,N_21454);
nand U23509 (N_23509,N_20821,N_20457);
nand U23510 (N_23510,N_22089,N_20606);
xnor U23511 (N_23511,N_21728,N_20060);
xor U23512 (N_23512,N_21294,N_20397);
or U23513 (N_23513,N_20684,N_22495);
or U23514 (N_23514,N_21046,N_20251);
nand U23515 (N_23515,N_20564,N_20859);
nor U23516 (N_23516,N_21691,N_21870);
xnor U23517 (N_23517,N_20378,N_21453);
xnor U23518 (N_23518,N_21702,N_21923);
or U23519 (N_23519,N_22280,N_21071);
xor U23520 (N_23520,N_20945,N_21195);
nand U23521 (N_23521,N_20406,N_20339);
xnor U23522 (N_23522,N_20994,N_21700);
nor U23523 (N_23523,N_21061,N_20840);
nor U23524 (N_23524,N_20876,N_22424);
xor U23525 (N_23525,N_20040,N_22158);
nor U23526 (N_23526,N_21581,N_21627);
xor U23527 (N_23527,N_21604,N_21612);
xor U23528 (N_23528,N_20678,N_21532);
nor U23529 (N_23529,N_22024,N_22480);
and U23530 (N_23530,N_22034,N_22126);
nand U23531 (N_23531,N_20716,N_21228);
and U23532 (N_23532,N_21031,N_22066);
or U23533 (N_23533,N_20381,N_21548);
or U23534 (N_23534,N_20694,N_20039);
nand U23535 (N_23535,N_20158,N_21342);
xnor U23536 (N_23536,N_20367,N_21681);
and U23537 (N_23537,N_22483,N_20916);
nand U23538 (N_23538,N_21744,N_22153);
nand U23539 (N_23539,N_21646,N_22182);
nand U23540 (N_23540,N_21907,N_22287);
or U23541 (N_23541,N_20650,N_21202);
nor U23542 (N_23542,N_21387,N_21180);
nor U23543 (N_23543,N_20484,N_20046);
nand U23544 (N_23544,N_22135,N_22216);
nand U23545 (N_23545,N_20504,N_21529);
or U23546 (N_23546,N_20114,N_20723);
nor U23547 (N_23547,N_21842,N_20686);
or U23548 (N_23548,N_22303,N_20988);
or U23549 (N_23549,N_22136,N_22235);
or U23550 (N_23550,N_20161,N_20605);
nor U23551 (N_23551,N_20955,N_20781);
nand U23552 (N_23552,N_20145,N_21620);
and U23553 (N_23553,N_21404,N_22451);
or U23554 (N_23554,N_20688,N_21541);
or U23555 (N_23555,N_20074,N_21856);
or U23556 (N_23556,N_20482,N_21749);
or U23557 (N_23557,N_21005,N_22327);
nand U23558 (N_23558,N_21463,N_22421);
nand U23559 (N_23559,N_22036,N_21762);
and U23560 (N_23560,N_20438,N_20023);
or U23561 (N_23561,N_21493,N_20829);
or U23562 (N_23562,N_20634,N_21433);
and U23563 (N_23563,N_22433,N_22199);
or U23564 (N_23564,N_20085,N_20066);
nand U23565 (N_23565,N_21756,N_20455);
nor U23566 (N_23566,N_20692,N_22383);
nand U23567 (N_23567,N_20917,N_22318);
nand U23568 (N_23568,N_20430,N_21086);
or U23569 (N_23569,N_20869,N_21994);
nor U23570 (N_23570,N_21334,N_21112);
or U23571 (N_23571,N_22060,N_21758);
or U23572 (N_23572,N_22008,N_21459);
nor U23573 (N_23573,N_20159,N_20053);
xnor U23574 (N_23574,N_22408,N_20764);
xnor U23575 (N_23575,N_21293,N_21341);
nor U23576 (N_23576,N_21431,N_22386);
nand U23577 (N_23577,N_20803,N_20434);
or U23578 (N_23578,N_20741,N_20947);
xor U23579 (N_23579,N_21230,N_20395);
xnor U23580 (N_23580,N_20860,N_21767);
xnor U23581 (N_23581,N_21605,N_20125);
and U23582 (N_23582,N_21093,N_20903);
and U23583 (N_23583,N_21348,N_21146);
nand U23584 (N_23584,N_21029,N_21617);
and U23585 (N_23585,N_21380,N_22397);
or U23586 (N_23586,N_22205,N_21434);
nand U23587 (N_23587,N_22420,N_22348);
or U23588 (N_23588,N_20135,N_20528);
nand U23589 (N_23589,N_21367,N_21836);
xnor U23590 (N_23590,N_20246,N_21895);
xor U23591 (N_23591,N_21458,N_20111);
nor U23592 (N_23592,N_20543,N_22443);
or U23593 (N_23593,N_20461,N_21610);
xnor U23594 (N_23594,N_21545,N_21442);
or U23595 (N_23595,N_22050,N_21534);
and U23596 (N_23596,N_20807,N_22191);
and U23597 (N_23597,N_21999,N_22336);
nor U23598 (N_23598,N_21645,N_21972);
xnor U23599 (N_23599,N_21425,N_21316);
and U23600 (N_23600,N_22449,N_20344);
and U23601 (N_23601,N_21285,N_21440);
nor U23602 (N_23602,N_22363,N_20979);
xor U23603 (N_23603,N_21412,N_21407);
nor U23604 (N_23604,N_21260,N_21383);
and U23605 (N_23605,N_21054,N_21734);
or U23606 (N_23606,N_21752,N_21297);
nand U23607 (N_23607,N_20797,N_21116);
xnor U23608 (N_23608,N_20737,N_20007);
xor U23609 (N_23609,N_20780,N_20763);
or U23610 (N_23610,N_20582,N_21954);
nand U23611 (N_23611,N_22207,N_21349);
and U23612 (N_23612,N_20766,N_21705);
nand U23613 (N_23613,N_21221,N_20072);
nand U23614 (N_23614,N_20725,N_22021);
or U23615 (N_23615,N_20532,N_21661);
xor U23616 (N_23616,N_21017,N_20077);
and U23617 (N_23617,N_21696,N_20425);
nand U23618 (N_23618,N_20186,N_20967);
or U23619 (N_23619,N_22392,N_22238);
xnor U23620 (N_23620,N_21774,N_21649);
and U23621 (N_23621,N_21887,N_21389);
nor U23622 (N_23622,N_21191,N_22038);
xor U23623 (N_23623,N_20640,N_20355);
and U23624 (N_23624,N_22428,N_20266);
nor U23625 (N_23625,N_21687,N_21821);
xnor U23626 (N_23626,N_22251,N_21557);
and U23627 (N_23627,N_20743,N_22356);
nand U23628 (N_23628,N_22147,N_21184);
nand U23629 (N_23629,N_20292,N_21490);
or U23630 (N_23630,N_22241,N_21227);
nor U23631 (N_23631,N_21208,N_21707);
xnor U23632 (N_23632,N_21662,N_20256);
and U23633 (N_23633,N_20566,N_21331);
xor U23634 (N_23634,N_21144,N_20652);
xnor U23635 (N_23635,N_20387,N_22291);
nor U23636 (N_23636,N_20073,N_20089);
and U23637 (N_23637,N_21088,N_20848);
nand U23638 (N_23638,N_21519,N_22230);
nand U23639 (N_23639,N_21828,N_20130);
xor U23640 (N_23640,N_20919,N_20265);
xnor U23641 (N_23641,N_21746,N_21920);
nand U23642 (N_23642,N_22086,N_20558);
and U23643 (N_23643,N_22122,N_20237);
nor U23644 (N_23644,N_21674,N_21708);
and U23645 (N_23645,N_21760,N_22143);
xnor U23646 (N_23646,N_21639,N_21934);
xor U23647 (N_23647,N_21780,N_21219);
nor U23648 (N_23648,N_22006,N_21224);
nor U23649 (N_23649,N_20465,N_21580);
and U23650 (N_23650,N_22102,N_22221);
xnor U23651 (N_23651,N_22463,N_21302);
xor U23652 (N_23652,N_20391,N_20660);
nor U23653 (N_23653,N_20877,N_21063);
or U23654 (N_23654,N_20845,N_20142);
xnor U23655 (N_23655,N_21170,N_20196);
xnor U23656 (N_23656,N_20436,N_20320);
or U23657 (N_23657,N_20431,N_20117);
nor U23658 (N_23658,N_22416,N_22072);
or U23659 (N_23659,N_20727,N_20211);
xnor U23660 (N_23660,N_22412,N_20291);
xor U23661 (N_23661,N_20106,N_20312);
and U23662 (N_23662,N_20834,N_22274);
xor U23663 (N_23663,N_21967,N_22346);
nor U23664 (N_23664,N_21038,N_22290);
nor U23665 (N_23665,N_21099,N_21857);
or U23666 (N_23666,N_22252,N_21321);
or U23667 (N_23667,N_20071,N_21449);
or U23668 (N_23668,N_22085,N_21045);
and U23669 (N_23669,N_22178,N_20569);
xor U23670 (N_23670,N_21283,N_21820);
xnor U23671 (N_23671,N_22379,N_20838);
and U23672 (N_23672,N_22190,N_20913);
nand U23673 (N_23673,N_21212,N_20087);
and U23674 (N_23674,N_21369,N_21683);
nor U23675 (N_23675,N_21417,N_20376);
and U23676 (N_23676,N_21521,N_22120);
nand U23677 (N_23677,N_21713,N_22215);
or U23678 (N_23678,N_22155,N_20653);
nor U23679 (N_23679,N_22342,N_21916);
xor U23680 (N_23680,N_21218,N_21957);
nor U23681 (N_23681,N_20352,N_22485);
and U23682 (N_23682,N_21353,N_21254);
xor U23683 (N_23683,N_20204,N_22262);
nand U23684 (N_23684,N_22360,N_21527);
nor U23685 (N_23685,N_21273,N_20193);
nand U23686 (N_23686,N_22312,N_20974);
nor U23687 (N_23687,N_20181,N_21025);
or U23688 (N_23688,N_20811,N_20124);
and U23689 (N_23689,N_22194,N_20828);
nand U23690 (N_23690,N_20002,N_21085);
nand U23691 (N_23691,N_21811,N_20520);
or U23692 (N_23692,N_20373,N_22429);
nor U23693 (N_23693,N_21249,N_22297);
xnor U23694 (N_23694,N_20658,N_20553);
nor U23695 (N_23695,N_21816,N_21199);
nand U23696 (N_23696,N_20328,N_20245);
xnor U23697 (N_23697,N_20179,N_21215);
and U23698 (N_23698,N_21287,N_20301);
nand U23699 (N_23699,N_22438,N_20778);
nand U23700 (N_23700,N_21991,N_22142);
and U23701 (N_23701,N_20173,N_20667);
and U23702 (N_23702,N_20305,N_20970);
and U23703 (N_23703,N_22244,N_21806);
nand U23704 (N_23704,N_22263,N_20858);
and U23705 (N_23705,N_20614,N_21798);
or U23706 (N_23706,N_21436,N_21900);
and U23707 (N_23707,N_21443,N_21975);
nand U23708 (N_23708,N_20665,N_21986);
or U23709 (N_23709,N_21168,N_20689);
xor U23710 (N_23710,N_20402,N_21550);
nor U23711 (N_23711,N_20413,N_21222);
nor U23712 (N_23712,N_21777,N_21868);
nand U23713 (N_23713,N_22177,N_21435);
nand U23714 (N_23714,N_21860,N_20162);
and U23715 (N_23715,N_21508,N_21263);
xnor U23716 (N_23716,N_20827,N_21768);
and U23717 (N_23717,N_20441,N_22141);
nor U23718 (N_23718,N_21104,N_21372);
nand U23719 (N_23719,N_20949,N_20891);
nor U23720 (N_23720,N_22145,N_20407);
xor U23721 (N_23721,N_20706,N_21176);
xnor U23722 (N_23722,N_21850,N_20708);
and U23723 (N_23723,N_21925,N_20309);
or U23724 (N_23724,N_21996,N_22154);
xor U23725 (N_23725,N_20996,N_20018);
nand U23726 (N_23726,N_21952,N_21770);
or U23727 (N_23727,N_20170,N_21738);
nand U23728 (N_23728,N_21034,N_22214);
nor U23729 (N_23729,N_20770,N_20058);
and U23730 (N_23730,N_20899,N_21761);
xor U23731 (N_23731,N_21476,N_20386);
and U23732 (N_23732,N_20926,N_20636);
xnor U23733 (N_23733,N_20038,N_22256);
or U23734 (N_23734,N_20346,N_20783);
nand U23735 (N_23735,N_20578,N_22496);
and U23736 (N_23736,N_20808,N_22227);
nand U23737 (N_23737,N_21120,N_22459);
or U23738 (N_23738,N_21363,N_21472);
nand U23739 (N_23739,N_22125,N_21792);
xor U23740 (N_23740,N_20390,N_22452);
nand U23741 (N_23741,N_20392,N_20607);
nor U23742 (N_23742,N_21102,N_22293);
and U23743 (N_23743,N_20602,N_20788);
and U23744 (N_23744,N_22469,N_20017);
or U23745 (N_23745,N_20311,N_21606);
nor U23746 (N_23746,N_20281,N_20681);
xnor U23747 (N_23747,N_20886,N_22246);
or U23748 (N_23748,N_22115,N_21423);
or U23749 (N_23749,N_22127,N_20531);
nand U23750 (N_23750,N_21149,N_20438);
or U23751 (N_23751,N_20204,N_20448);
xnor U23752 (N_23752,N_20157,N_20747);
nand U23753 (N_23753,N_22366,N_21919);
nor U23754 (N_23754,N_22430,N_22145);
xor U23755 (N_23755,N_22198,N_22233);
and U23756 (N_23756,N_20072,N_22086);
nand U23757 (N_23757,N_20510,N_20701);
nand U23758 (N_23758,N_21959,N_20783);
nand U23759 (N_23759,N_22474,N_21794);
xor U23760 (N_23760,N_22251,N_21334);
or U23761 (N_23761,N_21613,N_20723);
or U23762 (N_23762,N_20062,N_20780);
and U23763 (N_23763,N_20517,N_21906);
or U23764 (N_23764,N_20960,N_20272);
and U23765 (N_23765,N_20469,N_22102);
and U23766 (N_23766,N_21217,N_20742);
and U23767 (N_23767,N_22133,N_20882);
xor U23768 (N_23768,N_22107,N_22462);
or U23769 (N_23769,N_20516,N_21420);
nor U23770 (N_23770,N_21281,N_20329);
nor U23771 (N_23771,N_20902,N_20105);
nand U23772 (N_23772,N_21495,N_20535);
xor U23773 (N_23773,N_20931,N_21521);
or U23774 (N_23774,N_21928,N_22482);
or U23775 (N_23775,N_21486,N_22094);
nand U23776 (N_23776,N_21817,N_21786);
nor U23777 (N_23777,N_20212,N_22294);
nor U23778 (N_23778,N_20168,N_21059);
and U23779 (N_23779,N_22482,N_20761);
and U23780 (N_23780,N_21783,N_21087);
xnor U23781 (N_23781,N_21494,N_21482);
or U23782 (N_23782,N_22379,N_22064);
xor U23783 (N_23783,N_21289,N_22401);
xnor U23784 (N_23784,N_21864,N_22305);
xor U23785 (N_23785,N_20843,N_20311);
xnor U23786 (N_23786,N_22227,N_21955);
xnor U23787 (N_23787,N_21992,N_20311);
xor U23788 (N_23788,N_22136,N_21612);
and U23789 (N_23789,N_20754,N_22299);
xnor U23790 (N_23790,N_22259,N_21105);
and U23791 (N_23791,N_21054,N_20530);
and U23792 (N_23792,N_20933,N_22332);
nand U23793 (N_23793,N_20519,N_21386);
and U23794 (N_23794,N_21485,N_22101);
and U23795 (N_23795,N_21344,N_22305);
or U23796 (N_23796,N_20595,N_20322);
nand U23797 (N_23797,N_21567,N_21953);
or U23798 (N_23798,N_21889,N_22490);
or U23799 (N_23799,N_21464,N_21253);
xor U23800 (N_23800,N_20955,N_21392);
and U23801 (N_23801,N_20938,N_21050);
and U23802 (N_23802,N_21075,N_22035);
or U23803 (N_23803,N_21030,N_21236);
nand U23804 (N_23804,N_20391,N_21305);
xnor U23805 (N_23805,N_21730,N_21739);
xor U23806 (N_23806,N_21603,N_21750);
nand U23807 (N_23807,N_21415,N_21580);
nor U23808 (N_23808,N_22490,N_22368);
nand U23809 (N_23809,N_20852,N_22421);
and U23810 (N_23810,N_22301,N_20109);
xor U23811 (N_23811,N_20763,N_20464);
and U23812 (N_23812,N_20824,N_22225);
nand U23813 (N_23813,N_20181,N_21731);
and U23814 (N_23814,N_22300,N_22251);
nor U23815 (N_23815,N_22159,N_20481);
and U23816 (N_23816,N_22068,N_21724);
nand U23817 (N_23817,N_21027,N_21289);
or U23818 (N_23818,N_20966,N_20050);
nor U23819 (N_23819,N_21427,N_20765);
or U23820 (N_23820,N_20595,N_21710);
and U23821 (N_23821,N_22311,N_20722);
or U23822 (N_23822,N_21747,N_21902);
or U23823 (N_23823,N_20639,N_20087);
nand U23824 (N_23824,N_20734,N_21874);
nand U23825 (N_23825,N_22203,N_20512);
nand U23826 (N_23826,N_22468,N_21543);
or U23827 (N_23827,N_20804,N_21443);
nand U23828 (N_23828,N_21366,N_20651);
xnor U23829 (N_23829,N_20182,N_20561);
nand U23830 (N_23830,N_20605,N_21143);
nand U23831 (N_23831,N_21255,N_20609);
and U23832 (N_23832,N_21919,N_21449);
nand U23833 (N_23833,N_20935,N_22242);
xor U23834 (N_23834,N_21220,N_21226);
and U23835 (N_23835,N_21595,N_20307);
and U23836 (N_23836,N_20726,N_21210);
xor U23837 (N_23837,N_20100,N_20826);
xnor U23838 (N_23838,N_20898,N_21794);
nor U23839 (N_23839,N_20883,N_21443);
or U23840 (N_23840,N_21425,N_21343);
nand U23841 (N_23841,N_20911,N_21449);
nor U23842 (N_23842,N_20782,N_21134);
or U23843 (N_23843,N_21035,N_21956);
and U23844 (N_23844,N_20840,N_20500);
nor U23845 (N_23845,N_21490,N_21516);
and U23846 (N_23846,N_22227,N_21316);
or U23847 (N_23847,N_21961,N_20926);
or U23848 (N_23848,N_20876,N_21696);
nand U23849 (N_23849,N_22495,N_20159);
nand U23850 (N_23850,N_22104,N_21898);
nor U23851 (N_23851,N_21029,N_20889);
nand U23852 (N_23852,N_21208,N_20996);
and U23853 (N_23853,N_21221,N_20874);
nor U23854 (N_23854,N_20108,N_20573);
nor U23855 (N_23855,N_20460,N_20852);
or U23856 (N_23856,N_20926,N_20063);
xnor U23857 (N_23857,N_21368,N_20218);
xor U23858 (N_23858,N_20059,N_21510);
nor U23859 (N_23859,N_20721,N_22089);
xnor U23860 (N_23860,N_20172,N_21476);
or U23861 (N_23861,N_21408,N_21905);
nand U23862 (N_23862,N_22217,N_20348);
nor U23863 (N_23863,N_20649,N_20910);
xor U23864 (N_23864,N_22363,N_21658);
and U23865 (N_23865,N_20584,N_21314);
nor U23866 (N_23866,N_20812,N_21660);
nor U23867 (N_23867,N_20476,N_20247);
nand U23868 (N_23868,N_22430,N_20058);
or U23869 (N_23869,N_21840,N_20090);
nand U23870 (N_23870,N_20833,N_21892);
nand U23871 (N_23871,N_20238,N_21857);
nor U23872 (N_23872,N_21312,N_21106);
nand U23873 (N_23873,N_20612,N_20277);
and U23874 (N_23874,N_21396,N_20631);
nor U23875 (N_23875,N_20289,N_21516);
xnor U23876 (N_23876,N_21477,N_20787);
xor U23877 (N_23877,N_22124,N_22248);
xor U23878 (N_23878,N_22245,N_20934);
and U23879 (N_23879,N_22264,N_22382);
nor U23880 (N_23880,N_20925,N_21821);
and U23881 (N_23881,N_21135,N_20091);
or U23882 (N_23882,N_20106,N_20564);
nand U23883 (N_23883,N_21299,N_21438);
xor U23884 (N_23884,N_20582,N_22311);
and U23885 (N_23885,N_22032,N_22335);
xor U23886 (N_23886,N_21828,N_20857);
and U23887 (N_23887,N_20985,N_21381);
xor U23888 (N_23888,N_22298,N_21726);
nor U23889 (N_23889,N_20058,N_20145);
nand U23890 (N_23890,N_21764,N_20858);
nor U23891 (N_23891,N_22164,N_20045);
nor U23892 (N_23892,N_20433,N_20783);
and U23893 (N_23893,N_20445,N_21489);
nor U23894 (N_23894,N_21036,N_22091);
nor U23895 (N_23895,N_20036,N_20104);
and U23896 (N_23896,N_20944,N_20480);
and U23897 (N_23897,N_20793,N_22128);
nand U23898 (N_23898,N_20025,N_21471);
nand U23899 (N_23899,N_21015,N_20184);
xnor U23900 (N_23900,N_22093,N_22011);
xnor U23901 (N_23901,N_21799,N_20303);
xor U23902 (N_23902,N_20452,N_21816);
and U23903 (N_23903,N_21693,N_21523);
nand U23904 (N_23904,N_20370,N_20584);
xnor U23905 (N_23905,N_21943,N_21132);
nand U23906 (N_23906,N_20031,N_20557);
or U23907 (N_23907,N_22395,N_21149);
nor U23908 (N_23908,N_22105,N_20337);
nor U23909 (N_23909,N_21240,N_20929);
and U23910 (N_23910,N_20767,N_20186);
or U23911 (N_23911,N_21654,N_21387);
or U23912 (N_23912,N_21951,N_22086);
or U23913 (N_23913,N_21798,N_20640);
nor U23914 (N_23914,N_22391,N_20165);
nor U23915 (N_23915,N_20449,N_21804);
or U23916 (N_23916,N_20141,N_20390);
nor U23917 (N_23917,N_21439,N_21742);
nor U23918 (N_23918,N_22158,N_22168);
nor U23919 (N_23919,N_22226,N_20634);
xor U23920 (N_23920,N_20731,N_21530);
or U23921 (N_23921,N_21591,N_21316);
nand U23922 (N_23922,N_20420,N_21543);
nor U23923 (N_23923,N_21836,N_21185);
nor U23924 (N_23924,N_21966,N_22449);
xnor U23925 (N_23925,N_21460,N_20001);
and U23926 (N_23926,N_22294,N_20582);
or U23927 (N_23927,N_21961,N_20228);
nor U23928 (N_23928,N_20824,N_21017);
and U23929 (N_23929,N_20498,N_21164);
and U23930 (N_23930,N_20788,N_20681);
and U23931 (N_23931,N_21826,N_20650);
or U23932 (N_23932,N_21087,N_20719);
nor U23933 (N_23933,N_22075,N_21996);
nand U23934 (N_23934,N_21736,N_20994);
xor U23935 (N_23935,N_20102,N_21865);
and U23936 (N_23936,N_22482,N_20463);
nand U23937 (N_23937,N_20995,N_21363);
xor U23938 (N_23938,N_20244,N_21752);
and U23939 (N_23939,N_22154,N_21020);
nand U23940 (N_23940,N_21782,N_21126);
nor U23941 (N_23941,N_22033,N_22148);
nand U23942 (N_23942,N_21595,N_21891);
or U23943 (N_23943,N_21658,N_21826);
xnor U23944 (N_23944,N_21684,N_20075);
nor U23945 (N_23945,N_20123,N_22020);
nand U23946 (N_23946,N_20591,N_20886);
and U23947 (N_23947,N_21499,N_20241);
xnor U23948 (N_23948,N_22142,N_21409);
or U23949 (N_23949,N_20070,N_21324);
and U23950 (N_23950,N_21265,N_21418);
xnor U23951 (N_23951,N_21083,N_20192);
or U23952 (N_23952,N_21916,N_21042);
xnor U23953 (N_23953,N_21090,N_21294);
or U23954 (N_23954,N_21784,N_21493);
or U23955 (N_23955,N_22444,N_22075);
or U23956 (N_23956,N_21895,N_20884);
and U23957 (N_23957,N_20051,N_22243);
and U23958 (N_23958,N_20694,N_22469);
or U23959 (N_23959,N_20920,N_20515);
or U23960 (N_23960,N_22491,N_22282);
and U23961 (N_23961,N_20296,N_22200);
xor U23962 (N_23962,N_22047,N_21079);
and U23963 (N_23963,N_21627,N_22184);
and U23964 (N_23964,N_21976,N_22230);
nor U23965 (N_23965,N_20581,N_21130);
or U23966 (N_23966,N_21129,N_22179);
and U23967 (N_23967,N_21906,N_20570);
or U23968 (N_23968,N_22006,N_21506);
and U23969 (N_23969,N_20602,N_22119);
nand U23970 (N_23970,N_20438,N_22449);
and U23971 (N_23971,N_21256,N_22438);
or U23972 (N_23972,N_20055,N_20685);
nand U23973 (N_23973,N_22397,N_21525);
nor U23974 (N_23974,N_22434,N_20897);
nand U23975 (N_23975,N_21734,N_20412);
nand U23976 (N_23976,N_21109,N_21698);
nand U23977 (N_23977,N_20225,N_21858);
nand U23978 (N_23978,N_21772,N_22303);
and U23979 (N_23979,N_22367,N_22258);
nand U23980 (N_23980,N_21785,N_21627);
nor U23981 (N_23981,N_20640,N_20362);
nand U23982 (N_23982,N_20825,N_20985);
xnor U23983 (N_23983,N_21397,N_22307);
xor U23984 (N_23984,N_21950,N_22131);
nand U23985 (N_23985,N_22402,N_21193);
xor U23986 (N_23986,N_20308,N_21749);
nor U23987 (N_23987,N_20844,N_20078);
nand U23988 (N_23988,N_21399,N_20202);
xor U23989 (N_23989,N_21846,N_22305);
or U23990 (N_23990,N_21880,N_21732);
nor U23991 (N_23991,N_21176,N_20649);
xor U23992 (N_23992,N_22254,N_21206);
or U23993 (N_23993,N_20853,N_21282);
and U23994 (N_23994,N_21407,N_21459);
or U23995 (N_23995,N_20669,N_21501);
xor U23996 (N_23996,N_20378,N_21069);
nand U23997 (N_23997,N_21250,N_21670);
or U23998 (N_23998,N_21221,N_21864);
nor U23999 (N_23999,N_21040,N_21428);
xor U24000 (N_24000,N_20143,N_21685);
xor U24001 (N_24001,N_20226,N_21869);
xnor U24002 (N_24002,N_22042,N_22068);
nand U24003 (N_24003,N_20280,N_21964);
xnor U24004 (N_24004,N_22050,N_20581);
or U24005 (N_24005,N_21928,N_21420);
or U24006 (N_24006,N_21455,N_21910);
xor U24007 (N_24007,N_20508,N_20566);
or U24008 (N_24008,N_20251,N_21157);
and U24009 (N_24009,N_20655,N_22172);
or U24010 (N_24010,N_22413,N_21262);
nand U24011 (N_24011,N_20505,N_20351);
nor U24012 (N_24012,N_20968,N_21574);
nand U24013 (N_24013,N_20005,N_21049);
nor U24014 (N_24014,N_22439,N_20171);
and U24015 (N_24015,N_20608,N_22439);
nand U24016 (N_24016,N_22158,N_20240);
xor U24017 (N_24017,N_22195,N_20693);
xor U24018 (N_24018,N_20197,N_21629);
and U24019 (N_24019,N_20533,N_20109);
xor U24020 (N_24020,N_22403,N_20034);
or U24021 (N_24021,N_20314,N_20856);
nand U24022 (N_24022,N_20737,N_21983);
and U24023 (N_24023,N_22497,N_21957);
xnor U24024 (N_24024,N_20878,N_22060);
xnor U24025 (N_24025,N_21749,N_22054);
nor U24026 (N_24026,N_21675,N_21114);
and U24027 (N_24027,N_22078,N_20108);
xor U24028 (N_24028,N_22043,N_20459);
xor U24029 (N_24029,N_20407,N_20269);
xor U24030 (N_24030,N_20266,N_20950);
or U24031 (N_24031,N_22060,N_21096);
and U24032 (N_24032,N_21702,N_20819);
nor U24033 (N_24033,N_21198,N_20619);
xor U24034 (N_24034,N_20608,N_21139);
nor U24035 (N_24035,N_20296,N_22197);
and U24036 (N_24036,N_21538,N_21129);
or U24037 (N_24037,N_20028,N_21721);
or U24038 (N_24038,N_21750,N_21475);
or U24039 (N_24039,N_20519,N_22321);
or U24040 (N_24040,N_21499,N_21543);
nor U24041 (N_24041,N_21981,N_21664);
nand U24042 (N_24042,N_20733,N_21616);
and U24043 (N_24043,N_21411,N_21639);
and U24044 (N_24044,N_20488,N_22373);
xor U24045 (N_24045,N_22423,N_20928);
nand U24046 (N_24046,N_22174,N_21288);
or U24047 (N_24047,N_21243,N_21573);
nor U24048 (N_24048,N_20687,N_20161);
xnor U24049 (N_24049,N_20889,N_20298);
nand U24050 (N_24050,N_20289,N_22273);
and U24051 (N_24051,N_21763,N_21893);
nand U24052 (N_24052,N_21152,N_21062);
or U24053 (N_24053,N_20891,N_20813);
and U24054 (N_24054,N_21367,N_22480);
nor U24055 (N_24055,N_22218,N_22425);
xnor U24056 (N_24056,N_20594,N_22009);
xor U24057 (N_24057,N_22201,N_20750);
xor U24058 (N_24058,N_20977,N_21475);
xnor U24059 (N_24059,N_20751,N_21666);
nor U24060 (N_24060,N_22001,N_22396);
nor U24061 (N_24061,N_20992,N_21411);
xnor U24062 (N_24062,N_20768,N_22404);
xnor U24063 (N_24063,N_21224,N_21016);
nor U24064 (N_24064,N_21028,N_22402);
nor U24065 (N_24065,N_21942,N_20912);
nand U24066 (N_24066,N_20711,N_21575);
nand U24067 (N_24067,N_20748,N_22104);
nand U24068 (N_24068,N_21254,N_22491);
xnor U24069 (N_24069,N_20947,N_20923);
xnor U24070 (N_24070,N_21980,N_22352);
nor U24071 (N_24071,N_21373,N_21515);
nor U24072 (N_24072,N_20075,N_21278);
or U24073 (N_24073,N_21786,N_22244);
nand U24074 (N_24074,N_21305,N_21449);
xor U24075 (N_24075,N_20840,N_20713);
and U24076 (N_24076,N_21800,N_21611);
nand U24077 (N_24077,N_20269,N_21569);
xnor U24078 (N_24078,N_22090,N_22447);
and U24079 (N_24079,N_22053,N_22231);
xnor U24080 (N_24080,N_20751,N_21323);
xor U24081 (N_24081,N_21019,N_21588);
xnor U24082 (N_24082,N_20193,N_20271);
nor U24083 (N_24083,N_20412,N_22079);
and U24084 (N_24084,N_20138,N_20076);
or U24085 (N_24085,N_20869,N_21596);
or U24086 (N_24086,N_22195,N_20999);
or U24087 (N_24087,N_20675,N_21023);
and U24088 (N_24088,N_21766,N_21785);
nor U24089 (N_24089,N_22217,N_20053);
or U24090 (N_24090,N_22064,N_20794);
or U24091 (N_24091,N_22204,N_20809);
or U24092 (N_24092,N_20613,N_21209);
xor U24093 (N_24093,N_21162,N_22259);
nor U24094 (N_24094,N_21182,N_21205);
nand U24095 (N_24095,N_21588,N_22219);
nand U24096 (N_24096,N_21907,N_20615);
nor U24097 (N_24097,N_21194,N_21149);
nor U24098 (N_24098,N_20333,N_20322);
and U24099 (N_24099,N_20917,N_20931);
nand U24100 (N_24100,N_21410,N_21574);
xor U24101 (N_24101,N_22454,N_20294);
and U24102 (N_24102,N_20468,N_21062);
and U24103 (N_24103,N_22178,N_22211);
or U24104 (N_24104,N_20783,N_21364);
and U24105 (N_24105,N_20830,N_21988);
and U24106 (N_24106,N_22062,N_21975);
or U24107 (N_24107,N_20450,N_21843);
nand U24108 (N_24108,N_22451,N_20316);
nand U24109 (N_24109,N_20289,N_20594);
and U24110 (N_24110,N_20382,N_20505);
xnor U24111 (N_24111,N_22475,N_22321);
nand U24112 (N_24112,N_21264,N_21068);
xor U24113 (N_24113,N_20707,N_20786);
nor U24114 (N_24114,N_21410,N_21038);
nand U24115 (N_24115,N_20582,N_21531);
nand U24116 (N_24116,N_20687,N_21839);
and U24117 (N_24117,N_20892,N_21453);
xor U24118 (N_24118,N_21083,N_21073);
or U24119 (N_24119,N_20937,N_21611);
nor U24120 (N_24120,N_21608,N_21929);
nand U24121 (N_24121,N_21324,N_21563);
xnor U24122 (N_24122,N_21391,N_22344);
nand U24123 (N_24123,N_21892,N_20143);
xor U24124 (N_24124,N_21395,N_22458);
xnor U24125 (N_24125,N_20891,N_20015);
nand U24126 (N_24126,N_21389,N_21275);
xor U24127 (N_24127,N_21451,N_21181);
nor U24128 (N_24128,N_22313,N_20453);
nor U24129 (N_24129,N_20445,N_20314);
and U24130 (N_24130,N_20107,N_21627);
xor U24131 (N_24131,N_21331,N_20505);
xor U24132 (N_24132,N_20947,N_20292);
and U24133 (N_24133,N_21642,N_20936);
nor U24134 (N_24134,N_20750,N_21590);
and U24135 (N_24135,N_20988,N_20867);
xnor U24136 (N_24136,N_21100,N_21216);
and U24137 (N_24137,N_20026,N_20984);
and U24138 (N_24138,N_20228,N_20396);
nor U24139 (N_24139,N_22278,N_21236);
nor U24140 (N_24140,N_20987,N_21724);
or U24141 (N_24141,N_22257,N_21009);
or U24142 (N_24142,N_20835,N_20615);
or U24143 (N_24143,N_21791,N_20049);
and U24144 (N_24144,N_20357,N_22245);
and U24145 (N_24145,N_20852,N_21331);
or U24146 (N_24146,N_22007,N_20171);
xnor U24147 (N_24147,N_21479,N_21392);
and U24148 (N_24148,N_21572,N_21820);
or U24149 (N_24149,N_20331,N_21592);
nor U24150 (N_24150,N_20199,N_20776);
and U24151 (N_24151,N_21452,N_21804);
nand U24152 (N_24152,N_21752,N_20626);
nand U24153 (N_24153,N_20652,N_20222);
xor U24154 (N_24154,N_20613,N_20142);
and U24155 (N_24155,N_20922,N_20916);
or U24156 (N_24156,N_20740,N_22397);
or U24157 (N_24157,N_20805,N_21718);
xnor U24158 (N_24158,N_20744,N_20834);
and U24159 (N_24159,N_20433,N_20690);
or U24160 (N_24160,N_21109,N_20893);
or U24161 (N_24161,N_20864,N_20915);
or U24162 (N_24162,N_21596,N_21156);
nand U24163 (N_24163,N_21605,N_21554);
xnor U24164 (N_24164,N_21428,N_22134);
and U24165 (N_24165,N_20879,N_20922);
nand U24166 (N_24166,N_20364,N_20601);
nand U24167 (N_24167,N_21730,N_20833);
nand U24168 (N_24168,N_21896,N_21517);
xor U24169 (N_24169,N_20702,N_20633);
or U24170 (N_24170,N_22487,N_20260);
nand U24171 (N_24171,N_22426,N_21827);
xor U24172 (N_24172,N_21072,N_21391);
nor U24173 (N_24173,N_20652,N_21882);
or U24174 (N_24174,N_21926,N_20494);
nor U24175 (N_24175,N_20983,N_20730);
or U24176 (N_24176,N_22444,N_20850);
or U24177 (N_24177,N_21382,N_20420);
and U24178 (N_24178,N_20193,N_22048);
or U24179 (N_24179,N_21535,N_22337);
nand U24180 (N_24180,N_21170,N_20390);
and U24181 (N_24181,N_22061,N_20919);
and U24182 (N_24182,N_21583,N_22314);
nand U24183 (N_24183,N_20985,N_20673);
or U24184 (N_24184,N_20893,N_20269);
nor U24185 (N_24185,N_21776,N_20736);
nor U24186 (N_24186,N_21854,N_21636);
xor U24187 (N_24187,N_22352,N_22263);
nor U24188 (N_24188,N_21601,N_20234);
nand U24189 (N_24189,N_21964,N_20663);
and U24190 (N_24190,N_20785,N_22398);
or U24191 (N_24191,N_20279,N_21250);
xor U24192 (N_24192,N_22465,N_21460);
or U24193 (N_24193,N_21724,N_22248);
xnor U24194 (N_24194,N_20735,N_20683);
nand U24195 (N_24195,N_21139,N_21622);
nand U24196 (N_24196,N_21835,N_21135);
xnor U24197 (N_24197,N_20704,N_22217);
xor U24198 (N_24198,N_21568,N_21217);
xor U24199 (N_24199,N_21518,N_20715);
xnor U24200 (N_24200,N_20684,N_22292);
nor U24201 (N_24201,N_21573,N_21750);
xor U24202 (N_24202,N_21658,N_21934);
nand U24203 (N_24203,N_20067,N_21981);
nand U24204 (N_24204,N_22138,N_20745);
xnor U24205 (N_24205,N_22383,N_20137);
and U24206 (N_24206,N_21373,N_21439);
or U24207 (N_24207,N_22178,N_22248);
xor U24208 (N_24208,N_20169,N_21478);
xor U24209 (N_24209,N_21222,N_21874);
and U24210 (N_24210,N_21101,N_22079);
xor U24211 (N_24211,N_21908,N_21901);
or U24212 (N_24212,N_21441,N_22067);
xor U24213 (N_24213,N_21702,N_21258);
nor U24214 (N_24214,N_20283,N_20911);
and U24215 (N_24215,N_21189,N_22308);
or U24216 (N_24216,N_21682,N_21961);
and U24217 (N_24217,N_21842,N_20242);
or U24218 (N_24218,N_20006,N_20305);
and U24219 (N_24219,N_20869,N_21932);
and U24220 (N_24220,N_20381,N_22300);
nor U24221 (N_24221,N_20426,N_22326);
nand U24222 (N_24222,N_21309,N_20592);
nor U24223 (N_24223,N_21808,N_20196);
and U24224 (N_24224,N_21888,N_20044);
and U24225 (N_24225,N_20571,N_22420);
or U24226 (N_24226,N_20350,N_21744);
nand U24227 (N_24227,N_20171,N_20515);
nand U24228 (N_24228,N_21835,N_22347);
nor U24229 (N_24229,N_20506,N_22340);
and U24230 (N_24230,N_22254,N_22413);
xor U24231 (N_24231,N_20546,N_21730);
nand U24232 (N_24232,N_21612,N_21092);
and U24233 (N_24233,N_22367,N_21506);
or U24234 (N_24234,N_21918,N_21710);
and U24235 (N_24235,N_21094,N_21616);
xnor U24236 (N_24236,N_20599,N_22323);
nor U24237 (N_24237,N_22460,N_20700);
or U24238 (N_24238,N_21042,N_20363);
nand U24239 (N_24239,N_21663,N_22363);
nor U24240 (N_24240,N_21745,N_21831);
nor U24241 (N_24241,N_21885,N_21136);
xor U24242 (N_24242,N_20837,N_20920);
nand U24243 (N_24243,N_21393,N_20752);
nand U24244 (N_24244,N_21015,N_20786);
xor U24245 (N_24245,N_20352,N_21079);
nand U24246 (N_24246,N_22296,N_20093);
xnor U24247 (N_24247,N_20878,N_22117);
and U24248 (N_24248,N_22019,N_21059);
nand U24249 (N_24249,N_20480,N_21462);
or U24250 (N_24250,N_22115,N_20751);
and U24251 (N_24251,N_21524,N_21210);
and U24252 (N_24252,N_20729,N_21220);
nor U24253 (N_24253,N_22021,N_20668);
nor U24254 (N_24254,N_21373,N_20620);
xnor U24255 (N_24255,N_20519,N_22312);
nand U24256 (N_24256,N_21213,N_20878);
nand U24257 (N_24257,N_22452,N_21922);
xor U24258 (N_24258,N_22002,N_22003);
and U24259 (N_24259,N_20080,N_20411);
xor U24260 (N_24260,N_21316,N_21526);
nor U24261 (N_24261,N_22065,N_21539);
xnor U24262 (N_24262,N_21220,N_21416);
or U24263 (N_24263,N_21746,N_21636);
nand U24264 (N_24264,N_22066,N_20691);
nor U24265 (N_24265,N_21680,N_22355);
nor U24266 (N_24266,N_21447,N_20775);
nand U24267 (N_24267,N_20093,N_22403);
or U24268 (N_24268,N_22365,N_22150);
nor U24269 (N_24269,N_21697,N_21975);
nand U24270 (N_24270,N_20686,N_22316);
and U24271 (N_24271,N_21475,N_20353);
nand U24272 (N_24272,N_20642,N_20456);
and U24273 (N_24273,N_20100,N_22402);
xnor U24274 (N_24274,N_21520,N_22312);
nor U24275 (N_24275,N_21925,N_22186);
or U24276 (N_24276,N_21035,N_21301);
xnor U24277 (N_24277,N_20153,N_21390);
nor U24278 (N_24278,N_20234,N_21191);
nor U24279 (N_24279,N_21608,N_22421);
and U24280 (N_24280,N_20553,N_21734);
or U24281 (N_24281,N_21367,N_21976);
nor U24282 (N_24282,N_20104,N_22161);
and U24283 (N_24283,N_20155,N_21246);
nand U24284 (N_24284,N_22303,N_20602);
or U24285 (N_24285,N_21390,N_21814);
nand U24286 (N_24286,N_22395,N_20761);
and U24287 (N_24287,N_20708,N_20510);
nor U24288 (N_24288,N_21855,N_20705);
or U24289 (N_24289,N_20006,N_20845);
or U24290 (N_24290,N_20687,N_21101);
or U24291 (N_24291,N_21120,N_21495);
xor U24292 (N_24292,N_22114,N_22461);
nor U24293 (N_24293,N_21182,N_21565);
xnor U24294 (N_24294,N_21537,N_22174);
nand U24295 (N_24295,N_20656,N_22181);
and U24296 (N_24296,N_21517,N_20736);
and U24297 (N_24297,N_20376,N_20894);
or U24298 (N_24298,N_22325,N_22467);
or U24299 (N_24299,N_21155,N_21540);
xnor U24300 (N_24300,N_20237,N_21924);
and U24301 (N_24301,N_20265,N_21182);
xnor U24302 (N_24302,N_21240,N_20683);
or U24303 (N_24303,N_20697,N_22086);
and U24304 (N_24304,N_21661,N_21549);
nor U24305 (N_24305,N_20375,N_21994);
nand U24306 (N_24306,N_21262,N_21767);
or U24307 (N_24307,N_21763,N_20561);
xor U24308 (N_24308,N_21055,N_22359);
and U24309 (N_24309,N_21543,N_20447);
nor U24310 (N_24310,N_21886,N_20585);
xnor U24311 (N_24311,N_22129,N_20760);
and U24312 (N_24312,N_22434,N_20572);
nor U24313 (N_24313,N_22397,N_22024);
nor U24314 (N_24314,N_20292,N_21053);
nor U24315 (N_24315,N_21388,N_20841);
and U24316 (N_24316,N_22022,N_22359);
xor U24317 (N_24317,N_21561,N_20200);
nor U24318 (N_24318,N_22310,N_21500);
nand U24319 (N_24319,N_20993,N_20344);
nand U24320 (N_24320,N_22301,N_21564);
and U24321 (N_24321,N_22297,N_20295);
and U24322 (N_24322,N_21373,N_21590);
or U24323 (N_24323,N_20079,N_20262);
nor U24324 (N_24324,N_20307,N_20244);
and U24325 (N_24325,N_22167,N_20387);
nand U24326 (N_24326,N_21762,N_20370);
nor U24327 (N_24327,N_20803,N_22023);
nor U24328 (N_24328,N_21201,N_20513);
or U24329 (N_24329,N_20611,N_20554);
or U24330 (N_24330,N_22407,N_20784);
xor U24331 (N_24331,N_20734,N_20790);
nor U24332 (N_24332,N_21184,N_20928);
and U24333 (N_24333,N_22413,N_21028);
xor U24334 (N_24334,N_20334,N_20470);
and U24335 (N_24335,N_22295,N_22178);
nand U24336 (N_24336,N_20717,N_20227);
nand U24337 (N_24337,N_21145,N_20851);
and U24338 (N_24338,N_20661,N_22132);
nand U24339 (N_24339,N_21685,N_21153);
xor U24340 (N_24340,N_20230,N_21118);
xnor U24341 (N_24341,N_21061,N_22380);
xor U24342 (N_24342,N_21443,N_20750);
nand U24343 (N_24343,N_21549,N_22175);
or U24344 (N_24344,N_21884,N_21094);
or U24345 (N_24345,N_20509,N_20093);
and U24346 (N_24346,N_20331,N_20741);
nor U24347 (N_24347,N_22057,N_20639);
xnor U24348 (N_24348,N_21872,N_21686);
xor U24349 (N_24349,N_21467,N_20483);
and U24350 (N_24350,N_21337,N_22302);
xnor U24351 (N_24351,N_20132,N_20751);
xor U24352 (N_24352,N_22045,N_20424);
nand U24353 (N_24353,N_22443,N_20444);
and U24354 (N_24354,N_21548,N_21560);
nor U24355 (N_24355,N_20466,N_21978);
nor U24356 (N_24356,N_20757,N_21806);
xnor U24357 (N_24357,N_21549,N_21122);
nor U24358 (N_24358,N_20105,N_22070);
and U24359 (N_24359,N_21387,N_22476);
nand U24360 (N_24360,N_20641,N_21117);
nand U24361 (N_24361,N_21509,N_21208);
nor U24362 (N_24362,N_21869,N_22132);
nand U24363 (N_24363,N_21439,N_20511);
or U24364 (N_24364,N_20901,N_21118);
or U24365 (N_24365,N_20576,N_21050);
nand U24366 (N_24366,N_22041,N_21985);
and U24367 (N_24367,N_22178,N_20336);
or U24368 (N_24368,N_21850,N_20135);
or U24369 (N_24369,N_20295,N_21848);
or U24370 (N_24370,N_22199,N_21326);
nand U24371 (N_24371,N_21762,N_21446);
nor U24372 (N_24372,N_21618,N_20293);
or U24373 (N_24373,N_20932,N_21599);
nand U24374 (N_24374,N_22208,N_21214);
nand U24375 (N_24375,N_21664,N_20203);
nor U24376 (N_24376,N_22270,N_22066);
nand U24377 (N_24377,N_21096,N_20408);
xor U24378 (N_24378,N_20129,N_21229);
xnor U24379 (N_24379,N_21169,N_20011);
xnor U24380 (N_24380,N_21366,N_20872);
nand U24381 (N_24381,N_21743,N_21551);
nand U24382 (N_24382,N_20176,N_21932);
xor U24383 (N_24383,N_21066,N_21977);
xor U24384 (N_24384,N_21377,N_21882);
nand U24385 (N_24385,N_22263,N_21430);
nor U24386 (N_24386,N_22164,N_20513);
nand U24387 (N_24387,N_20616,N_21055);
and U24388 (N_24388,N_21982,N_20798);
and U24389 (N_24389,N_20930,N_21918);
nor U24390 (N_24390,N_21832,N_20984);
xor U24391 (N_24391,N_20946,N_21533);
or U24392 (N_24392,N_21086,N_21284);
nor U24393 (N_24393,N_20127,N_21531);
xor U24394 (N_24394,N_21274,N_20374);
xnor U24395 (N_24395,N_20436,N_20868);
nand U24396 (N_24396,N_20632,N_21150);
and U24397 (N_24397,N_22165,N_21140);
or U24398 (N_24398,N_21691,N_22295);
or U24399 (N_24399,N_21679,N_20451);
nand U24400 (N_24400,N_22406,N_20493);
xnor U24401 (N_24401,N_21032,N_21093);
xor U24402 (N_24402,N_20860,N_20714);
and U24403 (N_24403,N_20730,N_22385);
or U24404 (N_24404,N_21760,N_20962);
nor U24405 (N_24405,N_20822,N_20448);
and U24406 (N_24406,N_20419,N_22346);
xor U24407 (N_24407,N_21700,N_20920);
xor U24408 (N_24408,N_21678,N_21675);
or U24409 (N_24409,N_21717,N_20713);
and U24410 (N_24410,N_21593,N_21600);
nor U24411 (N_24411,N_20709,N_20393);
nor U24412 (N_24412,N_21583,N_21205);
nor U24413 (N_24413,N_20985,N_20283);
nand U24414 (N_24414,N_22288,N_20234);
xnor U24415 (N_24415,N_21650,N_20107);
nor U24416 (N_24416,N_20325,N_20572);
or U24417 (N_24417,N_20686,N_22366);
nand U24418 (N_24418,N_21660,N_20337);
or U24419 (N_24419,N_21118,N_20473);
xor U24420 (N_24420,N_21184,N_21824);
or U24421 (N_24421,N_20955,N_20960);
xnor U24422 (N_24422,N_21549,N_20452);
nor U24423 (N_24423,N_20689,N_21954);
or U24424 (N_24424,N_20152,N_20438);
nor U24425 (N_24425,N_20926,N_21424);
xor U24426 (N_24426,N_21315,N_20032);
nor U24427 (N_24427,N_22369,N_20612);
nor U24428 (N_24428,N_21930,N_21688);
nand U24429 (N_24429,N_22109,N_20043);
nor U24430 (N_24430,N_20533,N_21251);
xnor U24431 (N_24431,N_21137,N_21694);
nand U24432 (N_24432,N_22439,N_21545);
or U24433 (N_24433,N_20704,N_20390);
xnor U24434 (N_24434,N_21351,N_22136);
nor U24435 (N_24435,N_21586,N_20500);
xor U24436 (N_24436,N_21155,N_21884);
and U24437 (N_24437,N_21548,N_21779);
nand U24438 (N_24438,N_22093,N_21481);
or U24439 (N_24439,N_21292,N_22336);
or U24440 (N_24440,N_20666,N_20278);
and U24441 (N_24441,N_20574,N_20021);
xor U24442 (N_24442,N_21945,N_21208);
and U24443 (N_24443,N_20724,N_22314);
or U24444 (N_24444,N_21481,N_20150);
xnor U24445 (N_24445,N_21602,N_20151);
nand U24446 (N_24446,N_22370,N_20474);
or U24447 (N_24447,N_22091,N_21788);
nand U24448 (N_24448,N_20588,N_20617);
and U24449 (N_24449,N_22473,N_20666);
nor U24450 (N_24450,N_20787,N_21825);
or U24451 (N_24451,N_20976,N_22361);
xor U24452 (N_24452,N_20903,N_21246);
nand U24453 (N_24453,N_22288,N_21241);
nor U24454 (N_24454,N_22360,N_21398);
or U24455 (N_24455,N_21367,N_20656);
and U24456 (N_24456,N_20296,N_20442);
nand U24457 (N_24457,N_20984,N_22198);
or U24458 (N_24458,N_22117,N_22373);
and U24459 (N_24459,N_22072,N_21226);
xor U24460 (N_24460,N_21129,N_20230);
xnor U24461 (N_24461,N_22210,N_20481);
and U24462 (N_24462,N_20774,N_21225);
xor U24463 (N_24463,N_22139,N_21478);
nand U24464 (N_24464,N_21912,N_20450);
or U24465 (N_24465,N_20167,N_21624);
xor U24466 (N_24466,N_20344,N_22104);
nand U24467 (N_24467,N_21875,N_20356);
nor U24468 (N_24468,N_22366,N_22028);
xor U24469 (N_24469,N_21810,N_21852);
xor U24470 (N_24470,N_22221,N_20052);
nand U24471 (N_24471,N_21727,N_22215);
or U24472 (N_24472,N_20875,N_21919);
xor U24473 (N_24473,N_21879,N_21859);
nand U24474 (N_24474,N_22289,N_20344);
nand U24475 (N_24475,N_20315,N_21584);
or U24476 (N_24476,N_20365,N_21445);
nand U24477 (N_24477,N_21513,N_21103);
or U24478 (N_24478,N_21701,N_21198);
nor U24479 (N_24479,N_20225,N_20821);
and U24480 (N_24480,N_21030,N_20372);
and U24481 (N_24481,N_21967,N_20161);
nand U24482 (N_24482,N_21151,N_21702);
xnor U24483 (N_24483,N_21417,N_20095);
or U24484 (N_24484,N_20626,N_22308);
or U24485 (N_24485,N_20457,N_21024);
xor U24486 (N_24486,N_21808,N_21697);
nor U24487 (N_24487,N_21023,N_20443);
nor U24488 (N_24488,N_21671,N_21677);
nand U24489 (N_24489,N_21073,N_22448);
nor U24490 (N_24490,N_22383,N_20013);
and U24491 (N_24491,N_20580,N_21045);
and U24492 (N_24492,N_22179,N_20012);
nand U24493 (N_24493,N_22191,N_20185);
xnor U24494 (N_24494,N_21208,N_21415);
or U24495 (N_24495,N_20018,N_20451);
and U24496 (N_24496,N_20344,N_20415);
nand U24497 (N_24497,N_22219,N_20637);
nor U24498 (N_24498,N_21601,N_22460);
or U24499 (N_24499,N_21716,N_20007);
nor U24500 (N_24500,N_20133,N_20401);
nand U24501 (N_24501,N_22408,N_22402);
and U24502 (N_24502,N_20210,N_22331);
nand U24503 (N_24503,N_21831,N_21094);
nand U24504 (N_24504,N_21057,N_20896);
and U24505 (N_24505,N_21258,N_20683);
nor U24506 (N_24506,N_21611,N_21580);
nand U24507 (N_24507,N_21620,N_20376);
and U24508 (N_24508,N_21900,N_20403);
nand U24509 (N_24509,N_20035,N_21706);
or U24510 (N_24510,N_22410,N_20630);
nor U24511 (N_24511,N_22415,N_21443);
nor U24512 (N_24512,N_22033,N_21113);
and U24513 (N_24513,N_20468,N_21277);
nand U24514 (N_24514,N_22111,N_21045);
or U24515 (N_24515,N_22432,N_21815);
and U24516 (N_24516,N_22272,N_20494);
xnor U24517 (N_24517,N_21845,N_20514);
or U24518 (N_24518,N_22056,N_21551);
xnor U24519 (N_24519,N_20716,N_21932);
or U24520 (N_24520,N_20248,N_20273);
nor U24521 (N_24521,N_21859,N_21719);
nand U24522 (N_24522,N_21059,N_21724);
nand U24523 (N_24523,N_21790,N_20182);
nor U24524 (N_24524,N_20065,N_22122);
xnor U24525 (N_24525,N_22367,N_22478);
xor U24526 (N_24526,N_20830,N_20531);
or U24527 (N_24527,N_22182,N_20067);
xor U24528 (N_24528,N_21196,N_20821);
xor U24529 (N_24529,N_20678,N_21090);
nor U24530 (N_24530,N_21702,N_21888);
xor U24531 (N_24531,N_22346,N_21078);
and U24532 (N_24532,N_21615,N_21132);
or U24533 (N_24533,N_20714,N_20523);
or U24534 (N_24534,N_20901,N_21502);
nand U24535 (N_24535,N_22139,N_20935);
nor U24536 (N_24536,N_20042,N_21478);
and U24537 (N_24537,N_20431,N_22051);
or U24538 (N_24538,N_21925,N_20758);
nand U24539 (N_24539,N_22124,N_22312);
or U24540 (N_24540,N_21030,N_20485);
xor U24541 (N_24541,N_20100,N_21590);
or U24542 (N_24542,N_21319,N_21390);
nor U24543 (N_24543,N_20624,N_20841);
or U24544 (N_24544,N_21262,N_21819);
xor U24545 (N_24545,N_22346,N_20114);
nand U24546 (N_24546,N_20698,N_22334);
nand U24547 (N_24547,N_21698,N_21573);
and U24548 (N_24548,N_21054,N_20156);
nand U24549 (N_24549,N_21899,N_21713);
nand U24550 (N_24550,N_20506,N_21300);
nor U24551 (N_24551,N_20415,N_22132);
nand U24552 (N_24552,N_20091,N_20543);
xnor U24553 (N_24553,N_22159,N_21253);
and U24554 (N_24554,N_22161,N_21730);
nand U24555 (N_24555,N_22040,N_20193);
nand U24556 (N_24556,N_20123,N_20373);
nor U24557 (N_24557,N_20596,N_20457);
nor U24558 (N_24558,N_22313,N_22110);
and U24559 (N_24559,N_20199,N_20124);
xor U24560 (N_24560,N_21629,N_22284);
or U24561 (N_24561,N_20497,N_22469);
nor U24562 (N_24562,N_22316,N_21548);
nand U24563 (N_24563,N_21066,N_21071);
nand U24564 (N_24564,N_20028,N_21863);
xnor U24565 (N_24565,N_20984,N_21587);
or U24566 (N_24566,N_21490,N_20104);
nor U24567 (N_24567,N_21611,N_20409);
or U24568 (N_24568,N_21429,N_21575);
xor U24569 (N_24569,N_21544,N_20883);
and U24570 (N_24570,N_21676,N_20677);
and U24571 (N_24571,N_20762,N_21984);
xnor U24572 (N_24572,N_21774,N_20284);
or U24573 (N_24573,N_20770,N_21774);
nor U24574 (N_24574,N_20034,N_20623);
nor U24575 (N_24575,N_20931,N_22289);
nand U24576 (N_24576,N_22033,N_21465);
nand U24577 (N_24577,N_21478,N_21169);
or U24578 (N_24578,N_21902,N_20999);
or U24579 (N_24579,N_20957,N_21464);
and U24580 (N_24580,N_22470,N_21445);
or U24581 (N_24581,N_21420,N_22417);
nand U24582 (N_24582,N_20936,N_20500);
nand U24583 (N_24583,N_22464,N_20049);
xor U24584 (N_24584,N_21767,N_21935);
nand U24585 (N_24585,N_21673,N_21747);
xor U24586 (N_24586,N_21387,N_20339);
or U24587 (N_24587,N_21781,N_21581);
nand U24588 (N_24588,N_20613,N_21707);
nand U24589 (N_24589,N_20838,N_22270);
or U24590 (N_24590,N_21870,N_20284);
and U24591 (N_24591,N_21707,N_22313);
or U24592 (N_24592,N_20520,N_22470);
nor U24593 (N_24593,N_20870,N_20564);
nor U24594 (N_24594,N_21169,N_20823);
nand U24595 (N_24595,N_20095,N_22336);
nor U24596 (N_24596,N_20060,N_20268);
nor U24597 (N_24597,N_20278,N_20178);
nor U24598 (N_24598,N_20316,N_21502);
xnor U24599 (N_24599,N_21688,N_20393);
xor U24600 (N_24600,N_21380,N_22104);
and U24601 (N_24601,N_22275,N_21645);
xnor U24602 (N_24602,N_21051,N_20931);
nor U24603 (N_24603,N_22191,N_20510);
xor U24604 (N_24604,N_20464,N_20463);
nor U24605 (N_24605,N_21911,N_20253);
xnor U24606 (N_24606,N_22131,N_21330);
nor U24607 (N_24607,N_21085,N_21212);
nand U24608 (N_24608,N_21471,N_21487);
xor U24609 (N_24609,N_20310,N_22257);
nor U24610 (N_24610,N_21650,N_20968);
and U24611 (N_24611,N_21018,N_20862);
nand U24612 (N_24612,N_21292,N_21699);
xnor U24613 (N_24613,N_21295,N_20446);
and U24614 (N_24614,N_21669,N_21656);
and U24615 (N_24615,N_20885,N_20305);
or U24616 (N_24616,N_21385,N_21599);
xor U24617 (N_24617,N_21867,N_20994);
nand U24618 (N_24618,N_20959,N_21342);
or U24619 (N_24619,N_21270,N_20822);
nor U24620 (N_24620,N_21254,N_20828);
nor U24621 (N_24621,N_20478,N_20615);
nand U24622 (N_24622,N_21305,N_20561);
nor U24623 (N_24623,N_22422,N_21385);
or U24624 (N_24624,N_21090,N_22416);
xor U24625 (N_24625,N_21642,N_21306);
nor U24626 (N_24626,N_22251,N_20632);
xor U24627 (N_24627,N_22106,N_21745);
xnor U24628 (N_24628,N_21825,N_20740);
nand U24629 (N_24629,N_20655,N_20915);
or U24630 (N_24630,N_21783,N_20440);
xnor U24631 (N_24631,N_22454,N_20188);
nand U24632 (N_24632,N_20578,N_20105);
or U24633 (N_24633,N_21632,N_22449);
or U24634 (N_24634,N_20949,N_20580);
nand U24635 (N_24635,N_20429,N_21674);
xnor U24636 (N_24636,N_20997,N_21771);
xnor U24637 (N_24637,N_21432,N_21352);
or U24638 (N_24638,N_22162,N_22136);
or U24639 (N_24639,N_22105,N_20122);
nor U24640 (N_24640,N_21913,N_20590);
and U24641 (N_24641,N_21751,N_20690);
xor U24642 (N_24642,N_21489,N_21279);
nor U24643 (N_24643,N_21778,N_21161);
or U24644 (N_24644,N_20904,N_21990);
xor U24645 (N_24645,N_20898,N_21559);
or U24646 (N_24646,N_21139,N_20495);
and U24647 (N_24647,N_21015,N_20560);
xor U24648 (N_24648,N_20075,N_21223);
and U24649 (N_24649,N_20215,N_20005);
or U24650 (N_24650,N_21242,N_20989);
nor U24651 (N_24651,N_21130,N_21151);
nor U24652 (N_24652,N_22408,N_20033);
nand U24653 (N_24653,N_21964,N_22254);
nor U24654 (N_24654,N_22141,N_20609);
and U24655 (N_24655,N_20542,N_20166);
nor U24656 (N_24656,N_20415,N_20855);
xnor U24657 (N_24657,N_20091,N_22068);
nand U24658 (N_24658,N_20618,N_20507);
nor U24659 (N_24659,N_20679,N_20090);
or U24660 (N_24660,N_20014,N_20488);
and U24661 (N_24661,N_20448,N_20329);
or U24662 (N_24662,N_21911,N_21445);
or U24663 (N_24663,N_21110,N_21316);
nand U24664 (N_24664,N_21409,N_20518);
and U24665 (N_24665,N_21949,N_21952);
xnor U24666 (N_24666,N_21880,N_21665);
nand U24667 (N_24667,N_21648,N_21827);
nand U24668 (N_24668,N_20963,N_22130);
nand U24669 (N_24669,N_21649,N_21750);
nand U24670 (N_24670,N_22472,N_21276);
and U24671 (N_24671,N_21586,N_22451);
xnor U24672 (N_24672,N_20226,N_20892);
nor U24673 (N_24673,N_22179,N_20377);
xor U24674 (N_24674,N_22135,N_20366);
or U24675 (N_24675,N_21039,N_20188);
xnor U24676 (N_24676,N_21027,N_21038);
xor U24677 (N_24677,N_21804,N_20381);
and U24678 (N_24678,N_21856,N_21618);
xnor U24679 (N_24679,N_21369,N_22373);
or U24680 (N_24680,N_21708,N_21804);
nand U24681 (N_24681,N_20140,N_21358);
nand U24682 (N_24682,N_22092,N_21640);
or U24683 (N_24683,N_21757,N_20693);
xnor U24684 (N_24684,N_21270,N_21247);
or U24685 (N_24685,N_20384,N_20194);
nand U24686 (N_24686,N_21510,N_22406);
or U24687 (N_24687,N_22235,N_21170);
nor U24688 (N_24688,N_21530,N_20456);
or U24689 (N_24689,N_22171,N_20298);
or U24690 (N_24690,N_20340,N_20075);
nand U24691 (N_24691,N_21286,N_20137);
nand U24692 (N_24692,N_21694,N_20848);
or U24693 (N_24693,N_21978,N_21166);
and U24694 (N_24694,N_20146,N_20386);
xnor U24695 (N_24695,N_20547,N_22268);
xnor U24696 (N_24696,N_21040,N_21814);
nor U24697 (N_24697,N_22471,N_21087);
xnor U24698 (N_24698,N_22385,N_20299);
or U24699 (N_24699,N_21774,N_20041);
nand U24700 (N_24700,N_20252,N_20456);
and U24701 (N_24701,N_20651,N_22319);
nor U24702 (N_24702,N_21577,N_20355);
nand U24703 (N_24703,N_20333,N_20008);
nand U24704 (N_24704,N_21341,N_20222);
nand U24705 (N_24705,N_22319,N_20051);
or U24706 (N_24706,N_20399,N_21085);
xor U24707 (N_24707,N_20380,N_20676);
nor U24708 (N_24708,N_21381,N_21889);
and U24709 (N_24709,N_22283,N_20211);
or U24710 (N_24710,N_21074,N_21156);
or U24711 (N_24711,N_20273,N_22492);
xnor U24712 (N_24712,N_20878,N_21818);
and U24713 (N_24713,N_20790,N_22464);
nor U24714 (N_24714,N_21474,N_20186);
nand U24715 (N_24715,N_21824,N_20989);
xnor U24716 (N_24716,N_22386,N_20090);
or U24717 (N_24717,N_21188,N_21505);
and U24718 (N_24718,N_22350,N_20417);
nor U24719 (N_24719,N_20091,N_22039);
and U24720 (N_24720,N_20144,N_21175);
nor U24721 (N_24721,N_21869,N_22394);
nor U24722 (N_24722,N_22247,N_20118);
nor U24723 (N_24723,N_21326,N_22401);
and U24724 (N_24724,N_20467,N_21430);
and U24725 (N_24725,N_21385,N_21655);
nor U24726 (N_24726,N_22313,N_20282);
nor U24727 (N_24727,N_21968,N_20649);
and U24728 (N_24728,N_21087,N_21193);
or U24729 (N_24729,N_21847,N_20391);
xor U24730 (N_24730,N_22426,N_20149);
xor U24731 (N_24731,N_20171,N_20624);
and U24732 (N_24732,N_22287,N_20220);
xnor U24733 (N_24733,N_21252,N_21553);
nand U24734 (N_24734,N_21294,N_22224);
nor U24735 (N_24735,N_21439,N_21172);
nor U24736 (N_24736,N_20030,N_20047);
xor U24737 (N_24737,N_21547,N_21640);
and U24738 (N_24738,N_21124,N_20934);
nand U24739 (N_24739,N_21627,N_20192);
and U24740 (N_24740,N_20048,N_22241);
or U24741 (N_24741,N_21999,N_20629);
xor U24742 (N_24742,N_21005,N_22311);
and U24743 (N_24743,N_22476,N_20199);
nand U24744 (N_24744,N_21342,N_20134);
or U24745 (N_24745,N_21809,N_22471);
nand U24746 (N_24746,N_21394,N_20609);
xor U24747 (N_24747,N_21868,N_21615);
and U24748 (N_24748,N_20980,N_22329);
nand U24749 (N_24749,N_20492,N_20761);
and U24750 (N_24750,N_20866,N_21005);
and U24751 (N_24751,N_20395,N_21619);
xnor U24752 (N_24752,N_21243,N_21259);
xnor U24753 (N_24753,N_20745,N_20589);
or U24754 (N_24754,N_20622,N_20350);
nand U24755 (N_24755,N_21176,N_20489);
and U24756 (N_24756,N_21219,N_21202);
nor U24757 (N_24757,N_21790,N_20193);
nor U24758 (N_24758,N_21316,N_21207);
nor U24759 (N_24759,N_20506,N_20871);
or U24760 (N_24760,N_21373,N_22097);
nand U24761 (N_24761,N_22131,N_20481);
nand U24762 (N_24762,N_20092,N_20678);
nor U24763 (N_24763,N_22191,N_22425);
and U24764 (N_24764,N_21406,N_20366);
xor U24765 (N_24765,N_20272,N_21915);
nand U24766 (N_24766,N_20236,N_21239);
and U24767 (N_24767,N_21549,N_21485);
nor U24768 (N_24768,N_21915,N_21109);
and U24769 (N_24769,N_20514,N_21959);
nand U24770 (N_24770,N_21093,N_21686);
or U24771 (N_24771,N_20778,N_21167);
and U24772 (N_24772,N_21965,N_20840);
or U24773 (N_24773,N_20471,N_21685);
nor U24774 (N_24774,N_22126,N_20484);
nor U24775 (N_24775,N_21914,N_22284);
and U24776 (N_24776,N_20905,N_21477);
and U24777 (N_24777,N_21141,N_22304);
nor U24778 (N_24778,N_20648,N_20295);
or U24779 (N_24779,N_20779,N_20310);
nor U24780 (N_24780,N_22344,N_20733);
xor U24781 (N_24781,N_20319,N_22415);
and U24782 (N_24782,N_22394,N_22448);
nand U24783 (N_24783,N_21485,N_22124);
and U24784 (N_24784,N_21334,N_20375);
nor U24785 (N_24785,N_20723,N_21898);
nor U24786 (N_24786,N_20647,N_22201);
or U24787 (N_24787,N_21096,N_22003);
nor U24788 (N_24788,N_20568,N_21035);
nor U24789 (N_24789,N_21409,N_20011);
xnor U24790 (N_24790,N_20045,N_20040);
xor U24791 (N_24791,N_20804,N_22049);
and U24792 (N_24792,N_21656,N_22244);
or U24793 (N_24793,N_22397,N_20922);
nor U24794 (N_24794,N_20892,N_22427);
xor U24795 (N_24795,N_20181,N_22223);
or U24796 (N_24796,N_20515,N_20650);
and U24797 (N_24797,N_21721,N_22284);
and U24798 (N_24798,N_22057,N_20688);
nor U24799 (N_24799,N_20452,N_21075);
and U24800 (N_24800,N_21328,N_20365);
nor U24801 (N_24801,N_22498,N_20417);
xnor U24802 (N_24802,N_21455,N_20538);
nand U24803 (N_24803,N_21761,N_21360);
nand U24804 (N_24804,N_20667,N_20792);
and U24805 (N_24805,N_20982,N_21357);
or U24806 (N_24806,N_21883,N_21816);
nor U24807 (N_24807,N_21641,N_21706);
and U24808 (N_24808,N_21588,N_21030);
or U24809 (N_24809,N_22042,N_21952);
xnor U24810 (N_24810,N_20939,N_21952);
and U24811 (N_24811,N_22381,N_20861);
nor U24812 (N_24812,N_21322,N_21479);
and U24813 (N_24813,N_21841,N_22198);
or U24814 (N_24814,N_22399,N_21746);
and U24815 (N_24815,N_20520,N_20974);
nand U24816 (N_24816,N_21559,N_21314);
and U24817 (N_24817,N_20544,N_22191);
and U24818 (N_24818,N_21870,N_21906);
nor U24819 (N_24819,N_21321,N_22316);
xor U24820 (N_24820,N_20738,N_20145);
xnor U24821 (N_24821,N_21669,N_21954);
nand U24822 (N_24822,N_21594,N_21998);
or U24823 (N_24823,N_21279,N_20597);
nor U24824 (N_24824,N_21554,N_21847);
xnor U24825 (N_24825,N_22406,N_21236);
nand U24826 (N_24826,N_21295,N_20508);
nor U24827 (N_24827,N_21394,N_21463);
or U24828 (N_24828,N_20295,N_20349);
and U24829 (N_24829,N_22208,N_21670);
nand U24830 (N_24830,N_20791,N_21542);
xnor U24831 (N_24831,N_21316,N_21563);
nand U24832 (N_24832,N_21957,N_21921);
or U24833 (N_24833,N_22370,N_22043);
nand U24834 (N_24834,N_20797,N_22149);
nor U24835 (N_24835,N_20166,N_22482);
and U24836 (N_24836,N_20450,N_22389);
nor U24837 (N_24837,N_21246,N_21274);
nand U24838 (N_24838,N_22159,N_21797);
nand U24839 (N_24839,N_20274,N_22335);
nor U24840 (N_24840,N_22065,N_21548);
or U24841 (N_24841,N_22397,N_20691);
xor U24842 (N_24842,N_20414,N_21046);
and U24843 (N_24843,N_22303,N_20631);
xnor U24844 (N_24844,N_20545,N_21598);
xor U24845 (N_24845,N_21729,N_20481);
and U24846 (N_24846,N_20645,N_20494);
and U24847 (N_24847,N_20352,N_21606);
or U24848 (N_24848,N_20597,N_21612);
and U24849 (N_24849,N_20254,N_20178);
or U24850 (N_24850,N_21748,N_21051);
or U24851 (N_24851,N_21908,N_20063);
nand U24852 (N_24852,N_20192,N_21023);
and U24853 (N_24853,N_22039,N_20107);
nand U24854 (N_24854,N_21827,N_21928);
xnor U24855 (N_24855,N_21592,N_21878);
nor U24856 (N_24856,N_21921,N_21131);
or U24857 (N_24857,N_21980,N_21721);
xnor U24858 (N_24858,N_20369,N_22210);
nand U24859 (N_24859,N_20317,N_21974);
nand U24860 (N_24860,N_21340,N_21027);
nor U24861 (N_24861,N_21998,N_20131);
xor U24862 (N_24862,N_20813,N_21131);
nand U24863 (N_24863,N_22008,N_20690);
nand U24864 (N_24864,N_21157,N_22103);
nor U24865 (N_24865,N_22137,N_20815);
or U24866 (N_24866,N_20226,N_21480);
nand U24867 (N_24867,N_21157,N_21175);
or U24868 (N_24868,N_20074,N_20244);
xor U24869 (N_24869,N_20748,N_20504);
nand U24870 (N_24870,N_22014,N_21399);
or U24871 (N_24871,N_21465,N_21344);
and U24872 (N_24872,N_22037,N_21950);
or U24873 (N_24873,N_22115,N_20396);
and U24874 (N_24874,N_20102,N_21737);
nand U24875 (N_24875,N_20796,N_20056);
or U24876 (N_24876,N_20578,N_22330);
nand U24877 (N_24877,N_20008,N_22016);
xor U24878 (N_24878,N_21683,N_21449);
nand U24879 (N_24879,N_22274,N_20262);
and U24880 (N_24880,N_21184,N_20863);
nand U24881 (N_24881,N_20893,N_21420);
nand U24882 (N_24882,N_22249,N_20914);
nand U24883 (N_24883,N_22471,N_22079);
xor U24884 (N_24884,N_21178,N_21946);
and U24885 (N_24885,N_20252,N_20636);
xor U24886 (N_24886,N_20802,N_20463);
nand U24887 (N_24887,N_20583,N_20710);
nand U24888 (N_24888,N_20958,N_21071);
and U24889 (N_24889,N_20937,N_21441);
nand U24890 (N_24890,N_21764,N_22451);
or U24891 (N_24891,N_22486,N_20793);
xnor U24892 (N_24892,N_21240,N_21024);
xor U24893 (N_24893,N_20824,N_21385);
nand U24894 (N_24894,N_20326,N_20835);
and U24895 (N_24895,N_21127,N_20561);
nand U24896 (N_24896,N_22203,N_22389);
nand U24897 (N_24897,N_21727,N_20537);
nand U24898 (N_24898,N_20988,N_20880);
and U24899 (N_24899,N_20169,N_21604);
or U24900 (N_24900,N_21720,N_22141);
nand U24901 (N_24901,N_20826,N_21138);
nand U24902 (N_24902,N_20353,N_21347);
nor U24903 (N_24903,N_20066,N_21626);
nand U24904 (N_24904,N_20288,N_20603);
nand U24905 (N_24905,N_20420,N_20103);
or U24906 (N_24906,N_20882,N_20126);
nor U24907 (N_24907,N_21623,N_21184);
or U24908 (N_24908,N_22489,N_21757);
and U24909 (N_24909,N_21449,N_22488);
and U24910 (N_24910,N_21160,N_21083);
nand U24911 (N_24911,N_22072,N_22029);
nand U24912 (N_24912,N_21165,N_20894);
nor U24913 (N_24913,N_22348,N_21055);
and U24914 (N_24914,N_21219,N_20514);
nand U24915 (N_24915,N_21961,N_21839);
and U24916 (N_24916,N_21666,N_20342);
xor U24917 (N_24917,N_22373,N_21110);
nor U24918 (N_24918,N_21724,N_20755);
nor U24919 (N_24919,N_20878,N_21031);
or U24920 (N_24920,N_22156,N_20992);
or U24921 (N_24921,N_21189,N_20351);
or U24922 (N_24922,N_20618,N_21563);
nor U24923 (N_24923,N_20221,N_22028);
and U24924 (N_24924,N_20178,N_21583);
xor U24925 (N_24925,N_22020,N_21868);
or U24926 (N_24926,N_21357,N_21049);
and U24927 (N_24927,N_21172,N_20734);
nor U24928 (N_24928,N_20076,N_22434);
nor U24929 (N_24929,N_21646,N_22494);
or U24930 (N_24930,N_20172,N_21185);
xnor U24931 (N_24931,N_22429,N_20545);
nand U24932 (N_24932,N_20777,N_22310);
or U24933 (N_24933,N_20267,N_21564);
xnor U24934 (N_24934,N_21887,N_21864);
nand U24935 (N_24935,N_20822,N_20090);
nor U24936 (N_24936,N_21337,N_21075);
xnor U24937 (N_24937,N_21465,N_22424);
nor U24938 (N_24938,N_21658,N_20504);
nand U24939 (N_24939,N_22446,N_22258);
nor U24940 (N_24940,N_20319,N_21935);
and U24941 (N_24941,N_20103,N_20483);
nor U24942 (N_24942,N_21143,N_20377);
nand U24943 (N_24943,N_21983,N_20822);
nor U24944 (N_24944,N_20942,N_20134);
or U24945 (N_24945,N_22306,N_22242);
nand U24946 (N_24946,N_20747,N_20828);
and U24947 (N_24947,N_21257,N_21249);
nor U24948 (N_24948,N_20444,N_20800);
nand U24949 (N_24949,N_21120,N_22384);
and U24950 (N_24950,N_20236,N_20069);
nor U24951 (N_24951,N_21966,N_21715);
nor U24952 (N_24952,N_20103,N_20764);
or U24953 (N_24953,N_22047,N_22218);
nand U24954 (N_24954,N_20575,N_21127);
xor U24955 (N_24955,N_22398,N_21551);
xor U24956 (N_24956,N_22407,N_20199);
nand U24957 (N_24957,N_20873,N_22181);
xor U24958 (N_24958,N_20710,N_22352);
xnor U24959 (N_24959,N_20249,N_22188);
xor U24960 (N_24960,N_21812,N_20198);
nand U24961 (N_24961,N_20589,N_21977);
nor U24962 (N_24962,N_20689,N_21864);
or U24963 (N_24963,N_21973,N_20962);
nor U24964 (N_24964,N_20167,N_22007);
nor U24965 (N_24965,N_21294,N_20258);
or U24966 (N_24966,N_20196,N_21237);
or U24967 (N_24967,N_20533,N_20187);
or U24968 (N_24968,N_21848,N_20570);
xnor U24969 (N_24969,N_20962,N_20292);
xor U24970 (N_24970,N_22185,N_22291);
nor U24971 (N_24971,N_20413,N_20746);
nor U24972 (N_24972,N_20645,N_21743);
and U24973 (N_24973,N_20020,N_20053);
xor U24974 (N_24974,N_21140,N_20199);
or U24975 (N_24975,N_21106,N_22452);
or U24976 (N_24976,N_22143,N_20189);
and U24977 (N_24977,N_21061,N_22312);
or U24978 (N_24978,N_20597,N_21075);
nand U24979 (N_24979,N_21918,N_21196);
nor U24980 (N_24980,N_22369,N_20255);
nor U24981 (N_24981,N_20140,N_21134);
or U24982 (N_24982,N_20024,N_21584);
xnor U24983 (N_24983,N_21823,N_21012);
xor U24984 (N_24984,N_21450,N_20002);
or U24985 (N_24985,N_20026,N_22356);
nor U24986 (N_24986,N_21562,N_22263);
and U24987 (N_24987,N_21308,N_22306);
nor U24988 (N_24988,N_22400,N_22071);
and U24989 (N_24989,N_21772,N_21744);
or U24990 (N_24990,N_21291,N_20044);
or U24991 (N_24991,N_22063,N_22470);
and U24992 (N_24992,N_21125,N_20083);
nor U24993 (N_24993,N_20208,N_20928);
xor U24994 (N_24994,N_20776,N_22296);
or U24995 (N_24995,N_20015,N_21002);
or U24996 (N_24996,N_20169,N_22276);
nand U24997 (N_24997,N_21341,N_20654);
nand U24998 (N_24998,N_21501,N_21434);
nand U24999 (N_24999,N_21591,N_22272);
or UO_0 (O_0,N_23551,N_23089);
xor UO_1 (O_1,N_23149,N_22758);
and UO_2 (O_2,N_23530,N_23348);
xnor UO_3 (O_3,N_24279,N_24282);
and UO_4 (O_4,N_22879,N_23343);
nand UO_5 (O_5,N_23346,N_23376);
nand UO_6 (O_6,N_23693,N_24806);
or UO_7 (O_7,N_23688,N_24639);
xor UO_8 (O_8,N_23023,N_23528);
nand UO_9 (O_9,N_22885,N_24109);
xnor UO_10 (O_10,N_24140,N_24718);
nand UO_11 (O_11,N_22853,N_23807);
nand UO_12 (O_12,N_23709,N_22617);
nor UO_13 (O_13,N_23483,N_23587);
nand UO_14 (O_14,N_23972,N_24356);
xor UO_15 (O_15,N_23162,N_24375);
nor UO_16 (O_16,N_24829,N_23355);
and UO_17 (O_17,N_24599,N_23990);
or UO_18 (O_18,N_22654,N_22888);
nor UO_19 (O_19,N_24251,N_22965);
nor UO_20 (O_20,N_22823,N_24208);
xnor UO_21 (O_21,N_22928,N_24107);
nand UO_22 (O_22,N_23529,N_23466);
xor UO_23 (O_23,N_24555,N_23536);
xor UO_24 (O_24,N_22726,N_24573);
or UO_25 (O_25,N_24200,N_22933);
or UO_26 (O_26,N_23007,N_23690);
and UO_27 (O_27,N_23632,N_24483);
nor UO_28 (O_28,N_24582,N_24930);
and UO_29 (O_29,N_24754,N_22652);
nor UO_30 (O_30,N_23431,N_23758);
xnor UO_31 (O_31,N_24874,N_23264);
and UO_32 (O_32,N_23054,N_24393);
nand UO_33 (O_33,N_22880,N_24996);
and UO_34 (O_34,N_22956,N_22760);
nand UO_35 (O_35,N_24454,N_23438);
and UO_36 (O_36,N_22532,N_24605);
xor UO_37 (O_37,N_22741,N_24537);
xnor UO_38 (O_38,N_23887,N_24481);
nand UO_39 (O_39,N_23952,N_23523);
and UO_40 (O_40,N_23961,N_23595);
and UO_41 (O_41,N_23907,N_24931);
nand UO_42 (O_42,N_23527,N_24296);
nor UO_43 (O_43,N_24530,N_23055);
nor UO_44 (O_44,N_24390,N_24765);
nor UO_45 (O_45,N_24065,N_22775);
and UO_46 (O_46,N_22680,N_23967);
xor UO_47 (O_47,N_24699,N_23652);
xnor UO_48 (O_48,N_24774,N_22649);
xnor UO_49 (O_49,N_24170,N_23039);
nor UO_50 (O_50,N_22552,N_23666);
nand UO_51 (O_51,N_23925,N_24244);
or UO_52 (O_52,N_23391,N_24805);
and UO_53 (O_53,N_22924,N_24321);
nor UO_54 (O_54,N_22980,N_24852);
and UO_55 (O_55,N_23881,N_24482);
and UO_56 (O_56,N_23778,N_22650);
xnor UO_57 (O_57,N_24882,N_24717);
nor UO_58 (O_58,N_23463,N_24928);
nor UO_59 (O_59,N_23368,N_23286);
nor UO_60 (O_60,N_23626,N_22867);
nor UO_61 (O_61,N_24948,N_24617);
or UO_62 (O_62,N_22651,N_23775);
and UO_63 (O_63,N_22539,N_23507);
nor UO_64 (O_64,N_24411,N_22819);
nor UO_65 (O_65,N_23899,N_24712);
nor UO_66 (O_66,N_24516,N_22629);
nand UO_67 (O_67,N_23697,N_24383);
and UO_68 (O_68,N_23012,N_23442);
nor UO_69 (O_69,N_24893,N_23160);
or UO_70 (O_70,N_24377,N_23405);
nand UO_71 (O_71,N_23969,N_24804);
nand UO_72 (O_72,N_24091,N_23737);
xor UO_73 (O_73,N_22546,N_23426);
and UO_74 (O_74,N_23201,N_23640);
xnor UO_75 (O_75,N_24263,N_23742);
or UO_76 (O_76,N_23924,N_22585);
and UO_77 (O_77,N_24402,N_23494);
nor UO_78 (O_78,N_24694,N_23156);
and UO_79 (O_79,N_22923,N_23784);
and UO_80 (O_80,N_22902,N_22643);
and UO_81 (O_81,N_23402,N_23103);
xor UO_82 (O_82,N_23075,N_24194);
and UO_83 (O_83,N_23322,N_22661);
and UO_84 (O_84,N_24843,N_24205);
nand UO_85 (O_85,N_23733,N_22663);
or UO_86 (O_86,N_24775,N_23830);
or UO_87 (O_87,N_22524,N_22542);
xor UO_88 (O_88,N_24461,N_23216);
or UO_89 (O_89,N_24380,N_23128);
or UO_90 (O_90,N_23844,N_24837);
xor UO_91 (O_91,N_23304,N_23735);
nor UO_92 (O_92,N_22863,N_22891);
or UO_93 (O_93,N_24048,N_23866);
nor UO_94 (O_94,N_24836,N_22547);
or UO_95 (O_95,N_22765,N_22844);
or UO_96 (O_96,N_23829,N_24651);
xor UO_97 (O_97,N_24723,N_24795);
and UO_98 (O_98,N_24011,N_24325);
xor UO_99 (O_99,N_22779,N_23325);
or UO_100 (O_100,N_23892,N_23454);
and UO_101 (O_101,N_22845,N_23239);
nand UO_102 (O_102,N_24565,N_23479);
or UO_103 (O_103,N_23612,N_22852);
or UO_104 (O_104,N_24221,N_23058);
xor UO_105 (O_105,N_23817,N_23085);
xnor UO_106 (O_106,N_24185,N_22857);
xnor UO_107 (O_107,N_22747,N_22721);
xor UO_108 (O_108,N_24871,N_22623);
and UO_109 (O_109,N_23407,N_23918);
or UO_110 (O_110,N_22789,N_24070);
and UO_111 (O_111,N_22517,N_23281);
nand UO_112 (O_112,N_23123,N_24112);
xnor UO_113 (O_113,N_23379,N_24297);
nor UO_114 (O_114,N_23436,N_24157);
and UO_115 (O_115,N_23364,N_24105);
and UO_116 (O_116,N_23300,N_23041);
nor UO_117 (O_117,N_24577,N_24252);
or UO_118 (O_118,N_24755,N_22785);
nand UO_119 (O_119,N_24389,N_22575);
nand UO_120 (O_120,N_24035,N_22809);
nand UO_121 (O_121,N_24624,N_24067);
nor UO_122 (O_122,N_22782,N_23589);
or UO_123 (O_123,N_24448,N_23982);
xor UO_124 (O_124,N_23674,N_23511);
nor UO_125 (O_125,N_23766,N_23414);
and UO_126 (O_126,N_24036,N_22755);
xnor UO_127 (O_127,N_22712,N_24691);
nor UO_128 (O_128,N_24658,N_24143);
xor UO_129 (O_129,N_24751,N_23113);
and UO_130 (O_130,N_23077,N_23739);
or UO_131 (O_131,N_22770,N_24972);
nand UO_132 (O_132,N_23799,N_22806);
and UO_133 (O_133,N_23771,N_24769);
nand UO_134 (O_134,N_24058,N_22574);
and UO_135 (O_135,N_24258,N_22884);
nor UO_136 (O_136,N_24367,N_24951);
and UO_137 (O_137,N_23657,N_24172);
nand UO_138 (O_138,N_23471,N_24523);
nand UO_139 (O_139,N_22903,N_23986);
nor UO_140 (O_140,N_24696,N_23221);
nor UO_141 (O_141,N_22694,N_24436);
and UO_142 (O_142,N_22508,N_24929);
and UO_143 (O_143,N_22949,N_24584);
xnor UO_144 (O_144,N_22757,N_22679);
nand UO_145 (O_145,N_24120,N_23649);
and UO_146 (O_146,N_23100,N_24669);
and UO_147 (O_147,N_22826,N_23382);
nor UO_148 (O_148,N_22696,N_24895);
xnor UO_149 (O_149,N_22776,N_23352);
xnor UO_150 (O_150,N_24273,N_22930);
or UO_151 (O_151,N_23010,N_24098);
and UO_152 (O_152,N_22750,N_24809);
or UO_153 (O_153,N_24322,N_22571);
or UO_154 (O_154,N_23171,N_22876);
or UO_155 (O_155,N_24462,N_23219);
or UO_156 (O_156,N_23013,N_23552);
xor UO_157 (O_157,N_23340,N_22787);
xnor UO_158 (O_158,N_23137,N_23499);
or UO_159 (O_159,N_24469,N_24018);
xnor UO_160 (O_160,N_24864,N_22892);
nor UO_161 (O_161,N_23412,N_24417);
or UO_162 (O_162,N_24731,N_22934);
nand UO_163 (O_163,N_23531,N_23490);
or UO_164 (O_164,N_24222,N_23234);
and UO_165 (O_165,N_22786,N_23290);
and UO_166 (O_166,N_22973,N_22536);
xnor UO_167 (O_167,N_24434,N_24333);
and UO_168 (O_168,N_22725,N_24927);
and UO_169 (O_169,N_23107,N_23823);
and UO_170 (O_170,N_22894,N_23026);
xnor UO_171 (O_171,N_22794,N_24026);
and UO_172 (O_172,N_23440,N_24772);
or UO_173 (O_173,N_24733,N_24368);
nand UO_174 (O_174,N_23195,N_24202);
or UO_175 (O_175,N_24568,N_23413);
xor UO_176 (O_176,N_23548,N_22904);
nor UO_177 (O_177,N_24032,N_22506);
xnor UO_178 (O_178,N_23298,N_24165);
or UO_179 (O_179,N_23549,N_23331);
and UO_180 (O_180,N_23679,N_23940);
nor UO_181 (O_181,N_23247,N_24014);
nand UO_182 (O_182,N_24196,N_23152);
and UO_183 (O_183,N_23028,N_22516);
or UO_184 (O_184,N_23522,N_23524);
xor UO_185 (O_185,N_24862,N_23995);
or UO_186 (O_186,N_23683,N_24618);
nand UO_187 (O_187,N_23453,N_24101);
xnor UO_188 (O_188,N_23890,N_23339);
nand UO_189 (O_189,N_23064,N_24231);
nand UO_190 (O_190,N_24062,N_23947);
nand UO_191 (O_191,N_24802,N_24596);
nand UO_192 (O_192,N_23199,N_23804);
nand UO_193 (O_193,N_23916,N_24726);
or UO_194 (O_194,N_24515,N_22865);
nand UO_195 (O_195,N_23648,N_22735);
nand UO_196 (O_196,N_23689,N_23896);
nand UO_197 (O_197,N_24697,N_22579);
nand UO_198 (O_198,N_24089,N_24053);
or UO_199 (O_199,N_24442,N_23747);
nor UO_200 (O_200,N_24281,N_23257);
and UO_201 (O_201,N_23808,N_22607);
xor UO_202 (O_202,N_24647,N_24936);
nand UO_203 (O_203,N_23143,N_24817);
and UO_204 (O_204,N_23083,N_22983);
xnor UO_205 (O_205,N_22957,N_23744);
xnor UO_206 (O_206,N_22591,N_24486);
or UO_207 (O_207,N_24267,N_24746);
or UO_208 (O_208,N_23224,N_24496);
nor UO_209 (O_209,N_24005,N_23682);
and UO_210 (O_210,N_23606,N_23713);
nor UO_211 (O_211,N_23717,N_24665);
nor UO_212 (O_212,N_23686,N_24635);
nor UO_213 (O_213,N_22642,N_23711);
nor UO_214 (O_214,N_24518,N_24360);
nand UO_215 (O_215,N_24791,N_24787);
and UO_216 (O_216,N_22702,N_23313);
or UO_217 (O_217,N_23932,N_22893);
or UO_218 (O_218,N_24077,N_23669);
nor UO_219 (O_219,N_23585,N_23870);
xnor UO_220 (O_220,N_22715,N_23335);
xor UO_221 (O_221,N_23024,N_24752);
and UO_222 (O_222,N_24569,N_23545);
or UO_223 (O_223,N_23477,N_22946);
and UO_224 (O_224,N_22985,N_24145);
nand UO_225 (O_225,N_24685,N_22821);
and UO_226 (O_226,N_23147,N_24234);
xor UO_227 (O_227,N_23299,N_24578);
xnor UO_228 (O_228,N_23349,N_22703);
or UO_229 (O_229,N_24447,N_24896);
nor UO_230 (O_230,N_23242,N_24198);
nand UO_231 (O_231,N_24302,N_23462);
nor UO_232 (O_232,N_24766,N_23588);
xnor UO_233 (O_233,N_24920,N_24855);
and UO_234 (O_234,N_22850,N_24484);
nand UO_235 (O_235,N_22995,N_24060);
nor UO_236 (O_236,N_24338,N_23743);
nor UO_237 (O_237,N_24400,N_22534);
nor UO_238 (O_238,N_23213,N_22831);
nor UO_239 (O_239,N_23333,N_24501);
nand UO_240 (O_240,N_24277,N_24293);
xor UO_241 (O_241,N_23228,N_22753);
or UO_242 (O_242,N_23929,N_22667);
xor UO_243 (O_243,N_23037,N_24667);
or UO_244 (O_244,N_24676,N_24668);
nand UO_245 (O_245,N_23303,N_24068);
nand UO_246 (O_246,N_24937,N_23989);
and UO_247 (O_247,N_24092,N_23190);
nand UO_248 (O_248,N_24689,N_22635);
and UO_249 (O_249,N_23501,N_24917);
nand UO_250 (O_250,N_23517,N_24227);
or UO_251 (O_251,N_24275,N_23678);
and UO_252 (O_252,N_23187,N_23610);
nor UO_253 (O_253,N_22645,N_23819);
nor UO_254 (O_254,N_24419,N_23814);
nor UO_255 (O_255,N_22996,N_23192);
and UO_256 (O_256,N_24315,N_23293);
nor UO_257 (O_257,N_22837,N_22616);
xor UO_258 (O_258,N_23035,N_24261);
nor UO_259 (O_259,N_22628,N_24406);
nor UO_260 (O_260,N_24810,N_23279);
and UO_261 (O_261,N_22916,N_24283);
xor UO_262 (O_262,N_24660,N_22793);
nand UO_263 (O_263,N_23473,N_24716);
and UO_264 (O_264,N_23435,N_23197);
nand UO_265 (O_265,N_24040,N_24362);
xor UO_266 (O_266,N_22962,N_24246);
and UO_267 (O_267,N_24798,N_24575);
nand UO_268 (O_268,N_24099,N_24865);
nor UO_269 (O_269,N_22736,N_23305);
or UO_270 (O_270,N_23820,N_23757);
nand UO_271 (O_271,N_23812,N_24888);
nand UO_272 (O_272,N_23984,N_23145);
and UO_273 (O_273,N_23205,N_23810);
nor UO_274 (O_274,N_24834,N_23960);
and UO_275 (O_275,N_24151,N_23425);
and UO_276 (O_276,N_24816,N_23267);
nand UO_277 (O_277,N_23939,N_24870);
nand UO_278 (O_278,N_23127,N_24211);
nor UO_279 (O_279,N_22593,N_23136);
and UO_280 (O_280,N_24385,N_23353);
nor UO_281 (O_281,N_23115,N_23895);
xnor UO_282 (O_282,N_23868,N_23575);
nor UO_283 (O_283,N_22769,N_23356);
and UO_284 (O_284,N_22937,N_23445);
nand UO_285 (O_285,N_23594,N_24264);
nand UO_286 (O_286,N_22711,N_23596);
or UO_287 (O_287,N_23667,N_23066);
and UO_288 (O_288,N_22739,N_23470);
or UO_289 (O_289,N_23122,N_24045);
xor UO_290 (O_290,N_24813,N_24858);
and UO_291 (O_291,N_23794,N_23558);
and UO_292 (O_292,N_23577,N_22588);
or UO_293 (O_293,N_23306,N_24922);
or UO_294 (O_294,N_24800,N_24104);
or UO_295 (O_295,N_23334,N_24916);
nand UO_296 (O_296,N_23297,N_24294);
xnor UO_297 (O_297,N_22917,N_23973);
and UO_298 (O_298,N_24373,N_24585);
xnor UO_299 (O_299,N_24973,N_22706);
nor UO_300 (O_300,N_23447,N_24298);
and UO_301 (O_301,N_23618,N_24978);
and UO_302 (O_302,N_23276,N_23371);
nand UO_303 (O_303,N_24892,N_23319);
xor UO_304 (O_304,N_23120,N_23639);
or UO_305 (O_305,N_23601,N_23991);
or UO_306 (O_306,N_23110,N_24576);
or UO_307 (O_307,N_22567,N_23033);
and UO_308 (O_308,N_23394,N_24452);
nor UO_309 (O_309,N_24108,N_23354);
or UO_310 (O_310,N_22801,N_24729);
nor UO_311 (O_311,N_24184,N_24342);
nor UO_312 (O_312,N_22655,N_24134);
xor UO_313 (O_313,N_24027,N_23229);
and UO_314 (O_314,N_23624,N_24397);
and UO_315 (O_315,N_23998,N_23395);
xnor UO_316 (O_316,N_24705,N_23316);
and UO_317 (O_317,N_23602,N_23900);
and UO_318 (O_318,N_22570,N_22841);
nor UO_319 (O_319,N_23863,N_24768);
nor UO_320 (O_320,N_23519,N_23392);
or UO_321 (O_321,N_24012,N_24290);
or UO_322 (O_322,N_24080,N_23148);
nand UO_323 (O_323,N_24890,N_22685);
nor UO_324 (O_324,N_24631,N_24842);
nor UO_325 (O_325,N_24875,N_22781);
nor UO_326 (O_326,N_22900,N_23498);
nor UO_327 (O_327,N_24431,N_24079);
nor UO_328 (O_328,N_24331,N_22615);
nor UO_329 (O_329,N_24144,N_23439);
nor UO_330 (O_330,N_22859,N_24409);
nand UO_331 (O_331,N_24097,N_24270);
or UO_332 (O_332,N_23203,N_24921);
xnor UO_333 (O_333,N_24629,N_24586);
nand UO_334 (O_334,N_23954,N_24081);
or UO_335 (O_335,N_24849,N_23614);
nand UO_336 (O_336,N_24472,N_24103);
nor UO_337 (O_337,N_22960,N_24102);
xnor UO_338 (O_338,N_24295,N_23167);
xnor UO_339 (O_339,N_23034,N_23897);
and UO_340 (O_340,N_24821,N_24158);
xnor UO_341 (O_341,N_23036,N_24509);
nor UO_342 (O_342,N_22862,N_24028);
or UO_343 (O_343,N_24478,N_22535);
or UO_344 (O_344,N_23877,N_23084);
or UO_345 (O_345,N_24621,N_24460);
nand UO_346 (O_346,N_24259,N_23755);
nand UO_347 (O_347,N_23788,N_23792);
xnor UO_348 (O_348,N_24055,N_23104);
nand UO_349 (O_349,N_24756,N_22691);
nand UO_350 (O_350,N_23225,N_24812);
and UO_351 (O_351,N_24680,N_22873);
nor UO_352 (O_352,N_24487,N_23637);
xor UO_353 (O_353,N_23159,N_22871);
or UO_354 (O_354,N_23262,N_23038);
or UO_355 (O_355,N_22919,N_22732);
nand UO_356 (O_356,N_23106,N_22503);
nor UO_357 (O_357,N_24525,N_23361);
nor UO_358 (O_358,N_24789,N_22662);
xor UO_359 (O_359,N_23537,N_24828);
nor UO_360 (O_360,N_23783,N_24815);
nand UO_361 (O_361,N_24300,N_24709);
xor UO_362 (O_362,N_22901,N_24632);
nor UO_363 (O_363,N_24316,N_24220);
or UO_364 (O_364,N_24991,N_24894);
nor UO_365 (O_365,N_22827,N_22676);
xnor UO_366 (O_366,N_22825,N_24790);
or UO_367 (O_367,N_23324,N_24507);
nand UO_368 (O_368,N_23902,N_23288);
or UO_369 (O_369,N_22564,N_24350);
nand UO_370 (O_370,N_23806,N_23941);
nand UO_371 (O_371,N_24713,N_24745);
nand UO_372 (O_372,N_23375,N_22689);
and UO_373 (O_373,N_24637,N_24784);
xor UO_374 (O_374,N_24044,N_23600);
nor UO_375 (O_375,N_24136,N_22625);
xnor UO_376 (O_376,N_24952,N_24470);
nor UO_377 (O_377,N_24612,N_24418);
nand UO_378 (O_378,N_23000,N_24223);
and UO_379 (O_379,N_24913,N_22563);
nand UO_380 (O_380,N_22745,N_23226);
xnor UO_381 (O_381,N_24513,N_24173);
nand UO_382 (O_382,N_23980,N_24857);
and UO_383 (O_383,N_22843,N_24638);
xor UO_384 (O_384,N_24663,N_24544);
or UO_385 (O_385,N_23621,N_23046);
nand UO_386 (O_386,N_24702,N_24910);
or UO_387 (O_387,N_23605,N_22800);
xnor UO_388 (O_388,N_24410,N_24859);
or UO_389 (O_389,N_24620,N_24649);
and UO_390 (O_390,N_24132,N_23144);
xnor UO_391 (O_391,N_24840,N_24778);
nor UO_392 (O_392,N_23419,N_23428);
and UO_393 (O_393,N_24734,N_24796);
xor UO_394 (O_394,N_22521,N_23119);
or UO_395 (O_395,N_24161,N_23503);
xor UO_396 (O_396,N_24823,N_23323);
xnor UO_397 (O_397,N_22815,N_23702);
and UO_398 (O_398,N_23381,N_23401);
nand UO_399 (O_399,N_24116,N_24381);
xnor UO_400 (O_400,N_23164,N_23211);
nand UO_401 (O_401,N_24695,N_23047);
or UO_402 (O_402,N_23846,N_23117);
or UO_403 (O_403,N_22587,N_23853);
nand UO_404 (O_404,N_22999,N_24391);
xor UO_405 (O_405,N_22874,N_23665);
nand UO_406 (O_406,N_24566,N_23574);
xor UO_407 (O_407,N_23663,N_22773);
nor UO_408 (O_408,N_23749,N_23158);
or UO_409 (O_409,N_23315,N_24940);
and UO_410 (O_410,N_24572,N_24762);
nand UO_411 (O_411,N_22899,N_23268);
nand UO_412 (O_412,N_22622,N_22979);
and UO_413 (O_413,N_23030,N_22584);
and UO_414 (O_414,N_23931,N_23096);
xnor UO_415 (O_415,N_24054,N_24529);
xor UO_416 (O_416,N_24959,N_24289);
and UO_417 (O_417,N_23327,N_24312);
xor UO_418 (O_418,N_24947,N_23485);
xnor UO_419 (O_419,N_23712,N_23701);
xor UO_420 (O_420,N_23831,N_24063);
nand UO_421 (O_421,N_22577,N_22633);
or UO_422 (O_422,N_24480,N_23206);
and UO_423 (O_423,N_24477,N_23732);
xor UO_424 (O_424,N_22849,N_24590);
and UO_425 (O_425,N_23176,N_23597);
or UO_426 (O_426,N_24379,N_23975);
nor UO_427 (O_427,N_24394,N_23977);
nor UO_428 (O_428,N_24899,N_23911);
nor UO_429 (O_429,N_22795,N_23328);
xor UO_430 (O_430,N_24979,N_23563);
and UO_431 (O_431,N_23072,N_22935);
or UO_432 (O_432,N_23180,N_24962);
xnor UO_433 (O_433,N_23849,N_24994);
xnor UO_434 (O_434,N_23027,N_24992);
or UO_435 (O_435,N_23468,N_24628);
or UO_436 (O_436,N_23525,N_22986);
or UO_437 (O_437,N_24412,N_23920);
xnor UO_438 (O_438,N_23111,N_23389);
xnor UO_439 (O_439,N_23884,N_22566);
or UO_440 (O_440,N_24623,N_24847);
xnor UO_441 (O_441,N_23001,N_23150);
nand UO_442 (O_442,N_24110,N_22549);
nor UO_443 (O_443,N_23151,N_23223);
or UO_444 (O_444,N_22969,N_22614);
nand UO_445 (O_445,N_23646,N_24912);
and UO_446 (O_446,N_24341,N_24583);
nor UO_447 (O_447,N_23329,N_24239);
and UO_448 (O_448,N_22820,N_23198);
nor UO_449 (O_449,N_23273,N_23488);
xor UO_450 (O_450,N_24127,N_22648);
nor UO_451 (O_451,N_23876,N_22505);
nor UO_452 (O_452,N_23252,N_22955);
and UO_453 (O_453,N_23214,N_22610);
and UO_454 (O_454,N_24182,N_22783);
or UO_455 (O_455,N_23173,N_22520);
nand UO_456 (O_456,N_23196,N_24985);
and UO_457 (O_457,N_23764,N_24682);
nor UO_458 (O_458,N_23782,N_23664);
or UO_459 (O_459,N_24711,N_24771);
xor UO_460 (O_460,N_23358,N_24958);
and UO_461 (O_461,N_24451,N_23094);
nand UO_462 (O_462,N_22784,N_23271);
nor UO_463 (O_463,N_24384,N_24288);
or UO_464 (O_464,N_23917,N_23889);
xor UO_465 (O_465,N_24210,N_23759);
nand UO_466 (O_466,N_24963,N_22778);
nand UO_467 (O_467,N_23641,N_22641);
xnor UO_468 (O_468,N_24183,N_22941);
and UO_469 (O_469,N_24650,N_24681);
nand UO_470 (O_470,N_24904,N_24494);
nor UO_471 (O_471,N_24266,N_23175);
xnor UO_472 (O_472,N_23769,N_23933);
and UO_473 (O_473,N_24944,N_24464);
or UO_474 (O_474,N_24309,N_22525);
xor UO_475 (O_475,N_23584,N_22818);
and UO_476 (O_476,N_24057,N_23133);
xor UO_477 (O_477,N_23177,N_23613);
nor UO_478 (O_478,N_23811,N_22762);
nor UO_479 (O_479,N_24861,N_24953);
nor UO_480 (O_480,N_24614,N_23512);
or UO_481 (O_481,N_23922,N_24788);
nor UO_482 (O_482,N_23822,N_24589);
nand UO_483 (O_483,N_23533,N_22981);
nand UO_484 (O_484,N_22541,N_24925);
nand UO_485 (O_485,N_24317,N_24401);
and UO_486 (O_486,N_24508,N_24616);
or UO_487 (O_487,N_24207,N_23891);
or UO_488 (O_488,N_24708,N_24492);
nor UO_489 (O_489,N_23056,N_24056);
xor UO_490 (O_490,N_24491,N_24588);
or UO_491 (O_491,N_23694,N_22522);
xnor UO_492 (O_492,N_24797,N_23475);
or UO_493 (O_493,N_24898,N_24678);
or UO_494 (O_494,N_23386,N_23586);
nor UO_495 (O_495,N_23894,N_24719);
nand UO_496 (O_496,N_23018,N_22742);
nand UO_497 (O_497,N_23248,N_24533);
nand UO_498 (O_498,N_22713,N_23979);
xor UO_499 (O_499,N_22814,N_23815);
nor UO_500 (O_500,N_23653,N_24113);
and UO_501 (O_501,N_24126,N_24688);
and UO_502 (O_502,N_22734,N_24560);
xnor UO_503 (O_503,N_24886,N_22848);
nor UO_504 (O_504,N_22710,N_23675);
or UO_505 (O_505,N_22692,N_24945);
nand UO_506 (O_506,N_22988,N_23948);
nor UO_507 (O_507,N_22945,N_23179);
or UO_508 (O_508,N_22510,N_22994);
and UO_509 (O_509,N_23882,N_23629);
and UO_510 (O_510,N_22513,N_24909);
nor UO_511 (O_511,N_23504,N_23859);
xnor UO_512 (O_512,N_23581,N_24520);
nand UO_513 (O_513,N_24030,N_23341);
and UO_514 (O_514,N_22936,N_22519);
nand UO_515 (O_515,N_24824,N_23723);
xnor UO_516 (O_516,N_24982,N_23710);
xor UO_517 (O_517,N_24939,N_24655);
nand UO_518 (O_518,N_24420,N_24757);
and UO_519 (O_519,N_23400,N_22529);
and UO_520 (O_520,N_23818,N_23032);
and UO_521 (O_521,N_23677,N_24167);
nor UO_522 (O_522,N_24354,N_24814);
xor UO_523 (O_523,N_24066,N_24807);
xnor UO_524 (O_524,N_23193,N_24343);
or UO_525 (O_525,N_22716,N_24670);
and UO_526 (O_526,N_24274,N_23858);
nor UO_527 (O_527,N_22683,N_24352);
and UO_528 (O_528,N_23295,N_22611);
and UO_529 (O_529,N_24869,N_24303);
nand UO_530 (O_530,N_23235,N_22630);
or UO_531 (O_531,N_22840,N_22976);
xnor UO_532 (O_532,N_24998,N_23244);
nor UO_533 (O_533,N_23108,N_23893);
xnor UO_534 (O_534,N_24114,N_23114);
xor UO_535 (O_535,N_24744,N_24522);
and UO_536 (O_536,N_22772,N_22523);
xnor UO_537 (O_537,N_24794,N_24128);
and UO_538 (O_538,N_23970,N_23185);
nor UO_539 (O_539,N_23542,N_23307);
nor UO_540 (O_540,N_22653,N_23074);
xnor UO_541 (O_541,N_23828,N_23603);
nand UO_542 (O_542,N_24247,N_23050);
nand UO_543 (O_543,N_24100,N_24233);
nor UO_544 (O_544,N_24094,N_23457);
nand UO_545 (O_545,N_22723,N_23446);
and UO_546 (O_546,N_23671,N_23964);
xnor UO_547 (O_547,N_23555,N_23153);
and UO_548 (O_548,N_23418,N_24218);
nor UO_549 (O_549,N_24811,N_23182);
xor UO_550 (O_550,N_24272,N_24485);
or UO_551 (O_551,N_22504,N_24701);
nand UO_552 (O_552,N_24698,N_22816);
and UO_553 (O_553,N_22974,N_24162);
or UO_554 (O_554,N_22752,N_23999);
and UO_555 (O_555,N_22686,N_23025);
and UO_556 (O_556,N_23057,N_24465);
nor UO_557 (O_557,N_22599,N_24934);
nand UO_558 (O_558,N_23209,N_23350);
and UO_559 (O_559,N_23014,N_24064);
nand UO_560 (O_560,N_24195,N_24881);
and UO_561 (O_561,N_23140,N_23443);
nand UO_562 (O_562,N_23885,N_24493);
xnor UO_563 (O_563,N_22586,N_23746);
or UO_564 (O_564,N_24388,N_23538);
or UO_565 (O_565,N_23043,N_22911);
nor UO_566 (O_566,N_23741,N_23310);
nand UO_567 (O_567,N_22606,N_22834);
and UO_568 (O_568,N_23727,N_22687);
nand UO_569 (O_569,N_22731,N_22856);
xor UO_570 (O_570,N_23467,N_23130);
and UO_571 (O_571,N_24376,N_23091);
nor UO_572 (O_572,N_24935,N_24301);
or UO_573 (O_573,N_24137,N_24538);
nand UO_574 (O_574,N_23843,N_24511);
xnor UO_575 (O_575,N_23070,N_24084);
and UO_576 (O_576,N_23554,N_24201);
nor UO_577 (O_577,N_22951,N_24117);
nand UO_578 (O_578,N_24178,N_23730);
or UO_579 (O_579,N_24610,N_23342);
nor UO_580 (O_580,N_24730,N_22639);
or UO_581 (O_581,N_23856,N_23178);
xor UO_582 (O_582,N_24353,N_22500);
and UO_583 (O_583,N_24832,N_24603);
or UO_584 (O_584,N_23487,N_22557);
and UO_585 (O_585,N_23236,N_23189);
and UO_586 (O_586,N_22927,N_24276);
nand UO_587 (O_587,N_23274,N_24125);
and UO_588 (O_588,N_23053,N_22963);
or UO_589 (O_589,N_24361,N_22763);
xor UO_590 (O_590,N_22507,N_23420);
nor UO_591 (O_591,N_23230,N_24265);
and UO_592 (O_592,N_24009,N_23672);
and UO_593 (O_593,N_23966,N_24372);
xor UO_594 (O_594,N_24031,N_22569);
nand UO_595 (O_595,N_23655,N_23905);
nor UO_596 (O_596,N_22601,N_23169);
and UO_597 (O_597,N_24122,N_22560);
xor UO_598 (O_598,N_23816,N_22515);
nor UO_599 (O_599,N_22670,N_24327);
xnor UO_600 (O_600,N_23718,N_24407);
or UO_601 (O_601,N_24160,N_23790);
nand UO_602 (O_602,N_23166,N_23874);
nand UO_603 (O_603,N_22637,N_24232);
and UO_604 (O_604,N_23097,N_23559);
nor UO_605 (O_605,N_23330,N_23714);
nand UO_606 (O_606,N_24786,N_23550);
and UO_607 (O_607,N_22993,N_23797);
or UO_608 (O_608,N_23765,N_22939);
xnor UO_609 (O_609,N_24911,N_23388);
nor UO_610 (O_610,N_23497,N_24396);
and UO_611 (O_611,N_23284,N_23852);
xor UO_612 (O_612,N_23285,N_23101);
nand UO_613 (O_613,N_23851,N_24019);
nand UO_614 (O_614,N_24186,N_24311);
xor UO_615 (O_615,N_23093,N_23194);
or UO_616 (O_616,N_23928,N_23565);
xnor UO_617 (O_617,N_22699,N_24332);
nor UO_618 (O_618,N_24278,N_24374);
nand UO_619 (O_619,N_23069,N_24918);
xnor UO_620 (O_620,N_22913,N_23345);
and UO_621 (O_621,N_24506,N_23146);
nor UO_622 (O_622,N_23578,N_23029);
xor UO_623 (O_623,N_24720,N_23875);
and UO_624 (O_624,N_23832,N_24328);
nand UO_625 (O_625,N_22920,N_23243);
or UO_626 (O_626,N_22830,N_23781);
nor UO_627 (O_627,N_23780,N_24770);
or UO_628 (O_628,N_23842,N_23553);
and UO_629 (O_629,N_23452,N_24831);
nand UO_630 (O_630,N_23684,N_24554);
and UO_631 (O_631,N_23738,N_24826);
nor UO_632 (O_632,N_23374,N_24348);
or UO_633 (O_633,N_22527,N_23955);
nand UO_634 (O_634,N_24524,N_23919);
and UO_635 (O_635,N_23636,N_24602);
nand UO_636 (O_636,N_23872,N_23065);
nor UO_637 (O_637,N_24887,N_24366);
or UO_638 (O_638,N_23390,N_22697);
nor UO_639 (O_639,N_23410,N_23609);
and UO_640 (O_640,N_24010,N_23910);
or UO_641 (O_641,N_23857,N_24753);
nand UO_642 (O_642,N_22627,N_22688);
or UO_643 (O_643,N_22526,N_23841);
xnor UO_644 (O_644,N_24033,N_23720);
or UO_645 (O_645,N_22678,N_24474);
xnor UO_646 (O_646,N_22597,N_22774);
and UO_647 (O_647,N_24883,N_23576);
xnor UO_648 (O_648,N_24078,N_23415);
nand UO_649 (O_649,N_23593,N_24075);
nand UO_650 (O_650,N_23434,N_23351);
nand UO_651 (O_651,N_24987,N_22727);
or UO_652 (O_652,N_24355,N_23957);
xnor UO_653 (O_653,N_23662,N_24335);
xnor UO_654 (O_654,N_23992,N_24435);
nor UO_655 (O_655,N_22501,N_22640);
xnor UO_656 (O_656,N_23021,N_23628);
xor UO_657 (O_657,N_23867,N_22668);
and UO_658 (O_658,N_22953,N_22847);
nand UO_659 (O_659,N_24155,N_24715);
or UO_660 (O_660,N_24129,N_24001);
and UO_661 (O_661,N_24241,N_24193);
nand UO_662 (O_662,N_22604,N_24683);
or UO_663 (O_663,N_24086,N_23493);
xnor UO_664 (O_664,N_24243,N_24250);
nand UO_665 (O_665,N_22987,N_23927);
or UO_666 (O_666,N_23016,N_24499);
and UO_667 (O_667,N_23945,N_22748);
xnor UO_668 (O_668,N_24449,N_24532);
nor UO_669 (O_669,N_22554,N_22537);
xor UO_670 (O_670,N_23432,N_24652);
or UO_671 (O_671,N_23040,N_24986);
xor UO_672 (O_672,N_24497,N_24848);
xor UO_673 (O_673,N_23520,N_23650);
or UO_674 (O_674,N_23118,N_24721);
nor UO_675 (O_675,N_24269,N_22910);
and UO_676 (O_676,N_24725,N_24471);
nand UO_677 (O_677,N_23854,N_24236);
xor UO_678 (O_678,N_23076,N_23482);
xor UO_679 (O_679,N_23068,N_22798);
and UO_680 (O_680,N_23569,N_22858);
and UO_681 (O_681,N_22908,N_23125);
nand UO_682 (O_682,N_22878,N_23777);
and UO_683 (O_683,N_22984,N_22675);
xor UO_684 (O_684,N_24641,N_24286);
nand UO_685 (O_685,N_23474,N_22756);
nand UO_686 (O_686,N_23269,N_24850);
nor UO_687 (O_687,N_22644,N_24395);
or UO_688 (O_688,N_23988,N_23862);
xnor UO_689 (O_689,N_22802,N_24013);
nor UO_690 (O_690,N_23082,N_23800);
or UO_691 (O_691,N_22718,N_24844);
and UO_692 (O_692,N_24181,N_22851);
xor UO_693 (O_693,N_23833,N_24408);
and UO_694 (O_694,N_22562,N_24622);
or UO_695 (O_695,N_24310,N_23855);
nand UO_696 (O_696,N_24285,N_22817);
xnor UO_697 (O_697,N_23616,N_22573);
and UO_698 (O_698,N_22624,N_22958);
or UO_699 (O_699,N_23959,N_24868);
nand UO_700 (O_700,N_24004,N_22583);
nor UO_701 (O_701,N_24889,N_24463);
xor UO_702 (O_702,N_23864,N_24037);
nand UO_703 (O_703,N_24906,N_24106);
nor UO_704 (O_704,N_24307,N_22719);
and UO_705 (O_705,N_24989,N_24627);
and UO_706 (O_706,N_23170,N_23560);
or UO_707 (O_707,N_23956,N_24046);
nand UO_708 (O_708,N_22854,N_23921);
nand UO_709 (O_709,N_23708,N_24710);
xor UO_710 (O_710,N_23756,N_23936);
nor UO_711 (O_711,N_23253,N_22990);
xnor UO_712 (O_712,N_23261,N_24642);
nand UO_713 (O_713,N_24405,N_24433);
and UO_714 (O_714,N_24432,N_23699);
or UO_715 (O_715,N_24743,N_23745);
nand UO_716 (O_716,N_23978,N_23004);
nor UO_717 (O_717,N_22509,N_24153);
or UO_718 (O_718,N_23706,N_23102);
xor UO_719 (O_719,N_23008,N_23985);
xnor UO_720 (O_720,N_24592,N_22511);
xor UO_721 (O_721,N_22530,N_23062);
xor UO_722 (O_722,N_23338,N_23987);
or UO_723 (O_723,N_24597,N_23617);
nor UO_724 (O_724,N_24230,N_24799);
nor UO_725 (O_725,N_24932,N_24154);
or UO_726 (O_726,N_23321,N_24500);
nand UO_727 (O_727,N_24147,N_24007);
nor UO_728 (O_728,N_22555,N_24159);
or UO_729 (O_729,N_22898,N_23272);
and UO_730 (O_730,N_23417,N_24690);
nand UO_731 (O_731,N_23935,N_24228);
and UO_732 (O_732,N_23809,N_23993);
nand UO_733 (O_733,N_22565,N_22982);
and UO_734 (O_734,N_24021,N_22589);
and UO_735 (O_735,N_23680,N_23044);
and UO_736 (O_736,N_23456,N_23208);
nand UO_737 (O_737,N_23080,N_24564);
xnor UO_738 (O_738,N_24581,N_23045);
or UO_739 (O_739,N_22780,N_24439);
nor UO_740 (O_740,N_23962,N_24133);
nand UO_741 (O_741,N_24398,N_23700);
nor UO_742 (O_742,N_23753,N_22531);
and UO_743 (O_743,N_23620,N_24071);
or UO_744 (O_744,N_24679,N_24245);
or UO_745 (O_745,N_24539,N_23455);
nor UO_746 (O_746,N_24504,N_23622);
and UO_747 (O_747,N_24562,N_23378);
nand UO_748 (O_748,N_24598,N_23347);
nor UO_749 (O_749,N_24336,N_24946);
xor UO_750 (O_750,N_24924,N_23761);
nor UO_751 (O_751,N_23063,N_24072);
nand UO_752 (O_752,N_24337,N_24319);
or UO_753 (O_753,N_24841,N_23638);
xnor UO_754 (O_754,N_24801,N_22886);
xnor UO_755 (O_755,N_24257,N_24659);
xor UO_756 (O_756,N_23562,N_23656);
and UO_757 (O_757,N_24526,N_22609);
nor UO_758 (O_758,N_22728,N_22553);
nor UO_759 (O_759,N_22842,N_23059);
xnor UO_760 (O_760,N_22626,N_22620);
and UO_761 (O_761,N_23052,N_23731);
and UO_762 (O_762,N_23383,N_23767);
and UO_763 (O_763,N_22666,N_23258);
nand UO_764 (O_764,N_22634,N_23791);
and UO_765 (O_765,N_23532,N_23478);
and UO_766 (O_766,N_23661,N_23514);
and UO_767 (O_767,N_24489,N_23266);
and UO_768 (O_768,N_24908,N_23526);
or UO_769 (O_769,N_24287,N_23309);
or UO_770 (O_770,N_23996,N_24706);
or UO_771 (O_771,N_23399,N_24119);
nor UO_772 (O_772,N_22512,N_22991);
xnor UO_773 (O_773,N_23406,N_22695);
and UO_774 (O_774,N_24965,N_23789);
xnor UO_775 (O_775,N_23188,N_22998);
nand UO_776 (O_776,N_23698,N_24141);
or UO_777 (O_777,N_24051,N_24880);
nand UO_778 (O_778,N_24860,N_22673);
nor UO_779 (O_779,N_22805,N_24253);
and UO_780 (O_780,N_24838,N_24878);
or UO_781 (O_781,N_22558,N_24557);
and UO_782 (O_782,N_24541,N_22877);
nand UO_783 (O_783,N_24192,N_24061);
nor UO_784 (O_784,N_24124,N_23020);
or UO_785 (O_785,N_24975,N_23202);
or UO_786 (O_786,N_24422,N_22613);
nand UO_787 (O_787,N_24648,N_24866);
nor UO_788 (O_788,N_23729,N_24226);
and UO_789 (O_789,N_24262,N_23500);
and UO_790 (O_790,N_23580,N_24677);
nor UO_791 (O_791,N_24964,N_23949);
nor UO_792 (O_792,N_24115,N_24950);
and UO_793 (O_793,N_24510,N_24846);
or UO_794 (O_794,N_24473,N_23691);
xnor UO_795 (O_795,N_22636,N_22907);
and UO_796 (O_796,N_23424,N_24853);
nor UO_797 (O_797,N_23186,N_24015);
and UO_798 (O_798,N_23233,N_22698);
or UO_799 (O_799,N_23458,N_24867);
nand UO_800 (O_800,N_24625,N_24644);
xor UO_801 (O_801,N_24087,N_24291);
or UO_802 (O_802,N_24248,N_24613);
nor UO_803 (O_803,N_22931,N_24550);
or UO_804 (O_804,N_23901,N_23088);
nor UO_805 (O_805,N_24142,N_24314);
xnor UO_806 (O_806,N_24741,N_24467);
xor UO_807 (O_807,N_22790,N_23496);
nand UO_808 (O_808,N_23019,N_23734);
xor UO_809 (O_809,N_24457,N_24425);
and UO_810 (O_810,N_24399,N_24856);
xor UO_811 (O_811,N_23212,N_24700);
and UO_812 (O_812,N_23908,N_22822);
xor UO_813 (O_813,N_24299,N_22714);
and UO_814 (O_814,N_24579,N_23903);
xor UO_815 (O_815,N_24654,N_23573);
nand UO_816 (O_816,N_24540,N_23944);
and UO_817 (O_817,N_23131,N_24549);
or UO_818 (O_818,N_23615,N_24038);
or UO_819 (O_819,N_23567,N_22869);
or UO_820 (O_820,N_23591,N_24271);
nand UO_821 (O_821,N_22777,N_23480);
or UO_822 (O_822,N_23878,N_24334);
xnor UO_823 (O_823,N_22647,N_22855);
and UO_824 (O_824,N_24763,N_23465);
nand UO_825 (O_825,N_24249,N_23839);
and UO_826 (O_826,N_23484,N_24966);
nand UO_827 (O_827,N_23009,N_23311);
nand UO_828 (O_828,N_23518,N_23472);
nand UO_829 (O_829,N_23363,N_24558);
xnor UO_830 (O_830,N_22918,N_24156);
xor UO_831 (O_831,N_24073,N_22681);
nand UO_832 (O_832,N_23509,N_22950);
xnor UO_833 (O_833,N_24961,N_24008);
nand UO_834 (O_834,N_23370,N_24988);
and UO_835 (O_835,N_24661,N_24176);
or UO_836 (O_836,N_23326,N_24029);
xnor UO_837 (O_837,N_23942,N_24313);
or UO_838 (O_838,N_23486,N_24459);
xor UO_839 (O_839,N_22514,N_24739);
xor UO_840 (O_840,N_24242,N_24703);
or UO_841 (O_841,N_23748,N_22883);
nor UO_842 (O_842,N_22605,N_23994);
xor UO_843 (O_843,N_23564,N_24926);
xnor UO_844 (O_844,N_23464,N_24949);
or UO_845 (O_845,N_23515,N_22767);
and UO_846 (O_846,N_23696,N_24851);
and UO_847 (O_847,N_22674,N_24561);
xor UO_848 (O_848,N_24839,N_24371);
or UO_849 (O_849,N_24601,N_23191);
nand UO_850 (O_850,N_23377,N_24955);
nor UO_851 (O_851,N_23291,N_24587);
or UO_852 (O_852,N_24545,N_22972);
nand UO_853 (O_853,N_23135,N_22612);
and UO_854 (O_854,N_24052,N_23280);
nor UO_855 (O_855,N_24197,N_23909);
xor UO_856 (O_856,N_22959,N_23129);
or UO_857 (O_857,N_23508,N_22664);
xor UO_858 (O_858,N_24490,N_23098);
nand UO_859 (O_859,N_23695,N_22811);
and UO_860 (O_860,N_23215,N_24535);
nor UO_861 (O_861,N_24039,N_23566);
nor UO_862 (O_862,N_24971,N_24326);
and UO_863 (O_863,N_23222,N_23850);
xnor UO_864 (O_864,N_22669,N_23660);
xor UO_865 (O_865,N_23275,N_23751);
nand UO_866 (O_866,N_23250,N_24131);
nor UO_867 (O_867,N_22518,N_22659);
nor UO_868 (O_868,N_22568,N_23703);
nor UO_869 (O_869,N_23259,N_22621);
nor UO_870 (O_870,N_23571,N_24984);
xor UO_871 (O_871,N_24954,N_24704);
nor UO_872 (O_872,N_24450,N_23017);
nand UO_873 (O_873,N_23301,N_22975);
or UO_874 (O_874,N_23155,N_23302);
or UO_875 (O_875,N_22846,N_22997);
nand UO_876 (O_876,N_24189,N_22572);
and UO_877 (O_877,N_24445,N_24488);
nand UO_878 (O_878,N_22646,N_23642);
nor UO_879 (O_879,N_23687,N_23461);
and UO_880 (O_880,N_24822,N_22968);
nor UO_881 (O_881,N_23296,N_23965);
or UO_882 (O_882,N_23451,N_23930);
xnor UO_883 (O_883,N_24392,N_22977);
or UO_884 (O_884,N_24724,N_24609);
nand UO_885 (O_885,N_24606,N_22870);
nand UO_886 (O_886,N_23681,N_23635);
nand UO_887 (O_887,N_23218,N_24345);
and UO_888 (O_888,N_23154,N_24594);
and UO_889 (O_889,N_22693,N_23547);
or UO_890 (O_890,N_24897,N_23535);
or UO_891 (O_891,N_23824,N_24370);
and UO_892 (O_892,N_23002,N_24580);
and UO_893 (O_893,N_24968,N_24750);
xor UO_894 (O_894,N_23716,N_23200);
xor UO_895 (O_895,N_22544,N_22828);
xor UO_896 (O_896,N_23366,N_24437);
nor UO_897 (O_897,N_24758,N_22875);
nand UO_898 (O_898,N_22799,N_24351);
xnor UO_899 (O_899,N_22730,N_23848);
nand UO_900 (O_900,N_23099,N_23668);
nand UO_901 (O_901,N_24320,N_24923);
nand UO_902 (O_902,N_23448,N_23914);
and UO_903 (O_903,N_22744,N_22708);
nor UO_904 (O_904,N_22733,N_22890);
nor UO_905 (O_905,N_23599,N_24542);
nand UO_906 (O_906,N_23802,N_24498);
nand UO_907 (O_907,N_22749,N_23923);
nor UO_908 (O_908,N_23409,N_22603);
or UO_909 (O_909,N_22971,N_24416);
nor UO_910 (O_910,N_22970,N_23938);
or UO_911 (O_911,N_22835,N_22812);
nor UO_912 (O_912,N_24803,N_24737);
nor UO_913 (O_913,N_24020,N_24468);
or UO_914 (O_914,N_23071,N_23255);
xnor UO_915 (O_915,N_23079,N_22720);
xor UO_916 (O_916,N_23249,N_22895);
nand UO_917 (O_917,N_24876,N_23337);
nand UO_918 (O_918,N_23898,N_24684);
xor UO_919 (O_919,N_24551,N_23105);
nor UO_920 (O_920,N_23314,N_24686);
xnor UO_921 (O_921,N_24415,N_22740);
nand UO_922 (O_922,N_24085,N_24017);
nor UO_923 (O_923,N_24707,N_23502);
and UO_924 (O_924,N_22889,N_23061);
nor UO_925 (O_925,N_24495,N_24306);
and UO_926 (O_926,N_24329,N_24782);
nand UO_927 (O_927,N_23254,N_24254);
and UO_928 (O_928,N_24139,N_24349);
or UO_929 (O_929,N_23692,N_24854);
or UO_930 (O_930,N_23707,N_23590);
or UO_931 (O_931,N_23879,N_23915);
xor UO_932 (O_932,N_22824,N_22940);
and UO_933 (O_933,N_23583,N_23231);
or UO_934 (O_934,N_24833,N_22882);
nand UO_935 (O_935,N_23847,N_23634);
and UO_936 (O_936,N_22533,N_24990);
nor UO_937 (O_937,N_24779,N_24969);
nand UO_938 (O_938,N_24571,N_22961);
xor UO_939 (O_939,N_22751,N_24773);
nor UO_940 (O_940,N_24179,N_24776);
or UO_941 (O_941,N_24025,N_24528);
and UO_942 (O_942,N_24121,N_24213);
and UO_943 (O_943,N_24475,N_22743);
and UO_944 (O_944,N_24727,N_24212);
or UO_945 (O_945,N_23060,N_24456);
or UO_946 (O_946,N_23513,N_22540);
or UO_947 (O_947,N_23633,N_24003);
or UO_948 (O_948,N_22665,N_24479);
nor UO_949 (O_949,N_24292,N_24792);
xnor UO_950 (O_950,N_23845,N_22944);
nor UO_951 (O_951,N_23631,N_24111);
or UO_952 (O_952,N_23109,N_23003);
or UO_953 (O_953,N_22864,N_23049);
or UO_954 (O_954,N_23871,N_22915);
xor UO_955 (O_955,N_24933,N_24305);
and UO_956 (O_956,N_22906,N_23762);
and UO_957 (O_957,N_24002,N_23095);
xnor UO_958 (O_958,N_23367,N_23568);
and UO_959 (O_959,N_22921,N_22594);
or UO_960 (O_960,N_24096,N_22912);
nor UO_961 (O_961,N_24268,N_23495);
nor UO_962 (O_962,N_24981,N_24076);
nor UO_963 (O_963,N_22788,N_23736);
nand UO_964 (O_964,N_23676,N_24818);
and UO_965 (O_965,N_24203,N_24382);
xor UO_966 (O_966,N_24175,N_24956);
nor UO_967 (O_967,N_24235,N_24430);
xor UO_968 (O_968,N_24404,N_22768);
nor UO_969 (O_969,N_23643,N_23521);
nand UO_970 (O_970,N_24548,N_24476);
or UO_971 (O_971,N_23081,N_24206);
and UO_972 (O_972,N_24748,N_23132);
xor UO_973 (O_973,N_22619,N_24793);
xnor UO_974 (O_974,N_23217,N_24093);
and UO_975 (O_975,N_23116,N_23429);
nand UO_976 (O_976,N_23489,N_22929);
xor UO_977 (O_977,N_22657,N_24090);
nand UO_978 (O_978,N_22914,N_23332);
xor UO_979 (O_979,N_22729,N_22598);
nand UO_980 (O_980,N_23579,N_23861);
nor UO_981 (O_981,N_23481,N_23785);
nor UO_982 (O_982,N_22707,N_22808);
xor UO_983 (O_983,N_23670,N_24118);
nor UO_984 (O_984,N_23237,N_24000);
nor UO_985 (O_985,N_22705,N_23838);
or UO_986 (O_986,N_24006,N_23570);
xnor UO_987 (O_987,N_24595,N_23015);
or UO_988 (O_988,N_24191,N_23270);
or UO_989 (O_989,N_24148,N_23207);
or UO_990 (O_990,N_23997,N_24692);
nor UO_991 (O_991,N_22797,N_24216);
xnor UO_992 (O_992,N_24024,N_23090);
or UO_993 (O_993,N_24041,N_23786);
nand UO_994 (O_994,N_23912,N_23673);
xnor UO_995 (O_995,N_22704,N_23369);
or UO_996 (O_996,N_23773,N_24344);
nor UO_997 (O_997,N_22737,N_23411);
or UO_998 (O_998,N_24204,N_23372);
nand UO_999 (O_999,N_23067,N_22700);
xnor UO_1000 (O_1000,N_24225,N_23139);
nand UO_1001 (O_1001,N_22660,N_22803);
and UO_1002 (O_1002,N_22551,N_24543);
nor UO_1003 (O_1003,N_24088,N_24403);
xnor UO_1004 (O_1004,N_24138,N_23344);
and UO_1005 (O_1005,N_24169,N_24215);
or UO_1006 (O_1006,N_24593,N_23408);
or UO_1007 (O_1007,N_23768,N_24229);
and UO_1008 (O_1008,N_23444,N_24152);
nand UO_1009 (O_1009,N_24619,N_22631);
or UO_1010 (O_1010,N_22602,N_24761);
xor UO_1011 (O_1011,N_24877,N_23934);
or UO_1012 (O_1012,N_22925,N_23805);
xnor UO_1013 (O_1013,N_24357,N_24905);
xor UO_1014 (O_1014,N_23582,N_23865);
or UO_1015 (O_1015,N_23950,N_23142);
or UO_1016 (O_1016,N_24608,N_23238);
xnor UO_1017 (O_1017,N_22722,N_24323);
nor UO_1018 (O_1018,N_24884,N_24657);
nand UO_1019 (O_1019,N_24256,N_23834);
or UO_1020 (O_1020,N_24574,N_24069);
nand UO_1021 (O_1021,N_24664,N_22796);
and UO_1022 (O_1022,N_23825,N_23292);
xor UO_1023 (O_1023,N_22596,N_23608);
or UO_1024 (O_1024,N_24240,N_23627);
nand UO_1025 (O_1025,N_24238,N_23240);
nand UO_1026 (O_1026,N_24600,N_22658);
nand UO_1027 (O_1027,N_24559,N_24903);
nor UO_1028 (O_1028,N_23726,N_24671);
nand UO_1029 (O_1029,N_24942,N_22709);
and UO_1030 (O_1030,N_24378,N_23625);
xnor UO_1031 (O_1031,N_23385,N_23813);
nand UO_1032 (O_1032,N_24993,N_24427);
and UO_1033 (O_1033,N_24237,N_22738);
and UO_1034 (O_1034,N_24123,N_24974);
or UO_1035 (O_1035,N_23951,N_23449);
xor UO_1036 (O_1036,N_24666,N_23835);
nand UO_1037 (O_1037,N_24736,N_23953);
and UO_1038 (O_1038,N_23396,N_23793);
nand UO_1039 (O_1039,N_24885,N_24527);
xor UO_1040 (O_1040,N_24845,N_23138);
nand UO_1041 (O_1041,N_23943,N_24426);
or UO_1042 (O_1042,N_23557,N_24536);
nor UO_1043 (O_1043,N_23277,N_23232);
or UO_1044 (O_1044,N_24034,N_22764);
nor UO_1045 (O_1045,N_23630,N_23357);
or UO_1046 (O_1046,N_23705,N_23441);
or UO_1047 (O_1047,N_24304,N_23556);
nand UO_1048 (O_1048,N_22717,N_24180);
nand UO_1049 (O_1049,N_24749,N_22881);
xnor UO_1050 (O_1050,N_24764,N_23546);
or UO_1051 (O_1051,N_23880,N_24997);
xnor UO_1052 (O_1052,N_24514,N_23976);
or UO_1053 (O_1053,N_24819,N_22866);
and UO_1054 (O_1054,N_23946,N_23750);
or UO_1055 (O_1055,N_23774,N_23728);
and UO_1056 (O_1056,N_24901,N_23163);
nand UO_1057 (O_1057,N_23715,N_24505);
or UO_1058 (O_1058,N_24164,N_22545);
xnor UO_1059 (O_1059,N_24049,N_23263);
xnor UO_1060 (O_1060,N_23042,N_22766);
nand UO_1061 (O_1061,N_23869,N_23183);
or UO_1062 (O_1062,N_22836,N_24732);
and UO_1063 (O_1063,N_24016,N_24387);
and UO_1064 (O_1064,N_23397,N_23644);
xnor UO_1065 (O_1065,N_24873,N_23510);
or UO_1066 (O_1066,N_23541,N_23645);
and UO_1067 (O_1067,N_24330,N_24872);
xor UO_1068 (O_1068,N_24458,N_23860);
and UO_1069 (O_1069,N_24149,N_23658);
nor UO_1070 (O_1070,N_23174,N_23763);
nor UO_1071 (O_1071,N_23659,N_24646);
and UO_1072 (O_1072,N_24611,N_24938);
nor UO_1073 (O_1073,N_22672,N_24553);
or UO_1074 (O_1074,N_24050,N_23172);
or UO_1075 (O_1075,N_24970,N_22943);
nand UO_1076 (O_1076,N_22618,N_23124);
xnor UO_1077 (O_1077,N_23317,N_23798);
or UO_1078 (O_1078,N_24640,N_24177);
or UO_1079 (O_1079,N_23416,N_24150);
and UO_1080 (O_1080,N_23607,N_22838);
and UO_1081 (O_1081,N_22922,N_22528);
nor UO_1082 (O_1082,N_22833,N_23722);
nand UO_1083 (O_1083,N_22550,N_24742);
or UO_1084 (O_1084,N_22581,N_24531);
or UO_1085 (O_1085,N_24747,N_23421);
and UO_1086 (O_1086,N_24907,N_22548);
or UO_1087 (O_1087,N_23754,N_22832);
nor UO_1088 (O_1088,N_24095,N_23380);
and UO_1089 (O_1089,N_24636,N_23772);
nand UO_1090 (O_1090,N_24517,N_23359);
xnor UO_1091 (O_1091,N_23427,N_24780);
xnor UO_1092 (O_1092,N_22502,N_24339);
nand UO_1093 (O_1093,N_23821,N_24634);
nor UO_1094 (O_1094,N_23604,N_22992);
nor UO_1095 (O_1095,N_24760,N_22872);
nor UO_1096 (O_1096,N_23787,N_24662);
or UO_1097 (O_1097,N_24219,N_23906);
nor UO_1098 (O_1098,N_22887,N_22682);
or UO_1099 (O_1099,N_24453,N_24340);
xor UO_1100 (O_1100,N_23265,N_24424);
and UO_1101 (O_1101,N_23210,N_23450);
nor UO_1102 (O_1102,N_22896,N_22556);
xor UO_1103 (O_1103,N_23592,N_24643);
or UO_1104 (O_1104,N_23051,N_22684);
nand UO_1105 (O_1105,N_23958,N_23181);
nor UO_1106 (O_1106,N_24943,N_23752);
nand UO_1107 (O_1107,N_24941,N_23827);
nand UO_1108 (O_1108,N_22905,N_24022);
xor UO_1109 (O_1109,N_24759,N_22938);
nand UO_1110 (O_1110,N_23251,N_24174);
nand UO_1111 (O_1111,N_24879,N_22978);
and UO_1112 (O_1112,N_24386,N_23422);
and UO_1113 (O_1113,N_22632,N_24674);
and UO_1114 (O_1114,N_23005,N_22926);
or UO_1115 (O_1115,N_23245,N_22561);
xor UO_1116 (O_1116,N_24547,N_24633);
or UO_1117 (O_1117,N_23078,N_24429);
nor UO_1118 (O_1118,N_22582,N_23048);
xnor UO_1119 (O_1119,N_23505,N_23320);
xor UO_1120 (O_1120,N_24863,N_23161);
nand UO_1121 (O_1121,N_22829,N_23572);
nor UO_1122 (O_1122,N_22967,N_23318);
nand UO_1123 (O_1123,N_22576,N_22909);
nor UO_1124 (O_1124,N_23360,N_24438);
or UO_1125 (O_1125,N_24446,N_23157);
nand UO_1126 (O_1126,N_24687,N_23795);
and UO_1127 (O_1127,N_24983,N_23282);
nand UO_1128 (O_1128,N_23837,N_22543);
or UO_1129 (O_1129,N_24556,N_24047);
xnor UO_1130 (O_1130,N_23492,N_22807);
nand UO_1131 (O_1131,N_24199,N_24214);
or UO_1132 (O_1132,N_23459,N_24059);
or UO_1133 (O_1133,N_23423,N_22746);
nand UO_1134 (O_1134,N_24735,N_24146);
and UO_1135 (O_1135,N_23283,N_23516);
nand UO_1136 (O_1136,N_23260,N_22861);
or UO_1137 (O_1137,N_23112,N_24645);
or UO_1138 (O_1138,N_24260,N_23087);
or UO_1139 (O_1139,N_24977,N_23460);
nor UO_1140 (O_1140,N_23403,N_23544);
nand UO_1141 (O_1141,N_24767,N_23022);
and UO_1142 (O_1142,N_23886,N_23491);
nor UO_1143 (O_1143,N_22600,N_23006);
xor UO_1144 (O_1144,N_22580,N_23365);
and UO_1145 (O_1145,N_24369,N_23937);
and UO_1146 (O_1146,N_22897,N_24919);
and UO_1147 (O_1147,N_23312,N_23963);
or UO_1148 (O_1148,N_22948,N_24783);
xnor UO_1149 (O_1149,N_24255,N_24441);
or UO_1150 (O_1150,N_24546,N_24324);
nand UO_1151 (O_1151,N_24423,N_23373);
nor UO_1152 (O_1152,N_22608,N_22868);
xor UO_1153 (O_1153,N_23888,N_23540);
nor UO_1154 (O_1154,N_23168,N_23654);
xnor UO_1155 (O_1155,N_24672,N_24363);
nand UO_1156 (O_1156,N_23704,N_24607);
nand UO_1157 (O_1157,N_23803,N_22952);
nand UO_1158 (O_1158,N_24519,N_24563);
and UO_1159 (O_1159,N_24673,N_23719);
xor UO_1160 (O_1160,N_24346,N_23623);
and UO_1161 (O_1161,N_24914,N_22954);
xor UO_1162 (O_1162,N_23534,N_23308);
nand UO_1163 (O_1163,N_24825,N_23883);
and UO_1164 (O_1164,N_24714,N_23539);
nor UO_1165 (O_1165,N_24365,N_23256);
nand UO_1166 (O_1166,N_22947,N_23430);
or UO_1167 (O_1167,N_23561,N_23031);
and UO_1168 (O_1168,N_24722,N_23227);
or UO_1169 (O_1169,N_24999,N_24960);
or UO_1170 (O_1170,N_24421,N_22964);
xnor UO_1171 (O_1171,N_24043,N_23740);
xnor UO_1172 (O_1172,N_24163,N_24785);
or UO_1173 (O_1173,N_24675,N_24187);
xnor UO_1174 (O_1174,N_24414,N_24808);
nor UO_1175 (O_1175,N_24552,N_23393);
or UO_1176 (O_1176,N_24364,N_24023);
xnor UO_1177 (O_1177,N_23779,N_22656);
or UO_1178 (O_1178,N_23092,N_24168);
nor UO_1179 (O_1179,N_24630,N_23836);
or UO_1180 (O_1180,N_22804,N_23433);
nor UO_1181 (O_1181,N_23776,N_23134);
nor UO_1182 (O_1182,N_24777,N_23725);
xor UO_1183 (O_1183,N_24957,N_24915);
or UO_1184 (O_1184,N_22942,N_24042);
nand UO_1185 (O_1185,N_24615,N_23241);
and UO_1186 (O_1186,N_24188,N_23543);
nand UO_1187 (O_1187,N_23184,N_24413);
nor UO_1188 (O_1188,N_23278,N_24728);
xnor UO_1189 (O_1189,N_23796,N_23974);
or UO_1190 (O_1190,N_24318,N_24995);
or UO_1191 (O_1191,N_23971,N_23611);
xnor UO_1192 (O_1192,N_23840,N_24209);
nand UO_1193 (O_1193,N_24166,N_24444);
xor UO_1194 (O_1194,N_23437,N_22559);
nor UO_1195 (O_1195,N_24781,N_22590);
nand UO_1196 (O_1196,N_23469,N_24591);
nor UO_1197 (O_1197,N_24428,N_24130);
nor UO_1198 (O_1198,N_23165,N_24503);
xor UO_1199 (O_1199,N_24521,N_23246);
nor UO_1200 (O_1200,N_24358,N_24308);
nor UO_1201 (O_1201,N_22771,N_22792);
or UO_1202 (O_1202,N_24835,N_22810);
nor UO_1203 (O_1203,N_22932,N_24900);
or UO_1204 (O_1204,N_23724,N_24502);
or UO_1205 (O_1205,N_22592,N_23294);
nor UO_1206 (O_1206,N_23404,N_24740);
nor UO_1207 (O_1207,N_24626,N_23141);
or UO_1208 (O_1208,N_22538,N_23926);
nor UO_1209 (O_1209,N_23011,N_22595);
or UO_1210 (O_1210,N_22677,N_24976);
nor UO_1211 (O_1211,N_23968,N_24359);
or UO_1212 (O_1212,N_24738,N_24534);
or UO_1213 (O_1213,N_23506,N_23760);
and UO_1214 (O_1214,N_23647,N_22839);
xor UO_1215 (O_1215,N_24135,N_22638);
nor UO_1216 (O_1216,N_24656,N_24224);
nand UO_1217 (O_1217,N_22578,N_23220);
and UO_1218 (O_1218,N_24827,N_23721);
or UO_1219 (O_1219,N_23398,N_23598);
xnor UO_1220 (O_1220,N_23126,N_23801);
or UO_1221 (O_1221,N_23913,N_22813);
nand UO_1222 (O_1222,N_24171,N_23476);
xnor UO_1223 (O_1223,N_23826,N_22791);
and UO_1224 (O_1224,N_23981,N_22759);
or UO_1225 (O_1225,N_24082,N_24284);
nor UO_1226 (O_1226,N_24967,N_24653);
xnor UO_1227 (O_1227,N_22724,N_23073);
or UO_1228 (O_1228,N_22671,N_23362);
or UO_1229 (O_1229,N_24980,N_24570);
or UO_1230 (O_1230,N_22701,N_23336);
nor UO_1231 (O_1231,N_23685,N_23770);
xor UO_1232 (O_1232,N_22989,N_23651);
or UO_1233 (O_1233,N_23204,N_24902);
nand UO_1234 (O_1234,N_24074,N_23086);
nand UO_1235 (O_1235,N_23384,N_22966);
and UO_1236 (O_1236,N_24891,N_22860);
or UO_1237 (O_1237,N_23619,N_24693);
or UO_1238 (O_1238,N_22690,N_24820);
or UO_1239 (O_1239,N_23983,N_23904);
and UO_1240 (O_1240,N_24830,N_22754);
nand UO_1241 (O_1241,N_24440,N_23121);
and UO_1242 (O_1242,N_24443,N_24190);
or UO_1243 (O_1243,N_23287,N_24512);
nand UO_1244 (O_1244,N_23873,N_24567);
and UO_1245 (O_1245,N_24455,N_23289);
and UO_1246 (O_1246,N_24217,N_22761);
xor UO_1247 (O_1247,N_24466,N_24280);
xnor UO_1248 (O_1248,N_24083,N_23387);
nor UO_1249 (O_1249,N_24604,N_24347);
nand UO_1250 (O_1250,N_24287,N_23295);
and UO_1251 (O_1251,N_24440,N_24515);
nor UO_1252 (O_1252,N_24760,N_24406);
and UO_1253 (O_1253,N_22611,N_22962);
or UO_1254 (O_1254,N_23005,N_23270);
nand UO_1255 (O_1255,N_24589,N_24201);
or UO_1256 (O_1256,N_24855,N_22907);
and UO_1257 (O_1257,N_22841,N_22572);
nand UO_1258 (O_1258,N_23060,N_23897);
or UO_1259 (O_1259,N_24949,N_22881);
nand UO_1260 (O_1260,N_23923,N_24466);
nand UO_1261 (O_1261,N_23409,N_23975);
nor UO_1262 (O_1262,N_24463,N_23284);
and UO_1263 (O_1263,N_23167,N_22803);
nand UO_1264 (O_1264,N_24359,N_24200);
nor UO_1265 (O_1265,N_23579,N_23886);
nor UO_1266 (O_1266,N_24792,N_24304);
xnor UO_1267 (O_1267,N_24408,N_23665);
xor UO_1268 (O_1268,N_22749,N_23566);
xnor UO_1269 (O_1269,N_24139,N_24987);
or UO_1270 (O_1270,N_22534,N_24394);
nand UO_1271 (O_1271,N_23486,N_23824);
and UO_1272 (O_1272,N_24224,N_24688);
xnor UO_1273 (O_1273,N_24531,N_23246);
nand UO_1274 (O_1274,N_24324,N_23714);
or UO_1275 (O_1275,N_24665,N_23704);
nor UO_1276 (O_1276,N_23706,N_22985);
or UO_1277 (O_1277,N_23730,N_22620);
nor UO_1278 (O_1278,N_23370,N_24719);
xor UO_1279 (O_1279,N_22654,N_23752);
nand UO_1280 (O_1280,N_23898,N_24202);
or UO_1281 (O_1281,N_24874,N_22811);
or UO_1282 (O_1282,N_23321,N_22635);
xnor UO_1283 (O_1283,N_24985,N_24622);
nor UO_1284 (O_1284,N_24409,N_24643);
xnor UO_1285 (O_1285,N_22589,N_24863);
or UO_1286 (O_1286,N_24954,N_23598);
and UO_1287 (O_1287,N_24206,N_22854);
or UO_1288 (O_1288,N_24545,N_22602);
nor UO_1289 (O_1289,N_24197,N_23416);
nor UO_1290 (O_1290,N_23538,N_23405);
nor UO_1291 (O_1291,N_24475,N_24737);
xor UO_1292 (O_1292,N_22514,N_24742);
and UO_1293 (O_1293,N_23872,N_24132);
and UO_1294 (O_1294,N_24894,N_23310);
and UO_1295 (O_1295,N_24093,N_23129);
nor UO_1296 (O_1296,N_24519,N_22854);
nand UO_1297 (O_1297,N_24704,N_24101);
xnor UO_1298 (O_1298,N_22804,N_23910);
nor UO_1299 (O_1299,N_23979,N_24077);
nand UO_1300 (O_1300,N_23695,N_22535);
xnor UO_1301 (O_1301,N_22609,N_23453);
nand UO_1302 (O_1302,N_23138,N_22864);
nand UO_1303 (O_1303,N_23224,N_23221);
xor UO_1304 (O_1304,N_23784,N_23335);
nor UO_1305 (O_1305,N_24219,N_23079);
xor UO_1306 (O_1306,N_24015,N_23604);
nand UO_1307 (O_1307,N_22773,N_23588);
nor UO_1308 (O_1308,N_23972,N_24286);
and UO_1309 (O_1309,N_24407,N_24387);
and UO_1310 (O_1310,N_23900,N_23380);
nor UO_1311 (O_1311,N_22583,N_24931);
nor UO_1312 (O_1312,N_24743,N_22881);
or UO_1313 (O_1313,N_22714,N_24169);
nand UO_1314 (O_1314,N_23972,N_23528);
nor UO_1315 (O_1315,N_23948,N_24086);
nand UO_1316 (O_1316,N_23715,N_23639);
or UO_1317 (O_1317,N_23216,N_22665);
nor UO_1318 (O_1318,N_23664,N_23213);
and UO_1319 (O_1319,N_24031,N_24508);
xnor UO_1320 (O_1320,N_23618,N_24393);
and UO_1321 (O_1321,N_23132,N_23177);
nand UO_1322 (O_1322,N_23537,N_22756);
nand UO_1323 (O_1323,N_23886,N_23782);
or UO_1324 (O_1324,N_23610,N_23218);
nand UO_1325 (O_1325,N_23679,N_24878);
nand UO_1326 (O_1326,N_22765,N_23837);
nand UO_1327 (O_1327,N_24411,N_23787);
xnor UO_1328 (O_1328,N_22582,N_23355);
or UO_1329 (O_1329,N_23617,N_24539);
and UO_1330 (O_1330,N_23859,N_23140);
and UO_1331 (O_1331,N_22584,N_24101);
or UO_1332 (O_1332,N_23462,N_24108);
xor UO_1333 (O_1333,N_23250,N_23161);
or UO_1334 (O_1334,N_24260,N_22568);
nand UO_1335 (O_1335,N_23545,N_24703);
nand UO_1336 (O_1336,N_23808,N_24304);
nor UO_1337 (O_1337,N_23879,N_23056);
nor UO_1338 (O_1338,N_24644,N_22815);
xor UO_1339 (O_1339,N_22632,N_24497);
nand UO_1340 (O_1340,N_23758,N_23480);
and UO_1341 (O_1341,N_24135,N_24473);
nor UO_1342 (O_1342,N_24123,N_23704);
xor UO_1343 (O_1343,N_24967,N_23733);
nor UO_1344 (O_1344,N_22839,N_24040);
or UO_1345 (O_1345,N_24487,N_24702);
nand UO_1346 (O_1346,N_23921,N_23806);
nand UO_1347 (O_1347,N_24645,N_24174);
nand UO_1348 (O_1348,N_24477,N_24822);
and UO_1349 (O_1349,N_22846,N_22939);
nor UO_1350 (O_1350,N_23563,N_22877);
nor UO_1351 (O_1351,N_24682,N_24088);
or UO_1352 (O_1352,N_24979,N_24358);
and UO_1353 (O_1353,N_22892,N_24969);
or UO_1354 (O_1354,N_24432,N_24565);
nand UO_1355 (O_1355,N_23812,N_23684);
nor UO_1356 (O_1356,N_23808,N_23121);
nor UO_1357 (O_1357,N_23008,N_23989);
or UO_1358 (O_1358,N_24921,N_24407);
xor UO_1359 (O_1359,N_23957,N_24973);
nor UO_1360 (O_1360,N_23267,N_24808);
or UO_1361 (O_1361,N_24767,N_22620);
nor UO_1362 (O_1362,N_23943,N_23215);
and UO_1363 (O_1363,N_22645,N_23494);
nand UO_1364 (O_1364,N_24002,N_24926);
and UO_1365 (O_1365,N_24184,N_24503);
xnor UO_1366 (O_1366,N_23805,N_22998);
nand UO_1367 (O_1367,N_23135,N_23656);
xnor UO_1368 (O_1368,N_23335,N_22916);
nand UO_1369 (O_1369,N_24575,N_24110);
and UO_1370 (O_1370,N_23123,N_24660);
nor UO_1371 (O_1371,N_23801,N_24181);
nor UO_1372 (O_1372,N_22981,N_24752);
or UO_1373 (O_1373,N_24004,N_24649);
xor UO_1374 (O_1374,N_24304,N_23837);
nand UO_1375 (O_1375,N_22659,N_24313);
and UO_1376 (O_1376,N_23716,N_23451);
nand UO_1377 (O_1377,N_22943,N_24229);
xor UO_1378 (O_1378,N_22727,N_24207);
xor UO_1379 (O_1379,N_24504,N_23137);
or UO_1380 (O_1380,N_23059,N_24875);
xor UO_1381 (O_1381,N_24018,N_23264);
nor UO_1382 (O_1382,N_23305,N_24886);
or UO_1383 (O_1383,N_23157,N_24059);
or UO_1384 (O_1384,N_24180,N_23342);
and UO_1385 (O_1385,N_23959,N_24311);
xnor UO_1386 (O_1386,N_22989,N_24326);
or UO_1387 (O_1387,N_24450,N_24532);
nor UO_1388 (O_1388,N_24088,N_24710);
xor UO_1389 (O_1389,N_22609,N_24177);
or UO_1390 (O_1390,N_24997,N_23274);
or UO_1391 (O_1391,N_24265,N_23319);
nand UO_1392 (O_1392,N_24610,N_23967);
nand UO_1393 (O_1393,N_22606,N_23268);
or UO_1394 (O_1394,N_23312,N_24584);
xnor UO_1395 (O_1395,N_24638,N_22673);
xor UO_1396 (O_1396,N_22955,N_24131);
or UO_1397 (O_1397,N_23677,N_24758);
nand UO_1398 (O_1398,N_24124,N_23433);
nor UO_1399 (O_1399,N_23301,N_22570);
or UO_1400 (O_1400,N_24530,N_24388);
xor UO_1401 (O_1401,N_23928,N_24485);
xnor UO_1402 (O_1402,N_24725,N_22876);
or UO_1403 (O_1403,N_23673,N_23853);
and UO_1404 (O_1404,N_23106,N_24399);
nand UO_1405 (O_1405,N_24263,N_23172);
or UO_1406 (O_1406,N_23896,N_23361);
and UO_1407 (O_1407,N_23828,N_23094);
nand UO_1408 (O_1408,N_22715,N_24203);
xnor UO_1409 (O_1409,N_23860,N_22648);
or UO_1410 (O_1410,N_23151,N_23633);
xnor UO_1411 (O_1411,N_23756,N_24590);
and UO_1412 (O_1412,N_23476,N_24050);
xor UO_1413 (O_1413,N_23713,N_23024);
xor UO_1414 (O_1414,N_23281,N_24757);
or UO_1415 (O_1415,N_23300,N_23638);
nand UO_1416 (O_1416,N_24959,N_23137);
xor UO_1417 (O_1417,N_23518,N_24613);
and UO_1418 (O_1418,N_23072,N_23776);
or UO_1419 (O_1419,N_22819,N_23954);
nor UO_1420 (O_1420,N_24259,N_23618);
nor UO_1421 (O_1421,N_22645,N_23543);
nand UO_1422 (O_1422,N_23465,N_22846);
nand UO_1423 (O_1423,N_22828,N_23066);
or UO_1424 (O_1424,N_23788,N_24910);
or UO_1425 (O_1425,N_23100,N_24737);
or UO_1426 (O_1426,N_23465,N_24173);
or UO_1427 (O_1427,N_23649,N_23178);
and UO_1428 (O_1428,N_23883,N_24919);
and UO_1429 (O_1429,N_23470,N_23306);
xnor UO_1430 (O_1430,N_24210,N_22625);
or UO_1431 (O_1431,N_23509,N_24309);
and UO_1432 (O_1432,N_22965,N_24281);
and UO_1433 (O_1433,N_23113,N_22892);
or UO_1434 (O_1434,N_23303,N_24778);
nor UO_1435 (O_1435,N_24977,N_22903);
nor UO_1436 (O_1436,N_23940,N_23270);
and UO_1437 (O_1437,N_24711,N_24831);
or UO_1438 (O_1438,N_23010,N_22847);
or UO_1439 (O_1439,N_22949,N_23555);
nor UO_1440 (O_1440,N_22599,N_24391);
nand UO_1441 (O_1441,N_24502,N_23203);
nor UO_1442 (O_1442,N_23085,N_23880);
xnor UO_1443 (O_1443,N_23363,N_23788);
nor UO_1444 (O_1444,N_23431,N_24359);
xor UO_1445 (O_1445,N_24991,N_24849);
or UO_1446 (O_1446,N_23343,N_23156);
or UO_1447 (O_1447,N_23117,N_23194);
xor UO_1448 (O_1448,N_24351,N_23793);
or UO_1449 (O_1449,N_24236,N_23843);
and UO_1450 (O_1450,N_23793,N_24069);
nand UO_1451 (O_1451,N_22954,N_23692);
nand UO_1452 (O_1452,N_22977,N_23290);
nand UO_1453 (O_1453,N_23174,N_24685);
nor UO_1454 (O_1454,N_24933,N_23456);
xor UO_1455 (O_1455,N_24310,N_24136);
and UO_1456 (O_1456,N_23625,N_24073);
xnor UO_1457 (O_1457,N_23811,N_23884);
nand UO_1458 (O_1458,N_23340,N_23271);
nand UO_1459 (O_1459,N_24866,N_23643);
and UO_1460 (O_1460,N_24212,N_22523);
and UO_1461 (O_1461,N_23600,N_23123);
nand UO_1462 (O_1462,N_24043,N_22598);
or UO_1463 (O_1463,N_23937,N_22896);
nor UO_1464 (O_1464,N_24808,N_24297);
xnor UO_1465 (O_1465,N_23646,N_22766);
or UO_1466 (O_1466,N_24304,N_23492);
xor UO_1467 (O_1467,N_24352,N_23535);
xnor UO_1468 (O_1468,N_23801,N_23979);
and UO_1469 (O_1469,N_24415,N_23727);
and UO_1470 (O_1470,N_24552,N_23324);
nand UO_1471 (O_1471,N_24510,N_24292);
nand UO_1472 (O_1472,N_22923,N_23990);
nor UO_1473 (O_1473,N_24779,N_24683);
nand UO_1474 (O_1474,N_24847,N_24610);
or UO_1475 (O_1475,N_23573,N_24605);
and UO_1476 (O_1476,N_23756,N_23757);
nor UO_1477 (O_1477,N_23740,N_24031);
xnor UO_1478 (O_1478,N_23416,N_24375);
nor UO_1479 (O_1479,N_23141,N_24245);
nand UO_1480 (O_1480,N_23724,N_23195);
or UO_1481 (O_1481,N_24059,N_23172);
nor UO_1482 (O_1482,N_23988,N_24447);
and UO_1483 (O_1483,N_23158,N_24613);
nor UO_1484 (O_1484,N_24639,N_24977);
or UO_1485 (O_1485,N_24031,N_24017);
nand UO_1486 (O_1486,N_23869,N_24986);
nor UO_1487 (O_1487,N_24266,N_24340);
nor UO_1488 (O_1488,N_24298,N_23297);
or UO_1489 (O_1489,N_23098,N_22702);
nor UO_1490 (O_1490,N_23838,N_24193);
or UO_1491 (O_1491,N_24990,N_24984);
or UO_1492 (O_1492,N_23734,N_24136);
xnor UO_1493 (O_1493,N_23940,N_23315);
nor UO_1494 (O_1494,N_24234,N_23786);
nor UO_1495 (O_1495,N_24040,N_24859);
or UO_1496 (O_1496,N_23335,N_24401);
or UO_1497 (O_1497,N_22562,N_22995);
nor UO_1498 (O_1498,N_23363,N_22582);
or UO_1499 (O_1499,N_24736,N_23996);
and UO_1500 (O_1500,N_23412,N_22741);
nand UO_1501 (O_1501,N_24135,N_22685);
nor UO_1502 (O_1502,N_24384,N_24203);
nor UO_1503 (O_1503,N_24242,N_24923);
xnor UO_1504 (O_1504,N_23469,N_22555);
and UO_1505 (O_1505,N_23117,N_23346);
nor UO_1506 (O_1506,N_22637,N_23897);
xor UO_1507 (O_1507,N_24795,N_23248);
or UO_1508 (O_1508,N_23562,N_23244);
and UO_1509 (O_1509,N_22518,N_22786);
nor UO_1510 (O_1510,N_24943,N_22670);
xnor UO_1511 (O_1511,N_23320,N_23349);
xnor UO_1512 (O_1512,N_23831,N_24428);
or UO_1513 (O_1513,N_24195,N_22932);
nand UO_1514 (O_1514,N_22836,N_24121);
and UO_1515 (O_1515,N_23222,N_24910);
or UO_1516 (O_1516,N_24638,N_22804);
nand UO_1517 (O_1517,N_23188,N_24336);
nand UO_1518 (O_1518,N_24616,N_23370);
and UO_1519 (O_1519,N_23713,N_23248);
nor UO_1520 (O_1520,N_23400,N_23795);
nor UO_1521 (O_1521,N_24943,N_23690);
and UO_1522 (O_1522,N_23987,N_23507);
xnor UO_1523 (O_1523,N_23487,N_22920);
nor UO_1524 (O_1524,N_23244,N_23128);
nand UO_1525 (O_1525,N_24036,N_23757);
and UO_1526 (O_1526,N_23780,N_23473);
nand UO_1527 (O_1527,N_22635,N_23618);
xor UO_1528 (O_1528,N_24333,N_24331);
nor UO_1529 (O_1529,N_23837,N_22738);
and UO_1530 (O_1530,N_24129,N_22660);
nor UO_1531 (O_1531,N_22595,N_23661);
nand UO_1532 (O_1532,N_24783,N_23684);
or UO_1533 (O_1533,N_22720,N_23809);
nor UO_1534 (O_1534,N_24410,N_24777);
nor UO_1535 (O_1535,N_22852,N_23526);
nor UO_1536 (O_1536,N_23836,N_23056);
nand UO_1537 (O_1537,N_23018,N_24735);
and UO_1538 (O_1538,N_22848,N_22931);
nand UO_1539 (O_1539,N_23497,N_22613);
nor UO_1540 (O_1540,N_24763,N_22576);
or UO_1541 (O_1541,N_23149,N_22548);
nor UO_1542 (O_1542,N_24201,N_22609);
xnor UO_1543 (O_1543,N_22959,N_24417);
xor UO_1544 (O_1544,N_22596,N_23076);
and UO_1545 (O_1545,N_23073,N_23096);
nor UO_1546 (O_1546,N_23193,N_22675);
nor UO_1547 (O_1547,N_24049,N_23616);
or UO_1548 (O_1548,N_24428,N_23194);
xnor UO_1549 (O_1549,N_24939,N_24096);
and UO_1550 (O_1550,N_23641,N_23607);
and UO_1551 (O_1551,N_24815,N_23438);
nand UO_1552 (O_1552,N_24682,N_22645);
xor UO_1553 (O_1553,N_23212,N_24481);
nor UO_1554 (O_1554,N_24858,N_24270);
or UO_1555 (O_1555,N_23929,N_23755);
nor UO_1556 (O_1556,N_22950,N_22560);
xor UO_1557 (O_1557,N_23354,N_23873);
nor UO_1558 (O_1558,N_23981,N_24683);
and UO_1559 (O_1559,N_23455,N_24389);
nand UO_1560 (O_1560,N_24259,N_23297);
nand UO_1561 (O_1561,N_23240,N_24535);
and UO_1562 (O_1562,N_24926,N_24818);
nor UO_1563 (O_1563,N_23999,N_24459);
or UO_1564 (O_1564,N_23988,N_24270);
and UO_1565 (O_1565,N_22994,N_24587);
and UO_1566 (O_1566,N_23879,N_24666);
and UO_1567 (O_1567,N_23582,N_23410);
xnor UO_1568 (O_1568,N_23365,N_23960);
or UO_1569 (O_1569,N_24349,N_23396);
or UO_1570 (O_1570,N_23657,N_23752);
or UO_1571 (O_1571,N_23647,N_22954);
nand UO_1572 (O_1572,N_23164,N_24654);
or UO_1573 (O_1573,N_23609,N_22683);
nand UO_1574 (O_1574,N_24175,N_23324);
nand UO_1575 (O_1575,N_24025,N_22578);
nand UO_1576 (O_1576,N_24896,N_23783);
or UO_1577 (O_1577,N_24958,N_24882);
nor UO_1578 (O_1578,N_23261,N_23821);
xor UO_1579 (O_1579,N_23406,N_24144);
or UO_1580 (O_1580,N_22702,N_24434);
and UO_1581 (O_1581,N_22819,N_23562);
or UO_1582 (O_1582,N_22517,N_22773);
nand UO_1583 (O_1583,N_23961,N_22937);
xnor UO_1584 (O_1584,N_23602,N_23591);
or UO_1585 (O_1585,N_22560,N_24195);
nor UO_1586 (O_1586,N_22905,N_22878);
or UO_1587 (O_1587,N_24303,N_23655);
xnor UO_1588 (O_1588,N_22521,N_23533);
nor UO_1589 (O_1589,N_22699,N_24532);
nand UO_1590 (O_1590,N_22774,N_24217);
and UO_1591 (O_1591,N_23567,N_24546);
or UO_1592 (O_1592,N_22990,N_24145);
nor UO_1593 (O_1593,N_24117,N_24713);
and UO_1594 (O_1594,N_24321,N_22690);
nand UO_1595 (O_1595,N_23835,N_22530);
xnor UO_1596 (O_1596,N_23308,N_23504);
xor UO_1597 (O_1597,N_23984,N_24159);
or UO_1598 (O_1598,N_22881,N_23503);
nor UO_1599 (O_1599,N_23636,N_23475);
and UO_1600 (O_1600,N_24960,N_24526);
nor UO_1601 (O_1601,N_24439,N_23333);
xor UO_1602 (O_1602,N_23351,N_23226);
and UO_1603 (O_1603,N_23712,N_24080);
or UO_1604 (O_1604,N_24776,N_23547);
and UO_1605 (O_1605,N_23957,N_22956);
xnor UO_1606 (O_1606,N_24917,N_22671);
nand UO_1607 (O_1607,N_24527,N_24040);
and UO_1608 (O_1608,N_22969,N_24766);
xnor UO_1609 (O_1609,N_22866,N_22736);
or UO_1610 (O_1610,N_23185,N_24072);
xnor UO_1611 (O_1611,N_24694,N_24744);
and UO_1612 (O_1612,N_24808,N_24129);
or UO_1613 (O_1613,N_23682,N_24158);
and UO_1614 (O_1614,N_23392,N_23668);
nor UO_1615 (O_1615,N_23046,N_23317);
nand UO_1616 (O_1616,N_24548,N_24472);
nand UO_1617 (O_1617,N_24770,N_24469);
nand UO_1618 (O_1618,N_22794,N_23332);
or UO_1619 (O_1619,N_24731,N_22847);
nand UO_1620 (O_1620,N_24580,N_23579);
or UO_1621 (O_1621,N_24060,N_23839);
nand UO_1622 (O_1622,N_22814,N_23217);
or UO_1623 (O_1623,N_23444,N_23429);
and UO_1624 (O_1624,N_24078,N_23008);
xor UO_1625 (O_1625,N_24566,N_24074);
xnor UO_1626 (O_1626,N_24162,N_24109);
nor UO_1627 (O_1627,N_24961,N_24224);
nor UO_1628 (O_1628,N_23385,N_22770);
or UO_1629 (O_1629,N_24472,N_24364);
or UO_1630 (O_1630,N_24761,N_23389);
or UO_1631 (O_1631,N_23842,N_22906);
nand UO_1632 (O_1632,N_23611,N_23247);
or UO_1633 (O_1633,N_24914,N_23621);
or UO_1634 (O_1634,N_22521,N_23888);
and UO_1635 (O_1635,N_24303,N_23363);
nand UO_1636 (O_1636,N_22654,N_24723);
nor UO_1637 (O_1637,N_24726,N_24445);
xor UO_1638 (O_1638,N_22993,N_22852);
xnor UO_1639 (O_1639,N_24557,N_24439);
nand UO_1640 (O_1640,N_24292,N_23648);
nor UO_1641 (O_1641,N_22550,N_22783);
nand UO_1642 (O_1642,N_23375,N_22915);
nor UO_1643 (O_1643,N_24555,N_24435);
or UO_1644 (O_1644,N_23445,N_24326);
nor UO_1645 (O_1645,N_23916,N_22975);
nand UO_1646 (O_1646,N_24518,N_23182);
or UO_1647 (O_1647,N_22825,N_22805);
nand UO_1648 (O_1648,N_23763,N_22717);
or UO_1649 (O_1649,N_23253,N_24165);
or UO_1650 (O_1650,N_23146,N_23828);
nor UO_1651 (O_1651,N_23931,N_24504);
nand UO_1652 (O_1652,N_23045,N_24060);
nor UO_1653 (O_1653,N_23569,N_23391);
or UO_1654 (O_1654,N_23306,N_22552);
nor UO_1655 (O_1655,N_22699,N_24884);
nor UO_1656 (O_1656,N_22792,N_22822);
and UO_1657 (O_1657,N_23835,N_23651);
and UO_1658 (O_1658,N_24523,N_23549);
or UO_1659 (O_1659,N_22642,N_24341);
nand UO_1660 (O_1660,N_24076,N_23343);
or UO_1661 (O_1661,N_24736,N_23752);
and UO_1662 (O_1662,N_23697,N_22673);
and UO_1663 (O_1663,N_24755,N_24319);
xnor UO_1664 (O_1664,N_23484,N_22708);
or UO_1665 (O_1665,N_23515,N_24643);
and UO_1666 (O_1666,N_24118,N_24590);
and UO_1667 (O_1667,N_24933,N_23443);
and UO_1668 (O_1668,N_24686,N_24102);
nor UO_1669 (O_1669,N_23400,N_22898);
nand UO_1670 (O_1670,N_22522,N_23111);
nor UO_1671 (O_1671,N_23093,N_23004);
and UO_1672 (O_1672,N_23380,N_23518);
nor UO_1673 (O_1673,N_24914,N_24194);
nand UO_1674 (O_1674,N_24299,N_24048);
nand UO_1675 (O_1675,N_23047,N_24838);
nor UO_1676 (O_1676,N_23683,N_24718);
and UO_1677 (O_1677,N_23046,N_24942);
nand UO_1678 (O_1678,N_23561,N_23343);
and UO_1679 (O_1679,N_23209,N_24451);
and UO_1680 (O_1680,N_22536,N_24586);
or UO_1681 (O_1681,N_23015,N_23206);
nand UO_1682 (O_1682,N_23281,N_23315);
nand UO_1683 (O_1683,N_24160,N_24510);
xnor UO_1684 (O_1684,N_23239,N_24931);
xor UO_1685 (O_1685,N_24974,N_24119);
nor UO_1686 (O_1686,N_24960,N_22578);
or UO_1687 (O_1687,N_24474,N_24017);
and UO_1688 (O_1688,N_22872,N_22551);
and UO_1689 (O_1689,N_23532,N_24885);
xnor UO_1690 (O_1690,N_23941,N_23347);
nand UO_1691 (O_1691,N_22931,N_24698);
nor UO_1692 (O_1692,N_22775,N_23928);
xnor UO_1693 (O_1693,N_24257,N_22644);
nor UO_1694 (O_1694,N_23329,N_23161);
nor UO_1695 (O_1695,N_24813,N_23587);
xor UO_1696 (O_1696,N_22688,N_24555);
nand UO_1697 (O_1697,N_22981,N_22895);
nor UO_1698 (O_1698,N_23797,N_23512);
nand UO_1699 (O_1699,N_23881,N_22641);
xnor UO_1700 (O_1700,N_23369,N_22554);
nor UO_1701 (O_1701,N_22982,N_22648);
xor UO_1702 (O_1702,N_24779,N_24419);
xnor UO_1703 (O_1703,N_23512,N_22560);
and UO_1704 (O_1704,N_24634,N_24587);
and UO_1705 (O_1705,N_24439,N_24934);
or UO_1706 (O_1706,N_23732,N_23165);
or UO_1707 (O_1707,N_24670,N_23213);
xor UO_1708 (O_1708,N_23737,N_24398);
and UO_1709 (O_1709,N_24934,N_24346);
and UO_1710 (O_1710,N_23198,N_23930);
and UO_1711 (O_1711,N_22685,N_23271);
and UO_1712 (O_1712,N_23363,N_22874);
nand UO_1713 (O_1713,N_22540,N_24085);
nand UO_1714 (O_1714,N_22934,N_22603);
or UO_1715 (O_1715,N_23502,N_23096);
or UO_1716 (O_1716,N_22504,N_24890);
nand UO_1717 (O_1717,N_23562,N_23181);
nor UO_1718 (O_1718,N_22805,N_23249);
nand UO_1719 (O_1719,N_24164,N_23076);
xor UO_1720 (O_1720,N_22739,N_22505);
or UO_1721 (O_1721,N_23424,N_24069);
xor UO_1722 (O_1722,N_23389,N_24877);
or UO_1723 (O_1723,N_23476,N_24077);
xnor UO_1724 (O_1724,N_24498,N_22937);
xnor UO_1725 (O_1725,N_23960,N_24945);
nand UO_1726 (O_1726,N_22961,N_23244);
or UO_1727 (O_1727,N_23359,N_23374);
xor UO_1728 (O_1728,N_23005,N_23090);
nor UO_1729 (O_1729,N_23247,N_24428);
and UO_1730 (O_1730,N_23017,N_24822);
or UO_1731 (O_1731,N_22525,N_23683);
and UO_1732 (O_1732,N_24002,N_22736);
nor UO_1733 (O_1733,N_22816,N_23052);
nand UO_1734 (O_1734,N_22734,N_22737);
or UO_1735 (O_1735,N_24854,N_23609);
nor UO_1736 (O_1736,N_24523,N_22917);
and UO_1737 (O_1737,N_23437,N_24572);
nor UO_1738 (O_1738,N_22944,N_23451);
xor UO_1739 (O_1739,N_24386,N_23652);
or UO_1740 (O_1740,N_24768,N_23734);
nor UO_1741 (O_1741,N_22773,N_24534);
and UO_1742 (O_1742,N_23146,N_23840);
nor UO_1743 (O_1743,N_23256,N_22543);
and UO_1744 (O_1744,N_23276,N_24629);
xor UO_1745 (O_1745,N_24330,N_24515);
xor UO_1746 (O_1746,N_24597,N_23536);
nor UO_1747 (O_1747,N_24734,N_24903);
nor UO_1748 (O_1748,N_22557,N_24124);
xnor UO_1749 (O_1749,N_24657,N_24419);
or UO_1750 (O_1750,N_23122,N_24237);
nand UO_1751 (O_1751,N_22855,N_23960);
or UO_1752 (O_1752,N_22767,N_23428);
xnor UO_1753 (O_1753,N_23918,N_22532);
nand UO_1754 (O_1754,N_24838,N_24723);
or UO_1755 (O_1755,N_22878,N_22936);
and UO_1756 (O_1756,N_22634,N_23713);
nor UO_1757 (O_1757,N_23792,N_22852);
and UO_1758 (O_1758,N_24113,N_24495);
or UO_1759 (O_1759,N_23382,N_24891);
or UO_1760 (O_1760,N_23688,N_22613);
and UO_1761 (O_1761,N_22795,N_24938);
xnor UO_1762 (O_1762,N_22541,N_24417);
nor UO_1763 (O_1763,N_22580,N_22862);
xnor UO_1764 (O_1764,N_23950,N_22919);
nand UO_1765 (O_1765,N_24674,N_24435);
nor UO_1766 (O_1766,N_23264,N_24460);
nor UO_1767 (O_1767,N_23395,N_23503);
or UO_1768 (O_1768,N_23398,N_23563);
or UO_1769 (O_1769,N_24358,N_24465);
xor UO_1770 (O_1770,N_24260,N_24181);
and UO_1771 (O_1771,N_23729,N_22824);
nor UO_1772 (O_1772,N_24808,N_23569);
nand UO_1773 (O_1773,N_23571,N_24048);
or UO_1774 (O_1774,N_24642,N_24066);
and UO_1775 (O_1775,N_24300,N_23355);
and UO_1776 (O_1776,N_23964,N_23912);
nand UO_1777 (O_1777,N_22513,N_23569);
or UO_1778 (O_1778,N_23007,N_24697);
xor UO_1779 (O_1779,N_24614,N_24925);
xor UO_1780 (O_1780,N_24344,N_23775);
nor UO_1781 (O_1781,N_24397,N_23399);
nor UO_1782 (O_1782,N_23011,N_23522);
xnor UO_1783 (O_1783,N_22609,N_23125);
nor UO_1784 (O_1784,N_22783,N_22571);
and UO_1785 (O_1785,N_24258,N_23829);
nand UO_1786 (O_1786,N_24129,N_23239);
xor UO_1787 (O_1787,N_23507,N_22922);
or UO_1788 (O_1788,N_22563,N_22876);
xor UO_1789 (O_1789,N_22954,N_22608);
nand UO_1790 (O_1790,N_24378,N_24194);
or UO_1791 (O_1791,N_24314,N_24137);
or UO_1792 (O_1792,N_23327,N_23197);
nand UO_1793 (O_1793,N_24218,N_22527);
or UO_1794 (O_1794,N_23995,N_22671);
nand UO_1795 (O_1795,N_24623,N_22569);
xor UO_1796 (O_1796,N_24196,N_24310);
and UO_1797 (O_1797,N_23592,N_24073);
and UO_1798 (O_1798,N_22754,N_24541);
and UO_1799 (O_1799,N_24069,N_23713);
and UO_1800 (O_1800,N_24563,N_23824);
xnor UO_1801 (O_1801,N_22811,N_24719);
xor UO_1802 (O_1802,N_23913,N_22753);
or UO_1803 (O_1803,N_24376,N_24160);
or UO_1804 (O_1804,N_24195,N_22686);
and UO_1805 (O_1805,N_23780,N_23757);
and UO_1806 (O_1806,N_23565,N_22791);
xnor UO_1807 (O_1807,N_24910,N_24155);
and UO_1808 (O_1808,N_24370,N_24844);
and UO_1809 (O_1809,N_23113,N_23826);
xor UO_1810 (O_1810,N_22718,N_23240);
nor UO_1811 (O_1811,N_22920,N_23507);
nand UO_1812 (O_1812,N_23529,N_24044);
nor UO_1813 (O_1813,N_23888,N_22995);
or UO_1814 (O_1814,N_22827,N_24752);
nor UO_1815 (O_1815,N_24390,N_23676);
and UO_1816 (O_1816,N_23061,N_22931);
xnor UO_1817 (O_1817,N_24477,N_23813);
xor UO_1818 (O_1818,N_24306,N_24118);
xnor UO_1819 (O_1819,N_22753,N_23888);
or UO_1820 (O_1820,N_23147,N_24970);
nor UO_1821 (O_1821,N_24144,N_24634);
nor UO_1822 (O_1822,N_22800,N_23233);
nand UO_1823 (O_1823,N_23586,N_24515);
or UO_1824 (O_1824,N_24522,N_23612);
and UO_1825 (O_1825,N_22665,N_23812);
or UO_1826 (O_1826,N_23450,N_24246);
or UO_1827 (O_1827,N_23411,N_24921);
xnor UO_1828 (O_1828,N_23127,N_24337);
xnor UO_1829 (O_1829,N_23322,N_23708);
nand UO_1830 (O_1830,N_23263,N_24142);
or UO_1831 (O_1831,N_24852,N_23965);
nand UO_1832 (O_1832,N_24591,N_24358);
or UO_1833 (O_1833,N_24419,N_24772);
xnor UO_1834 (O_1834,N_24932,N_24601);
or UO_1835 (O_1835,N_23436,N_23468);
nor UO_1836 (O_1836,N_24086,N_24264);
and UO_1837 (O_1837,N_24496,N_23365);
or UO_1838 (O_1838,N_24307,N_23571);
xnor UO_1839 (O_1839,N_23751,N_24727);
nor UO_1840 (O_1840,N_24451,N_23029);
nor UO_1841 (O_1841,N_22872,N_23851);
nand UO_1842 (O_1842,N_24546,N_22683);
xor UO_1843 (O_1843,N_24522,N_24619);
and UO_1844 (O_1844,N_22742,N_22927);
nor UO_1845 (O_1845,N_23592,N_23244);
xnor UO_1846 (O_1846,N_24148,N_22652);
and UO_1847 (O_1847,N_23568,N_24855);
and UO_1848 (O_1848,N_24200,N_24144);
and UO_1849 (O_1849,N_24939,N_23857);
and UO_1850 (O_1850,N_22945,N_24262);
or UO_1851 (O_1851,N_23425,N_22662);
nand UO_1852 (O_1852,N_23278,N_22602);
nor UO_1853 (O_1853,N_22775,N_23873);
nand UO_1854 (O_1854,N_23208,N_24161);
nor UO_1855 (O_1855,N_23426,N_24300);
xor UO_1856 (O_1856,N_24982,N_23874);
or UO_1857 (O_1857,N_22950,N_24835);
xor UO_1858 (O_1858,N_23544,N_24921);
or UO_1859 (O_1859,N_24820,N_23792);
xnor UO_1860 (O_1860,N_24764,N_23669);
or UO_1861 (O_1861,N_24982,N_24986);
xor UO_1862 (O_1862,N_22857,N_24215);
or UO_1863 (O_1863,N_22877,N_24793);
nor UO_1864 (O_1864,N_24077,N_22917);
or UO_1865 (O_1865,N_24885,N_24791);
and UO_1866 (O_1866,N_24321,N_23935);
or UO_1867 (O_1867,N_24773,N_23851);
or UO_1868 (O_1868,N_23436,N_24467);
or UO_1869 (O_1869,N_23481,N_23008);
xor UO_1870 (O_1870,N_24395,N_22828);
nor UO_1871 (O_1871,N_24159,N_23590);
nor UO_1872 (O_1872,N_24648,N_23667);
or UO_1873 (O_1873,N_23314,N_22657);
or UO_1874 (O_1874,N_22589,N_24974);
or UO_1875 (O_1875,N_24294,N_22757);
and UO_1876 (O_1876,N_23899,N_24180);
nand UO_1877 (O_1877,N_24975,N_23241);
xnor UO_1878 (O_1878,N_24224,N_24412);
xnor UO_1879 (O_1879,N_23234,N_24165);
or UO_1880 (O_1880,N_23189,N_24404);
and UO_1881 (O_1881,N_24470,N_22598);
xnor UO_1882 (O_1882,N_23711,N_23497);
and UO_1883 (O_1883,N_23174,N_24243);
and UO_1884 (O_1884,N_23940,N_23227);
or UO_1885 (O_1885,N_22903,N_24577);
and UO_1886 (O_1886,N_22623,N_23539);
xnor UO_1887 (O_1887,N_24468,N_24984);
nand UO_1888 (O_1888,N_22709,N_23371);
nor UO_1889 (O_1889,N_22867,N_24951);
xor UO_1890 (O_1890,N_23271,N_22700);
nor UO_1891 (O_1891,N_24149,N_24972);
nor UO_1892 (O_1892,N_24966,N_24529);
nand UO_1893 (O_1893,N_22579,N_22797);
or UO_1894 (O_1894,N_23635,N_24228);
and UO_1895 (O_1895,N_23725,N_24244);
nor UO_1896 (O_1896,N_24257,N_22666);
xor UO_1897 (O_1897,N_24466,N_24099);
and UO_1898 (O_1898,N_23264,N_23355);
xor UO_1899 (O_1899,N_23057,N_24019);
and UO_1900 (O_1900,N_23658,N_24252);
xnor UO_1901 (O_1901,N_24449,N_24443);
or UO_1902 (O_1902,N_23086,N_23911);
nand UO_1903 (O_1903,N_22928,N_23829);
and UO_1904 (O_1904,N_24328,N_24620);
xor UO_1905 (O_1905,N_24882,N_23077);
nand UO_1906 (O_1906,N_24317,N_24327);
nor UO_1907 (O_1907,N_24120,N_22685);
nand UO_1908 (O_1908,N_24195,N_23656);
nor UO_1909 (O_1909,N_24698,N_23274);
and UO_1910 (O_1910,N_23913,N_24602);
nor UO_1911 (O_1911,N_24840,N_24808);
xor UO_1912 (O_1912,N_23204,N_24616);
or UO_1913 (O_1913,N_23130,N_24814);
nor UO_1914 (O_1914,N_23933,N_24896);
nand UO_1915 (O_1915,N_24428,N_23783);
xnor UO_1916 (O_1916,N_22714,N_23087);
xor UO_1917 (O_1917,N_23288,N_24914);
xor UO_1918 (O_1918,N_22640,N_24014);
or UO_1919 (O_1919,N_23736,N_23062);
xor UO_1920 (O_1920,N_22803,N_24580);
xor UO_1921 (O_1921,N_23218,N_23043);
xnor UO_1922 (O_1922,N_22594,N_24083);
or UO_1923 (O_1923,N_24875,N_24283);
or UO_1924 (O_1924,N_24034,N_24578);
nand UO_1925 (O_1925,N_22906,N_23435);
nand UO_1926 (O_1926,N_23817,N_24646);
nand UO_1927 (O_1927,N_23066,N_23496);
or UO_1928 (O_1928,N_24462,N_22669);
nor UO_1929 (O_1929,N_23566,N_23697);
and UO_1930 (O_1930,N_24489,N_24912);
xor UO_1931 (O_1931,N_23984,N_23251);
xor UO_1932 (O_1932,N_23090,N_23821);
or UO_1933 (O_1933,N_23979,N_24549);
nor UO_1934 (O_1934,N_23047,N_23316);
xnor UO_1935 (O_1935,N_23267,N_24838);
and UO_1936 (O_1936,N_24643,N_22787);
and UO_1937 (O_1937,N_23366,N_24383);
nor UO_1938 (O_1938,N_22872,N_22967);
xor UO_1939 (O_1939,N_24927,N_22865);
xnor UO_1940 (O_1940,N_24468,N_23943);
or UO_1941 (O_1941,N_22894,N_24705);
xor UO_1942 (O_1942,N_23183,N_24272);
nand UO_1943 (O_1943,N_23780,N_24802);
and UO_1944 (O_1944,N_24695,N_24161);
xor UO_1945 (O_1945,N_24320,N_24660);
or UO_1946 (O_1946,N_23492,N_22599);
xor UO_1947 (O_1947,N_22846,N_23420);
nand UO_1948 (O_1948,N_23168,N_24121);
xor UO_1949 (O_1949,N_23713,N_23069);
or UO_1950 (O_1950,N_24602,N_24217);
nand UO_1951 (O_1951,N_24819,N_24708);
or UO_1952 (O_1952,N_23310,N_24981);
xor UO_1953 (O_1953,N_23030,N_22717);
and UO_1954 (O_1954,N_23780,N_22994);
or UO_1955 (O_1955,N_22812,N_22625);
nand UO_1956 (O_1956,N_23091,N_24608);
or UO_1957 (O_1957,N_24298,N_24414);
nand UO_1958 (O_1958,N_23318,N_24359);
xnor UO_1959 (O_1959,N_23693,N_24251);
and UO_1960 (O_1960,N_24468,N_22682);
and UO_1961 (O_1961,N_23252,N_23001);
nor UO_1962 (O_1962,N_24559,N_22529);
and UO_1963 (O_1963,N_22627,N_23468);
nor UO_1964 (O_1964,N_24297,N_24997);
nand UO_1965 (O_1965,N_24139,N_24025);
and UO_1966 (O_1966,N_24624,N_22507);
xnor UO_1967 (O_1967,N_23299,N_24830);
nand UO_1968 (O_1968,N_24494,N_23799);
nor UO_1969 (O_1969,N_24548,N_24186);
nand UO_1970 (O_1970,N_24803,N_24393);
xnor UO_1971 (O_1971,N_24426,N_24627);
or UO_1972 (O_1972,N_24148,N_24333);
nor UO_1973 (O_1973,N_23039,N_23384);
and UO_1974 (O_1974,N_24503,N_23267);
nor UO_1975 (O_1975,N_23007,N_22703);
or UO_1976 (O_1976,N_23472,N_24742);
or UO_1977 (O_1977,N_24351,N_22810);
xor UO_1978 (O_1978,N_22565,N_24259);
nand UO_1979 (O_1979,N_24076,N_23512);
or UO_1980 (O_1980,N_23856,N_24880);
or UO_1981 (O_1981,N_23137,N_22956);
nor UO_1982 (O_1982,N_23769,N_24118);
nor UO_1983 (O_1983,N_24800,N_24009);
nor UO_1984 (O_1984,N_24307,N_24762);
and UO_1985 (O_1985,N_24471,N_22631);
nor UO_1986 (O_1986,N_22968,N_23637);
nand UO_1987 (O_1987,N_24196,N_24961);
nand UO_1988 (O_1988,N_24585,N_24721);
xor UO_1989 (O_1989,N_24341,N_24969);
nor UO_1990 (O_1990,N_23984,N_22632);
xor UO_1991 (O_1991,N_22561,N_23785);
or UO_1992 (O_1992,N_23331,N_24222);
and UO_1993 (O_1993,N_24185,N_23700);
nand UO_1994 (O_1994,N_22902,N_24517);
xnor UO_1995 (O_1995,N_24731,N_24269);
and UO_1996 (O_1996,N_23251,N_23743);
or UO_1997 (O_1997,N_22775,N_24139);
or UO_1998 (O_1998,N_23651,N_22864);
and UO_1999 (O_1999,N_24253,N_23651);
xnor UO_2000 (O_2000,N_24609,N_23188);
and UO_2001 (O_2001,N_23904,N_23497);
or UO_2002 (O_2002,N_24264,N_22545);
xnor UO_2003 (O_2003,N_23716,N_24081);
xnor UO_2004 (O_2004,N_24143,N_24289);
and UO_2005 (O_2005,N_22722,N_23406);
nand UO_2006 (O_2006,N_23213,N_23524);
nand UO_2007 (O_2007,N_23789,N_23614);
and UO_2008 (O_2008,N_24823,N_23515);
or UO_2009 (O_2009,N_23041,N_22661);
nand UO_2010 (O_2010,N_24998,N_22981);
and UO_2011 (O_2011,N_24075,N_23452);
and UO_2012 (O_2012,N_22505,N_24767);
xnor UO_2013 (O_2013,N_22564,N_23212);
nand UO_2014 (O_2014,N_24392,N_23570);
or UO_2015 (O_2015,N_24975,N_23892);
xor UO_2016 (O_2016,N_24583,N_22538);
or UO_2017 (O_2017,N_23441,N_22576);
xnor UO_2018 (O_2018,N_23697,N_24184);
nor UO_2019 (O_2019,N_23361,N_22985);
or UO_2020 (O_2020,N_22661,N_22595);
nor UO_2021 (O_2021,N_23161,N_24974);
xnor UO_2022 (O_2022,N_24088,N_22939);
nand UO_2023 (O_2023,N_23736,N_24949);
nand UO_2024 (O_2024,N_22713,N_24508);
nand UO_2025 (O_2025,N_23114,N_23169);
nor UO_2026 (O_2026,N_24669,N_24371);
or UO_2027 (O_2027,N_22853,N_22598);
nand UO_2028 (O_2028,N_23311,N_24318);
xor UO_2029 (O_2029,N_22721,N_23398);
and UO_2030 (O_2030,N_23620,N_23596);
or UO_2031 (O_2031,N_24237,N_23275);
xor UO_2032 (O_2032,N_23405,N_23667);
and UO_2033 (O_2033,N_24188,N_24360);
and UO_2034 (O_2034,N_23095,N_23936);
or UO_2035 (O_2035,N_22995,N_23191);
nor UO_2036 (O_2036,N_23475,N_24888);
xor UO_2037 (O_2037,N_23871,N_24836);
xor UO_2038 (O_2038,N_22970,N_23556);
xnor UO_2039 (O_2039,N_24453,N_23441);
and UO_2040 (O_2040,N_22582,N_24051);
and UO_2041 (O_2041,N_23382,N_23355);
or UO_2042 (O_2042,N_23192,N_24878);
nor UO_2043 (O_2043,N_23993,N_24272);
xor UO_2044 (O_2044,N_24424,N_22792);
nand UO_2045 (O_2045,N_23549,N_22607);
nand UO_2046 (O_2046,N_23964,N_24935);
and UO_2047 (O_2047,N_22861,N_23348);
nor UO_2048 (O_2048,N_24375,N_23314);
and UO_2049 (O_2049,N_23439,N_22764);
or UO_2050 (O_2050,N_22613,N_22950);
xnor UO_2051 (O_2051,N_24530,N_22875);
nor UO_2052 (O_2052,N_24496,N_23722);
nand UO_2053 (O_2053,N_24923,N_24415);
and UO_2054 (O_2054,N_23142,N_23655);
nand UO_2055 (O_2055,N_24089,N_23914);
or UO_2056 (O_2056,N_24501,N_22634);
nor UO_2057 (O_2057,N_24091,N_23184);
xor UO_2058 (O_2058,N_22667,N_24633);
or UO_2059 (O_2059,N_24402,N_23282);
nor UO_2060 (O_2060,N_22888,N_24840);
nand UO_2061 (O_2061,N_22786,N_24621);
xnor UO_2062 (O_2062,N_23226,N_24002);
nor UO_2063 (O_2063,N_22531,N_24378);
xor UO_2064 (O_2064,N_22925,N_22951);
or UO_2065 (O_2065,N_23246,N_22942);
nand UO_2066 (O_2066,N_24395,N_24760);
and UO_2067 (O_2067,N_22705,N_24453);
nor UO_2068 (O_2068,N_23395,N_22942);
nor UO_2069 (O_2069,N_23531,N_24804);
and UO_2070 (O_2070,N_23061,N_23032);
nand UO_2071 (O_2071,N_24030,N_24742);
and UO_2072 (O_2072,N_24730,N_24433);
nand UO_2073 (O_2073,N_22639,N_24254);
nand UO_2074 (O_2074,N_24432,N_23962);
and UO_2075 (O_2075,N_22848,N_24683);
xor UO_2076 (O_2076,N_24902,N_24762);
nor UO_2077 (O_2077,N_24720,N_23732);
and UO_2078 (O_2078,N_24865,N_23611);
nor UO_2079 (O_2079,N_23438,N_24279);
nand UO_2080 (O_2080,N_24324,N_23754);
xnor UO_2081 (O_2081,N_22586,N_24413);
xor UO_2082 (O_2082,N_24698,N_24916);
xnor UO_2083 (O_2083,N_23359,N_24972);
and UO_2084 (O_2084,N_23142,N_23448);
xnor UO_2085 (O_2085,N_23357,N_22788);
nor UO_2086 (O_2086,N_22677,N_22798);
xnor UO_2087 (O_2087,N_24963,N_24381);
and UO_2088 (O_2088,N_22845,N_24737);
nand UO_2089 (O_2089,N_24184,N_24407);
nand UO_2090 (O_2090,N_22749,N_22754);
or UO_2091 (O_2091,N_24116,N_22654);
nand UO_2092 (O_2092,N_23930,N_24144);
or UO_2093 (O_2093,N_22622,N_23379);
nand UO_2094 (O_2094,N_23779,N_24802);
nor UO_2095 (O_2095,N_24225,N_24631);
xnor UO_2096 (O_2096,N_24626,N_24229);
xnor UO_2097 (O_2097,N_23150,N_23336);
nor UO_2098 (O_2098,N_24385,N_23731);
and UO_2099 (O_2099,N_23392,N_23169);
nor UO_2100 (O_2100,N_24282,N_22824);
or UO_2101 (O_2101,N_24892,N_23119);
xnor UO_2102 (O_2102,N_24894,N_24680);
xnor UO_2103 (O_2103,N_23032,N_24686);
or UO_2104 (O_2104,N_24145,N_23333);
or UO_2105 (O_2105,N_22850,N_22994);
nor UO_2106 (O_2106,N_24543,N_23715);
nor UO_2107 (O_2107,N_24118,N_22762);
nand UO_2108 (O_2108,N_23041,N_24509);
xnor UO_2109 (O_2109,N_22867,N_24725);
and UO_2110 (O_2110,N_22857,N_24820);
or UO_2111 (O_2111,N_22669,N_23985);
or UO_2112 (O_2112,N_24350,N_22573);
and UO_2113 (O_2113,N_22613,N_24668);
nand UO_2114 (O_2114,N_23246,N_23153);
xor UO_2115 (O_2115,N_22736,N_23009);
nor UO_2116 (O_2116,N_23099,N_23986);
nand UO_2117 (O_2117,N_23270,N_22528);
or UO_2118 (O_2118,N_24417,N_23946);
and UO_2119 (O_2119,N_22735,N_24470);
nand UO_2120 (O_2120,N_24315,N_24254);
xor UO_2121 (O_2121,N_23101,N_24289);
and UO_2122 (O_2122,N_22594,N_23160);
xor UO_2123 (O_2123,N_24380,N_24383);
and UO_2124 (O_2124,N_22529,N_23233);
and UO_2125 (O_2125,N_23330,N_23550);
xnor UO_2126 (O_2126,N_24450,N_22898);
and UO_2127 (O_2127,N_23261,N_24674);
or UO_2128 (O_2128,N_23840,N_24365);
nor UO_2129 (O_2129,N_22663,N_22542);
nor UO_2130 (O_2130,N_24809,N_24617);
nor UO_2131 (O_2131,N_24840,N_24076);
nor UO_2132 (O_2132,N_24496,N_22920);
nand UO_2133 (O_2133,N_24429,N_22682);
nand UO_2134 (O_2134,N_23664,N_24760);
or UO_2135 (O_2135,N_22779,N_23636);
or UO_2136 (O_2136,N_23014,N_22810);
or UO_2137 (O_2137,N_23790,N_23443);
nor UO_2138 (O_2138,N_22545,N_24091);
nor UO_2139 (O_2139,N_24942,N_24556);
or UO_2140 (O_2140,N_23930,N_22790);
nor UO_2141 (O_2141,N_24176,N_22845);
or UO_2142 (O_2142,N_24634,N_22589);
nor UO_2143 (O_2143,N_24355,N_24994);
nand UO_2144 (O_2144,N_23927,N_23278);
and UO_2145 (O_2145,N_23826,N_23551);
and UO_2146 (O_2146,N_24331,N_23455);
and UO_2147 (O_2147,N_23837,N_23414);
or UO_2148 (O_2148,N_24815,N_22990);
or UO_2149 (O_2149,N_23834,N_22655);
nor UO_2150 (O_2150,N_23651,N_24278);
and UO_2151 (O_2151,N_22975,N_23593);
nor UO_2152 (O_2152,N_23415,N_24701);
nand UO_2153 (O_2153,N_24970,N_22895);
nand UO_2154 (O_2154,N_23248,N_24127);
and UO_2155 (O_2155,N_22870,N_24897);
nor UO_2156 (O_2156,N_23169,N_24198);
or UO_2157 (O_2157,N_24794,N_24230);
and UO_2158 (O_2158,N_22769,N_24674);
xnor UO_2159 (O_2159,N_24504,N_22630);
nor UO_2160 (O_2160,N_23776,N_24045);
nand UO_2161 (O_2161,N_24420,N_22836);
or UO_2162 (O_2162,N_24635,N_24881);
xnor UO_2163 (O_2163,N_24771,N_24017);
or UO_2164 (O_2164,N_24514,N_23241);
or UO_2165 (O_2165,N_22975,N_23666);
and UO_2166 (O_2166,N_24325,N_24319);
or UO_2167 (O_2167,N_24664,N_24409);
nand UO_2168 (O_2168,N_24260,N_23391);
xor UO_2169 (O_2169,N_24542,N_24220);
nand UO_2170 (O_2170,N_23751,N_23197);
nor UO_2171 (O_2171,N_23158,N_24933);
nand UO_2172 (O_2172,N_23924,N_24905);
and UO_2173 (O_2173,N_23204,N_23833);
nand UO_2174 (O_2174,N_24842,N_24905);
nand UO_2175 (O_2175,N_24677,N_24791);
nor UO_2176 (O_2176,N_24075,N_23407);
and UO_2177 (O_2177,N_23822,N_23962);
and UO_2178 (O_2178,N_24619,N_24066);
nand UO_2179 (O_2179,N_24276,N_22979);
nor UO_2180 (O_2180,N_23979,N_22739);
and UO_2181 (O_2181,N_24338,N_22777);
xnor UO_2182 (O_2182,N_24795,N_23251);
xnor UO_2183 (O_2183,N_24094,N_23293);
nand UO_2184 (O_2184,N_24908,N_24054);
nand UO_2185 (O_2185,N_24612,N_23329);
nor UO_2186 (O_2186,N_23733,N_22685);
and UO_2187 (O_2187,N_23391,N_23411);
nor UO_2188 (O_2188,N_22722,N_24780);
and UO_2189 (O_2189,N_23030,N_24176);
nor UO_2190 (O_2190,N_24424,N_24156);
and UO_2191 (O_2191,N_24074,N_23440);
nand UO_2192 (O_2192,N_24197,N_22561);
nand UO_2193 (O_2193,N_24064,N_23382);
nor UO_2194 (O_2194,N_23862,N_22554);
xnor UO_2195 (O_2195,N_23649,N_24842);
and UO_2196 (O_2196,N_24469,N_22518);
nor UO_2197 (O_2197,N_23702,N_23869);
xor UO_2198 (O_2198,N_23279,N_24278);
nor UO_2199 (O_2199,N_24936,N_23527);
and UO_2200 (O_2200,N_23470,N_23632);
nor UO_2201 (O_2201,N_23603,N_22576);
xor UO_2202 (O_2202,N_24395,N_24021);
and UO_2203 (O_2203,N_24146,N_23121);
nor UO_2204 (O_2204,N_23300,N_22998);
xor UO_2205 (O_2205,N_23918,N_24335);
or UO_2206 (O_2206,N_24794,N_23766);
xor UO_2207 (O_2207,N_22919,N_23612);
nand UO_2208 (O_2208,N_23302,N_23050);
nor UO_2209 (O_2209,N_23797,N_24076);
and UO_2210 (O_2210,N_22527,N_23074);
nor UO_2211 (O_2211,N_24060,N_23888);
and UO_2212 (O_2212,N_22925,N_24589);
nor UO_2213 (O_2213,N_23858,N_23939);
xnor UO_2214 (O_2214,N_24231,N_23539);
nor UO_2215 (O_2215,N_24589,N_23675);
nor UO_2216 (O_2216,N_23692,N_24430);
xor UO_2217 (O_2217,N_22576,N_22686);
and UO_2218 (O_2218,N_22870,N_23381);
and UO_2219 (O_2219,N_24826,N_24106);
nor UO_2220 (O_2220,N_23584,N_24055);
and UO_2221 (O_2221,N_24676,N_23738);
nand UO_2222 (O_2222,N_24008,N_22530);
nor UO_2223 (O_2223,N_23186,N_23461);
nand UO_2224 (O_2224,N_24528,N_23725);
xnor UO_2225 (O_2225,N_24526,N_23744);
nor UO_2226 (O_2226,N_22978,N_23364);
nand UO_2227 (O_2227,N_22840,N_23973);
nand UO_2228 (O_2228,N_23520,N_24165);
or UO_2229 (O_2229,N_24599,N_23162);
or UO_2230 (O_2230,N_24441,N_24522);
or UO_2231 (O_2231,N_22811,N_23526);
and UO_2232 (O_2232,N_24285,N_23587);
or UO_2233 (O_2233,N_23806,N_23825);
or UO_2234 (O_2234,N_24480,N_23062);
and UO_2235 (O_2235,N_24447,N_23310);
or UO_2236 (O_2236,N_24670,N_23565);
nor UO_2237 (O_2237,N_23717,N_23716);
and UO_2238 (O_2238,N_23521,N_24140);
and UO_2239 (O_2239,N_24627,N_23581);
or UO_2240 (O_2240,N_22861,N_22536);
or UO_2241 (O_2241,N_24186,N_22724);
nand UO_2242 (O_2242,N_22768,N_23011);
xnor UO_2243 (O_2243,N_24445,N_22766);
xor UO_2244 (O_2244,N_24429,N_23274);
nor UO_2245 (O_2245,N_23441,N_22877);
nor UO_2246 (O_2246,N_22774,N_23961);
or UO_2247 (O_2247,N_24044,N_24026);
and UO_2248 (O_2248,N_24849,N_24788);
nand UO_2249 (O_2249,N_22660,N_22602);
xnor UO_2250 (O_2250,N_22800,N_23741);
xor UO_2251 (O_2251,N_24910,N_24472);
xor UO_2252 (O_2252,N_24424,N_23035);
nor UO_2253 (O_2253,N_22707,N_24578);
and UO_2254 (O_2254,N_24841,N_24577);
nor UO_2255 (O_2255,N_22511,N_24243);
xor UO_2256 (O_2256,N_24066,N_22977);
or UO_2257 (O_2257,N_23094,N_23235);
nor UO_2258 (O_2258,N_23598,N_24569);
nand UO_2259 (O_2259,N_23451,N_23934);
and UO_2260 (O_2260,N_23949,N_23913);
and UO_2261 (O_2261,N_23090,N_23485);
and UO_2262 (O_2262,N_24429,N_23424);
nor UO_2263 (O_2263,N_23080,N_23677);
or UO_2264 (O_2264,N_22708,N_24361);
nand UO_2265 (O_2265,N_23254,N_24616);
xnor UO_2266 (O_2266,N_22952,N_24350);
and UO_2267 (O_2267,N_24649,N_24574);
nand UO_2268 (O_2268,N_23170,N_23709);
nor UO_2269 (O_2269,N_23383,N_24962);
nand UO_2270 (O_2270,N_23117,N_23210);
or UO_2271 (O_2271,N_23553,N_23367);
nor UO_2272 (O_2272,N_24121,N_23244);
or UO_2273 (O_2273,N_22959,N_24099);
nor UO_2274 (O_2274,N_23062,N_23549);
or UO_2275 (O_2275,N_22562,N_22797);
nand UO_2276 (O_2276,N_24838,N_23309);
or UO_2277 (O_2277,N_23244,N_23905);
nor UO_2278 (O_2278,N_23489,N_22822);
xnor UO_2279 (O_2279,N_22943,N_23265);
nand UO_2280 (O_2280,N_24294,N_24110);
or UO_2281 (O_2281,N_23389,N_23392);
and UO_2282 (O_2282,N_22612,N_23033);
nand UO_2283 (O_2283,N_23797,N_23673);
nor UO_2284 (O_2284,N_22668,N_22699);
nor UO_2285 (O_2285,N_22799,N_23384);
nand UO_2286 (O_2286,N_22847,N_23699);
xor UO_2287 (O_2287,N_24776,N_23727);
and UO_2288 (O_2288,N_23945,N_24259);
nand UO_2289 (O_2289,N_23118,N_23902);
xor UO_2290 (O_2290,N_23182,N_22927);
nand UO_2291 (O_2291,N_23100,N_24405);
nor UO_2292 (O_2292,N_23453,N_22656);
nand UO_2293 (O_2293,N_23260,N_24745);
nand UO_2294 (O_2294,N_23145,N_22797);
or UO_2295 (O_2295,N_23376,N_24633);
xnor UO_2296 (O_2296,N_23867,N_24617);
and UO_2297 (O_2297,N_24994,N_24864);
nand UO_2298 (O_2298,N_24543,N_24440);
or UO_2299 (O_2299,N_23608,N_23448);
xor UO_2300 (O_2300,N_23465,N_23420);
nand UO_2301 (O_2301,N_24118,N_23295);
nor UO_2302 (O_2302,N_24524,N_24257);
or UO_2303 (O_2303,N_24727,N_24643);
or UO_2304 (O_2304,N_22871,N_24028);
nor UO_2305 (O_2305,N_24564,N_24402);
nand UO_2306 (O_2306,N_22735,N_22878);
nand UO_2307 (O_2307,N_22552,N_24436);
or UO_2308 (O_2308,N_23659,N_24788);
or UO_2309 (O_2309,N_23474,N_23865);
or UO_2310 (O_2310,N_24920,N_22708);
nand UO_2311 (O_2311,N_23040,N_24441);
xor UO_2312 (O_2312,N_22572,N_23906);
and UO_2313 (O_2313,N_22993,N_22698);
nor UO_2314 (O_2314,N_23663,N_23063);
nand UO_2315 (O_2315,N_23343,N_22903);
or UO_2316 (O_2316,N_23922,N_23608);
nand UO_2317 (O_2317,N_22584,N_24881);
nor UO_2318 (O_2318,N_24517,N_24042);
and UO_2319 (O_2319,N_22990,N_23046);
nand UO_2320 (O_2320,N_24356,N_22703);
and UO_2321 (O_2321,N_22654,N_23018);
nor UO_2322 (O_2322,N_23041,N_23708);
nor UO_2323 (O_2323,N_24123,N_22629);
nor UO_2324 (O_2324,N_22507,N_24646);
nand UO_2325 (O_2325,N_23453,N_22643);
nor UO_2326 (O_2326,N_22692,N_24617);
xnor UO_2327 (O_2327,N_24317,N_23129);
nor UO_2328 (O_2328,N_23684,N_22981);
nor UO_2329 (O_2329,N_24361,N_22994);
nand UO_2330 (O_2330,N_23229,N_22528);
xor UO_2331 (O_2331,N_24206,N_24072);
xnor UO_2332 (O_2332,N_23092,N_23242);
nand UO_2333 (O_2333,N_23800,N_24647);
nand UO_2334 (O_2334,N_24818,N_23802);
and UO_2335 (O_2335,N_22747,N_24675);
and UO_2336 (O_2336,N_24930,N_23333);
nand UO_2337 (O_2337,N_23908,N_24677);
and UO_2338 (O_2338,N_24772,N_23157);
and UO_2339 (O_2339,N_23017,N_23952);
nor UO_2340 (O_2340,N_24560,N_24657);
and UO_2341 (O_2341,N_24472,N_23051);
nand UO_2342 (O_2342,N_23949,N_23009);
nand UO_2343 (O_2343,N_23218,N_24292);
nand UO_2344 (O_2344,N_23930,N_24063);
xnor UO_2345 (O_2345,N_22751,N_24432);
or UO_2346 (O_2346,N_24563,N_23692);
and UO_2347 (O_2347,N_23753,N_23727);
xor UO_2348 (O_2348,N_22829,N_22686);
nor UO_2349 (O_2349,N_23432,N_23676);
nor UO_2350 (O_2350,N_22782,N_24770);
nand UO_2351 (O_2351,N_24930,N_22783);
xnor UO_2352 (O_2352,N_22858,N_22753);
or UO_2353 (O_2353,N_23204,N_23437);
and UO_2354 (O_2354,N_22639,N_22540);
and UO_2355 (O_2355,N_24670,N_24253);
and UO_2356 (O_2356,N_24105,N_24449);
nand UO_2357 (O_2357,N_22592,N_23394);
nor UO_2358 (O_2358,N_24558,N_22565);
and UO_2359 (O_2359,N_24938,N_24467);
xnor UO_2360 (O_2360,N_23726,N_23366);
nor UO_2361 (O_2361,N_23707,N_24920);
nor UO_2362 (O_2362,N_24497,N_24265);
or UO_2363 (O_2363,N_24816,N_24163);
xnor UO_2364 (O_2364,N_24999,N_23948);
nor UO_2365 (O_2365,N_22727,N_23934);
nand UO_2366 (O_2366,N_22573,N_23571);
xnor UO_2367 (O_2367,N_23279,N_24332);
xnor UO_2368 (O_2368,N_23319,N_22819);
or UO_2369 (O_2369,N_23956,N_23523);
or UO_2370 (O_2370,N_24730,N_22920);
nand UO_2371 (O_2371,N_24224,N_24953);
and UO_2372 (O_2372,N_22917,N_23056);
xnor UO_2373 (O_2373,N_24747,N_23440);
xnor UO_2374 (O_2374,N_23167,N_24598);
and UO_2375 (O_2375,N_24547,N_24532);
nor UO_2376 (O_2376,N_24879,N_24137);
nand UO_2377 (O_2377,N_22565,N_24116);
xnor UO_2378 (O_2378,N_24443,N_24400);
or UO_2379 (O_2379,N_24805,N_24556);
or UO_2380 (O_2380,N_23084,N_24889);
or UO_2381 (O_2381,N_22746,N_23392);
or UO_2382 (O_2382,N_23616,N_23430);
or UO_2383 (O_2383,N_22688,N_24362);
nand UO_2384 (O_2384,N_24123,N_24626);
and UO_2385 (O_2385,N_22534,N_24937);
nor UO_2386 (O_2386,N_23245,N_23112);
or UO_2387 (O_2387,N_24211,N_24888);
or UO_2388 (O_2388,N_23403,N_23473);
or UO_2389 (O_2389,N_24822,N_24679);
nor UO_2390 (O_2390,N_24482,N_22951);
and UO_2391 (O_2391,N_23610,N_22835);
and UO_2392 (O_2392,N_24009,N_23103);
and UO_2393 (O_2393,N_22847,N_23368);
or UO_2394 (O_2394,N_24201,N_24051);
nand UO_2395 (O_2395,N_23055,N_23410);
or UO_2396 (O_2396,N_22566,N_23373);
or UO_2397 (O_2397,N_23580,N_22508);
xnor UO_2398 (O_2398,N_24994,N_23354);
and UO_2399 (O_2399,N_23197,N_24526);
nand UO_2400 (O_2400,N_23109,N_24147);
xnor UO_2401 (O_2401,N_23980,N_23383);
nand UO_2402 (O_2402,N_24769,N_24029);
nor UO_2403 (O_2403,N_24131,N_24397);
or UO_2404 (O_2404,N_24987,N_24283);
nand UO_2405 (O_2405,N_24237,N_24323);
and UO_2406 (O_2406,N_23476,N_24296);
nand UO_2407 (O_2407,N_23506,N_23975);
nand UO_2408 (O_2408,N_24632,N_24978);
nor UO_2409 (O_2409,N_23541,N_22696);
xnor UO_2410 (O_2410,N_24190,N_23460);
or UO_2411 (O_2411,N_23986,N_22625);
xor UO_2412 (O_2412,N_22530,N_24639);
and UO_2413 (O_2413,N_23786,N_22612);
nand UO_2414 (O_2414,N_24939,N_23323);
or UO_2415 (O_2415,N_23688,N_23220);
or UO_2416 (O_2416,N_24315,N_24581);
xnor UO_2417 (O_2417,N_24254,N_23014);
xor UO_2418 (O_2418,N_23111,N_23163);
or UO_2419 (O_2419,N_23222,N_24156);
and UO_2420 (O_2420,N_22550,N_24126);
and UO_2421 (O_2421,N_23684,N_24889);
nor UO_2422 (O_2422,N_24501,N_24675);
and UO_2423 (O_2423,N_23664,N_24218);
nor UO_2424 (O_2424,N_24267,N_22873);
xor UO_2425 (O_2425,N_23150,N_22683);
xor UO_2426 (O_2426,N_23337,N_23583);
xor UO_2427 (O_2427,N_23081,N_24439);
xor UO_2428 (O_2428,N_23599,N_24671);
or UO_2429 (O_2429,N_23414,N_23768);
nand UO_2430 (O_2430,N_24320,N_22832);
or UO_2431 (O_2431,N_24712,N_22933);
nor UO_2432 (O_2432,N_22547,N_24162);
xnor UO_2433 (O_2433,N_24630,N_24368);
xnor UO_2434 (O_2434,N_24313,N_23666);
xnor UO_2435 (O_2435,N_24675,N_23861);
nand UO_2436 (O_2436,N_23699,N_22929);
nand UO_2437 (O_2437,N_24045,N_24641);
and UO_2438 (O_2438,N_23276,N_22620);
nand UO_2439 (O_2439,N_23051,N_23294);
xor UO_2440 (O_2440,N_23202,N_22870);
xor UO_2441 (O_2441,N_24056,N_22946);
or UO_2442 (O_2442,N_23051,N_24238);
and UO_2443 (O_2443,N_23846,N_24682);
xor UO_2444 (O_2444,N_24631,N_24726);
xnor UO_2445 (O_2445,N_22961,N_22729);
or UO_2446 (O_2446,N_23590,N_24506);
xnor UO_2447 (O_2447,N_23261,N_24986);
nand UO_2448 (O_2448,N_24096,N_24570);
or UO_2449 (O_2449,N_24845,N_22993);
and UO_2450 (O_2450,N_24643,N_23243);
or UO_2451 (O_2451,N_24926,N_23697);
nand UO_2452 (O_2452,N_23090,N_23648);
nor UO_2453 (O_2453,N_24507,N_24304);
xnor UO_2454 (O_2454,N_23008,N_22727);
and UO_2455 (O_2455,N_24136,N_22631);
or UO_2456 (O_2456,N_24286,N_22604);
or UO_2457 (O_2457,N_24259,N_24816);
nor UO_2458 (O_2458,N_23403,N_22725);
nand UO_2459 (O_2459,N_24794,N_24117);
or UO_2460 (O_2460,N_23960,N_23581);
nor UO_2461 (O_2461,N_23058,N_24012);
or UO_2462 (O_2462,N_23468,N_24192);
xnor UO_2463 (O_2463,N_24905,N_22809);
xnor UO_2464 (O_2464,N_24525,N_22505);
xor UO_2465 (O_2465,N_22639,N_24493);
nand UO_2466 (O_2466,N_23369,N_23020);
xnor UO_2467 (O_2467,N_24757,N_23163);
xnor UO_2468 (O_2468,N_24116,N_24865);
or UO_2469 (O_2469,N_23934,N_24977);
xor UO_2470 (O_2470,N_22678,N_22604);
nor UO_2471 (O_2471,N_23200,N_23536);
nand UO_2472 (O_2472,N_24047,N_24169);
nand UO_2473 (O_2473,N_24978,N_24271);
nor UO_2474 (O_2474,N_24335,N_22911);
nor UO_2475 (O_2475,N_23232,N_23781);
or UO_2476 (O_2476,N_24724,N_24498);
and UO_2477 (O_2477,N_22670,N_24262);
and UO_2478 (O_2478,N_22551,N_24646);
xnor UO_2479 (O_2479,N_22984,N_22702);
nor UO_2480 (O_2480,N_24170,N_23584);
nand UO_2481 (O_2481,N_24456,N_24505);
nor UO_2482 (O_2482,N_22630,N_23256);
and UO_2483 (O_2483,N_23370,N_22612);
and UO_2484 (O_2484,N_23109,N_23460);
nor UO_2485 (O_2485,N_22615,N_24462);
nor UO_2486 (O_2486,N_24648,N_23600);
xnor UO_2487 (O_2487,N_24055,N_23806);
nor UO_2488 (O_2488,N_24854,N_24469);
nand UO_2489 (O_2489,N_23522,N_24121);
or UO_2490 (O_2490,N_24202,N_24587);
nand UO_2491 (O_2491,N_23605,N_24326);
nand UO_2492 (O_2492,N_23960,N_24288);
and UO_2493 (O_2493,N_22864,N_23155);
nand UO_2494 (O_2494,N_23818,N_23520);
nor UO_2495 (O_2495,N_24338,N_23594);
or UO_2496 (O_2496,N_24234,N_23484);
or UO_2497 (O_2497,N_24512,N_23708);
nand UO_2498 (O_2498,N_22803,N_23964);
xnor UO_2499 (O_2499,N_24394,N_22635);
nand UO_2500 (O_2500,N_23290,N_24164);
nand UO_2501 (O_2501,N_24437,N_23954);
nor UO_2502 (O_2502,N_22708,N_24317);
or UO_2503 (O_2503,N_24283,N_23122);
nand UO_2504 (O_2504,N_24025,N_22514);
nor UO_2505 (O_2505,N_23127,N_23730);
nand UO_2506 (O_2506,N_24718,N_24058);
and UO_2507 (O_2507,N_23350,N_22577);
or UO_2508 (O_2508,N_22707,N_22772);
and UO_2509 (O_2509,N_23932,N_23386);
nand UO_2510 (O_2510,N_22709,N_23370);
nor UO_2511 (O_2511,N_24811,N_24644);
or UO_2512 (O_2512,N_23110,N_22508);
nor UO_2513 (O_2513,N_22707,N_23876);
and UO_2514 (O_2514,N_24182,N_24976);
xor UO_2515 (O_2515,N_23957,N_23691);
and UO_2516 (O_2516,N_22651,N_23852);
xnor UO_2517 (O_2517,N_23549,N_22751);
and UO_2518 (O_2518,N_23744,N_23063);
and UO_2519 (O_2519,N_23021,N_24551);
nor UO_2520 (O_2520,N_24105,N_23454);
nand UO_2521 (O_2521,N_22849,N_23909);
and UO_2522 (O_2522,N_23100,N_23399);
nand UO_2523 (O_2523,N_23614,N_24787);
or UO_2524 (O_2524,N_23884,N_23928);
or UO_2525 (O_2525,N_23384,N_23179);
nand UO_2526 (O_2526,N_23348,N_24185);
nor UO_2527 (O_2527,N_22512,N_23134);
and UO_2528 (O_2528,N_23482,N_23888);
nand UO_2529 (O_2529,N_24238,N_23329);
or UO_2530 (O_2530,N_22978,N_24318);
nor UO_2531 (O_2531,N_22989,N_24385);
or UO_2532 (O_2532,N_24864,N_22839);
xor UO_2533 (O_2533,N_23036,N_24475);
nor UO_2534 (O_2534,N_22623,N_23886);
or UO_2535 (O_2535,N_23420,N_24281);
nor UO_2536 (O_2536,N_24854,N_23546);
or UO_2537 (O_2537,N_24955,N_23347);
xnor UO_2538 (O_2538,N_22894,N_23328);
nor UO_2539 (O_2539,N_23879,N_23081);
or UO_2540 (O_2540,N_23269,N_24223);
and UO_2541 (O_2541,N_24053,N_22757);
or UO_2542 (O_2542,N_23146,N_24891);
nor UO_2543 (O_2543,N_24544,N_23773);
or UO_2544 (O_2544,N_24518,N_23017);
nand UO_2545 (O_2545,N_24891,N_23438);
or UO_2546 (O_2546,N_22613,N_24924);
or UO_2547 (O_2547,N_22924,N_22829);
and UO_2548 (O_2548,N_22703,N_23875);
nand UO_2549 (O_2549,N_24370,N_23174);
or UO_2550 (O_2550,N_24454,N_23899);
or UO_2551 (O_2551,N_22996,N_24656);
and UO_2552 (O_2552,N_24544,N_24208);
nand UO_2553 (O_2553,N_24837,N_24635);
or UO_2554 (O_2554,N_23648,N_24339);
or UO_2555 (O_2555,N_24128,N_23797);
nand UO_2556 (O_2556,N_22609,N_24639);
nor UO_2557 (O_2557,N_23158,N_22646);
nand UO_2558 (O_2558,N_24168,N_24418);
nand UO_2559 (O_2559,N_22507,N_24818);
nor UO_2560 (O_2560,N_22644,N_22859);
nor UO_2561 (O_2561,N_23460,N_23363);
nand UO_2562 (O_2562,N_23509,N_22783);
xor UO_2563 (O_2563,N_24457,N_24911);
nand UO_2564 (O_2564,N_24349,N_24490);
xnor UO_2565 (O_2565,N_24480,N_22917);
nor UO_2566 (O_2566,N_24083,N_24684);
and UO_2567 (O_2567,N_24800,N_24237);
xnor UO_2568 (O_2568,N_24985,N_22719);
nand UO_2569 (O_2569,N_23083,N_24087);
and UO_2570 (O_2570,N_23119,N_23573);
and UO_2571 (O_2571,N_23942,N_23825);
nor UO_2572 (O_2572,N_24878,N_22540);
or UO_2573 (O_2573,N_24460,N_23631);
and UO_2574 (O_2574,N_23817,N_23548);
and UO_2575 (O_2575,N_22662,N_24129);
xnor UO_2576 (O_2576,N_23798,N_23473);
nor UO_2577 (O_2577,N_23542,N_24589);
or UO_2578 (O_2578,N_24385,N_23569);
or UO_2579 (O_2579,N_23442,N_23834);
xor UO_2580 (O_2580,N_23518,N_23623);
or UO_2581 (O_2581,N_23679,N_23073);
xor UO_2582 (O_2582,N_24137,N_24646);
or UO_2583 (O_2583,N_24329,N_22676);
or UO_2584 (O_2584,N_23834,N_23895);
nand UO_2585 (O_2585,N_23197,N_24423);
and UO_2586 (O_2586,N_23325,N_24907);
or UO_2587 (O_2587,N_23523,N_24143);
nor UO_2588 (O_2588,N_22817,N_22694);
xnor UO_2589 (O_2589,N_24239,N_23618);
nand UO_2590 (O_2590,N_23138,N_24438);
nand UO_2591 (O_2591,N_22609,N_24088);
xor UO_2592 (O_2592,N_23480,N_24401);
or UO_2593 (O_2593,N_22834,N_24268);
and UO_2594 (O_2594,N_23447,N_24822);
nor UO_2595 (O_2595,N_24319,N_23110);
or UO_2596 (O_2596,N_22748,N_23878);
xnor UO_2597 (O_2597,N_24447,N_24067);
or UO_2598 (O_2598,N_24068,N_24462);
or UO_2599 (O_2599,N_23105,N_24906);
nand UO_2600 (O_2600,N_23602,N_22709);
nor UO_2601 (O_2601,N_23916,N_22565);
nand UO_2602 (O_2602,N_22608,N_24758);
nand UO_2603 (O_2603,N_23822,N_24024);
and UO_2604 (O_2604,N_23769,N_24267);
nand UO_2605 (O_2605,N_24473,N_23598);
xnor UO_2606 (O_2606,N_22566,N_23382);
nor UO_2607 (O_2607,N_22943,N_24938);
nor UO_2608 (O_2608,N_23525,N_23583);
nand UO_2609 (O_2609,N_23762,N_22707);
or UO_2610 (O_2610,N_24013,N_24208);
or UO_2611 (O_2611,N_23878,N_23535);
and UO_2612 (O_2612,N_24660,N_23527);
nand UO_2613 (O_2613,N_24481,N_23739);
nand UO_2614 (O_2614,N_23218,N_24847);
nand UO_2615 (O_2615,N_22708,N_24556);
nand UO_2616 (O_2616,N_24866,N_24211);
nand UO_2617 (O_2617,N_23806,N_24439);
or UO_2618 (O_2618,N_23105,N_24678);
nor UO_2619 (O_2619,N_22540,N_23736);
nand UO_2620 (O_2620,N_23451,N_24451);
nor UO_2621 (O_2621,N_23739,N_24052);
nor UO_2622 (O_2622,N_23602,N_24231);
nor UO_2623 (O_2623,N_23068,N_23150);
nor UO_2624 (O_2624,N_23728,N_23529);
and UO_2625 (O_2625,N_23768,N_24442);
xnor UO_2626 (O_2626,N_24672,N_24949);
and UO_2627 (O_2627,N_24477,N_24788);
nor UO_2628 (O_2628,N_23441,N_23190);
and UO_2629 (O_2629,N_22562,N_23663);
nor UO_2630 (O_2630,N_24479,N_23879);
or UO_2631 (O_2631,N_24179,N_23906);
nand UO_2632 (O_2632,N_23846,N_22761);
nor UO_2633 (O_2633,N_23983,N_22572);
nor UO_2634 (O_2634,N_23007,N_23539);
or UO_2635 (O_2635,N_23460,N_22516);
and UO_2636 (O_2636,N_22660,N_22597);
nor UO_2637 (O_2637,N_23610,N_23343);
nor UO_2638 (O_2638,N_23612,N_24371);
xnor UO_2639 (O_2639,N_23900,N_22576);
or UO_2640 (O_2640,N_23989,N_23316);
xor UO_2641 (O_2641,N_22621,N_23362);
or UO_2642 (O_2642,N_23444,N_23689);
xnor UO_2643 (O_2643,N_24940,N_22536);
or UO_2644 (O_2644,N_23541,N_24100);
or UO_2645 (O_2645,N_23095,N_23276);
or UO_2646 (O_2646,N_22812,N_22763);
nand UO_2647 (O_2647,N_24637,N_24106);
nor UO_2648 (O_2648,N_24558,N_23509);
nand UO_2649 (O_2649,N_23375,N_23125);
and UO_2650 (O_2650,N_24802,N_24410);
or UO_2651 (O_2651,N_23472,N_23495);
nor UO_2652 (O_2652,N_22994,N_22641);
nand UO_2653 (O_2653,N_22762,N_24495);
xnor UO_2654 (O_2654,N_24277,N_24596);
or UO_2655 (O_2655,N_22921,N_23705);
and UO_2656 (O_2656,N_24282,N_23040);
nor UO_2657 (O_2657,N_23911,N_24226);
and UO_2658 (O_2658,N_24737,N_22985);
and UO_2659 (O_2659,N_22846,N_23130);
nand UO_2660 (O_2660,N_23712,N_23926);
nor UO_2661 (O_2661,N_24344,N_24104);
and UO_2662 (O_2662,N_24125,N_24640);
or UO_2663 (O_2663,N_24879,N_24838);
xor UO_2664 (O_2664,N_23882,N_24228);
nand UO_2665 (O_2665,N_24924,N_23682);
or UO_2666 (O_2666,N_23229,N_23526);
and UO_2667 (O_2667,N_22834,N_22902);
nand UO_2668 (O_2668,N_22711,N_22820);
and UO_2669 (O_2669,N_24588,N_24982);
or UO_2670 (O_2670,N_23717,N_22773);
xnor UO_2671 (O_2671,N_23701,N_23852);
xnor UO_2672 (O_2672,N_23618,N_22681);
nand UO_2673 (O_2673,N_23586,N_24220);
nor UO_2674 (O_2674,N_24175,N_24847);
or UO_2675 (O_2675,N_23143,N_23887);
xor UO_2676 (O_2676,N_24676,N_23790);
nand UO_2677 (O_2677,N_24635,N_23561);
nor UO_2678 (O_2678,N_23785,N_24777);
and UO_2679 (O_2679,N_23485,N_24439);
nand UO_2680 (O_2680,N_23876,N_24377);
xor UO_2681 (O_2681,N_23106,N_24543);
xnor UO_2682 (O_2682,N_24811,N_24632);
or UO_2683 (O_2683,N_22531,N_23694);
xor UO_2684 (O_2684,N_24417,N_23218);
or UO_2685 (O_2685,N_24305,N_22603);
xnor UO_2686 (O_2686,N_22731,N_24822);
xor UO_2687 (O_2687,N_23328,N_24827);
and UO_2688 (O_2688,N_23475,N_22627);
xor UO_2689 (O_2689,N_23468,N_23632);
or UO_2690 (O_2690,N_24488,N_24678);
or UO_2691 (O_2691,N_24842,N_23900);
nand UO_2692 (O_2692,N_24336,N_24117);
and UO_2693 (O_2693,N_23091,N_24606);
xor UO_2694 (O_2694,N_24646,N_23291);
or UO_2695 (O_2695,N_23076,N_23733);
and UO_2696 (O_2696,N_23414,N_24834);
nand UO_2697 (O_2697,N_24179,N_23136);
and UO_2698 (O_2698,N_23134,N_23426);
nand UO_2699 (O_2699,N_24887,N_24601);
xor UO_2700 (O_2700,N_24213,N_23901);
nor UO_2701 (O_2701,N_23548,N_24386);
nand UO_2702 (O_2702,N_24015,N_24061);
xnor UO_2703 (O_2703,N_23607,N_24499);
xnor UO_2704 (O_2704,N_23224,N_24360);
nand UO_2705 (O_2705,N_24989,N_24749);
nor UO_2706 (O_2706,N_24370,N_24455);
nand UO_2707 (O_2707,N_23239,N_23550);
nor UO_2708 (O_2708,N_23540,N_24900);
nand UO_2709 (O_2709,N_24400,N_24709);
xor UO_2710 (O_2710,N_23510,N_24018);
and UO_2711 (O_2711,N_22820,N_22937);
or UO_2712 (O_2712,N_23614,N_24931);
nand UO_2713 (O_2713,N_24005,N_24755);
nor UO_2714 (O_2714,N_23815,N_22663);
xnor UO_2715 (O_2715,N_23335,N_23587);
and UO_2716 (O_2716,N_23431,N_23166);
nor UO_2717 (O_2717,N_24233,N_23151);
nand UO_2718 (O_2718,N_22747,N_22565);
nor UO_2719 (O_2719,N_23796,N_24760);
or UO_2720 (O_2720,N_24418,N_23549);
or UO_2721 (O_2721,N_24588,N_24530);
or UO_2722 (O_2722,N_23198,N_24944);
xor UO_2723 (O_2723,N_23976,N_24316);
and UO_2724 (O_2724,N_23142,N_24809);
nand UO_2725 (O_2725,N_23507,N_24574);
nand UO_2726 (O_2726,N_24606,N_24554);
and UO_2727 (O_2727,N_23702,N_23059);
or UO_2728 (O_2728,N_24253,N_23447);
xnor UO_2729 (O_2729,N_23033,N_23197);
nand UO_2730 (O_2730,N_24136,N_24950);
nand UO_2731 (O_2731,N_24492,N_24560);
and UO_2732 (O_2732,N_23654,N_23947);
xor UO_2733 (O_2733,N_23639,N_22915);
xnor UO_2734 (O_2734,N_24089,N_24147);
xnor UO_2735 (O_2735,N_23724,N_24455);
xnor UO_2736 (O_2736,N_23178,N_23820);
or UO_2737 (O_2737,N_24459,N_24042);
or UO_2738 (O_2738,N_24201,N_22882);
and UO_2739 (O_2739,N_22653,N_24740);
or UO_2740 (O_2740,N_24919,N_22845);
nor UO_2741 (O_2741,N_23904,N_23822);
nand UO_2742 (O_2742,N_23953,N_23903);
or UO_2743 (O_2743,N_22772,N_23346);
nand UO_2744 (O_2744,N_24234,N_24460);
xor UO_2745 (O_2745,N_23880,N_24696);
or UO_2746 (O_2746,N_24046,N_23520);
nor UO_2747 (O_2747,N_24188,N_24514);
xnor UO_2748 (O_2748,N_24225,N_24047);
xor UO_2749 (O_2749,N_23588,N_24147);
xor UO_2750 (O_2750,N_23871,N_23539);
or UO_2751 (O_2751,N_23126,N_24869);
nor UO_2752 (O_2752,N_24771,N_24666);
nand UO_2753 (O_2753,N_24042,N_24770);
and UO_2754 (O_2754,N_23756,N_22538);
and UO_2755 (O_2755,N_23483,N_22760);
nand UO_2756 (O_2756,N_23877,N_23273);
and UO_2757 (O_2757,N_23608,N_23291);
or UO_2758 (O_2758,N_24210,N_24846);
and UO_2759 (O_2759,N_22979,N_22814);
nand UO_2760 (O_2760,N_22819,N_24740);
nand UO_2761 (O_2761,N_24278,N_24416);
or UO_2762 (O_2762,N_24884,N_22697);
xnor UO_2763 (O_2763,N_24637,N_22690);
xnor UO_2764 (O_2764,N_24010,N_24593);
nand UO_2765 (O_2765,N_22979,N_24229);
or UO_2766 (O_2766,N_23882,N_23219);
nor UO_2767 (O_2767,N_22703,N_24809);
or UO_2768 (O_2768,N_23157,N_23173);
nand UO_2769 (O_2769,N_23867,N_23460);
nor UO_2770 (O_2770,N_24066,N_23912);
nand UO_2771 (O_2771,N_22997,N_23173);
xnor UO_2772 (O_2772,N_22755,N_23115);
and UO_2773 (O_2773,N_23953,N_23813);
xnor UO_2774 (O_2774,N_24061,N_24123);
xor UO_2775 (O_2775,N_24380,N_23832);
xor UO_2776 (O_2776,N_24368,N_23415);
and UO_2777 (O_2777,N_22555,N_23203);
nand UO_2778 (O_2778,N_22621,N_24915);
or UO_2779 (O_2779,N_23249,N_24457);
and UO_2780 (O_2780,N_23269,N_24178);
or UO_2781 (O_2781,N_23963,N_24407);
nand UO_2782 (O_2782,N_23986,N_22939);
nand UO_2783 (O_2783,N_23445,N_24706);
and UO_2784 (O_2784,N_24551,N_23220);
or UO_2785 (O_2785,N_23899,N_23960);
xor UO_2786 (O_2786,N_23056,N_24880);
nor UO_2787 (O_2787,N_24940,N_23611);
nand UO_2788 (O_2788,N_24756,N_24641);
nor UO_2789 (O_2789,N_24167,N_22680);
or UO_2790 (O_2790,N_22945,N_23489);
or UO_2791 (O_2791,N_23954,N_22882);
xor UO_2792 (O_2792,N_23422,N_23687);
nand UO_2793 (O_2793,N_22623,N_22660);
or UO_2794 (O_2794,N_24463,N_23321);
nor UO_2795 (O_2795,N_23611,N_23366);
xnor UO_2796 (O_2796,N_24819,N_23430);
and UO_2797 (O_2797,N_22605,N_22532);
and UO_2798 (O_2798,N_22653,N_23219);
and UO_2799 (O_2799,N_22728,N_24995);
and UO_2800 (O_2800,N_24702,N_23183);
xor UO_2801 (O_2801,N_22969,N_23836);
nand UO_2802 (O_2802,N_24907,N_24489);
and UO_2803 (O_2803,N_22988,N_24849);
xor UO_2804 (O_2804,N_24744,N_22771);
xnor UO_2805 (O_2805,N_23922,N_23535);
nor UO_2806 (O_2806,N_24030,N_24833);
and UO_2807 (O_2807,N_22887,N_23463);
or UO_2808 (O_2808,N_22594,N_22802);
nor UO_2809 (O_2809,N_23398,N_23577);
and UO_2810 (O_2810,N_22541,N_24432);
and UO_2811 (O_2811,N_22902,N_24870);
or UO_2812 (O_2812,N_22944,N_23438);
nor UO_2813 (O_2813,N_22742,N_24094);
xnor UO_2814 (O_2814,N_24545,N_23532);
nor UO_2815 (O_2815,N_23088,N_23030);
and UO_2816 (O_2816,N_23805,N_23414);
and UO_2817 (O_2817,N_23968,N_23093);
or UO_2818 (O_2818,N_23023,N_24194);
nand UO_2819 (O_2819,N_22829,N_24421);
nor UO_2820 (O_2820,N_23230,N_23166);
nand UO_2821 (O_2821,N_23749,N_24311);
nand UO_2822 (O_2822,N_23815,N_24677);
xor UO_2823 (O_2823,N_23751,N_23126);
or UO_2824 (O_2824,N_23943,N_24592);
nand UO_2825 (O_2825,N_23055,N_22592);
nand UO_2826 (O_2826,N_24300,N_22973);
and UO_2827 (O_2827,N_24105,N_24089);
xor UO_2828 (O_2828,N_23014,N_23284);
or UO_2829 (O_2829,N_24874,N_24621);
nor UO_2830 (O_2830,N_24769,N_23286);
or UO_2831 (O_2831,N_24662,N_22576);
xor UO_2832 (O_2832,N_23970,N_24762);
nor UO_2833 (O_2833,N_22981,N_22654);
and UO_2834 (O_2834,N_23623,N_23267);
nand UO_2835 (O_2835,N_22580,N_24172);
or UO_2836 (O_2836,N_24615,N_24845);
and UO_2837 (O_2837,N_24113,N_24465);
or UO_2838 (O_2838,N_23332,N_23430);
xnor UO_2839 (O_2839,N_24267,N_24834);
nand UO_2840 (O_2840,N_23740,N_23049);
nand UO_2841 (O_2841,N_23891,N_23538);
or UO_2842 (O_2842,N_23430,N_24916);
nor UO_2843 (O_2843,N_23599,N_23386);
nor UO_2844 (O_2844,N_23636,N_23631);
or UO_2845 (O_2845,N_23277,N_23472);
nor UO_2846 (O_2846,N_24851,N_23746);
nand UO_2847 (O_2847,N_23122,N_24968);
and UO_2848 (O_2848,N_24536,N_23863);
and UO_2849 (O_2849,N_23031,N_22523);
nand UO_2850 (O_2850,N_23972,N_23886);
or UO_2851 (O_2851,N_24980,N_23557);
nand UO_2852 (O_2852,N_23978,N_22978);
xnor UO_2853 (O_2853,N_22903,N_24891);
and UO_2854 (O_2854,N_23617,N_23578);
nor UO_2855 (O_2855,N_22835,N_24456);
and UO_2856 (O_2856,N_24822,N_24796);
nand UO_2857 (O_2857,N_24150,N_24574);
or UO_2858 (O_2858,N_22802,N_24921);
and UO_2859 (O_2859,N_22686,N_22683);
nand UO_2860 (O_2860,N_23938,N_23018);
and UO_2861 (O_2861,N_22615,N_23862);
or UO_2862 (O_2862,N_24000,N_23309);
nor UO_2863 (O_2863,N_24859,N_24836);
and UO_2864 (O_2864,N_24173,N_22503);
nor UO_2865 (O_2865,N_22700,N_23162);
nor UO_2866 (O_2866,N_23706,N_23339);
nor UO_2867 (O_2867,N_22905,N_23726);
nor UO_2868 (O_2868,N_23507,N_24849);
and UO_2869 (O_2869,N_22802,N_23865);
nand UO_2870 (O_2870,N_23613,N_23777);
xor UO_2871 (O_2871,N_24844,N_22786);
nor UO_2872 (O_2872,N_23397,N_24984);
and UO_2873 (O_2873,N_23392,N_23568);
xnor UO_2874 (O_2874,N_23509,N_23859);
or UO_2875 (O_2875,N_24772,N_23714);
or UO_2876 (O_2876,N_24126,N_24635);
nor UO_2877 (O_2877,N_24961,N_24401);
nand UO_2878 (O_2878,N_23838,N_24595);
and UO_2879 (O_2879,N_24746,N_24526);
and UO_2880 (O_2880,N_23063,N_24362);
nor UO_2881 (O_2881,N_22882,N_24042);
nor UO_2882 (O_2882,N_22570,N_23093);
and UO_2883 (O_2883,N_24050,N_23297);
nand UO_2884 (O_2884,N_22926,N_24162);
xnor UO_2885 (O_2885,N_24312,N_23345);
nor UO_2886 (O_2886,N_23201,N_23251);
and UO_2887 (O_2887,N_22782,N_24277);
nor UO_2888 (O_2888,N_22981,N_23874);
or UO_2889 (O_2889,N_24312,N_23255);
xor UO_2890 (O_2890,N_23222,N_24680);
xor UO_2891 (O_2891,N_23953,N_23515);
xor UO_2892 (O_2892,N_22695,N_24461);
nand UO_2893 (O_2893,N_24921,N_22856);
nor UO_2894 (O_2894,N_24759,N_24076);
nand UO_2895 (O_2895,N_23053,N_23862);
nor UO_2896 (O_2896,N_22764,N_24731);
and UO_2897 (O_2897,N_23769,N_23680);
nor UO_2898 (O_2898,N_24622,N_24355);
nor UO_2899 (O_2899,N_22726,N_24404);
and UO_2900 (O_2900,N_22630,N_23053);
nand UO_2901 (O_2901,N_23108,N_23950);
nor UO_2902 (O_2902,N_22579,N_23634);
and UO_2903 (O_2903,N_24258,N_23012);
nand UO_2904 (O_2904,N_23243,N_22869);
nand UO_2905 (O_2905,N_22852,N_24670);
and UO_2906 (O_2906,N_23409,N_24004);
and UO_2907 (O_2907,N_24753,N_22933);
nor UO_2908 (O_2908,N_24582,N_22616);
xor UO_2909 (O_2909,N_22746,N_24179);
or UO_2910 (O_2910,N_24210,N_24145);
and UO_2911 (O_2911,N_23121,N_22972);
or UO_2912 (O_2912,N_23072,N_24334);
nor UO_2913 (O_2913,N_24213,N_24987);
and UO_2914 (O_2914,N_23388,N_22794);
and UO_2915 (O_2915,N_24508,N_24696);
or UO_2916 (O_2916,N_24928,N_24623);
and UO_2917 (O_2917,N_24452,N_23888);
nor UO_2918 (O_2918,N_22919,N_24898);
or UO_2919 (O_2919,N_24804,N_23745);
nor UO_2920 (O_2920,N_24754,N_24614);
nand UO_2921 (O_2921,N_23462,N_24270);
or UO_2922 (O_2922,N_24465,N_24693);
nand UO_2923 (O_2923,N_24572,N_23542);
nand UO_2924 (O_2924,N_22821,N_23332);
xor UO_2925 (O_2925,N_22913,N_22977);
and UO_2926 (O_2926,N_23220,N_24245);
and UO_2927 (O_2927,N_23055,N_23832);
xor UO_2928 (O_2928,N_24423,N_24574);
nand UO_2929 (O_2929,N_23728,N_23674);
nand UO_2930 (O_2930,N_24968,N_22803);
nand UO_2931 (O_2931,N_23776,N_23600);
nand UO_2932 (O_2932,N_24841,N_23620);
nand UO_2933 (O_2933,N_22981,N_22909);
xor UO_2934 (O_2934,N_24943,N_24730);
xnor UO_2935 (O_2935,N_24280,N_23644);
and UO_2936 (O_2936,N_24479,N_23010);
and UO_2937 (O_2937,N_24731,N_24863);
nor UO_2938 (O_2938,N_23743,N_22860);
nand UO_2939 (O_2939,N_24801,N_23639);
or UO_2940 (O_2940,N_23691,N_23001);
nor UO_2941 (O_2941,N_23081,N_24593);
and UO_2942 (O_2942,N_23363,N_23250);
xor UO_2943 (O_2943,N_24777,N_24494);
nand UO_2944 (O_2944,N_22750,N_23029);
nand UO_2945 (O_2945,N_23325,N_24756);
nor UO_2946 (O_2946,N_24118,N_23868);
or UO_2947 (O_2947,N_23705,N_23303);
nand UO_2948 (O_2948,N_22888,N_24237);
nand UO_2949 (O_2949,N_24514,N_24504);
nand UO_2950 (O_2950,N_23417,N_23549);
and UO_2951 (O_2951,N_23225,N_23284);
xnor UO_2952 (O_2952,N_24808,N_24003);
nand UO_2953 (O_2953,N_24281,N_24669);
xnor UO_2954 (O_2954,N_23784,N_24323);
or UO_2955 (O_2955,N_23931,N_24599);
xor UO_2956 (O_2956,N_23565,N_23292);
nand UO_2957 (O_2957,N_23746,N_23183);
nor UO_2958 (O_2958,N_23587,N_24360);
and UO_2959 (O_2959,N_24576,N_23187);
xnor UO_2960 (O_2960,N_22657,N_23149);
and UO_2961 (O_2961,N_24415,N_22817);
or UO_2962 (O_2962,N_22848,N_24471);
nor UO_2963 (O_2963,N_24168,N_23231);
nand UO_2964 (O_2964,N_23554,N_24147);
and UO_2965 (O_2965,N_24871,N_23574);
and UO_2966 (O_2966,N_23072,N_23450);
nand UO_2967 (O_2967,N_22914,N_24257);
xnor UO_2968 (O_2968,N_24759,N_23263);
or UO_2969 (O_2969,N_24732,N_24690);
nand UO_2970 (O_2970,N_24016,N_23328);
xor UO_2971 (O_2971,N_24383,N_24255);
or UO_2972 (O_2972,N_23892,N_22569);
and UO_2973 (O_2973,N_23887,N_24444);
nand UO_2974 (O_2974,N_23628,N_24144);
nand UO_2975 (O_2975,N_22530,N_22909);
and UO_2976 (O_2976,N_23783,N_23623);
xnor UO_2977 (O_2977,N_22981,N_22589);
or UO_2978 (O_2978,N_24045,N_23207);
xor UO_2979 (O_2979,N_22844,N_23897);
xor UO_2980 (O_2980,N_22819,N_24435);
or UO_2981 (O_2981,N_23485,N_24569);
nand UO_2982 (O_2982,N_24756,N_23879);
nor UO_2983 (O_2983,N_22995,N_24187);
or UO_2984 (O_2984,N_24445,N_22686);
xnor UO_2985 (O_2985,N_22874,N_23224);
xor UO_2986 (O_2986,N_24511,N_24081);
nor UO_2987 (O_2987,N_24769,N_24585);
xor UO_2988 (O_2988,N_23740,N_23632);
and UO_2989 (O_2989,N_23037,N_23501);
xor UO_2990 (O_2990,N_24758,N_23157);
or UO_2991 (O_2991,N_24210,N_23338);
and UO_2992 (O_2992,N_24239,N_22982);
nand UO_2993 (O_2993,N_22668,N_23409);
or UO_2994 (O_2994,N_24389,N_23698);
nor UO_2995 (O_2995,N_24303,N_24524);
and UO_2996 (O_2996,N_22811,N_23916);
or UO_2997 (O_2997,N_24909,N_22651);
and UO_2998 (O_2998,N_23604,N_23376);
nand UO_2999 (O_2999,N_22655,N_24178);
endmodule