module basic_1000_10000_1500_4_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_909,In_497);
nor U1 (N_1,In_983,In_487);
or U2 (N_2,In_163,In_486);
nor U3 (N_3,In_600,In_534);
or U4 (N_4,In_561,In_799);
or U5 (N_5,In_133,In_918);
or U6 (N_6,In_504,In_851);
and U7 (N_7,In_44,In_228);
or U8 (N_8,In_858,In_149);
or U9 (N_9,In_20,In_307);
nor U10 (N_10,In_996,In_246);
nand U11 (N_11,In_308,In_71);
nor U12 (N_12,In_256,In_452);
nor U13 (N_13,In_578,In_88);
nor U14 (N_14,In_984,In_939);
nor U15 (N_15,In_377,In_105);
or U16 (N_16,In_310,In_813);
nand U17 (N_17,In_570,In_254);
nand U18 (N_18,In_782,In_533);
nor U19 (N_19,In_510,In_325);
or U20 (N_20,In_917,In_949);
and U21 (N_21,In_746,In_962);
nor U22 (N_22,In_936,In_740);
nor U23 (N_23,In_944,In_340);
nor U24 (N_24,In_395,In_480);
nor U25 (N_25,In_147,In_502);
nand U26 (N_26,In_950,In_37);
and U27 (N_27,In_836,In_47);
nor U28 (N_28,In_104,In_679);
or U29 (N_29,In_328,In_172);
or U30 (N_30,In_542,In_16);
nand U31 (N_31,In_733,In_579);
nand U32 (N_32,In_439,In_346);
and U33 (N_33,In_192,In_882);
nand U34 (N_34,In_258,In_139);
nor U35 (N_35,In_519,In_273);
nor U36 (N_36,In_287,In_198);
nand U37 (N_37,In_576,In_0);
nand U38 (N_38,In_165,In_194);
and U39 (N_39,In_134,In_176);
and U40 (N_40,In_577,In_370);
xnor U41 (N_41,In_634,In_831);
xnor U42 (N_42,In_787,In_922);
or U43 (N_43,In_619,In_976);
nand U44 (N_44,In_343,In_801);
or U45 (N_45,In_613,In_617);
or U46 (N_46,In_415,In_568);
or U47 (N_47,In_540,In_276);
or U48 (N_48,In_771,In_249);
or U49 (N_49,In_441,In_896);
and U50 (N_50,In_349,In_51);
or U51 (N_51,In_825,In_253);
nand U52 (N_52,In_34,In_775);
nor U53 (N_53,In_436,In_989);
or U54 (N_54,In_709,In_162);
nor U55 (N_55,In_943,In_523);
or U56 (N_56,In_803,In_695);
or U57 (N_57,In_424,In_868);
nor U58 (N_58,In_505,In_394);
or U59 (N_59,In_814,In_95);
and U60 (N_60,In_969,In_443);
or U61 (N_61,In_379,In_83);
nor U62 (N_62,In_604,In_530);
or U63 (N_63,In_947,In_649);
and U64 (N_64,In_602,In_699);
or U65 (N_65,In_509,In_442);
or U66 (N_66,In_376,In_68);
and U67 (N_67,In_419,In_365);
and U68 (N_68,In_437,In_304);
nand U69 (N_69,In_333,In_206);
xnor U70 (N_70,In_400,In_60);
nor U71 (N_71,In_218,In_496);
or U72 (N_72,In_555,In_214);
nand U73 (N_73,In_190,In_942);
nand U74 (N_74,In_352,In_375);
nor U75 (N_75,In_824,In_702);
or U76 (N_76,In_76,In_627);
nor U77 (N_77,In_636,In_488);
or U78 (N_78,In_418,In_946);
and U79 (N_79,In_914,In_168);
nor U80 (N_80,In_716,In_562);
or U81 (N_81,In_200,In_433);
or U82 (N_82,In_120,In_770);
nor U83 (N_83,In_977,In_475);
nand U84 (N_84,In_238,In_817);
or U85 (N_85,In_675,In_887);
or U86 (N_86,In_351,In_177);
and U87 (N_87,In_131,In_390);
or U88 (N_88,In_109,In_591);
and U89 (N_89,In_654,In_148);
nand U90 (N_90,In_466,In_151);
nor U91 (N_91,In_528,In_678);
nand U92 (N_92,In_313,In_317);
nor U93 (N_93,In_311,In_669);
nor U94 (N_94,In_335,In_687);
nand U95 (N_95,In_762,In_220);
nand U96 (N_96,In_889,In_369);
and U97 (N_97,In_141,In_181);
and U98 (N_98,In_75,In_387);
nor U99 (N_99,In_684,In_144);
nand U100 (N_100,In_30,In_558);
and U101 (N_101,In_143,In_430);
or U102 (N_102,In_598,In_324);
nor U103 (N_103,In_638,In_535);
and U104 (N_104,In_284,In_671);
and U105 (N_105,In_462,In_900);
or U106 (N_106,In_501,In_221);
or U107 (N_107,In_92,In_551);
nand U108 (N_108,In_404,In_897);
nand U109 (N_109,In_987,In_538);
nand U110 (N_110,In_802,In_696);
nor U111 (N_111,In_268,In_211);
and U112 (N_112,In_145,In_137);
and U113 (N_113,In_848,In_507);
nand U114 (N_114,In_880,In_903);
and U115 (N_115,In_512,In_783);
or U116 (N_116,In_715,In_648);
or U117 (N_117,In_719,In_315);
or U118 (N_118,In_626,In_477);
nor U119 (N_119,In_64,In_749);
and U120 (N_120,In_590,In_291);
nand U121 (N_121,In_658,In_691);
and U122 (N_122,In_411,In_22);
nor U123 (N_123,In_881,In_854);
nor U124 (N_124,In_189,In_718);
and U125 (N_125,In_99,In_393);
or U126 (N_126,In_864,In_61);
or U127 (N_127,In_457,In_757);
or U128 (N_128,In_845,In_237);
nor U129 (N_129,In_282,In_999);
nand U130 (N_130,In_330,In_549);
and U131 (N_131,In_605,In_859);
nor U132 (N_132,In_642,In_456);
nand U133 (N_133,In_130,In_96);
and U134 (N_134,In_266,In_403);
nor U135 (N_135,In_731,In_809);
or U136 (N_136,In_263,In_650);
nand U137 (N_137,In_724,In_117);
or U138 (N_138,In_853,In_589);
or U139 (N_139,In_378,In_791);
and U140 (N_140,In_705,In_884);
nor U141 (N_141,In_170,In_837);
or U142 (N_142,In_520,In_839);
and U143 (N_143,In_612,In_132);
nand U144 (N_144,In_753,In_416);
or U145 (N_145,In_861,In_847);
or U146 (N_146,In_17,In_662);
or U147 (N_147,In_574,In_532);
and U148 (N_148,In_472,In_656);
and U149 (N_149,In_511,In_855);
and U150 (N_150,In_24,In_832);
or U151 (N_151,In_913,In_111);
or U152 (N_152,In_763,In_469);
nand U153 (N_153,In_123,In_85);
nand U154 (N_154,In_40,In_524);
and U155 (N_155,In_660,In_153);
or U156 (N_156,In_150,In_157);
nand U157 (N_157,In_710,In_86);
or U158 (N_158,In_923,In_956);
and U159 (N_159,In_478,In_657);
and U160 (N_160,In_384,In_385);
or U161 (N_161,In_810,In_309);
nor U162 (N_162,In_87,In_828);
nand U163 (N_163,In_713,In_197);
nor U164 (N_164,In_916,In_780);
or U165 (N_165,In_793,In_635);
or U166 (N_166,In_128,In_727);
or U167 (N_167,In_166,In_907);
nand U168 (N_168,In_222,In_171);
nor U169 (N_169,In_615,In_664);
or U170 (N_170,In_28,In_643);
nor U171 (N_171,In_54,In_259);
or U172 (N_172,In_722,In_483);
or U173 (N_173,In_373,In_371);
or U174 (N_174,In_863,In_611);
nand U175 (N_175,In_167,In_21);
and U176 (N_176,In_464,In_103);
nor U177 (N_177,In_547,In_618);
and U178 (N_178,In_750,In_525);
nand U179 (N_179,In_630,In_788);
and U180 (N_180,In_894,In_14);
or U181 (N_181,In_169,In_930);
and U182 (N_182,In_794,In_732);
nor U183 (N_183,In_712,In_53);
xnor U184 (N_184,In_427,In_739);
nor U185 (N_185,In_119,In_758);
and U186 (N_186,In_790,In_931);
nand U187 (N_187,In_700,In_46);
or U188 (N_188,In_431,In_676);
and U189 (N_189,In_10,In_647);
nand U190 (N_190,In_711,In_322);
nor U191 (N_191,In_777,In_596);
or U192 (N_192,In_429,In_65);
and U193 (N_193,In_125,In_216);
nand U194 (N_194,In_215,In_633);
and U195 (N_195,In_734,In_760);
nand U196 (N_196,In_808,In_986);
and U197 (N_197,In_18,In_693);
nand U198 (N_198,In_932,In_797);
nand U199 (N_199,In_970,In_666);
and U200 (N_200,In_632,In_721);
or U201 (N_201,In_629,In_892);
nor U202 (N_202,In_331,In_826);
and U203 (N_203,In_821,In_955);
nand U204 (N_204,In_232,In_689);
and U205 (N_205,In_280,In_529);
nor U206 (N_206,In_108,In_954);
nor U207 (N_207,In_895,In_468);
nor U208 (N_208,In_252,In_481);
or U209 (N_209,In_42,In_267);
and U210 (N_210,In_901,In_624);
and U211 (N_211,In_292,In_982);
or U212 (N_212,In_514,In_101);
or U213 (N_213,In_467,In_364);
and U214 (N_214,In_849,In_607);
nand U215 (N_215,In_243,In_332);
or U216 (N_216,In_455,In_623);
nor U217 (N_217,In_703,In_495);
nor U218 (N_218,In_417,In_186);
nor U219 (N_219,In_78,In_7);
and U220 (N_220,In_645,In_893);
or U221 (N_221,In_816,In_743);
nand U222 (N_222,In_992,In_935);
nor U223 (N_223,In_960,In_122);
and U224 (N_224,In_339,In_257);
or U225 (N_225,In_798,In_806);
nor U226 (N_226,In_846,In_730);
or U227 (N_227,In_326,In_334);
nand U228 (N_228,In_386,In_871);
and U229 (N_229,In_432,In_536);
nand U230 (N_230,In_242,In_142);
and U231 (N_231,In_974,In_911);
nand U232 (N_232,In_36,In_616);
nor U233 (N_233,In_840,In_174);
and U234 (N_234,In_91,In_637);
nor U235 (N_235,In_250,In_73);
or U236 (N_236,In_569,In_245);
or U237 (N_237,In_856,In_460);
nand U238 (N_238,In_476,In_751);
nand U239 (N_239,In_571,In_508);
nand U240 (N_240,In_873,In_941);
or U241 (N_241,In_230,In_708);
nand U242 (N_242,In_227,In_236);
nand U243 (N_243,In_398,In_207);
nor U244 (N_244,In_952,In_354);
nand U245 (N_245,In_203,In_97);
nand U246 (N_246,In_875,In_644);
and U247 (N_247,In_513,In_359);
nor U248 (N_248,In_926,In_792);
nor U249 (N_249,In_920,In_585);
and U250 (N_250,In_725,In_565);
nand U251 (N_251,In_231,In_164);
nor U252 (N_252,In_422,In_885);
xor U253 (N_253,In_973,In_659);
or U254 (N_254,In_233,In_77);
and U255 (N_255,In_193,In_518);
nand U256 (N_256,In_517,In_318);
nor U257 (N_257,In_539,In_870);
or U258 (N_258,In_420,In_736);
nand U259 (N_259,In_912,In_209);
and U260 (N_260,In_599,In_631);
nand U261 (N_261,In_902,In_444);
nor U262 (N_262,In_556,In_680);
nand U263 (N_263,In_473,In_426);
or U264 (N_264,In_672,In_500);
or U265 (N_265,In_158,In_503);
nand U266 (N_266,In_776,In_668);
nor U267 (N_267,In_552,In_557);
nor U268 (N_268,In_779,In_191);
and U269 (N_269,In_906,In_541);
nor U270 (N_270,In_360,In_872);
or U271 (N_271,In_819,In_597);
and U272 (N_272,In_405,In_298);
or U273 (N_273,In_964,In_247);
or U274 (N_274,In_625,In_124);
and U275 (N_275,In_723,In_261);
and U276 (N_276,In_592,In_670);
nor U277 (N_277,In_959,In_41);
nand U278 (N_278,In_82,In_127);
and U279 (N_279,In_6,In_448);
nor U280 (N_280,In_835,In_219);
or U281 (N_281,In_12,In_260);
and U282 (N_282,In_23,In_115);
nor U283 (N_283,In_971,In_929);
nor U284 (N_284,In_179,In_274);
nand U285 (N_285,In_240,In_62);
and U286 (N_286,In_766,In_159);
nor U287 (N_287,In_651,In_301);
and U288 (N_288,In_58,In_412);
nor U289 (N_289,In_747,In_434);
nand U290 (N_290,In_126,In_640);
and U291 (N_291,In_320,In_686);
nor U292 (N_292,In_321,In_842);
or U293 (N_293,In_327,In_471);
and U294 (N_294,In_957,In_720);
nand U295 (N_295,In_288,In_494);
nand U296 (N_296,In_31,In_294);
nor U297 (N_297,In_463,In_217);
or U298 (N_298,In_990,In_66);
or U299 (N_299,In_161,In_239);
nor U300 (N_300,In_402,In_756);
nor U301 (N_301,In_899,In_754);
or U302 (N_302,In_515,In_449);
nor U303 (N_303,In_934,In_305);
or U304 (N_304,In_204,In_362);
or U305 (N_305,In_614,In_347);
or U306 (N_306,In_993,In_474);
or U307 (N_307,In_554,In_461);
nand U308 (N_308,In_714,In_366);
nor U309 (N_309,In_271,In_805);
nand U310 (N_310,In_641,In_823);
and U311 (N_311,In_800,In_586);
nor U312 (N_312,In_414,In_188);
and U313 (N_313,In_685,In_620);
nor U314 (N_314,In_898,In_564);
nand U315 (N_315,In_963,In_269);
and U316 (N_316,In_453,In_933);
nor U317 (N_317,In_652,In_70);
nor U318 (N_318,In_178,In_69);
nor U319 (N_319,In_303,In_94);
or U320 (N_320,In_818,In_363);
and U321 (N_321,In_891,In_761);
or U322 (N_322,In_234,In_583);
and U323 (N_323,In_290,In_812);
and U324 (N_324,In_910,In_768);
and U325 (N_325,In_811,In_752);
nor U326 (N_326,In_735,In_850);
nor U327 (N_327,In_100,In_965);
nand U328 (N_328,In_544,In_865);
and U329 (N_329,In_195,In_961);
nand U330 (N_330,In_994,In_380);
and U331 (N_331,In_878,In_559);
nand U332 (N_332,In_833,In_183);
and U333 (N_333,In_458,In_350);
or U334 (N_334,In_278,In_820);
or U335 (N_335,In_726,In_498);
nor U336 (N_336,In_52,In_49);
or U337 (N_337,In_692,In_226);
nand U338 (N_338,In_830,In_396);
nand U339 (N_339,In_694,In_81);
nand U340 (N_340,In_84,In_829);
nor U341 (N_341,In_212,In_603);
nor U342 (N_342,In_673,In_784);
or U343 (N_343,In_201,In_265);
nand U344 (N_344,In_187,In_606);
and U345 (N_345,In_285,In_862);
and U346 (N_346,In_927,In_815);
xor U347 (N_347,In_796,In_857);
nand U348 (N_348,In_581,In_948);
or U349 (N_349,In_667,In_2);
nor U350 (N_350,In_136,In_459);
nor U351 (N_351,In_275,In_154);
nor U352 (N_352,In_866,In_838);
nand U353 (N_353,In_300,In_925);
nor U354 (N_354,In_665,In_272);
or U355 (N_355,In_56,In_470);
nand U356 (N_356,In_406,In_213);
and U357 (N_357,In_286,In_546);
nor U358 (N_358,In_35,In_527);
or U359 (N_359,In_492,In_399);
nand U360 (N_360,In_223,In_423);
nand U361 (N_361,In_755,In_450);
nand U362 (N_362,In_646,In_80);
or U363 (N_363,In_341,In_114);
nand U364 (N_364,In_852,In_877);
and U365 (N_365,In_876,In_608);
or U366 (N_366,In_277,In_663);
and U367 (N_367,In_372,In_224);
xor U368 (N_368,In_4,In_834);
nor U369 (N_369,In_410,In_921);
nor U370 (N_370,In_182,In_314);
or U371 (N_371,In_19,In_804);
or U372 (N_372,In_407,In_281);
nand U373 (N_373,In_33,In_451);
and U374 (N_374,In_593,In_297);
or U375 (N_375,In_25,In_937);
or U376 (N_376,In_681,In_381);
nand U377 (N_377,In_421,In_655);
nor U378 (N_378,In_594,In_958);
or U379 (N_379,In_368,In_844);
or U380 (N_380,In_90,In_382);
nand U381 (N_381,In_924,In_940);
nor U382 (N_382,In_336,In_184);
and U383 (N_383,In_118,In_353);
nand U384 (N_384,In_361,In_391);
and U385 (N_385,In_778,In_595);
nand U386 (N_386,In_706,In_786);
nand U387 (N_387,In_388,In_156);
or U388 (N_388,In_742,In_244);
and U389 (N_389,In_822,In_553);
and U390 (N_390,In_584,In_32);
nor U391 (N_391,In_582,In_262);
or U392 (N_392,In_409,In_116);
and U393 (N_393,In_11,In_57);
nand U394 (N_394,In_919,In_180);
xor U395 (N_395,In_697,In_435);
or U396 (N_396,In_93,In_785);
nand U397 (N_397,In_698,In_208);
nand U398 (N_398,In_628,In_867);
nor U399 (N_399,In_79,In_26);
and U400 (N_400,In_255,In_516);
nor U401 (N_401,In_428,In_356);
nand U402 (N_402,In_972,In_338);
nor U403 (N_403,In_979,In_425);
nand U404 (N_404,In_563,In_928);
nor U405 (N_405,In_489,In_1);
or U406 (N_406,In_202,In_745);
or U407 (N_407,In_323,In_107);
nand U408 (N_408,In_102,In_639);
nor U409 (N_409,In_572,In_454);
nand U410 (N_410,In_953,In_843);
nor U411 (N_411,In_357,In_175);
and U412 (N_412,In_344,In_485);
and U413 (N_413,In_446,In_879);
or U414 (N_414,In_991,In_38);
nor U415 (N_415,In_789,In_827);
nand U416 (N_416,In_438,In_938);
nand U417 (N_417,In_270,In_146);
and U418 (N_418,In_767,In_358);
nand U419 (N_419,In_205,In_521);
nand U420 (N_420,In_759,In_841);
nor U421 (N_421,In_550,In_774);
or U422 (N_422,In_748,In_342);
and U423 (N_423,In_975,In_264);
or U424 (N_424,In_110,In_674);
nor U425 (N_425,In_465,In_522);
nor U426 (N_426,In_988,In_329);
nand U427 (N_427,In_199,In_383);
nor U428 (N_428,In_5,In_293);
nor U429 (N_429,In_951,In_3);
nor U430 (N_430,In_355,In_886);
nand U431 (N_431,In_401,In_447);
nor U432 (N_432,In_765,In_241);
nor U433 (N_433,In_499,In_43);
and U434 (N_434,In_588,In_140);
and U435 (N_435,In_279,In_869);
nand U436 (N_436,In_560,In_690);
nand U437 (N_437,In_9,In_661);
nand U438 (N_438,In_883,In_980);
nor U439 (N_439,In_995,In_601);
nor U440 (N_440,In_138,In_537);
xnor U441 (N_441,In_543,In_737);
and U442 (N_442,In_580,In_29);
and U443 (N_443,In_55,In_235);
and U444 (N_444,In_945,In_337);
and U445 (N_445,In_729,In_704);
nor U446 (N_446,In_707,In_860);
and U447 (N_447,In_967,In_50);
or U448 (N_448,In_13,In_67);
nor U449 (N_449,In_160,In_196);
nand U450 (N_450,In_978,In_59);
nor U451 (N_451,In_981,In_573);
and U452 (N_452,In_985,In_389);
or U453 (N_453,In_997,In_769);
or U454 (N_454,In_306,In_781);
xor U455 (N_455,In_345,In_807);
and U456 (N_456,In_738,In_319);
nand U457 (N_457,In_374,In_98);
nor U458 (N_458,In_155,In_408);
and U459 (N_459,In_121,In_609);
nor U460 (N_460,In_283,In_744);
or U461 (N_461,In_295,In_717);
or U462 (N_462,In_251,In_72);
nand U463 (N_463,In_15,In_968);
or U464 (N_464,In_210,In_185);
and U465 (N_465,In_482,In_45);
nor U466 (N_466,In_915,In_484);
nand U467 (N_467,In_225,In_229);
or U468 (N_468,In_113,In_367);
or U469 (N_469,In_621,In_587);
and U470 (N_470,In_129,In_302);
nand U471 (N_471,In_772,In_567);
and U472 (N_472,In_566,In_998);
or U473 (N_473,In_173,In_63);
nand U474 (N_474,In_112,In_413);
nor U475 (N_475,In_677,In_106);
nor U476 (N_476,In_728,In_312);
nand U477 (N_477,In_888,In_39);
nand U478 (N_478,In_27,In_506);
or U479 (N_479,In_890,In_135);
and U480 (N_480,In_74,In_48);
nand U481 (N_481,In_490,In_653);
and U482 (N_482,In_622,In_688);
nand U483 (N_483,In_905,In_545);
or U484 (N_484,In_89,In_741);
nand U485 (N_485,In_904,In_764);
and U486 (N_486,In_531,In_248);
nand U487 (N_487,In_682,In_289);
nand U488 (N_488,In_874,In_479);
nand U489 (N_489,In_526,In_348);
nand U490 (N_490,In_152,In_795);
nand U491 (N_491,In_908,In_575);
nor U492 (N_492,In_397,In_773);
or U493 (N_493,In_392,In_701);
nand U494 (N_494,In_296,In_440);
and U495 (N_495,In_610,In_299);
or U496 (N_496,In_548,In_8);
and U497 (N_497,In_966,In_683);
nand U498 (N_498,In_493,In_445);
or U499 (N_499,In_491,In_316);
nand U500 (N_500,In_109,In_606);
nand U501 (N_501,In_19,In_669);
nor U502 (N_502,In_459,In_643);
and U503 (N_503,In_171,In_451);
nor U504 (N_504,In_141,In_803);
or U505 (N_505,In_422,In_802);
and U506 (N_506,In_25,In_665);
nor U507 (N_507,In_786,In_724);
nor U508 (N_508,In_164,In_21);
nor U509 (N_509,In_320,In_67);
or U510 (N_510,In_953,In_521);
nand U511 (N_511,In_234,In_482);
nand U512 (N_512,In_957,In_915);
or U513 (N_513,In_84,In_942);
and U514 (N_514,In_347,In_288);
or U515 (N_515,In_855,In_868);
and U516 (N_516,In_383,In_985);
nand U517 (N_517,In_23,In_785);
or U518 (N_518,In_695,In_878);
nand U519 (N_519,In_673,In_504);
nor U520 (N_520,In_509,In_32);
nand U521 (N_521,In_342,In_325);
and U522 (N_522,In_608,In_563);
nor U523 (N_523,In_253,In_324);
or U524 (N_524,In_745,In_703);
nor U525 (N_525,In_415,In_243);
nor U526 (N_526,In_858,In_807);
or U527 (N_527,In_548,In_33);
and U528 (N_528,In_222,In_880);
and U529 (N_529,In_395,In_786);
or U530 (N_530,In_719,In_813);
nand U531 (N_531,In_423,In_771);
nand U532 (N_532,In_522,In_766);
nor U533 (N_533,In_209,In_267);
or U534 (N_534,In_889,In_434);
nand U535 (N_535,In_415,In_822);
or U536 (N_536,In_134,In_49);
nand U537 (N_537,In_550,In_991);
nand U538 (N_538,In_5,In_239);
and U539 (N_539,In_498,In_8);
or U540 (N_540,In_91,In_553);
nand U541 (N_541,In_119,In_90);
and U542 (N_542,In_350,In_554);
or U543 (N_543,In_914,In_668);
or U544 (N_544,In_272,In_247);
or U545 (N_545,In_680,In_555);
nor U546 (N_546,In_227,In_697);
nor U547 (N_547,In_2,In_587);
or U548 (N_548,In_561,In_115);
nand U549 (N_549,In_783,In_380);
and U550 (N_550,In_348,In_482);
nor U551 (N_551,In_728,In_795);
nor U552 (N_552,In_649,In_298);
nor U553 (N_553,In_118,In_567);
or U554 (N_554,In_597,In_780);
nand U555 (N_555,In_378,In_704);
nor U556 (N_556,In_403,In_893);
or U557 (N_557,In_860,In_148);
nor U558 (N_558,In_347,In_858);
and U559 (N_559,In_775,In_628);
nand U560 (N_560,In_956,In_333);
and U561 (N_561,In_755,In_684);
or U562 (N_562,In_912,In_204);
or U563 (N_563,In_292,In_30);
nor U564 (N_564,In_608,In_830);
and U565 (N_565,In_592,In_576);
nor U566 (N_566,In_408,In_22);
nor U567 (N_567,In_131,In_713);
or U568 (N_568,In_276,In_903);
and U569 (N_569,In_621,In_471);
and U570 (N_570,In_3,In_962);
nor U571 (N_571,In_714,In_840);
nor U572 (N_572,In_342,In_538);
or U573 (N_573,In_945,In_482);
nand U574 (N_574,In_750,In_997);
or U575 (N_575,In_264,In_840);
nand U576 (N_576,In_853,In_803);
nor U577 (N_577,In_475,In_89);
nand U578 (N_578,In_120,In_435);
nand U579 (N_579,In_153,In_596);
nand U580 (N_580,In_279,In_844);
or U581 (N_581,In_512,In_649);
or U582 (N_582,In_940,In_800);
nand U583 (N_583,In_23,In_222);
nor U584 (N_584,In_224,In_594);
and U585 (N_585,In_747,In_575);
nor U586 (N_586,In_580,In_969);
nand U587 (N_587,In_905,In_234);
nand U588 (N_588,In_305,In_958);
xnor U589 (N_589,In_580,In_784);
and U590 (N_590,In_392,In_913);
nor U591 (N_591,In_157,In_822);
and U592 (N_592,In_513,In_223);
nor U593 (N_593,In_459,In_412);
or U594 (N_594,In_989,In_223);
or U595 (N_595,In_677,In_93);
and U596 (N_596,In_593,In_304);
nand U597 (N_597,In_931,In_22);
or U598 (N_598,In_135,In_130);
or U599 (N_599,In_659,In_585);
or U600 (N_600,In_189,In_334);
or U601 (N_601,In_161,In_663);
nor U602 (N_602,In_609,In_647);
and U603 (N_603,In_991,In_136);
or U604 (N_604,In_699,In_606);
and U605 (N_605,In_137,In_364);
nor U606 (N_606,In_848,In_43);
nand U607 (N_607,In_803,In_548);
nand U608 (N_608,In_990,In_502);
nor U609 (N_609,In_710,In_152);
nand U610 (N_610,In_527,In_53);
nor U611 (N_611,In_777,In_824);
and U612 (N_612,In_10,In_107);
or U613 (N_613,In_56,In_330);
nor U614 (N_614,In_963,In_549);
or U615 (N_615,In_306,In_448);
nor U616 (N_616,In_530,In_133);
and U617 (N_617,In_51,In_256);
or U618 (N_618,In_376,In_690);
nand U619 (N_619,In_4,In_196);
or U620 (N_620,In_301,In_189);
nand U621 (N_621,In_286,In_851);
and U622 (N_622,In_526,In_874);
nor U623 (N_623,In_325,In_574);
or U624 (N_624,In_320,In_58);
or U625 (N_625,In_803,In_362);
and U626 (N_626,In_611,In_150);
nand U627 (N_627,In_704,In_756);
nand U628 (N_628,In_953,In_719);
nand U629 (N_629,In_46,In_798);
nor U630 (N_630,In_761,In_509);
nor U631 (N_631,In_692,In_589);
and U632 (N_632,In_385,In_157);
and U633 (N_633,In_689,In_566);
or U634 (N_634,In_464,In_305);
and U635 (N_635,In_376,In_767);
nor U636 (N_636,In_943,In_0);
or U637 (N_637,In_169,In_259);
nor U638 (N_638,In_133,In_982);
or U639 (N_639,In_793,In_348);
or U640 (N_640,In_819,In_387);
or U641 (N_641,In_644,In_913);
and U642 (N_642,In_876,In_771);
nand U643 (N_643,In_986,In_663);
or U644 (N_644,In_986,In_695);
nor U645 (N_645,In_821,In_516);
nor U646 (N_646,In_764,In_43);
nor U647 (N_647,In_372,In_280);
and U648 (N_648,In_722,In_327);
nor U649 (N_649,In_171,In_346);
and U650 (N_650,In_492,In_199);
or U651 (N_651,In_774,In_984);
nand U652 (N_652,In_404,In_860);
or U653 (N_653,In_14,In_118);
or U654 (N_654,In_234,In_126);
nand U655 (N_655,In_549,In_0);
and U656 (N_656,In_304,In_557);
nor U657 (N_657,In_871,In_314);
or U658 (N_658,In_397,In_950);
or U659 (N_659,In_633,In_443);
nor U660 (N_660,In_699,In_903);
nand U661 (N_661,In_55,In_881);
and U662 (N_662,In_562,In_824);
nor U663 (N_663,In_862,In_441);
nand U664 (N_664,In_4,In_760);
or U665 (N_665,In_983,In_74);
or U666 (N_666,In_139,In_691);
nor U667 (N_667,In_773,In_301);
or U668 (N_668,In_230,In_311);
and U669 (N_669,In_69,In_563);
nor U670 (N_670,In_196,In_591);
or U671 (N_671,In_674,In_990);
and U672 (N_672,In_309,In_287);
or U673 (N_673,In_575,In_231);
nor U674 (N_674,In_96,In_122);
nor U675 (N_675,In_603,In_729);
nor U676 (N_676,In_243,In_596);
and U677 (N_677,In_743,In_186);
and U678 (N_678,In_21,In_852);
and U679 (N_679,In_812,In_868);
nand U680 (N_680,In_158,In_505);
and U681 (N_681,In_104,In_666);
nor U682 (N_682,In_738,In_199);
nor U683 (N_683,In_509,In_441);
nand U684 (N_684,In_733,In_906);
nand U685 (N_685,In_493,In_913);
nand U686 (N_686,In_453,In_114);
nor U687 (N_687,In_679,In_510);
or U688 (N_688,In_354,In_234);
nand U689 (N_689,In_602,In_944);
nor U690 (N_690,In_842,In_945);
and U691 (N_691,In_331,In_551);
nor U692 (N_692,In_239,In_244);
nand U693 (N_693,In_666,In_28);
or U694 (N_694,In_62,In_409);
or U695 (N_695,In_311,In_944);
and U696 (N_696,In_479,In_10);
nand U697 (N_697,In_247,In_112);
and U698 (N_698,In_634,In_22);
nand U699 (N_699,In_963,In_523);
nand U700 (N_700,In_145,In_228);
nand U701 (N_701,In_340,In_850);
nand U702 (N_702,In_100,In_647);
and U703 (N_703,In_46,In_71);
and U704 (N_704,In_427,In_829);
or U705 (N_705,In_936,In_682);
nor U706 (N_706,In_155,In_259);
and U707 (N_707,In_707,In_642);
nor U708 (N_708,In_884,In_380);
nor U709 (N_709,In_618,In_221);
nand U710 (N_710,In_9,In_515);
or U711 (N_711,In_165,In_731);
nand U712 (N_712,In_701,In_794);
nor U713 (N_713,In_161,In_778);
and U714 (N_714,In_228,In_160);
nand U715 (N_715,In_776,In_720);
or U716 (N_716,In_199,In_846);
nand U717 (N_717,In_482,In_504);
nand U718 (N_718,In_472,In_439);
nand U719 (N_719,In_169,In_765);
and U720 (N_720,In_352,In_515);
nor U721 (N_721,In_594,In_661);
or U722 (N_722,In_897,In_822);
nor U723 (N_723,In_570,In_547);
nor U724 (N_724,In_849,In_285);
or U725 (N_725,In_332,In_722);
or U726 (N_726,In_236,In_233);
nor U727 (N_727,In_307,In_294);
nand U728 (N_728,In_600,In_444);
or U729 (N_729,In_869,In_25);
nand U730 (N_730,In_859,In_950);
nand U731 (N_731,In_84,In_33);
or U732 (N_732,In_726,In_461);
and U733 (N_733,In_854,In_609);
nor U734 (N_734,In_373,In_957);
and U735 (N_735,In_610,In_94);
and U736 (N_736,In_890,In_3);
and U737 (N_737,In_948,In_322);
nand U738 (N_738,In_674,In_719);
and U739 (N_739,In_51,In_203);
or U740 (N_740,In_865,In_316);
nor U741 (N_741,In_87,In_554);
nand U742 (N_742,In_813,In_792);
or U743 (N_743,In_883,In_930);
and U744 (N_744,In_774,In_367);
or U745 (N_745,In_489,In_43);
nor U746 (N_746,In_347,In_29);
nand U747 (N_747,In_764,In_390);
and U748 (N_748,In_0,In_691);
nand U749 (N_749,In_770,In_972);
nor U750 (N_750,In_635,In_381);
xnor U751 (N_751,In_304,In_383);
or U752 (N_752,In_709,In_23);
or U753 (N_753,In_0,In_562);
and U754 (N_754,In_836,In_986);
nor U755 (N_755,In_190,In_407);
or U756 (N_756,In_121,In_519);
nand U757 (N_757,In_68,In_995);
and U758 (N_758,In_265,In_604);
or U759 (N_759,In_4,In_642);
nand U760 (N_760,In_393,In_818);
or U761 (N_761,In_595,In_636);
or U762 (N_762,In_554,In_727);
nor U763 (N_763,In_280,In_968);
or U764 (N_764,In_156,In_244);
nand U765 (N_765,In_236,In_316);
or U766 (N_766,In_316,In_670);
nand U767 (N_767,In_893,In_86);
nand U768 (N_768,In_233,In_975);
and U769 (N_769,In_925,In_670);
nor U770 (N_770,In_664,In_438);
nor U771 (N_771,In_133,In_551);
nor U772 (N_772,In_64,In_45);
and U773 (N_773,In_245,In_266);
nor U774 (N_774,In_759,In_147);
nor U775 (N_775,In_200,In_959);
and U776 (N_776,In_639,In_666);
nand U777 (N_777,In_417,In_385);
or U778 (N_778,In_711,In_190);
nor U779 (N_779,In_115,In_126);
or U780 (N_780,In_912,In_488);
xnor U781 (N_781,In_686,In_825);
nand U782 (N_782,In_903,In_23);
nor U783 (N_783,In_793,In_67);
and U784 (N_784,In_257,In_851);
or U785 (N_785,In_106,In_957);
or U786 (N_786,In_695,In_630);
and U787 (N_787,In_116,In_819);
nor U788 (N_788,In_935,In_959);
or U789 (N_789,In_948,In_63);
nand U790 (N_790,In_958,In_206);
or U791 (N_791,In_639,In_771);
nor U792 (N_792,In_123,In_348);
nand U793 (N_793,In_528,In_270);
and U794 (N_794,In_630,In_532);
or U795 (N_795,In_952,In_313);
or U796 (N_796,In_35,In_896);
or U797 (N_797,In_265,In_675);
and U798 (N_798,In_176,In_503);
nand U799 (N_799,In_719,In_273);
nand U800 (N_800,In_737,In_722);
or U801 (N_801,In_266,In_288);
nand U802 (N_802,In_926,In_155);
and U803 (N_803,In_217,In_509);
nor U804 (N_804,In_262,In_408);
nor U805 (N_805,In_591,In_736);
and U806 (N_806,In_22,In_892);
and U807 (N_807,In_708,In_303);
or U808 (N_808,In_494,In_858);
nand U809 (N_809,In_154,In_607);
or U810 (N_810,In_41,In_982);
nor U811 (N_811,In_239,In_603);
and U812 (N_812,In_83,In_151);
or U813 (N_813,In_792,In_324);
and U814 (N_814,In_584,In_699);
and U815 (N_815,In_563,In_735);
nand U816 (N_816,In_344,In_998);
nand U817 (N_817,In_526,In_89);
nand U818 (N_818,In_561,In_280);
and U819 (N_819,In_172,In_709);
nand U820 (N_820,In_216,In_537);
or U821 (N_821,In_678,In_702);
nand U822 (N_822,In_913,In_281);
nand U823 (N_823,In_530,In_935);
or U824 (N_824,In_441,In_832);
and U825 (N_825,In_647,In_539);
nand U826 (N_826,In_538,In_323);
nor U827 (N_827,In_924,In_464);
nand U828 (N_828,In_833,In_152);
and U829 (N_829,In_705,In_131);
nor U830 (N_830,In_921,In_978);
nor U831 (N_831,In_626,In_772);
and U832 (N_832,In_809,In_75);
or U833 (N_833,In_692,In_97);
nand U834 (N_834,In_47,In_343);
nand U835 (N_835,In_942,In_711);
or U836 (N_836,In_544,In_109);
and U837 (N_837,In_953,In_750);
and U838 (N_838,In_915,In_256);
or U839 (N_839,In_268,In_62);
nor U840 (N_840,In_211,In_908);
nor U841 (N_841,In_978,In_540);
nand U842 (N_842,In_519,In_906);
nand U843 (N_843,In_12,In_347);
nand U844 (N_844,In_438,In_172);
and U845 (N_845,In_480,In_974);
nand U846 (N_846,In_345,In_310);
and U847 (N_847,In_625,In_839);
or U848 (N_848,In_298,In_950);
and U849 (N_849,In_384,In_282);
nor U850 (N_850,In_660,In_822);
and U851 (N_851,In_410,In_402);
nand U852 (N_852,In_946,In_747);
nand U853 (N_853,In_719,In_793);
nor U854 (N_854,In_233,In_959);
nand U855 (N_855,In_804,In_461);
nor U856 (N_856,In_979,In_451);
and U857 (N_857,In_957,In_594);
nor U858 (N_858,In_987,In_51);
nor U859 (N_859,In_807,In_857);
nand U860 (N_860,In_439,In_742);
nand U861 (N_861,In_974,In_247);
and U862 (N_862,In_207,In_726);
or U863 (N_863,In_9,In_891);
nand U864 (N_864,In_526,In_98);
or U865 (N_865,In_324,In_119);
nand U866 (N_866,In_763,In_45);
or U867 (N_867,In_248,In_862);
nor U868 (N_868,In_245,In_430);
xnor U869 (N_869,In_292,In_103);
and U870 (N_870,In_767,In_514);
or U871 (N_871,In_935,In_904);
or U872 (N_872,In_762,In_694);
nor U873 (N_873,In_832,In_823);
or U874 (N_874,In_322,In_223);
xor U875 (N_875,In_181,In_765);
nand U876 (N_876,In_322,In_520);
and U877 (N_877,In_436,In_834);
and U878 (N_878,In_211,In_251);
nor U879 (N_879,In_800,In_460);
nor U880 (N_880,In_680,In_735);
or U881 (N_881,In_469,In_334);
or U882 (N_882,In_293,In_284);
nor U883 (N_883,In_853,In_647);
nand U884 (N_884,In_567,In_494);
nor U885 (N_885,In_183,In_710);
nor U886 (N_886,In_88,In_547);
and U887 (N_887,In_225,In_265);
nand U888 (N_888,In_450,In_301);
nand U889 (N_889,In_764,In_145);
nand U890 (N_890,In_467,In_447);
or U891 (N_891,In_320,In_45);
nand U892 (N_892,In_228,In_144);
nor U893 (N_893,In_929,In_182);
and U894 (N_894,In_744,In_181);
and U895 (N_895,In_591,In_36);
nand U896 (N_896,In_93,In_85);
or U897 (N_897,In_568,In_248);
or U898 (N_898,In_40,In_421);
or U899 (N_899,In_333,In_719);
nor U900 (N_900,In_900,In_455);
nand U901 (N_901,In_151,In_533);
nor U902 (N_902,In_317,In_876);
nand U903 (N_903,In_290,In_1);
and U904 (N_904,In_924,In_779);
or U905 (N_905,In_208,In_61);
and U906 (N_906,In_692,In_622);
nor U907 (N_907,In_151,In_939);
and U908 (N_908,In_702,In_455);
or U909 (N_909,In_532,In_170);
or U910 (N_910,In_100,In_779);
and U911 (N_911,In_633,In_915);
nand U912 (N_912,In_254,In_900);
and U913 (N_913,In_559,In_602);
or U914 (N_914,In_106,In_371);
or U915 (N_915,In_702,In_948);
or U916 (N_916,In_103,In_845);
and U917 (N_917,In_868,In_275);
nand U918 (N_918,In_665,In_715);
nor U919 (N_919,In_794,In_999);
or U920 (N_920,In_773,In_457);
or U921 (N_921,In_237,In_393);
and U922 (N_922,In_242,In_738);
or U923 (N_923,In_293,In_645);
and U924 (N_924,In_143,In_524);
or U925 (N_925,In_65,In_122);
nor U926 (N_926,In_613,In_994);
or U927 (N_927,In_779,In_585);
and U928 (N_928,In_901,In_865);
nand U929 (N_929,In_676,In_56);
nor U930 (N_930,In_296,In_95);
nand U931 (N_931,In_330,In_793);
nand U932 (N_932,In_669,In_93);
nor U933 (N_933,In_80,In_19);
nand U934 (N_934,In_84,In_529);
nand U935 (N_935,In_539,In_238);
nand U936 (N_936,In_238,In_250);
nor U937 (N_937,In_597,In_376);
nand U938 (N_938,In_332,In_95);
nor U939 (N_939,In_934,In_14);
nor U940 (N_940,In_207,In_547);
nand U941 (N_941,In_879,In_231);
or U942 (N_942,In_596,In_73);
and U943 (N_943,In_28,In_59);
or U944 (N_944,In_194,In_427);
and U945 (N_945,In_865,In_915);
nor U946 (N_946,In_891,In_510);
nor U947 (N_947,In_749,In_564);
or U948 (N_948,In_225,In_631);
or U949 (N_949,In_816,In_701);
or U950 (N_950,In_150,In_675);
nand U951 (N_951,In_457,In_408);
nand U952 (N_952,In_776,In_911);
nor U953 (N_953,In_891,In_915);
nor U954 (N_954,In_46,In_973);
and U955 (N_955,In_208,In_748);
nor U956 (N_956,In_891,In_286);
nand U957 (N_957,In_189,In_948);
or U958 (N_958,In_283,In_540);
and U959 (N_959,In_999,In_690);
nor U960 (N_960,In_106,In_743);
nor U961 (N_961,In_470,In_710);
and U962 (N_962,In_245,In_720);
nand U963 (N_963,In_249,In_845);
nor U964 (N_964,In_542,In_499);
or U965 (N_965,In_422,In_669);
nand U966 (N_966,In_460,In_6);
nand U967 (N_967,In_341,In_591);
nand U968 (N_968,In_801,In_41);
nand U969 (N_969,In_425,In_687);
nor U970 (N_970,In_250,In_351);
and U971 (N_971,In_365,In_703);
nor U972 (N_972,In_180,In_244);
nand U973 (N_973,In_871,In_49);
and U974 (N_974,In_445,In_988);
nand U975 (N_975,In_240,In_744);
nand U976 (N_976,In_405,In_24);
nor U977 (N_977,In_318,In_455);
xor U978 (N_978,In_449,In_983);
and U979 (N_979,In_996,In_516);
and U980 (N_980,In_593,In_152);
and U981 (N_981,In_63,In_650);
or U982 (N_982,In_28,In_874);
nand U983 (N_983,In_235,In_124);
nor U984 (N_984,In_39,In_899);
and U985 (N_985,In_239,In_294);
nand U986 (N_986,In_812,In_715);
nand U987 (N_987,In_505,In_103);
or U988 (N_988,In_418,In_479);
and U989 (N_989,In_704,In_648);
nand U990 (N_990,In_897,In_474);
nor U991 (N_991,In_192,In_863);
or U992 (N_992,In_52,In_362);
nand U993 (N_993,In_848,In_534);
and U994 (N_994,In_467,In_193);
nand U995 (N_995,In_68,In_893);
nand U996 (N_996,In_260,In_898);
xnor U997 (N_997,In_928,In_182);
or U998 (N_998,In_484,In_297);
nor U999 (N_999,In_992,In_795);
and U1000 (N_1000,In_623,In_244);
nor U1001 (N_1001,In_335,In_204);
nor U1002 (N_1002,In_784,In_66);
nand U1003 (N_1003,In_891,In_574);
nand U1004 (N_1004,In_716,In_127);
nand U1005 (N_1005,In_876,In_526);
or U1006 (N_1006,In_938,In_735);
nand U1007 (N_1007,In_4,In_576);
and U1008 (N_1008,In_506,In_571);
nand U1009 (N_1009,In_531,In_753);
nor U1010 (N_1010,In_894,In_806);
or U1011 (N_1011,In_530,In_494);
and U1012 (N_1012,In_360,In_279);
nor U1013 (N_1013,In_950,In_79);
nand U1014 (N_1014,In_928,In_469);
nor U1015 (N_1015,In_660,In_704);
and U1016 (N_1016,In_537,In_151);
or U1017 (N_1017,In_617,In_603);
nor U1018 (N_1018,In_659,In_600);
or U1019 (N_1019,In_776,In_297);
or U1020 (N_1020,In_302,In_989);
or U1021 (N_1021,In_168,In_119);
nand U1022 (N_1022,In_440,In_612);
and U1023 (N_1023,In_466,In_225);
and U1024 (N_1024,In_7,In_547);
nand U1025 (N_1025,In_265,In_879);
nand U1026 (N_1026,In_441,In_965);
nor U1027 (N_1027,In_683,In_635);
or U1028 (N_1028,In_216,In_282);
nand U1029 (N_1029,In_611,In_641);
and U1030 (N_1030,In_86,In_749);
or U1031 (N_1031,In_735,In_454);
nand U1032 (N_1032,In_988,In_517);
nand U1033 (N_1033,In_586,In_917);
nand U1034 (N_1034,In_230,In_250);
or U1035 (N_1035,In_940,In_663);
and U1036 (N_1036,In_740,In_317);
and U1037 (N_1037,In_324,In_246);
or U1038 (N_1038,In_739,In_451);
nand U1039 (N_1039,In_902,In_756);
and U1040 (N_1040,In_141,In_839);
and U1041 (N_1041,In_699,In_844);
nand U1042 (N_1042,In_766,In_122);
nor U1043 (N_1043,In_106,In_532);
nand U1044 (N_1044,In_381,In_60);
nor U1045 (N_1045,In_290,In_749);
and U1046 (N_1046,In_828,In_882);
nor U1047 (N_1047,In_350,In_634);
nor U1048 (N_1048,In_66,In_689);
nor U1049 (N_1049,In_117,In_931);
or U1050 (N_1050,In_280,In_712);
xnor U1051 (N_1051,In_16,In_718);
or U1052 (N_1052,In_915,In_284);
and U1053 (N_1053,In_163,In_0);
xor U1054 (N_1054,In_803,In_454);
nor U1055 (N_1055,In_428,In_313);
or U1056 (N_1056,In_932,In_489);
or U1057 (N_1057,In_982,In_589);
nor U1058 (N_1058,In_328,In_460);
nand U1059 (N_1059,In_300,In_43);
nand U1060 (N_1060,In_985,In_915);
or U1061 (N_1061,In_818,In_745);
nand U1062 (N_1062,In_549,In_620);
nor U1063 (N_1063,In_382,In_31);
and U1064 (N_1064,In_234,In_810);
and U1065 (N_1065,In_802,In_403);
nor U1066 (N_1066,In_712,In_197);
nand U1067 (N_1067,In_159,In_799);
or U1068 (N_1068,In_457,In_567);
or U1069 (N_1069,In_680,In_475);
and U1070 (N_1070,In_811,In_332);
or U1071 (N_1071,In_471,In_911);
and U1072 (N_1072,In_375,In_184);
and U1073 (N_1073,In_888,In_100);
and U1074 (N_1074,In_117,In_834);
nand U1075 (N_1075,In_129,In_343);
nor U1076 (N_1076,In_695,In_245);
nor U1077 (N_1077,In_512,In_391);
and U1078 (N_1078,In_239,In_854);
and U1079 (N_1079,In_417,In_698);
and U1080 (N_1080,In_716,In_382);
nor U1081 (N_1081,In_382,In_718);
or U1082 (N_1082,In_426,In_628);
or U1083 (N_1083,In_445,In_791);
nor U1084 (N_1084,In_216,In_340);
nand U1085 (N_1085,In_372,In_667);
nor U1086 (N_1086,In_514,In_487);
nor U1087 (N_1087,In_13,In_786);
nor U1088 (N_1088,In_885,In_225);
and U1089 (N_1089,In_427,In_353);
nand U1090 (N_1090,In_771,In_486);
and U1091 (N_1091,In_306,In_470);
or U1092 (N_1092,In_486,In_389);
nand U1093 (N_1093,In_53,In_664);
nand U1094 (N_1094,In_745,In_724);
or U1095 (N_1095,In_361,In_937);
or U1096 (N_1096,In_663,In_853);
nand U1097 (N_1097,In_739,In_971);
and U1098 (N_1098,In_674,In_770);
nand U1099 (N_1099,In_175,In_618);
or U1100 (N_1100,In_617,In_84);
nor U1101 (N_1101,In_217,In_632);
and U1102 (N_1102,In_392,In_627);
or U1103 (N_1103,In_793,In_851);
and U1104 (N_1104,In_788,In_443);
nor U1105 (N_1105,In_98,In_516);
xor U1106 (N_1106,In_705,In_100);
nor U1107 (N_1107,In_804,In_48);
and U1108 (N_1108,In_876,In_944);
nor U1109 (N_1109,In_324,In_809);
or U1110 (N_1110,In_725,In_541);
nor U1111 (N_1111,In_995,In_586);
or U1112 (N_1112,In_930,In_831);
or U1113 (N_1113,In_32,In_315);
nor U1114 (N_1114,In_271,In_672);
nand U1115 (N_1115,In_443,In_928);
nor U1116 (N_1116,In_267,In_810);
and U1117 (N_1117,In_41,In_961);
and U1118 (N_1118,In_982,In_706);
and U1119 (N_1119,In_808,In_917);
nand U1120 (N_1120,In_662,In_937);
and U1121 (N_1121,In_704,In_300);
nor U1122 (N_1122,In_418,In_263);
nor U1123 (N_1123,In_116,In_875);
and U1124 (N_1124,In_425,In_964);
nand U1125 (N_1125,In_522,In_955);
or U1126 (N_1126,In_365,In_746);
nor U1127 (N_1127,In_905,In_34);
and U1128 (N_1128,In_332,In_894);
nand U1129 (N_1129,In_657,In_475);
nor U1130 (N_1130,In_352,In_356);
and U1131 (N_1131,In_156,In_657);
and U1132 (N_1132,In_700,In_695);
nand U1133 (N_1133,In_681,In_551);
nor U1134 (N_1134,In_779,In_104);
and U1135 (N_1135,In_99,In_336);
and U1136 (N_1136,In_376,In_483);
nor U1137 (N_1137,In_22,In_840);
nand U1138 (N_1138,In_948,In_610);
nand U1139 (N_1139,In_161,In_800);
or U1140 (N_1140,In_305,In_144);
and U1141 (N_1141,In_69,In_107);
nand U1142 (N_1142,In_299,In_948);
nand U1143 (N_1143,In_670,In_575);
and U1144 (N_1144,In_275,In_899);
nor U1145 (N_1145,In_666,In_577);
or U1146 (N_1146,In_379,In_343);
and U1147 (N_1147,In_42,In_150);
nor U1148 (N_1148,In_753,In_932);
nand U1149 (N_1149,In_736,In_824);
or U1150 (N_1150,In_323,In_851);
nor U1151 (N_1151,In_840,In_891);
and U1152 (N_1152,In_396,In_679);
or U1153 (N_1153,In_663,In_74);
or U1154 (N_1154,In_163,In_831);
or U1155 (N_1155,In_843,In_628);
or U1156 (N_1156,In_198,In_329);
or U1157 (N_1157,In_365,In_932);
nand U1158 (N_1158,In_748,In_327);
or U1159 (N_1159,In_144,In_374);
nand U1160 (N_1160,In_105,In_473);
and U1161 (N_1161,In_314,In_283);
and U1162 (N_1162,In_343,In_800);
or U1163 (N_1163,In_25,In_591);
nand U1164 (N_1164,In_616,In_933);
nand U1165 (N_1165,In_719,In_222);
and U1166 (N_1166,In_723,In_10);
nand U1167 (N_1167,In_584,In_799);
and U1168 (N_1168,In_260,In_966);
and U1169 (N_1169,In_933,In_458);
nor U1170 (N_1170,In_300,In_881);
or U1171 (N_1171,In_479,In_765);
or U1172 (N_1172,In_128,In_950);
and U1173 (N_1173,In_594,In_325);
or U1174 (N_1174,In_463,In_223);
nor U1175 (N_1175,In_739,In_678);
nand U1176 (N_1176,In_336,In_881);
or U1177 (N_1177,In_247,In_682);
nand U1178 (N_1178,In_19,In_556);
nor U1179 (N_1179,In_528,In_596);
or U1180 (N_1180,In_731,In_135);
and U1181 (N_1181,In_626,In_499);
or U1182 (N_1182,In_158,In_460);
or U1183 (N_1183,In_1,In_973);
nor U1184 (N_1184,In_444,In_953);
nor U1185 (N_1185,In_707,In_418);
nand U1186 (N_1186,In_169,In_691);
or U1187 (N_1187,In_389,In_861);
nor U1188 (N_1188,In_997,In_954);
nand U1189 (N_1189,In_415,In_33);
or U1190 (N_1190,In_567,In_163);
nand U1191 (N_1191,In_608,In_571);
nor U1192 (N_1192,In_66,In_816);
and U1193 (N_1193,In_462,In_106);
and U1194 (N_1194,In_226,In_524);
nand U1195 (N_1195,In_472,In_308);
or U1196 (N_1196,In_620,In_404);
nor U1197 (N_1197,In_873,In_336);
nand U1198 (N_1198,In_149,In_76);
and U1199 (N_1199,In_751,In_767);
or U1200 (N_1200,In_829,In_213);
or U1201 (N_1201,In_416,In_254);
nand U1202 (N_1202,In_592,In_474);
nand U1203 (N_1203,In_502,In_900);
and U1204 (N_1204,In_164,In_184);
nor U1205 (N_1205,In_298,In_343);
or U1206 (N_1206,In_405,In_530);
nand U1207 (N_1207,In_90,In_185);
or U1208 (N_1208,In_451,In_15);
and U1209 (N_1209,In_222,In_560);
nor U1210 (N_1210,In_718,In_240);
and U1211 (N_1211,In_79,In_391);
or U1212 (N_1212,In_430,In_202);
or U1213 (N_1213,In_868,In_11);
nand U1214 (N_1214,In_810,In_263);
or U1215 (N_1215,In_607,In_786);
or U1216 (N_1216,In_189,In_390);
or U1217 (N_1217,In_674,In_219);
nand U1218 (N_1218,In_953,In_786);
and U1219 (N_1219,In_116,In_356);
and U1220 (N_1220,In_113,In_924);
nand U1221 (N_1221,In_667,In_646);
nand U1222 (N_1222,In_388,In_750);
nor U1223 (N_1223,In_945,In_119);
nand U1224 (N_1224,In_330,In_986);
or U1225 (N_1225,In_110,In_802);
or U1226 (N_1226,In_444,In_9);
or U1227 (N_1227,In_82,In_445);
or U1228 (N_1228,In_204,In_760);
nand U1229 (N_1229,In_329,In_943);
nand U1230 (N_1230,In_774,In_757);
nor U1231 (N_1231,In_416,In_226);
and U1232 (N_1232,In_582,In_55);
and U1233 (N_1233,In_990,In_474);
and U1234 (N_1234,In_208,In_994);
and U1235 (N_1235,In_28,In_677);
and U1236 (N_1236,In_732,In_285);
nand U1237 (N_1237,In_246,In_877);
nand U1238 (N_1238,In_147,In_500);
or U1239 (N_1239,In_47,In_978);
and U1240 (N_1240,In_968,In_162);
and U1241 (N_1241,In_523,In_21);
and U1242 (N_1242,In_498,In_806);
nand U1243 (N_1243,In_29,In_445);
xnor U1244 (N_1244,In_630,In_984);
nand U1245 (N_1245,In_304,In_255);
and U1246 (N_1246,In_239,In_208);
nand U1247 (N_1247,In_981,In_346);
nand U1248 (N_1248,In_557,In_387);
nand U1249 (N_1249,In_874,In_264);
nor U1250 (N_1250,In_163,In_614);
nand U1251 (N_1251,In_739,In_19);
or U1252 (N_1252,In_963,In_52);
or U1253 (N_1253,In_1,In_564);
nand U1254 (N_1254,In_729,In_280);
nor U1255 (N_1255,In_659,In_551);
and U1256 (N_1256,In_974,In_335);
and U1257 (N_1257,In_997,In_502);
or U1258 (N_1258,In_924,In_118);
nand U1259 (N_1259,In_751,In_451);
nor U1260 (N_1260,In_370,In_299);
nand U1261 (N_1261,In_176,In_472);
nand U1262 (N_1262,In_257,In_675);
nor U1263 (N_1263,In_254,In_259);
nor U1264 (N_1264,In_107,In_506);
and U1265 (N_1265,In_521,In_568);
nor U1266 (N_1266,In_585,In_957);
or U1267 (N_1267,In_190,In_801);
nor U1268 (N_1268,In_902,In_243);
nor U1269 (N_1269,In_875,In_79);
and U1270 (N_1270,In_890,In_514);
and U1271 (N_1271,In_810,In_37);
and U1272 (N_1272,In_620,In_743);
nor U1273 (N_1273,In_313,In_321);
or U1274 (N_1274,In_907,In_67);
and U1275 (N_1275,In_856,In_391);
nand U1276 (N_1276,In_231,In_936);
nand U1277 (N_1277,In_754,In_554);
or U1278 (N_1278,In_380,In_892);
or U1279 (N_1279,In_80,In_569);
and U1280 (N_1280,In_387,In_293);
nor U1281 (N_1281,In_65,In_332);
nor U1282 (N_1282,In_116,In_73);
nand U1283 (N_1283,In_415,In_341);
nor U1284 (N_1284,In_763,In_355);
or U1285 (N_1285,In_284,In_622);
nor U1286 (N_1286,In_428,In_7);
and U1287 (N_1287,In_174,In_973);
nand U1288 (N_1288,In_191,In_998);
or U1289 (N_1289,In_300,In_808);
and U1290 (N_1290,In_157,In_620);
nor U1291 (N_1291,In_531,In_752);
or U1292 (N_1292,In_829,In_287);
and U1293 (N_1293,In_634,In_540);
and U1294 (N_1294,In_911,In_570);
nand U1295 (N_1295,In_181,In_831);
nor U1296 (N_1296,In_199,In_435);
or U1297 (N_1297,In_136,In_943);
nand U1298 (N_1298,In_312,In_99);
nor U1299 (N_1299,In_545,In_623);
nor U1300 (N_1300,In_908,In_269);
or U1301 (N_1301,In_748,In_376);
and U1302 (N_1302,In_492,In_408);
or U1303 (N_1303,In_178,In_209);
nor U1304 (N_1304,In_577,In_467);
nand U1305 (N_1305,In_612,In_98);
or U1306 (N_1306,In_719,In_956);
nor U1307 (N_1307,In_688,In_209);
or U1308 (N_1308,In_464,In_71);
nand U1309 (N_1309,In_290,In_510);
nor U1310 (N_1310,In_794,In_159);
and U1311 (N_1311,In_551,In_579);
nand U1312 (N_1312,In_841,In_997);
or U1313 (N_1313,In_725,In_385);
or U1314 (N_1314,In_114,In_487);
nor U1315 (N_1315,In_773,In_532);
or U1316 (N_1316,In_203,In_109);
nand U1317 (N_1317,In_437,In_613);
or U1318 (N_1318,In_337,In_183);
and U1319 (N_1319,In_672,In_407);
xnor U1320 (N_1320,In_861,In_66);
nand U1321 (N_1321,In_36,In_47);
or U1322 (N_1322,In_43,In_880);
nor U1323 (N_1323,In_986,In_237);
nand U1324 (N_1324,In_648,In_836);
nor U1325 (N_1325,In_524,In_206);
nor U1326 (N_1326,In_696,In_484);
or U1327 (N_1327,In_149,In_317);
nand U1328 (N_1328,In_895,In_477);
or U1329 (N_1329,In_133,In_612);
nor U1330 (N_1330,In_483,In_514);
or U1331 (N_1331,In_104,In_471);
or U1332 (N_1332,In_615,In_439);
and U1333 (N_1333,In_5,In_220);
nor U1334 (N_1334,In_492,In_504);
and U1335 (N_1335,In_513,In_738);
or U1336 (N_1336,In_195,In_601);
nor U1337 (N_1337,In_872,In_653);
and U1338 (N_1338,In_430,In_815);
and U1339 (N_1339,In_609,In_76);
or U1340 (N_1340,In_635,In_943);
nor U1341 (N_1341,In_565,In_76);
or U1342 (N_1342,In_114,In_204);
nor U1343 (N_1343,In_764,In_86);
or U1344 (N_1344,In_39,In_40);
and U1345 (N_1345,In_891,In_449);
or U1346 (N_1346,In_812,In_645);
nor U1347 (N_1347,In_506,In_260);
or U1348 (N_1348,In_828,In_119);
and U1349 (N_1349,In_35,In_241);
nand U1350 (N_1350,In_990,In_651);
nand U1351 (N_1351,In_517,In_652);
or U1352 (N_1352,In_864,In_184);
and U1353 (N_1353,In_690,In_890);
and U1354 (N_1354,In_849,In_295);
or U1355 (N_1355,In_642,In_669);
nor U1356 (N_1356,In_667,In_805);
xor U1357 (N_1357,In_51,In_265);
nand U1358 (N_1358,In_771,In_963);
or U1359 (N_1359,In_599,In_666);
nand U1360 (N_1360,In_736,In_525);
nand U1361 (N_1361,In_422,In_133);
nor U1362 (N_1362,In_375,In_683);
and U1363 (N_1363,In_187,In_850);
nand U1364 (N_1364,In_206,In_925);
nand U1365 (N_1365,In_780,In_585);
and U1366 (N_1366,In_834,In_320);
nor U1367 (N_1367,In_203,In_20);
nor U1368 (N_1368,In_175,In_258);
or U1369 (N_1369,In_547,In_429);
nor U1370 (N_1370,In_276,In_986);
nor U1371 (N_1371,In_115,In_263);
or U1372 (N_1372,In_228,In_690);
nand U1373 (N_1373,In_246,In_372);
or U1374 (N_1374,In_128,In_105);
nor U1375 (N_1375,In_405,In_605);
or U1376 (N_1376,In_696,In_299);
nor U1377 (N_1377,In_42,In_820);
xnor U1378 (N_1378,In_242,In_697);
nor U1379 (N_1379,In_249,In_498);
or U1380 (N_1380,In_630,In_600);
or U1381 (N_1381,In_850,In_462);
nand U1382 (N_1382,In_57,In_281);
nor U1383 (N_1383,In_27,In_271);
nor U1384 (N_1384,In_757,In_352);
and U1385 (N_1385,In_540,In_964);
and U1386 (N_1386,In_177,In_315);
nand U1387 (N_1387,In_616,In_10);
or U1388 (N_1388,In_169,In_928);
nand U1389 (N_1389,In_837,In_754);
or U1390 (N_1390,In_436,In_858);
or U1391 (N_1391,In_512,In_39);
nand U1392 (N_1392,In_666,In_184);
or U1393 (N_1393,In_552,In_598);
nor U1394 (N_1394,In_462,In_879);
and U1395 (N_1395,In_477,In_202);
or U1396 (N_1396,In_277,In_622);
and U1397 (N_1397,In_958,In_14);
and U1398 (N_1398,In_692,In_112);
nand U1399 (N_1399,In_189,In_374);
nand U1400 (N_1400,In_338,In_989);
or U1401 (N_1401,In_908,In_698);
and U1402 (N_1402,In_281,In_837);
and U1403 (N_1403,In_404,In_664);
nor U1404 (N_1404,In_110,In_656);
and U1405 (N_1405,In_801,In_145);
or U1406 (N_1406,In_6,In_596);
and U1407 (N_1407,In_875,In_4);
nand U1408 (N_1408,In_941,In_493);
nand U1409 (N_1409,In_212,In_754);
nand U1410 (N_1410,In_584,In_852);
and U1411 (N_1411,In_107,In_753);
and U1412 (N_1412,In_273,In_204);
nor U1413 (N_1413,In_739,In_13);
nor U1414 (N_1414,In_514,In_113);
nor U1415 (N_1415,In_646,In_6);
nand U1416 (N_1416,In_222,In_351);
nand U1417 (N_1417,In_814,In_816);
nor U1418 (N_1418,In_672,In_746);
and U1419 (N_1419,In_13,In_846);
nand U1420 (N_1420,In_983,In_366);
nor U1421 (N_1421,In_269,In_506);
and U1422 (N_1422,In_942,In_563);
nand U1423 (N_1423,In_539,In_264);
nand U1424 (N_1424,In_599,In_976);
nor U1425 (N_1425,In_749,In_679);
nor U1426 (N_1426,In_883,In_116);
and U1427 (N_1427,In_525,In_360);
nor U1428 (N_1428,In_616,In_111);
nand U1429 (N_1429,In_746,In_526);
nor U1430 (N_1430,In_869,In_246);
nor U1431 (N_1431,In_883,In_364);
nor U1432 (N_1432,In_414,In_62);
nor U1433 (N_1433,In_137,In_464);
and U1434 (N_1434,In_692,In_160);
nor U1435 (N_1435,In_69,In_917);
and U1436 (N_1436,In_504,In_47);
nor U1437 (N_1437,In_185,In_774);
and U1438 (N_1438,In_656,In_911);
and U1439 (N_1439,In_901,In_43);
nor U1440 (N_1440,In_332,In_287);
and U1441 (N_1441,In_843,In_515);
and U1442 (N_1442,In_650,In_463);
or U1443 (N_1443,In_769,In_242);
nor U1444 (N_1444,In_137,In_457);
and U1445 (N_1445,In_176,In_522);
nor U1446 (N_1446,In_232,In_5);
nand U1447 (N_1447,In_256,In_551);
nand U1448 (N_1448,In_683,In_308);
nor U1449 (N_1449,In_193,In_98);
or U1450 (N_1450,In_53,In_498);
nor U1451 (N_1451,In_746,In_12);
nand U1452 (N_1452,In_890,In_320);
or U1453 (N_1453,In_735,In_458);
and U1454 (N_1454,In_840,In_872);
nand U1455 (N_1455,In_706,In_485);
and U1456 (N_1456,In_24,In_332);
or U1457 (N_1457,In_103,In_592);
nand U1458 (N_1458,In_704,In_711);
or U1459 (N_1459,In_87,In_174);
or U1460 (N_1460,In_636,In_373);
or U1461 (N_1461,In_836,In_161);
nand U1462 (N_1462,In_849,In_146);
nand U1463 (N_1463,In_798,In_526);
nor U1464 (N_1464,In_874,In_304);
nor U1465 (N_1465,In_259,In_353);
or U1466 (N_1466,In_348,In_372);
nor U1467 (N_1467,In_740,In_683);
nand U1468 (N_1468,In_224,In_964);
xnor U1469 (N_1469,In_273,In_432);
nand U1470 (N_1470,In_120,In_705);
nor U1471 (N_1471,In_747,In_214);
or U1472 (N_1472,In_905,In_29);
nand U1473 (N_1473,In_210,In_665);
or U1474 (N_1474,In_413,In_60);
or U1475 (N_1475,In_838,In_523);
and U1476 (N_1476,In_57,In_203);
nand U1477 (N_1477,In_532,In_750);
and U1478 (N_1478,In_158,In_806);
or U1479 (N_1479,In_812,In_961);
nand U1480 (N_1480,In_263,In_40);
nor U1481 (N_1481,In_824,In_371);
and U1482 (N_1482,In_788,In_513);
or U1483 (N_1483,In_130,In_11);
and U1484 (N_1484,In_389,In_999);
or U1485 (N_1485,In_126,In_825);
or U1486 (N_1486,In_115,In_602);
nor U1487 (N_1487,In_105,In_900);
or U1488 (N_1488,In_808,In_560);
nand U1489 (N_1489,In_624,In_860);
or U1490 (N_1490,In_729,In_550);
nand U1491 (N_1491,In_935,In_310);
nor U1492 (N_1492,In_263,In_189);
nor U1493 (N_1493,In_563,In_215);
nand U1494 (N_1494,In_177,In_529);
or U1495 (N_1495,In_363,In_81);
nand U1496 (N_1496,In_96,In_117);
nor U1497 (N_1497,In_202,In_444);
and U1498 (N_1498,In_405,In_531);
and U1499 (N_1499,In_892,In_977);
nor U1500 (N_1500,In_228,In_622);
nor U1501 (N_1501,In_307,In_587);
or U1502 (N_1502,In_928,In_130);
nor U1503 (N_1503,In_701,In_513);
nor U1504 (N_1504,In_519,In_552);
nand U1505 (N_1505,In_370,In_725);
nor U1506 (N_1506,In_348,In_545);
nand U1507 (N_1507,In_822,In_100);
nor U1508 (N_1508,In_102,In_663);
and U1509 (N_1509,In_17,In_219);
nor U1510 (N_1510,In_522,In_906);
or U1511 (N_1511,In_722,In_954);
nor U1512 (N_1512,In_331,In_24);
nand U1513 (N_1513,In_829,In_819);
or U1514 (N_1514,In_374,In_873);
or U1515 (N_1515,In_461,In_474);
nor U1516 (N_1516,In_657,In_735);
nor U1517 (N_1517,In_291,In_242);
nand U1518 (N_1518,In_26,In_435);
or U1519 (N_1519,In_337,In_776);
or U1520 (N_1520,In_112,In_245);
and U1521 (N_1521,In_682,In_365);
nand U1522 (N_1522,In_24,In_913);
nand U1523 (N_1523,In_920,In_350);
and U1524 (N_1524,In_59,In_226);
or U1525 (N_1525,In_332,In_623);
nand U1526 (N_1526,In_467,In_716);
and U1527 (N_1527,In_358,In_67);
and U1528 (N_1528,In_929,In_621);
or U1529 (N_1529,In_262,In_522);
nand U1530 (N_1530,In_859,In_31);
or U1531 (N_1531,In_494,In_49);
nand U1532 (N_1532,In_671,In_331);
nand U1533 (N_1533,In_702,In_803);
or U1534 (N_1534,In_364,In_461);
nor U1535 (N_1535,In_427,In_613);
nand U1536 (N_1536,In_903,In_160);
nand U1537 (N_1537,In_381,In_869);
xor U1538 (N_1538,In_336,In_501);
or U1539 (N_1539,In_932,In_973);
and U1540 (N_1540,In_748,In_309);
nor U1541 (N_1541,In_239,In_283);
nor U1542 (N_1542,In_630,In_680);
and U1543 (N_1543,In_511,In_217);
nand U1544 (N_1544,In_49,In_125);
nor U1545 (N_1545,In_438,In_327);
or U1546 (N_1546,In_319,In_447);
or U1547 (N_1547,In_302,In_281);
and U1548 (N_1548,In_472,In_801);
and U1549 (N_1549,In_986,In_931);
nand U1550 (N_1550,In_873,In_952);
and U1551 (N_1551,In_534,In_871);
nand U1552 (N_1552,In_384,In_327);
or U1553 (N_1553,In_812,In_935);
and U1554 (N_1554,In_390,In_920);
and U1555 (N_1555,In_550,In_917);
xor U1556 (N_1556,In_997,In_151);
or U1557 (N_1557,In_824,In_504);
nor U1558 (N_1558,In_637,In_173);
or U1559 (N_1559,In_27,In_230);
nor U1560 (N_1560,In_48,In_378);
nand U1561 (N_1561,In_253,In_845);
or U1562 (N_1562,In_781,In_789);
nor U1563 (N_1563,In_222,In_294);
nand U1564 (N_1564,In_315,In_724);
nor U1565 (N_1565,In_366,In_815);
or U1566 (N_1566,In_764,In_8);
nor U1567 (N_1567,In_959,In_526);
and U1568 (N_1568,In_279,In_701);
or U1569 (N_1569,In_262,In_472);
or U1570 (N_1570,In_915,In_272);
and U1571 (N_1571,In_878,In_267);
nand U1572 (N_1572,In_556,In_163);
nor U1573 (N_1573,In_35,In_935);
and U1574 (N_1574,In_983,In_306);
or U1575 (N_1575,In_869,In_698);
and U1576 (N_1576,In_814,In_632);
nor U1577 (N_1577,In_102,In_821);
and U1578 (N_1578,In_421,In_406);
or U1579 (N_1579,In_605,In_571);
nand U1580 (N_1580,In_700,In_143);
nand U1581 (N_1581,In_817,In_33);
nand U1582 (N_1582,In_243,In_655);
nand U1583 (N_1583,In_445,In_411);
nand U1584 (N_1584,In_273,In_28);
xor U1585 (N_1585,In_659,In_692);
nor U1586 (N_1586,In_917,In_358);
xor U1587 (N_1587,In_878,In_140);
nand U1588 (N_1588,In_290,In_561);
and U1589 (N_1589,In_521,In_372);
nor U1590 (N_1590,In_817,In_196);
and U1591 (N_1591,In_947,In_986);
and U1592 (N_1592,In_315,In_327);
nand U1593 (N_1593,In_259,In_14);
or U1594 (N_1594,In_941,In_232);
or U1595 (N_1595,In_713,In_642);
or U1596 (N_1596,In_49,In_444);
or U1597 (N_1597,In_231,In_431);
or U1598 (N_1598,In_596,In_958);
and U1599 (N_1599,In_409,In_170);
or U1600 (N_1600,In_977,In_316);
or U1601 (N_1601,In_561,In_888);
nand U1602 (N_1602,In_379,In_856);
nor U1603 (N_1603,In_274,In_83);
and U1604 (N_1604,In_705,In_376);
nand U1605 (N_1605,In_100,In_949);
or U1606 (N_1606,In_120,In_999);
nand U1607 (N_1607,In_877,In_204);
nor U1608 (N_1608,In_198,In_31);
and U1609 (N_1609,In_27,In_708);
nand U1610 (N_1610,In_744,In_804);
or U1611 (N_1611,In_869,In_856);
nand U1612 (N_1612,In_682,In_900);
or U1613 (N_1613,In_777,In_329);
nand U1614 (N_1614,In_34,In_661);
nand U1615 (N_1615,In_393,In_681);
and U1616 (N_1616,In_672,In_431);
nor U1617 (N_1617,In_669,In_425);
nand U1618 (N_1618,In_147,In_167);
or U1619 (N_1619,In_599,In_764);
and U1620 (N_1620,In_849,In_59);
and U1621 (N_1621,In_439,In_728);
nor U1622 (N_1622,In_635,In_339);
nor U1623 (N_1623,In_258,In_371);
nor U1624 (N_1624,In_734,In_125);
nand U1625 (N_1625,In_92,In_435);
and U1626 (N_1626,In_432,In_831);
or U1627 (N_1627,In_350,In_966);
nor U1628 (N_1628,In_868,In_122);
or U1629 (N_1629,In_976,In_412);
nand U1630 (N_1630,In_393,In_588);
nand U1631 (N_1631,In_721,In_735);
nor U1632 (N_1632,In_507,In_410);
and U1633 (N_1633,In_223,In_591);
and U1634 (N_1634,In_357,In_653);
and U1635 (N_1635,In_341,In_417);
nand U1636 (N_1636,In_468,In_846);
nor U1637 (N_1637,In_259,In_8);
nand U1638 (N_1638,In_662,In_658);
or U1639 (N_1639,In_606,In_242);
nor U1640 (N_1640,In_322,In_714);
or U1641 (N_1641,In_594,In_251);
and U1642 (N_1642,In_415,In_346);
and U1643 (N_1643,In_639,In_414);
nor U1644 (N_1644,In_878,In_526);
or U1645 (N_1645,In_501,In_591);
and U1646 (N_1646,In_798,In_615);
nor U1647 (N_1647,In_842,In_250);
or U1648 (N_1648,In_685,In_633);
and U1649 (N_1649,In_514,In_110);
nor U1650 (N_1650,In_709,In_658);
nor U1651 (N_1651,In_95,In_672);
nor U1652 (N_1652,In_673,In_927);
or U1653 (N_1653,In_893,In_693);
nor U1654 (N_1654,In_317,In_543);
nor U1655 (N_1655,In_495,In_840);
or U1656 (N_1656,In_479,In_297);
or U1657 (N_1657,In_373,In_869);
nor U1658 (N_1658,In_630,In_514);
nand U1659 (N_1659,In_895,In_620);
and U1660 (N_1660,In_738,In_991);
and U1661 (N_1661,In_506,In_809);
and U1662 (N_1662,In_550,In_357);
and U1663 (N_1663,In_638,In_933);
and U1664 (N_1664,In_97,In_961);
nor U1665 (N_1665,In_485,In_738);
nor U1666 (N_1666,In_496,In_446);
or U1667 (N_1667,In_57,In_464);
and U1668 (N_1668,In_827,In_702);
or U1669 (N_1669,In_724,In_621);
or U1670 (N_1670,In_132,In_344);
nand U1671 (N_1671,In_783,In_633);
and U1672 (N_1672,In_236,In_648);
or U1673 (N_1673,In_994,In_454);
nor U1674 (N_1674,In_460,In_31);
and U1675 (N_1675,In_178,In_500);
nand U1676 (N_1676,In_506,In_417);
or U1677 (N_1677,In_14,In_228);
nor U1678 (N_1678,In_797,In_617);
or U1679 (N_1679,In_975,In_678);
or U1680 (N_1680,In_612,In_334);
nor U1681 (N_1681,In_30,In_735);
nand U1682 (N_1682,In_631,In_63);
or U1683 (N_1683,In_94,In_764);
nor U1684 (N_1684,In_50,In_976);
and U1685 (N_1685,In_300,In_642);
nor U1686 (N_1686,In_430,In_557);
and U1687 (N_1687,In_180,In_192);
and U1688 (N_1688,In_909,In_531);
and U1689 (N_1689,In_667,In_416);
xor U1690 (N_1690,In_947,In_681);
or U1691 (N_1691,In_548,In_955);
nor U1692 (N_1692,In_284,In_17);
nand U1693 (N_1693,In_701,In_493);
nand U1694 (N_1694,In_752,In_843);
and U1695 (N_1695,In_566,In_562);
and U1696 (N_1696,In_701,In_277);
and U1697 (N_1697,In_976,In_648);
nand U1698 (N_1698,In_554,In_343);
nor U1699 (N_1699,In_544,In_259);
or U1700 (N_1700,In_140,In_984);
or U1701 (N_1701,In_249,In_737);
nand U1702 (N_1702,In_445,In_954);
or U1703 (N_1703,In_990,In_962);
and U1704 (N_1704,In_554,In_288);
and U1705 (N_1705,In_214,In_830);
or U1706 (N_1706,In_640,In_429);
or U1707 (N_1707,In_922,In_743);
and U1708 (N_1708,In_978,In_255);
nor U1709 (N_1709,In_468,In_148);
nand U1710 (N_1710,In_618,In_799);
nand U1711 (N_1711,In_960,In_632);
nor U1712 (N_1712,In_492,In_80);
and U1713 (N_1713,In_289,In_529);
nor U1714 (N_1714,In_101,In_562);
or U1715 (N_1715,In_291,In_862);
nor U1716 (N_1716,In_133,In_849);
and U1717 (N_1717,In_570,In_246);
nor U1718 (N_1718,In_254,In_878);
and U1719 (N_1719,In_607,In_82);
xnor U1720 (N_1720,In_966,In_227);
or U1721 (N_1721,In_485,In_912);
nand U1722 (N_1722,In_896,In_496);
or U1723 (N_1723,In_844,In_751);
nand U1724 (N_1724,In_75,In_411);
nor U1725 (N_1725,In_342,In_702);
nand U1726 (N_1726,In_328,In_401);
or U1727 (N_1727,In_937,In_96);
nor U1728 (N_1728,In_422,In_218);
xor U1729 (N_1729,In_488,In_458);
nor U1730 (N_1730,In_468,In_875);
nand U1731 (N_1731,In_498,In_432);
nor U1732 (N_1732,In_492,In_133);
and U1733 (N_1733,In_643,In_972);
nor U1734 (N_1734,In_599,In_560);
or U1735 (N_1735,In_588,In_945);
nor U1736 (N_1736,In_28,In_925);
nand U1737 (N_1737,In_315,In_610);
nand U1738 (N_1738,In_528,In_824);
nor U1739 (N_1739,In_507,In_157);
and U1740 (N_1740,In_745,In_450);
or U1741 (N_1741,In_455,In_128);
nor U1742 (N_1742,In_89,In_735);
and U1743 (N_1743,In_596,In_247);
or U1744 (N_1744,In_890,In_410);
or U1745 (N_1745,In_168,In_524);
or U1746 (N_1746,In_739,In_858);
and U1747 (N_1747,In_96,In_302);
nor U1748 (N_1748,In_65,In_149);
nor U1749 (N_1749,In_459,In_124);
and U1750 (N_1750,In_411,In_925);
or U1751 (N_1751,In_365,In_3);
nand U1752 (N_1752,In_406,In_89);
nor U1753 (N_1753,In_829,In_413);
nand U1754 (N_1754,In_374,In_439);
and U1755 (N_1755,In_305,In_179);
or U1756 (N_1756,In_36,In_367);
nor U1757 (N_1757,In_221,In_514);
nand U1758 (N_1758,In_924,In_467);
xor U1759 (N_1759,In_462,In_757);
nand U1760 (N_1760,In_311,In_278);
nand U1761 (N_1761,In_319,In_685);
or U1762 (N_1762,In_679,In_973);
and U1763 (N_1763,In_996,In_807);
or U1764 (N_1764,In_582,In_519);
or U1765 (N_1765,In_425,In_584);
or U1766 (N_1766,In_120,In_792);
nand U1767 (N_1767,In_976,In_745);
and U1768 (N_1768,In_852,In_38);
nand U1769 (N_1769,In_400,In_902);
and U1770 (N_1770,In_155,In_383);
and U1771 (N_1771,In_948,In_700);
and U1772 (N_1772,In_880,In_984);
nor U1773 (N_1773,In_642,In_803);
and U1774 (N_1774,In_549,In_136);
nor U1775 (N_1775,In_283,In_63);
nor U1776 (N_1776,In_643,In_441);
nor U1777 (N_1777,In_461,In_88);
nand U1778 (N_1778,In_915,In_513);
or U1779 (N_1779,In_66,In_605);
nor U1780 (N_1780,In_397,In_909);
nor U1781 (N_1781,In_189,In_46);
or U1782 (N_1782,In_396,In_913);
nand U1783 (N_1783,In_680,In_192);
nor U1784 (N_1784,In_426,In_129);
or U1785 (N_1785,In_59,In_870);
or U1786 (N_1786,In_674,In_804);
and U1787 (N_1787,In_894,In_239);
and U1788 (N_1788,In_548,In_819);
or U1789 (N_1789,In_752,In_240);
and U1790 (N_1790,In_605,In_155);
nor U1791 (N_1791,In_753,In_226);
nand U1792 (N_1792,In_633,In_819);
or U1793 (N_1793,In_485,In_38);
nor U1794 (N_1794,In_950,In_873);
nand U1795 (N_1795,In_63,In_933);
and U1796 (N_1796,In_628,In_377);
nor U1797 (N_1797,In_269,In_260);
nand U1798 (N_1798,In_140,In_172);
and U1799 (N_1799,In_380,In_111);
nor U1800 (N_1800,In_476,In_904);
nor U1801 (N_1801,In_368,In_529);
or U1802 (N_1802,In_657,In_207);
and U1803 (N_1803,In_874,In_501);
nor U1804 (N_1804,In_920,In_423);
or U1805 (N_1805,In_66,In_10);
xor U1806 (N_1806,In_205,In_204);
nand U1807 (N_1807,In_149,In_529);
or U1808 (N_1808,In_457,In_107);
nand U1809 (N_1809,In_358,In_686);
nor U1810 (N_1810,In_957,In_487);
and U1811 (N_1811,In_658,In_359);
nor U1812 (N_1812,In_286,In_947);
nor U1813 (N_1813,In_388,In_814);
and U1814 (N_1814,In_81,In_987);
or U1815 (N_1815,In_597,In_478);
nand U1816 (N_1816,In_771,In_120);
and U1817 (N_1817,In_702,In_81);
and U1818 (N_1818,In_577,In_451);
nor U1819 (N_1819,In_433,In_453);
nand U1820 (N_1820,In_946,In_478);
and U1821 (N_1821,In_601,In_424);
and U1822 (N_1822,In_426,In_808);
nor U1823 (N_1823,In_789,In_241);
and U1824 (N_1824,In_291,In_15);
or U1825 (N_1825,In_164,In_156);
and U1826 (N_1826,In_192,In_669);
or U1827 (N_1827,In_540,In_92);
or U1828 (N_1828,In_56,In_270);
nor U1829 (N_1829,In_512,In_631);
nand U1830 (N_1830,In_984,In_815);
nand U1831 (N_1831,In_719,In_637);
and U1832 (N_1832,In_776,In_68);
and U1833 (N_1833,In_529,In_888);
or U1834 (N_1834,In_874,In_476);
and U1835 (N_1835,In_612,In_192);
nand U1836 (N_1836,In_716,In_353);
nor U1837 (N_1837,In_363,In_654);
and U1838 (N_1838,In_694,In_146);
nand U1839 (N_1839,In_159,In_109);
nand U1840 (N_1840,In_538,In_365);
nor U1841 (N_1841,In_155,In_105);
or U1842 (N_1842,In_631,In_10);
nand U1843 (N_1843,In_25,In_451);
nor U1844 (N_1844,In_594,In_64);
and U1845 (N_1845,In_154,In_807);
nor U1846 (N_1846,In_521,In_104);
nand U1847 (N_1847,In_290,In_159);
or U1848 (N_1848,In_199,In_445);
nand U1849 (N_1849,In_838,In_949);
nor U1850 (N_1850,In_540,In_125);
or U1851 (N_1851,In_688,In_987);
or U1852 (N_1852,In_243,In_4);
and U1853 (N_1853,In_738,In_131);
nor U1854 (N_1854,In_150,In_962);
nor U1855 (N_1855,In_939,In_411);
or U1856 (N_1856,In_461,In_954);
nor U1857 (N_1857,In_521,In_240);
and U1858 (N_1858,In_275,In_206);
or U1859 (N_1859,In_898,In_280);
and U1860 (N_1860,In_554,In_357);
nand U1861 (N_1861,In_645,In_802);
nor U1862 (N_1862,In_718,In_278);
nand U1863 (N_1863,In_407,In_987);
nand U1864 (N_1864,In_860,In_307);
nor U1865 (N_1865,In_423,In_447);
nand U1866 (N_1866,In_978,In_284);
or U1867 (N_1867,In_2,In_798);
nor U1868 (N_1868,In_943,In_578);
and U1869 (N_1869,In_973,In_411);
nand U1870 (N_1870,In_366,In_929);
nand U1871 (N_1871,In_601,In_994);
and U1872 (N_1872,In_926,In_709);
nand U1873 (N_1873,In_1,In_404);
or U1874 (N_1874,In_817,In_214);
and U1875 (N_1875,In_831,In_11);
nor U1876 (N_1876,In_337,In_855);
and U1877 (N_1877,In_509,In_775);
and U1878 (N_1878,In_134,In_414);
and U1879 (N_1879,In_553,In_684);
nor U1880 (N_1880,In_78,In_905);
nor U1881 (N_1881,In_535,In_508);
nand U1882 (N_1882,In_952,In_718);
nand U1883 (N_1883,In_467,In_300);
or U1884 (N_1884,In_425,In_452);
and U1885 (N_1885,In_834,In_551);
and U1886 (N_1886,In_985,In_706);
and U1887 (N_1887,In_467,In_400);
and U1888 (N_1888,In_153,In_700);
nor U1889 (N_1889,In_473,In_887);
nand U1890 (N_1890,In_869,In_598);
nand U1891 (N_1891,In_257,In_747);
nand U1892 (N_1892,In_335,In_59);
or U1893 (N_1893,In_518,In_365);
and U1894 (N_1894,In_201,In_661);
nand U1895 (N_1895,In_674,In_252);
and U1896 (N_1896,In_518,In_828);
nand U1897 (N_1897,In_389,In_409);
nand U1898 (N_1898,In_164,In_97);
nor U1899 (N_1899,In_875,In_878);
and U1900 (N_1900,In_698,In_13);
or U1901 (N_1901,In_537,In_398);
or U1902 (N_1902,In_680,In_174);
nand U1903 (N_1903,In_5,In_428);
or U1904 (N_1904,In_246,In_426);
or U1905 (N_1905,In_851,In_894);
and U1906 (N_1906,In_759,In_788);
nor U1907 (N_1907,In_692,In_695);
nand U1908 (N_1908,In_904,In_923);
nor U1909 (N_1909,In_724,In_321);
nand U1910 (N_1910,In_874,In_584);
nor U1911 (N_1911,In_775,In_924);
nand U1912 (N_1912,In_252,In_335);
or U1913 (N_1913,In_428,In_961);
or U1914 (N_1914,In_356,In_145);
nand U1915 (N_1915,In_266,In_44);
or U1916 (N_1916,In_12,In_590);
nand U1917 (N_1917,In_797,In_402);
nor U1918 (N_1918,In_347,In_544);
or U1919 (N_1919,In_30,In_402);
or U1920 (N_1920,In_77,In_71);
nand U1921 (N_1921,In_193,In_437);
and U1922 (N_1922,In_868,In_439);
or U1923 (N_1923,In_599,In_694);
and U1924 (N_1924,In_86,In_661);
nand U1925 (N_1925,In_659,In_856);
and U1926 (N_1926,In_620,In_679);
or U1927 (N_1927,In_487,In_456);
nor U1928 (N_1928,In_44,In_587);
nand U1929 (N_1929,In_952,In_119);
and U1930 (N_1930,In_381,In_864);
and U1931 (N_1931,In_361,In_611);
nor U1932 (N_1932,In_392,In_246);
and U1933 (N_1933,In_444,In_812);
nor U1934 (N_1934,In_302,In_381);
nor U1935 (N_1935,In_544,In_908);
nor U1936 (N_1936,In_512,In_173);
nand U1937 (N_1937,In_228,In_772);
nor U1938 (N_1938,In_970,In_420);
or U1939 (N_1939,In_282,In_345);
nand U1940 (N_1940,In_73,In_318);
nand U1941 (N_1941,In_315,In_375);
nand U1942 (N_1942,In_228,In_261);
nor U1943 (N_1943,In_310,In_452);
and U1944 (N_1944,In_525,In_143);
and U1945 (N_1945,In_240,In_966);
and U1946 (N_1946,In_301,In_116);
nor U1947 (N_1947,In_419,In_332);
and U1948 (N_1948,In_73,In_447);
nor U1949 (N_1949,In_320,In_930);
nand U1950 (N_1950,In_272,In_737);
and U1951 (N_1951,In_162,In_348);
nand U1952 (N_1952,In_614,In_257);
nor U1953 (N_1953,In_310,In_327);
nor U1954 (N_1954,In_246,In_794);
or U1955 (N_1955,In_732,In_630);
nand U1956 (N_1956,In_603,In_435);
nor U1957 (N_1957,In_129,In_82);
and U1958 (N_1958,In_522,In_511);
or U1959 (N_1959,In_304,In_595);
or U1960 (N_1960,In_857,In_705);
nand U1961 (N_1961,In_616,In_599);
nand U1962 (N_1962,In_20,In_346);
or U1963 (N_1963,In_918,In_659);
or U1964 (N_1964,In_518,In_188);
or U1965 (N_1965,In_0,In_857);
nand U1966 (N_1966,In_370,In_863);
or U1967 (N_1967,In_298,In_823);
nor U1968 (N_1968,In_502,In_161);
nand U1969 (N_1969,In_586,In_135);
or U1970 (N_1970,In_22,In_400);
or U1971 (N_1971,In_107,In_870);
nand U1972 (N_1972,In_589,In_603);
nor U1973 (N_1973,In_694,In_302);
nand U1974 (N_1974,In_366,In_687);
nand U1975 (N_1975,In_281,In_60);
or U1976 (N_1976,In_299,In_86);
nand U1977 (N_1977,In_177,In_549);
or U1978 (N_1978,In_672,In_715);
or U1979 (N_1979,In_839,In_144);
xnor U1980 (N_1980,In_532,In_599);
or U1981 (N_1981,In_839,In_235);
nor U1982 (N_1982,In_714,In_576);
nor U1983 (N_1983,In_474,In_664);
and U1984 (N_1984,In_694,In_717);
or U1985 (N_1985,In_498,In_998);
nand U1986 (N_1986,In_650,In_530);
or U1987 (N_1987,In_806,In_779);
and U1988 (N_1988,In_684,In_628);
or U1989 (N_1989,In_388,In_236);
and U1990 (N_1990,In_465,In_105);
nor U1991 (N_1991,In_643,In_580);
or U1992 (N_1992,In_796,In_804);
nor U1993 (N_1993,In_888,In_947);
nand U1994 (N_1994,In_148,In_41);
nand U1995 (N_1995,In_672,In_850);
and U1996 (N_1996,In_51,In_7);
nor U1997 (N_1997,In_204,In_378);
and U1998 (N_1998,In_460,In_542);
and U1999 (N_1999,In_235,In_764);
or U2000 (N_2000,In_629,In_616);
nand U2001 (N_2001,In_477,In_249);
xnor U2002 (N_2002,In_409,In_567);
or U2003 (N_2003,In_774,In_132);
nor U2004 (N_2004,In_805,In_194);
nand U2005 (N_2005,In_244,In_523);
or U2006 (N_2006,In_998,In_386);
or U2007 (N_2007,In_754,In_440);
and U2008 (N_2008,In_890,In_363);
or U2009 (N_2009,In_725,In_821);
nor U2010 (N_2010,In_255,In_31);
and U2011 (N_2011,In_951,In_93);
xor U2012 (N_2012,In_611,In_11);
nor U2013 (N_2013,In_22,In_851);
and U2014 (N_2014,In_834,In_828);
and U2015 (N_2015,In_120,In_76);
nor U2016 (N_2016,In_304,In_453);
or U2017 (N_2017,In_514,In_461);
nand U2018 (N_2018,In_574,In_564);
and U2019 (N_2019,In_996,In_340);
nor U2020 (N_2020,In_938,In_48);
or U2021 (N_2021,In_250,In_931);
nor U2022 (N_2022,In_527,In_607);
and U2023 (N_2023,In_519,In_347);
and U2024 (N_2024,In_427,In_501);
nand U2025 (N_2025,In_412,In_794);
nand U2026 (N_2026,In_764,In_920);
nor U2027 (N_2027,In_822,In_429);
nor U2028 (N_2028,In_647,In_14);
nand U2029 (N_2029,In_558,In_135);
or U2030 (N_2030,In_139,In_456);
or U2031 (N_2031,In_944,In_727);
and U2032 (N_2032,In_399,In_364);
nand U2033 (N_2033,In_621,In_22);
and U2034 (N_2034,In_732,In_448);
nand U2035 (N_2035,In_915,In_605);
or U2036 (N_2036,In_693,In_933);
nand U2037 (N_2037,In_980,In_869);
or U2038 (N_2038,In_730,In_296);
and U2039 (N_2039,In_132,In_665);
nor U2040 (N_2040,In_26,In_316);
nor U2041 (N_2041,In_651,In_95);
and U2042 (N_2042,In_852,In_291);
or U2043 (N_2043,In_133,In_172);
and U2044 (N_2044,In_739,In_515);
nand U2045 (N_2045,In_631,In_509);
and U2046 (N_2046,In_170,In_143);
and U2047 (N_2047,In_356,In_713);
or U2048 (N_2048,In_910,In_987);
and U2049 (N_2049,In_581,In_326);
and U2050 (N_2050,In_273,In_974);
and U2051 (N_2051,In_524,In_285);
and U2052 (N_2052,In_398,In_410);
and U2053 (N_2053,In_684,In_70);
nor U2054 (N_2054,In_597,In_605);
nor U2055 (N_2055,In_211,In_52);
or U2056 (N_2056,In_389,In_922);
xor U2057 (N_2057,In_947,In_854);
nand U2058 (N_2058,In_480,In_297);
and U2059 (N_2059,In_180,In_183);
or U2060 (N_2060,In_781,In_855);
nor U2061 (N_2061,In_439,In_963);
or U2062 (N_2062,In_417,In_238);
nor U2063 (N_2063,In_660,In_497);
or U2064 (N_2064,In_976,In_299);
nor U2065 (N_2065,In_810,In_574);
nor U2066 (N_2066,In_591,In_306);
nand U2067 (N_2067,In_847,In_192);
nor U2068 (N_2068,In_172,In_811);
xor U2069 (N_2069,In_875,In_846);
nand U2070 (N_2070,In_684,In_746);
nand U2071 (N_2071,In_920,In_312);
or U2072 (N_2072,In_226,In_552);
and U2073 (N_2073,In_276,In_593);
and U2074 (N_2074,In_225,In_934);
or U2075 (N_2075,In_780,In_539);
or U2076 (N_2076,In_677,In_440);
or U2077 (N_2077,In_744,In_402);
or U2078 (N_2078,In_434,In_177);
nand U2079 (N_2079,In_27,In_188);
nor U2080 (N_2080,In_162,In_640);
nand U2081 (N_2081,In_536,In_952);
nand U2082 (N_2082,In_416,In_444);
or U2083 (N_2083,In_796,In_912);
nor U2084 (N_2084,In_633,In_963);
nand U2085 (N_2085,In_888,In_436);
nand U2086 (N_2086,In_312,In_575);
or U2087 (N_2087,In_616,In_419);
and U2088 (N_2088,In_994,In_618);
nor U2089 (N_2089,In_464,In_343);
nand U2090 (N_2090,In_386,In_345);
nand U2091 (N_2091,In_7,In_901);
or U2092 (N_2092,In_533,In_463);
or U2093 (N_2093,In_627,In_420);
or U2094 (N_2094,In_835,In_14);
or U2095 (N_2095,In_570,In_929);
nand U2096 (N_2096,In_570,In_119);
nor U2097 (N_2097,In_791,In_622);
or U2098 (N_2098,In_798,In_681);
nor U2099 (N_2099,In_349,In_981);
or U2100 (N_2100,In_409,In_365);
and U2101 (N_2101,In_34,In_921);
nand U2102 (N_2102,In_356,In_882);
or U2103 (N_2103,In_77,In_398);
and U2104 (N_2104,In_501,In_636);
or U2105 (N_2105,In_204,In_845);
nor U2106 (N_2106,In_903,In_419);
nor U2107 (N_2107,In_284,In_925);
and U2108 (N_2108,In_49,In_495);
or U2109 (N_2109,In_697,In_707);
nor U2110 (N_2110,In_860,In_206);
and U2111 (N_2111,In_291,In_841);
or U2112 (N_2112,In_947,In_70);
or U2113 (N_2113,In_141,In_755);
nor U2114 (N_2114,In_791,In_412);
and U2115 (N_2115,In_483,In_589);
nor U2116 (N_2116,In_397,In_885);
nor U2117 (N_2117,In_409,In_238);
or U2118 (N_2118,In_763,In_742);
nand U2119 (N_2119,In_555,In_570);
or U2120 (N_2120,In_851,In_647);
nor U2121 (N_2121,In_359,In_548);
nand U2122 (N_2122,In_459,In_919);
xor U2123 (N_2123,In_25,In_720);
nor U2124 (N_2124,In_712,In_276);
xnor U2125 (N_2125,In_717,In_766);
nand U2126 (N_2126,In_505,In_46);
or U2127 (N_2127,In_236,In_843);
nand U2128 (N_2128,In_751,In_574);
and U2129 (N_2129,In_8,In_541);
nand U2130 (N_2130,In_427,In_689);
nand U2131 (N_2131,In_893,In_59);
or U2132 (N_2132,In_544,In_19);
nand U2133 (N_2133,In_879,In_12);
nor U2134 (N_2134,In_66,In_401);
or U2135 (N_2135,In_226,In_87);
nor U2136 (N_2136,In_37,In_725);
nor U2137 (N_2137,In_240,In_465);
and U2138 (N_2138,In_731,In_315);
or U2139 (N_2139,In_969,In_47);
and U2140 (N_2140,In_844,In_8);
and U2141 (N_2141,In_900,In_116);
and U2142 (N_2142,In_562,In_202);
nand U2143 (N_2143,In_479,In_129);
nor U2144 (N_2144,In_723,In_852);
or U2145 (N_2145,In_97,In_775);
nor U2146 (N_2146,In_770,In_551);
nor U2147 (N_2147,In_105,In_40);
nand U2148 (N_2148,In_543,In_646);
nor U2149 (N_2149,In_122,In_211);
or U2150 (N_2150,In_82,In_128);
nor U2151 (N_2151,In_407,In_457);
nand U2152 (N_2152,In_857,In_162);
or U2153 (N_2153,In_659,In_488);
or U2154 (N_2154,In_264,In_933);
or U2155 (N_2155,In_231,In_846);
nor U2156 (N_2156,In_370,In_353);
and U2157 (N_2157,In_612,In_596);
or U2158 (N_2158,In_236,In_665);
nor U2159 (N_2159,In_162,In_527);
and U2160 (N_2160,In_236,In_170);
xnor U2161 (N_2161,In_102,In_738);
nor U2162 (N_2162,In_892,In_360);
and U2163 (N_2163,In_150,In_14);
nand U2164 (N_2164,In_422,In_788);
nor U2165 (N_2165,In_523,In_648);
nand U2166 (N_2166,In_897,In_91);
or U2167 (N_2167,In_323,In_223);
and U2168 (N_2168,In_241,In_100);
nand U2169 (N_2169,In_279,In_806);
nor U2170 (N_2170,In_384,In_321);
nor U2171 (N_2171,In_75,In_287);
nand U2172 (N_2172,In_534,In_460);
or U2173 (N_2173,In_538,In_930);
nor U2174 (N_2174,In_804,In_416);
or U2175 (N_2175,In_681,In_179);
nor U2176 (N_2176,In_870,In_71);
and U2177 (N_2177,In_295,In_349);
or U2178 (N_2178,In_170,In_945);
nor U2179 (N_2179,In_600,In_556);
and U2180 (N_2180,In_53,In_11);
and U2181 (N_2181,In_484,In_355);
and U2182 (N_2182,In_578,In_800);
and U2183 (N_2183,In_974,In_575);
or U2184 (N_2184,In_179,In_861);
and U2185 (N_2185,In_931,In_585);
or U2186 (N_2186,In_400,In_551);
nand U2187 (N_2187,In_152,In_210);
or U2188 (N_2188,In_624,In_444);
nor U2189 (N_2189,In_160,In_556);
nor U2190 (N_2190,In_408,In_673);
nor U2191 (N_2191,In_714,In_185);
nand U2192 (N_2192,In_474,In_654);
or U2193 (N_2193,In_409,In_873);
nor U2194 (N_2194,In_966,In_956);
or U2195 (N_2195,In_503,In_481);
and U2196 (N_2196,In_937,In_127);
nand U2197 (N_2197,In_984,In_676);
nand U2198 (N_2198,In_245,In_39);
nand U2199 (N_2199,In_734,In_660);
nor U2200 (N_2200,In_536,In_299);
nand U2201 (N_2201,In_973,In_998);
nand U2202 (N_2202,In_947,In_534);
and U2203 (N_2203,In_278,In_265);
and U2204 (N_2204,In_785,In_85);
or U2205 (N_2205,In_385,In_627);
or U2206 (N_2206,In_322,In_179);
nand U2207 (N_2207,In_890,In_735);
or U2208 (N_2208,In_580,In_811);
or U2209 (N_2209,In_270,In_162);
nand U2210 (N_2210,In_333,In_708);
and U2211 (N_2211,In_375,In_879);
or U2212 (N_2212,In_672,In_972);
or U2213 (N_2213,In_101,In_860);
and U2214 (N_2214,In_406,In_214);
and U2215 (N_2215,In_252,In_831);
nor U2216 (N_2216,In_455,In_33);
nor U2217 (N_2217,In_439,In_776);
nor U2218 (N_2218,In_289,In_133);
nand U2219 (N_2219,In_894,In_905);
nand U2220 (N_2220,In_972,In_293);
and U2221 (N_2221,In_316,In_163);
nor U2222 (N_2222,In_74,In_519);
and U2223 (N_2223,In_45,In_77);
nor U2224 (N_2224,In_957,In_711);
or U2225 (N_2225,In_773,In_712);
nand U2226 (N_2226,In_562,In_985);
nor U2227 (N_2227,In_362,In_923);
and U2228 (N_2228,In_762,In_462);
nor U2229 (N_2229,In_934,In_513);
or U2230 (N_2230,In_747,In_570);
or U2231 (N_2231,In_799,In_552);
nand U2232 (N_2232,In_57,In_605);
nor U2233 (N_2233,In_17,In_757);
nand U2234 (N_2234,In_975,In_11);
nand U2235 (N_2235,In_835,In_670);
or U2236 (N_2236,In_889,In_625);
nor U2237 (N_2237,In_134,In_361);
and U2238 (N_2238,In_453,In_588);
and U2239 (N_2239,In_220,In_897);
nor U2240 (N_2240,In_907,In_349);
nand U2241 (N_2241,In_689,In_893);
and U2242 (N_2242,In_470,In_286);
or U2243 (N_2243,In_127,In_291);
nor U2244 (N_2244,In_193,In_78);
nor U2245 (N_2245,In_752,In_64);
or U2246 (N_2246,In_598,In_492);
xnor U2247 (N_2247,In_132,In_289);
nor U2248 (N_2248,In_718,In_725);
nand U2249 (N_2249,In_624,In_868);
and U2250 (N_2250,In_824,In_922);
or U2251 (N_2251,In_377,In_79);
nor U2252 (N_2252,In_163,In_19);
and U2253 (N_2253,In_602,In_495);
nor U2254 (N_2254,In_954,In_505);
and U2255 (N_2255,In_909,In_933);
nor U2256 (N_2256,In_751,In_616);
and U2257 (N_2257,In_571,In_79);
or U2258 (N_2258,In_590,In_322);
nor U2259 (N_2259,In_800,In_63);
nor U2260 (N_2260,In_657,In_879);
or U2261 (N_2261,In_91,In_148);
nor U2262 (N_2262,In_338,In_322);
or U2263 (N_2263,In_868,In_206);
nor U2264 (N_2264,In_901,In_145);
and U2265 (N_2265,In_561,In_265);
nand U2266 (N_2266,In_649,In_202);
nor U2267 (N_2267,In_602,In_336);
and U2268 (N_2268,In_803,In_609);
nand U2269 (N_2269,In_675,In_488);
nand U2270 (N_2270,In_121,In_773);
nor U2271 (N_2271,In_216,In_594);
and U2272 (N_2272,In_358,In_724);
and U2273 (N_2273,In_835,In_154);
and U2274 (N_2274,In_506,In_885);
or U2275 (N_2275,In_571,In_289);
nand U2276 (N_2276,In_202,In_377);
nor U2277 (N_2277,In_728,In_222);
or U2278 (N_2278,In_868,In_741);
nor U2279 (N_2279,In_955,In_504);
nor U2280 (N_2280,In_390,In_126);
and U2281 (N_2281,In_790,In_594);
nor U2282 (N_2282,In_743,In_744);
nand U2283 (N_2283,In_966,In_536);
nor U2284 (N_2284,In_652,In_439);
nor U2285 (N_2285,In_568,In_879);
nand U2286 (N_2286,In_613,In_452);
or U2287 (N_2287,In_677,In_187);
and U2288 (N_2288,In_56,In_480);
nand U2289 (N_2289,In_508,In_194);
and U2290 (N_2290,In_551,In_370);
nand U2291 (N_2291,In_206,In_268);
or U2292 (N_2292,In_522,In_388);
nor U2293 (N_2293,In_872,In_946);
nand U2294 (N_2294,In_446,In_325);
nor U2295 (N_2295,In_776,In_508);
and U2296 (N_2296,In_65,In_403);
and U2297 (N_2297,In_879,In_165);
nand U2298 (N_2298,In_425,In_965);
nor U2299 (N_2299,In_273,In_439);
nand U2300 (N_2300,In_597,In_620);
nand U2301 (N_2301,In_822,In_5);
nand U2302 (N_2302,In_845,In_26);
xor U2303 (N_2303,In_103,In_967);
nor U2304 (N_2304,In_950,In_329);
and U2305 (N_2305,In_549,In_456);
and U2306 (N_2306,In_700,In_653);
or U2307 (N_2307,In_405,In_97);
and U2308 (N_2308,In_68,In_565);
nor U2309 (N_2309,In_560,In_993);
and U2310 (N_2310,In_36,In_486);
or U2311 (N_2311,In_558,In_946);
nor U2312 (N_2312,In_709,In_480);
nand U2313 (N_2313,In_890,In_989);
or U2314 (N_2314,In_727,In_634);
nor U2315 (N_2315,In_741,In_414);
nor U2316 (N_2316,In_120,In_698);
or U2317 (N_2317,In_926,In_382);
or U2318 (N_2318,In_504,In_642);
or U2319 (N_2319,In_999,In_880);
nand U2320 (N_2320,In_644,In_28);
nor U2321 (N_2321,In_648,In_886);
nor U2322 (N_2322,In_744,In_66);
nor U2323 (N_2323,In_644,In_665);
and U2324 (N_2324,In_875,In_794);
or U2325 (N_2325,In_726,In_779);
and U2326 (N_2326,In_865,In_226);
and U2327 (N_2327,In_68,In_662);
or U2328 (N_2328,In_542,In_347);
nand U2329 (N_2329,In_982,In_235);
or U2330 (N_2330,In_476,In_233);
and U2331 (N_2331,In_689,In_64);
and U2332 (N_2332,In_685,In_435);
nor U2333 (N_2333,In_207,In_605);
nor U2334 (N_2334,In_42,In_591);
and U2335 (N_2335,In_215,In_537);
nand U2336 (N_2336,In_128,In_158);
nand U2337 (N_2337,In_657,In_959);
and U2338 (N_2338,In_527,In_929);
and U2339 (N_2339,In_607,In_831);
nor U2340 (N_2340,In_707,In_910);
nor U2341 (N_2341,In_941,In_777);
nor U2342 (N_2342,In_319,In_583);
nor U2343 (N_2343,In_889,In_233);
nand U2344 (N_2344,In_394,In_576);
nor U2345 (N_2345,In_89,In_514);
and U2346 (N_2346,In_163,In_198);
nor U2347 (N_2347,In_175,In_26);
or U2348 (N_2348,In_781,In_209);
nor U2349 (N_2349,In_263,In_523);
or U2350 (N_2350,In_735,In_525);
or U2351 (N_2351,In_474,In_95);
nor U2352 (N_2352,In_326,In_944);
or U2353 (N_2353,In_714,In_566);
and U2354 (N_2354,In_702,In_141);
nor U2355 (N_2355,In_348,In_126);
or U2356 (N_2356,In_969,In_936);
or U2357 (N_2357,In_544,In_371);
or U2358 (N_2358,In_453,In_523);
xnor U2359 (N_2359,In_871,In_262);
and U2360 (N_2360,In_954,In_656);
nand U2361 (N_2361,In_579,In_999);
and U2362 (N_2362,In_428,In_976);
nor U2363 (N_2363,In_745,In_693);
and U2364 (N_2364,In_949,In_220);
or U2365 (N_2365,In_420,In_747);
nand U2366 (N_2366,In_708,In_62);
or U2367 (N_2367,In_369,In_854);
or U2368 (N_2368,In_105,In_103);
nor U2369 (N_2369,In_950,In_328);
and U2370 (N_2370,In_683,In_898);
nand U2371 (N_2371,In_182,In_219);
and U2372 (N_2372,In_966,In_94);
and U2373 (N_2373,In_132,In_709);
and U2374 (N_2374,In_228,In_68);
nor U2375 (N_2375,In_533,In_79);
nor U2376 (N_2376,In_765,In_859);
and U2377 (N_2377,In_305,In_135);
nand U2378 (N_2378,In_586,In_391);
and U2379 (N_2379,In_166,In_518);
and U2380 (N_2380,In_937,In_667);
and U2381 (N_2381,In_633,In_220);
or U2382 (N_2382,In_349,In_764);
and U2383 (N_2383,In_135,In_601);
and U2384 (N_2384,In_225,In_0);
nand U2385 (N_2385,In_568,In_691);
nor U2386 (N_2386,In_880,In_495);
or U2387 (N_2387,In_637,In_52);
nor U2388 (N_2388,In_78,In_917);
or U2389 (N_2389,In_587,In_855);
or U2390 (N_2390,In_294,In_164);
nor U2391 (N_2391,In_110,In_227);
and U2392 (N_2392,In_969,In_725);
or U2393 (N_2393,In_810,In_658);
nor U2394 (N_2394,In_633,In_769);
and U2395 (N_2395,In_625,In_945);
xor U2396 (N_2396,In_152,In_705);
and U2397 (N_2397,In_91,In_81);
and U2398 (N_2398,In_868,In_39);
nor U2399 (N_2399,In_177,In_663);
and U2400 (N_2400,In_844,In_982);
nand U2401 (N_2401,In_629,In_798);
and U2402 (N_2402,In_970,In_968);
or U2403 (N_2403,In_633,In_780);
or U2404 (N_2404,In_732,In_379);
nor U2405 (N_2405,In_500,In_570);
nor U2406 (N_2406,In_607,In_678);
and U2407 (N_2407,In_411,In_447);
or U2408 (N_2408,In_886,In_8);
nand U2409 (N_2409,In_431,In_126);
and U2410 (N_2410,In_548,In_208);
nor U2411 (N_2411,In_427,In_638);
and U2412 (N_2412,In_828,In_704);
and U2413 (N_2413,In_281,In_61);
and U2414 (N_2414,In_230,In_714);
nand U2415 (N_2415,In_685,In_656);
nand U2416 (N_2416,In_410,In_831);
nand U2417 (N_2417,In_264,In_84);
and U2418 (N_2418,In_909,In_555);
nand U2419 (N_2419,In_629,In_505);
or U2420 (N_2420,In_834,In_499);
and U2421 (N_2421,In_180,In_666);
nor U2422 (N_2422,In_476,In_887);
or U2423 (N_2423,In_438,In_444);
or U2424 (N_2424,In_995,In_325);
and U2425 (N_2425,In_665,In_549);
and U2426 (N_2426,In_431,In_226);
nand U2427 (N_2427,In_879,In_5);
nor U2428 (N_2428,In_531,In_751);
and U2429 (N_2429,In_853,In_914);
nor U2430 (N_2430,In_576,In_744);
and U2431 (N_2431,In_126,In_635);
and U2432 (N_2432,In_195,In_791);
and U2433 (N_2433,In_420,In_831);
and U2434 (N_2434,In_34,In_750);
and U2435 (N_2435,In_193,In_827);
nand U2436 (N_2436,In_208,In_310);
nand U2437 (N_2437,In_197,In_41);
nand U2438 (N_2438,In_568,In_868);
or U2439 (N_2439,In_783,In_728);
and U2440 (N_2440,In_985,In_594);
nand U2441 (N_2441,In_362,In_851);
and U2442 (N_2442,In_160,In_170);
or U2443 (N_2443,In_753,In_669);
or U2444 (N_2444,In_980,In_380);
or U2445 (N_2445,In_670,In_232);
and U2446 (N_2446,In_968,In_29);
nor U2447 (N_2447,In_583,In_702);
nor U2448 (N_2448,In_755,In_724);
and U2449 (N_2449,In_97,In_737);
nand U2450 (N_2450,In_534,In_233);
nor U2451 (N_2451,In_45,In_261);
nand U2452 (N_2452,In_810,In_678);
nand U2453 (N_2453,In_502,In_10);
and U2454 (N_2454,In_23,In_349);
or U2455 (N_2455,In_904,In_776);
and U2456 (N_2456,In_459,In_690);
xnor U2457 (N_2457,In_332,In_317);
nand U2458 (N_2458,In_278,In_384);
nor U2459 (N_2459,In_503,In_326);
nand U2460 (N_2460,In_999,In_923);
xnor U2461 (N_2461,In_226,In_745);
or U2462 (N_2462,In_604,In_557);
nor U2463 (N_2463,In_667,In_951);
or U2464 (N_2464,In_424,In_111);
or U2465 (N_2465,In_883,In_737);
nand U2466 (N_2466,In_550,In_969);
nand U2467 (N_2467,In_696,In_921);
nor U2468 (N_2468,In_299,In_401);
nand U2469 (N_2469,In_941,In_5);
nand U2470 (N_2470,In_343,In_768);
nor U2471 (N_2471,In_368,In_591);
nand U2472 (N_2472,In_792,In_560);
nand U2473 (N_2473,In_441,In_527);
or U2474 (N_2474,In_80,In_153);
and U2475 (N_2475,In_212,In_433);
xor U2476 (N_2476,In_543,In_426);
or U2477 (N_2477,In_677,In_759);
or U2478 (N_2478,In_770,In_415);
and U2479 (N_2479,In_418,In_550);
or U2480 (N_2480,In_732,In_333);
or U2481 (N_2481,In_244,In_106);
nand U2482 (N_2482,In_301,In_123);
nand U2483 (N_2483,In_11,In_980);
nor U2484 (N_2484,In_89,In_944);
or U2485 (N_2485,In_437,In_574);
nor U2486 (N_2486,In_487,In_577);
or U2487 (N_2487,In_372,In_278);
or U2488 (N_2488,In_940,In_260);
nor U2489 (N_2489,In_208,In_249);
nor U2490 (N_2490,In_718,In_564);
and U2491 (N_2491,In_292,In_654);
and U2492 (N_2492,In_910,In_744);
nor U2493 (N_2493,In_189,In_163);
nor U2494 (N_2494,In_247,In_137);
nor U2495 (N_2495,In_456,In_854);
nand U2496 (N_2496,In_53,In_497);
or U2497 (N_2497,In_64,In_227);
nand U2498 (N_2498,In_165,In_610);
and U2499 (N_2499,In_406,In_529);
or U2500 (N_2500,N_909,N_55);
xnor U2501 (N_2501,N_1832,N_2015);
nand U2502 (N_2502,N_741,N_361);
or U2503 (N_2503,N_1678,N_536);
and U2504 (N_2504,N_1479,N_1209);
nor U2505 (N_2505,N_141,N_1221);
and U2506 (N_2506,N_2234,N_870);
xnor U2507 (N_2507,N_320,N_2191);
or U2508 (N_2508,N_1421,N_1724);
nand U2509 (N_2509,N_1419,N_407);
and U2510 (N_2510,N_968,N_664);
nand U2511 (N_2511,N_1816,N_1723);
nand U2512 (N_2512,N_1972,N_1844);
nand U2513 (N_2513,N_1517,N_1606);
xor U2514 (N_2514,N_2039,N_2192);
nor U2515 (N_2515,N_47,N_610);
and U2516 (N_2516,N_148,N_1040);
or U2517 (N_2517,N_2346,N_1100);
and U2518 (N_2518,N_1371,N_744);
and U2519 (N_2519,N_1064,N_1049);
nor U2520 (N_2520,N_2443,N_1969);
or U2521 (N_2521,N_312,N_1516);
nand U2522 (N_2522,N_178,N_1171);
and U2523 (N_2523,N_2264,N_785);
and U2524 (N_2524,N_318,N_688);
nand U2525 (N_2525,N_1044,N_211);
nand U2526 (N_2526,N_1860,N_669);
or U2527 (N_2527,N_812,N_2085);
or U2528 (N_2528,N_1590,N_699);
or U2529 (N_2529,N_16,N_1332);
nand U2530 (N_2530,N_1938,N_2117);
nand U2531 (N_2531,N_2086,N_108);
nor U2532 (N_2532,N_1306,N_138);
nor U2533 (N_2533,N_74,N_1095);
nor U2534 (N_2534,N_535,N_1668);
nand U2535 (N_2535,N_1304,N_2054);
nor U2536 (N_2536,N_1900,N_853);
nor U2537 (N_2537,N_2223,N_1114);
and U2538 (N_2538,N_1030,N_1005);
nand U2539 (N_2539,N_1250,N_2017);
nor U2540 (N_2540,N_2103,N_1471);
or U2541 (N_2541,N_1023,N_1524);
or U2542 (N_2542,N_1999,N_991);
or U2543 (N_2543,N_2358,N_1817);
nor U2544 (N_2544,N_2477,N_1074);
or U2545 (N_2545,N_2309,N_1689);
and U2546 (N_2546,N_1249,N_2078);
nand U2547 (N_2547,N_1736,N_233);
or U2548 (N_2548,N_303,N_88);
or U2549 (N_2549,N_1592,N_949);
nand U2550 (N_2550,N_1499,N_1174);
and U2551 (N_2551,N_1807,N_366);
nand U2552 (N_2552,N_1551,N_1891);
and U2553 (N_2553,N_251,N_1641);
nand U2554 (N_2554,N_2450,N_1190);
nor U2555 (N_2555,N_90,N_477);
nand U2556 (N_2556,N_534,N_873);
and U2557 (N_2557,N_2132,N_564);
and U2558 (N_2558,N_2109,N_918);
nor U2559 (N_2559,N_2097,N_2025);
and U2560 (N_2560,N_866,N_2096);
and U2561 (N_2561,N_1895,N_2182);
nor U2562 (N_2562,N_1546,N_2059);
and U2563 (N_2563,N_1072,N_1191);
and U2564 (N_2564,N_1486,N_503);
and U2565 (N_2565,N_2325,N_1899);
and U2566 (N_2566,N_2475,N_1485);
or U2567 (N_2567,N_2471,N_2407);
nor U2568 (N_2568,N_1363,N_2386);
nand U2569 (N_2569,N_1926,N_1906);
nor U2570 (N_2570,N_422,N_618);
and U2571 (N_2571,N_1007,N_2359);
and U2572 (N_2572,N_1496,N_302);
and U2573 (N_2573,N_1520,N_983);
nor U2574 (N_2574,N_213,N_2008);
nand U2575 (N_2575,N_1697,N_2427);
or U2576 (N_2576,N_1772,N_624);
and U2577 (N_2577,N_2409,N_1324);
or U2578 (N_2578,N_293,N_379);
and U2579 (N_2579,N_735,N_1016);
and U2580 (N_2580,N_926,N_1967);
nor U2581 (N_2581,N_2490,N_329);
nand U2582 (N_2582,N_808,N_2076);
nor U2583 (N_2583,N_1734,N_2072);
and U2584 (N_2584,N_1325,N_1835);
nor U2585 (N_2585,N_1149,N_1033);
or U2586 (N_2586,N_638,N_523);
nand U2587 (N_2587,N_2499,N_1021);
xor U2588 (N_2588,N_364,N_925);
nor U2589 (N_2589,N_1168,N_520);
and U2590 (N_2590,N_572,N_1995);
or U2591 (N_2591,N_1583,N_892);
or U2592 (N_2592,N_869,N_2374);
and U2593 (N_2593,N_281,N_2379);
and U2594 (N_2594,N_1343,N_1236);
or U2595 (N_2595,N_1003,N_1718);
and U2596 (N_2596,N_201,N_1673);
and U2597 (N_2597,N_1271,N_2020);
nor U2598 (N_2598,N_2394,N_2058);
or U2599 (N_2599,N_1080,N_50);
or U2600 (N_2600,N_182,N_2043);
and U2601 (N_2601,N_758,N_1872);
nor U2602 (N_2602,N_444,N_1686);
and U2603 (N_2603,N_648,N_294);
nor U2604 (N_2604,N_448,N_1438);
nor U2605 (N_2605,N_2300,N_614);
nand U2606 (N_2606,N_1650,N_1894);
nand U2607 (N_2607,N_1411,N_2028);
or U2608 (N_2608,N_1317,N_1046);
xor U2609 (N_2609,N_969,N_1316);
nor U2610 (N_2610,N_418,N_929);
or U2611 (N_2611,N_224,N_159);
and U2612 (N_2612,N_982,N_2316);
or U2613 (N_2613,N_674,N_1312);
or U2614 (N_2614,N_1224,N_1982);
or U2615 (N_2615,N_1701,N_2202);
and U2616 (N_2616,N_537,N_1637);
nor U2617 (N_2617,N_501,N_2426);
xor U2618 (N_2618,N_1410,N_2460);
and U2619 (N_2619,N_867,N_1036);
nor U2620 (N_2620,N_31,N_1199);
or U2621 (N_2621,N_2495,N_401);
nand U2622 (N_2622,N_60,N_2153);
nand U2623 (N_2623,N_1071,N_2254);
nor U2624 (N_2624,N_2297,N_2380);
or U2625 (N_2625,N_1490,N_667);
or U2626 (N_2626,N_830,N_183);
nand U2627 (N_2627,N_1068,N_2046);
or U2628 (N_2628,N_1712,N_451);
nor U2629 (N_2629,N_194,N_166);
nand U2630 (N_2630,N_1179,N_557);
nand U2631 (N_2631,N_204,N_2229);
nor U2632 (N_2632,N_472,N_2323);
nand U2633 (N_2633,N_907,N_1243);
and U2634 (N_2634,N_894,N_1765);
or U2635 (N_2635,N_370,N_1276);
or U2636 (N_2636,N_247,N_615);
nand U2637 (N_2637,N_439,N_794);
and U2638 (N_2638,N_61,N_214);
nand U2639 (N_2639,N_41,N_2286);
or U2640 (N_2640,N_2494,N_945);
and U2641 (N_2641,N_1045,N_732);
or U2642 (N_2642,N_725,N_856);
nor U2643 (N_2643,N_1415,N_1245);
or U2644 (N_2644,N_642,N_298);
nor U2645 (N_2645,N_953,N_2142);
or U2646 (N_2646,N_2252,N_1795);
and U2647 (N_2647,N_1364,N_499);
xnor U2648 (N_2648,N_2240,N_2485);
nand U2649 (N_2649,N_554,N_415);
and U2650 (N_2650,N_2037,N_1634);
and U2651 (N_2651,N_475,N_162);
nand U2652 (N_2652,N_2023,N_193);
or U2653 (N_2653,N_1868,N_241);
and U2654 (N_2654,N_1349,N_510);
xor U2655 (N_2655,N_835,N_1735);
and U2656 (N_2656,N_643,N_286);
nor U2657 (N_2657,N_2127,N_2143);
or U2658 (N_2658,N_2051,N_1567);
and U2659 (N_2659,N_1941,N_124);
nand U2660 (N_2660,N_136,N_10);
or U2661 (N_2661,N_1210,N_2171);
nor U2662 (N_2662,N_2483,N_569);
or U2663 (N_2663,N_541,N_2404);
nor U2664 (N_2664,N_177,N_1172);
nand U2665 (N_2665,N_2105,N_1476);
or U2666 (N_2666,N_459,N_533);
nor U2667 (N_2667,N_2250,N_1561);
and U2668 (N_2668,N_649,N_2417);
and U2669 (N_2669,N_1764,N_2484);
and U2670 (N_2670,N_84,N_1949);
and U2671 (N_2671,N_1834,N_2188);
and U2672 (N_2672,N_2199,N_684);
nor U2673 (N_2673,N_2339,N_762);
or U2674 (N_2674,N_1408,N_728);
nor U2675 (N_2675,N_319,N_2470);
nor U2676 (N_2676,N_1144,N_1556);
and U2677 (N_2677,N_2355,N_2272);
xnor U2678 (N_2678,N_598,N_682);
or U2679 (N_2679,N_463,N_1060);
and U2680 (N_2680,N_2304,N_1744);
or U2681 (N_2681,N_2018,N_1915);
or U2682 (N_2682,N_2480,N_2243);
or U2683 (N_2683,N_553,N_2162);
nand U2684 (N_2684,N_1856,N_12);
and U2685 (N_2685,N_1288,N_1934);
and U2686 (N_2686,N_1390,N_1204);
nor U2687 (N_2687,N_2047,N_930);
or U2688 (N_2688,N_2486,N_1506);
or U2689 (N_2689,N_1294,N_1756);
nand U2690 (N_2690,N_186,N_1258);
or U2691 (N_2691,N_2137,N_726);
nand U2692 (N_2692,N_766,N_710);
nand U2693 (N_2693,N_230,N_81);
and U2694 (N_2694,N_469,N_2237);
nor U2695 (N_2695,N_252,N_1977);
or U2696 (N_2696,N_604,N_2381);
nand U2697 (N_2697,N_1162,N_1278);
or U2698 (N_2698,N_1921,N_36);
or U2699 (N_2699,N_279,N_952);
nand U2700 (N_2700,N_375,N_274);
nand U2701 (N_2701,N_1888,N_1383);
nand U2702 (N_2702,N_305,N_1388);
or U2703 (N_2703,N_2133,N_625);
and U2704 (N_2704,N_1051,N_2242);
or U2705 (N_2705,N_1008,N_482);
or U2706 (N_2706,N_849,N_378);
or U2707 (N_2707,N_2396,N_611);
nor U2708 (N_2708,N_1492,N_2282);
or U2709 (N_2709,N_1424,N_118);
and U2710 (N_2710,N_1662,N_2010);
nand U2711 (N_2711,N_33,N_2399);
and U2712 (N_2712,N_165,N_1035);
nand U2713 (N_2713,N_1439,N_2462);
and U2714 (N_2714,N_1629,N_2392);
nor U2715 (N_2715,N_1802,N_1851);
nor U2716 (N_2716,N_556,N_2126);
and U2717 (N_2717,N_1859,N_1176);
nor U2718 (N_2718,N_964,N_2000);
and U2719 (N_2719,N_357,N_635);
nand U2720 (N_2720,N_528,N_628);
and U2721 (N_2721,N_2401,N_244);
and U2722 (N_2722,N_2172,N_1960);
and U2723 (N_2723,N_2329,N_398);
nand U2724 (N_2724,N_46,N_215);
nor U2725 (N_2725,N_1061,N_217);
and U2726 (N_2726,N_511,N_462);
nand U2727 (N_2727,N_1283,N_683);
or U2728 (N_2728,N_955,N_923);
nand U2729 (N_2729,N_1804,N_1073);
nor U2730 (N_2730,N_546,N_23);
nor U2731 (N_2731,N_56,N_1548);
or U2732 (N_2732,N_2235,N_825);
nor U2733 (N_2733,N_2236,N_2040);
nand U2734 (N_2734,N_2418,N_2330);
or U2735 (N_2735,N_881,N_464);
nor U2736 (N_2736,N_1794,N_1671);
nor U2737 (N_2737,N_91,N_1335);
or U2738 (N_2738,N_1293,N_2413);
or U2739 (N_2739,N_1980,N_5);
nand U2740 (N_2740,N_325,N_587);
nor U2741 (N_2741,N_568,N_43);
and U2742 (N_2742,N_76,N_2310);
or U2743 (N_2743,N_2284,N_2122);
nand U2744 (N_2744,N_339,N_276);
and U2745 (N_2745,N_1790,N_1560);
nand U2746 (N_2746,N_2104,N_1993);
or U2747 (N_2747,N_2313,N_1867);
nand U2748 (N_2748,N_1882,N_1239);
nand U2749 (N_2749,N_59,N_1759);
and U2750 (N_2750,N_342,N_2004);
or U2751 (N_2751,N_496,N_752);
and U2752 (N_2752,N_509,N_863);
or U2753 (N_2753,N_1902,N_2148);
or U2754 (N_2754,N_1090,N_1848);
nand U2755 (N_2755,N_571,N_680);
and U2756 (N_2756,N_2301,N_1052);
or U2757 (N_2757,N_1836,N_54);
and U2758 (N_2758,N_486,N_2440);
nand U2759 (N_2759,N_2140,N_1550);
nor U2760 (N_2760,N_2389,N_153);
and U2761 (N_2761,N_2257,N_2263);
nor U2762 (N_2762,N_944,N_1101);
or U2763 (N_2763,N_282,N_2403);
and U2764 (N_2764,N_440,N_2449);
nor U2765 (N_2765,N_2273,N_310);
nand U2766 (N_2766,N_723,N_344);
and U2767 (N_2767,N_1357,N_1809);
nor U2768 (N_2768,N_2150,N_39);
nand U2769 (N_2769,N_35,N_990);
or U2770 (N_2770,N_1544,N_97);
or U2771 (N_2771,N_107,N_1392);
nand U2772 (N_2772,N_1373,N_2186);
or U2773 (N_2773,N_1400,N_1493);
nor U2774 (N_2774,N_714,N_1303);
nor U2775 (N_2775,N_295,N_2245);
nand U2776 (N_2776,N_701,N_268);
nand U2777 (N_2777,N_1473,N_1301);
or U2778 (N_2778,N_1922,N_784);
nor U2779 (N_2779,N_1495,N_961);
or U2780 (N_2780,N_2239,N_1222);
nand U2781 (N_2781,N_1311,N_271);
nand U2782 (N_2782,N_1394,N_210);
xnor U2783 (N_2783,N_1564,N_421);
and U2784 (N_2784,N_1553,N_103);
nor U2785 (N_2785,N_644,N_786);
nand U2786 (N_2786,N_872,N_1097);
and U2787 (N_2787,N_1793,N_1273);
nor U2788 (N_2788,N_1151,N_896);
nor U2789 (N_2789,N_1079,N_2084);
and U2790 (N_2790,N_542,N_2368);
nand U2791 (N_2791,N_309,N_2110);
nand U2792 (N_2792,N_2164,N_2168);
and U2793 (N_2793,N_678,N_780);
or U2794 (N_2794,N_1542,N_979);
or U2795 (N_2795,N_1808,N_629);
or U2796 (N_2796,N_1569,N_1092);
nand U2797 (N_2797,N_2479,N_1298);
and U2798 (N_2798,N_1990,N_670);
nor U2799 (N_2799,N_1015,N_363);
and U2800 (N_2800,N_1540,N_1070);
nand U2801 (N_2801,N_2094,N_489);
nor U2802 (N_2802,N_747,N_1050);
or U2803 (N_2803,N_1219,N_694);
or U2804 (N_2804,N_1720,N_527);
and U2805 (N_2805,N_1797,N_933);
nor U2806 (N_2806,N_1511,N_2189);
and U2807 (N_2807,N_592,N_2146);
or U2808 (N_2808,N_1633,N_1212);
xor U2809 (N_2809,N_1452,N_1164);
nor U2810 (N_2810,N_381,N_1346);
or U2811 (N_2811,N_1919,N_2038);
and U2812 (N_2812,N_284,N_150);
and U2813 (N_2813,N_878,N_2154);
and U2814 (N_2814,N_2217,N_1274);
nor U2815 (N_2815,N_842,N_1231);
and U2816 (N_2816,N_1541,N_1973);
nor U2817 (N_2817,N_1132,N_57);
nand U2818 (N_2818,N_919,N_1643);
nand U2819 (N_2819,N_1055,N_1063);
nand U2820 (N_2820,N_1806,N_538);
nand U2821 (N_2821,N_2241,N_597);
and U2822 (N_2822,N_1048,N_1351);
and U2823 (N_2823,N_2074,N_1375);
and U2824 (N_2824,N_994,N_2402);
nor U2825 (N_2825,N_1767,N_1896);
or U2826 (N_2826,N_770,N_1713);
or U2827 (N_2827,N_733,N_1122);
and U2828 (N_2828,N_1975,N_1255);
nand U2829 (N_2829,N_131,N_1126);
or U2830 (N_2830,N_1943,N_351);
or U2831 (N_2831,N_1710,N_2491);
nor U2832 (N_2832,N_651,N_2487);
and U2833 (N_2833,N_2002,N_2408);
nand U2834 (N_2834,N_2036,N_2395);
or U2835 (N_2835,N_973,N_754);
nor U2836 (N_2836,N_803,N_621);
and U2837 (N_2837,N_1321,N_17);
or U2838 (N_2838,N_142,N_704);
xnor U2839 (N_2839,N_601,N_1088);
and U2840 (N_2840,N_2466,N_291);
or U2841 (N_2841,N_2121,N_2388);
nand U2842 (N_2842,N_1200,N_703);
nor U2843 (N_2843,N_313,N_1109);
and U2844 (N_2844,N_876,N_1398);
nand U2845 (N_2845,N_2174,N_2071);
and U2846 (N_2846,N_1897,N_436);
nand U2847 (N_2847,N_646,N_1406);
or U2848 (N_2848,N_700,N_2152);
or U2849 (N_2849,N_2377,N_2033);
nor U2850 (N_2850,N_1676,N_1315);
or U2851 (N_2851,N_640,N_965);
nor U2852 (N_2852,N_345,N_169);
nand U2853 (N_2853,N_1205,N_1578);
nor U2854 (N_2854,N_1066,N_2414);
nor U2855 (N_2855,N_898,N_2442);
nand U2856 (N_2856,N_2412,N_709);
and U2857 (N_2857,N_2489,N_966);
nor U2858 (N_2858,N_1159,N_2014);
nor U2859 (N_2859,N_831,N_775);
nor U2860 (N_2860,N_1038,N_2225);
or U2861 (N_2861,N_1111,N_880);
and U2862 (N_2862,N_1874,N_1879);
nor U2863 (N_2863,N_393,N_340);
nand U2864 (N_2864,N_1218,N_137);
nor U2865 (N_2865,N_44,N_1956);
and U2866 (N_2866,N_1247,N_1773);
nand U2867 (N_2867,N_290,N_2361);
or U2868 (N_2868,N_696,N_299);
and U2869 (N_2869,N_995,N_2067);
or U2870 (N_2870,N_2276,N_1233);
or U2871 (N_2871,N_1024,N_1732);
nor U2872 (N_2872,N_1456,N_1427);
and U2873 (N_2873,N_1167,N_1730);
or U2874 (N_2874,N_253,N_539);
and U2875 (N_2875,N_1195,N_1057);
nor U2876 (N_2876,N_2131,N_2201);
nand U2877 (N_2877,N_396,N_2228);
nor U2878 (N_2878,N_2167,N_2093);
or U2879 (N_2879,N_788,N_1883);
or U2880 (N_2880,N_1491,N_1453);
or U2881 (N_2881,N_1370,N_1729);
nand U2882 (N_2882,N_374,N_2424);
nand U2883 (N_2883,N_2129,N_1534);
nor U2884 (N_2884,N_1535,N_1461);
and U2885 (N_2885,N_2367,N_1138);
or U2886 (N_2886,N_2344,N_117);
and U2887 (N_2887,N_630,N_782);
and U2888 (N_2888,N_481,N_2125);
and U2889 (N_2889,N_1314,N_2261);
nor U2890 (N_2890,N_425,N_2324);
and U2891 (N_2891,N_1620,N_1649);
or U2892 (N_2892,N_174,N_2342);
and U2893 (N_2893,N_1269,N_1465);
and U2894 (N_2894,N_2215,N_1876);
or U2895 (N_2895,N_1353,N_935);
or U2896 (N_2896,N_1225,N_2177);
xor U2897 (N_2897,N_388,N_2102);
and U2898 (N_2898,N_795,N_962);
and U2899 (N_2899,N_372,N_94);
nor U2900 (N_2900,N_1358,N_341);
and U2901 (N_2901,N_1474,N_1387);
nand U2902 (N_2902,N_1979,N_1839);
and U2903 (N_2903,N_2308,N_1158);
nand U2904 (N_2904,N_2351,N_792);
and U2905 (N_2905,N_473,N_225);
or U2906 (N_2906,N_2376,N_42);
nand U2907 (N_2907,N_1509,N_13);
nand U2908 (N_2908,N_2322,N_445);
or U2909 (N_2909,N_195,N_307);
or U2910 (N_2910,N_809,N_63);
and U2911 (N_2911,N_526,N_855);
nor U2912 (N_2912,N_200,N_1638);
or U2913 (N_2913,N_1340,N_921);
or U2914 (N_2914,N_1595,N_2317);
and U2915 (N_2915,N_2139,N_2283);
or U2916 (N_2916,N_2378,N_1426);
nor U2917 (N_2917,N_367,N_2292);
and U2918 (N_2918,N_358,N_1422);
or U2919 (N_2919,N_1266,N_517);
or U2920 (N_2920,N_1001,N_665);
and U2921 (N_2921,N_2218,N_978);
or U2922 (N_2922,N_1664,N_205);
and U2923 (N_2923,N_1572,N_1945);
or U2924 (N_2924,N_2472,N_1347);
nor U2925 (N_2925,N_765,N_330);
or U2926 (N_2926,N_2410,N_1589);
nor U2927 (N_2927,N_58,N_257);
nor U2928 (N_2928,N_1570,N_796);
and U2929 (N_2929,N_843,N_1536);
nand U2930 (N_2930,N_1531,N_206);
nand U2931 (N_2931,N_1965,N_2312);
nand U2932 (N_2932,N_963,N_2249);
nand U2933 (N_2933,N_1955,N_161);
or U2934 (N_2934,N_750,N_466);
and U2935 (N_2935,N_237,N_2269);
or U2936 (N_2936,N_1004,N_1418);
nand U2937 (N_2937,N_1870,N_851);
nand U2938 (N_2938,N_1705,N_2362);
and U2939 (N_2939,N_2198,N_327);
nand U2940 (N_2940,N_2482,N_52);
or U2941 (N_2941,N_404,N_2016);
xor U2942 (N_2942,N_1821,N_1268);
or U2943 (N_2943,N_1450,N_1291);
nor U2944 (N_2944,N_1157,N_2030);
nor U2945 (N_2945,N_164,N_1386);
nand U2946 (N_2946,N_1336,N_2256);
nor U2947 (N_2947,N_8,N_356);
nand U2948 (N_2948,N_2306,N_145);
nor U2949 (N_2949,N_685,N_1681);
nor U2950 (N_2950,N_347,N_1423);
nor U2951 (N_2951,N_127,N_1596);
nor U2952 (N_2952,N_810,N_838);
nor U2953 (N_2953,N_975,N_45);
or U2954 (N_2954,N_1295,N_1329);
nor U2955 (N_2955,N_829,N_987);
or U2956 (N_2956,N_560,N_260);
and U2957 (N_2957,N_981,N_111);
nand U2958 (N_2958,N_612,N_906);
nand U2959 (N_2959,N_68,N_191);
nand U2960 (N_2960,N_588,N_729);
and U2961 (N_2961,N_1402,N_1665);
or U2962 (N_2962,N_2405,N_811);
and U2963 (N_2963,N_1510,N_2247);
nor U2964 (N_2964,N_1555,N_460);
nor U2965 (N_2965,N_2314,N_1594);
and U2966 (N_2966,N_900,N_2145);
nor U2967 (N_2967,N_879,N_1573);
and U2968 (N_2968,N_751,N_2173);
or U2969 (N_2969,N_1263,N_755);
and U2970 (N_2970,N_1369,N_650);
nor U2971 (N_2971,N_1328,N_428);
and U2972 (N_2972,N_135,N_232);
nor U2973 (N_2973,N_2208,N_37);
and U2974 (N_2974,N_2034,N_1928);
or U2975 (N_2975,N_1580,N_1431);
and U2976 (N_2976,N_140,N_793);
nor U2977 (N_2977,N_2357,N_2348);
nand U2978 (N_2978,N_1103,N_1350);
or U2979 (N_2979,N_157,N_972);
nand U2980 (N_2980,N_1488,N_2387);
nand U2981 (N_2981,N_1339,N_852);
nand U2982 (N_2982,N_394,N_767);
and U2983 (N_2983,N_333,N_2406);
nand U2984 (N_2984,N_1500,N_1523);
and U2985 (N_2985,N_616,N_1841);
and U2986 (N_2986,N_1141,N_889);
nor U2987 (N_2987,N_2353,N_1568);
and U2988 (N_2988,N_1749,N_671);
or U2989 (N_2989,N_1796,N_1365);
nand U2990 (N_2990,N_483,N_218);
or U2991 (N_2991,N_1763,N_1933);
or U2992 (N_2992,N_673,N_1762);
and U2993 (N_2993,N_1672,N_2373);
nor U2994 (N_2994,N_1241,N_1611);
or U2995 (N_2995,N_2248,N_2013);
nand U2996 (N_2996,N_940,N_430);
and U2997 (N_2997,N_278,N_2032);
or U2998 (N_2998,N_1319,N_1711);
nor U2999 (N_2999,N_66,N_904);
or U3000 (N_3000,N_662,N_2463);
and U3001 (N_3001,N_2437,N_1942);
xnor U3002 (N_3002,N_2092,N_160);
and U3003 (N_3003,N_549,N_154);
or U3004 (N_3004,N_409,N_121);
or U3005 (N_3005,N_759,N_854);
nand U3006 (N_3006,N_304,N_653);
and U3007 (N_3007,N_1135,N_128);
nand U3008 (N_3008,N_2205,N_115);
and U3009 (N_3009,N_1147,N_1302);
and U3010 (N_3010,N_1521,N_822);
or U3011 (N_3011,N_1613,N_2327);
and U3012 (N_3012,N_1939,N_2400);
or U3013 (N_3013,N_2089,N_2082);
nand U3014 (N_3014,N_1626,N_1207);
and U3015 (N_3015,N_605,N_171);
and U3016 (N_3016,N_1805,N_986);
nand U3017 (N_3017,N_24,N_1320);
nor U3018 (N_3018,N_2343,N_1905);
xor U3019 (N_3019,N_2451,N_20);
nor U3020 (N_3020,N_1039,N_2183);
nand U3021 (N_3021,N_1012,N_816);
nand U3022 (N_3022,N_1522,N_779);
and U3023 (N_3023,N_753,N_2385);
or U3024 (N_3024,N_1475,N_1885);
and U3025 (N_3025,N_2098,N_529);
or U3026 (N_3026,N_1760,N_1916);
or U3027 (N_3027,N_2455,N_1498);
nand U3028 (N_3028,N_1997,N_1034);
and U3029 (N_3029,N_1690,N_864);
or U3030 (N_3030,N_1472,N_658);
or U3031 (N_3031,N_1670,N_1625);
nand U3032 (N_3032,N_941,N_657);
nand U3033 (N_3033,N_420,N_1920);
nand U3034 (N_3034,N_1624,N_1480);
or U3035 (N_3035,N_155,N_389);
nand U3036 (N_3036,N_577,N_2060);
or U3037 (N_3037,N_406,N_2492);
nor U3038 (N_3038,N_1525,N_1166);
or U3039 (N_3039,N_2302,N_2279);
nand U3040 (N_3040,N_1602,N_2433);
or U3041 (N_3041,N_262,N_637);
nor U3042 (N_3042,N_1047,N_936);
or U3043 (N_3043,N_1917,N_561);
nand U3044 (N_3044,N_1507,N_1947);
nor U3045 (N_3045,N_2001,N_73);
nor U3046 (N_3046,N_1133,N_1622);
or U3047 (N_3047,N_748,N_740);
or U3048 (N_3048,N_769,N_2114);
nor U3049 (N_3049,N_606,N_2195);
or U3050 (N_3050,N_2461,N_1177);
nand U3051 (N_3051,N_1429,N_116);
or U3052 (N_3052,N_1703,N_2444);
or U3053 (N_3053,N_273,N_1468);
and U3054 (N_3054,N_660,N_64);
or U3055 (N_3055,N_1505,N_819);
or U3056 (N_3056,N_661,N_806);
nand U3057 (N_3057,N_424,N_967);
nand U3058 (N_3058,N_40,N_1027);
or U3059 (N_3059,N_267,N_176);
nand U3060 (N_3060,N_1444,N_1441);
nand U3061 (N_3061,N_858,N_1186);
nor U3062 (N_3062,N_1214,N_300);
nor U3063 (N_3063,N_419,N_4);
nor U3064 (N_3064,N_1372,N_839);
and U3065 (N_3065,N_2285,N_1183);
and U3066 (N_3066,N_1069,N_603);
and U3067 (N_3067,N_708,N_1840);
nand U3068 (N_3068,N_1404,N_1675);
nor U3069 (N_3069,N_226,N_2035);
nor U3070 (N_3070,N_2147,N_1434);
and U3071 (N_3071,N_434,N_1009);
and U3072 (N_3072,N_1552,N_1238);
nand U3073 (N_3073,N_65,N_1175);
or U3074 (N_3074,N_681,N_452);
or U3075 (N_3075,N_435,N_2166);
nor U3076 (N_3076,N_959,N_738);
nand U3077 (N_3077,N_1484,N_992);
nand U3078 (N_3078,N_1827,N_1693);
or U3079 (N_3079,N_456,N_1850);
nor U3080 (N_3080,N_29,N_504);
nor U3081 (N_3081,N_1184,N_1612);
nor U3082 (N_3082,N_532,N_934);
nor U3083 (N_3083,N_2288,N_2298);
nor U3084 (N_3084,N_380,N_718);
and U3085 (N_3085,N_508,N_1615);
nand U3086 (N_3086,N_1076,N_1362);
nand U3087 (N_3087,N_882,N_1477);
nor U3088 (N_3088,N_1988,N_75);
and U3089 (N_3089,N_1102,N_173);
nand U3090 (N_3090,N_2419,N_2005);
nand U3091 (N_3091,N_1019,N_840);
nor U3092 (N_3092,N_1181,N_2022);
xor U3093 (N_3093,N_1285,N_1768);
or U3094 (N_3094,N_89,N_1246);
or U3095 (N_3095,N_875,N_326);
nor U3096 (N_3096,N_437,N_1748);
and U3097 (N_3097,N_1950,N_287);
nand U3098 (N_3098,N_1140,N_112);
and U3099 (N_3099,N_807,N_7);
nand U3100 (N_3100,N_1682,N_2439);
nor U3101 (N_3101,N_1296,N_296);
or U3102 (N_3102,N_619,N_515);
or U3103 (N_3103,N_1374,N_353);
or U3104 (N_3104,N_1774,N_1692);
or U3105 (N_3105,N_717,N_1547);
and U3106 (N_3106,N_2345,N_2119);
or U3107 (N_3107,N_1861,N_1907);
or U3108 (N_3108,N_147,N_2299);
nand U3109 (N_3109,N_1430,N_861);
and U3110 (N_3110,N_1989,N_2197);
and U3111 (N_3111,N_382,N_1694);
nor U3112 (N_3112,N_920,N_827);
nor U3113 (N_3113,N_847,N_332);
or U3114 (N_3114,N_2423,N_513);
nor U3115 (N_3115,N_911,N_1619);
or U3116 (N_3116,N_1978,N_1300);
or U3117 (N_3117,N_976,N_390);
or U3118 (N_3118,N_1725,N_168);
nor U3119 (N_3119,N_402,N_126);
nand U3120 (N_3120,N_1065,N_306);
nor U3121 (N_3121,N_1124,N_1259);
or U3122 (N_3122,N_2128,N_1341);
or U3123 (N_3123,N_1514,N_1952);
nor U3124 (N_3124,N_636,N_1110);
and U3125 (N_3125,N_1843,N_1944);
nor U3126 (N_3126,N_1537,N_1599);
nand U3127 (N_3127,N_1818,N_2438);
and U3128 (N_3128,N_1881,N_1931);
or U3129 (N_3129,N_1155,N_2422);
nand U3130 (N_3130,N_156,N_654);
and U3131 (N_3131,N_1337,N_1432);
nor U3132 (N_3132,N_1575,N_2333);
or U3133 (N_3133,N_512,N_1202);
nand U3134 (N_3134,N_100,N_1446);
nor U3135 (N_3135,N_652,N_540);
nor U3136 (N_3136,N_1313,N_245);
nor U3137 (N_3137,N_1152,N_1983);
and U3138 (N_3138,N_1728,N_413);
nor U3139 (N_3139,N_2227,N_2175);
and U3140 (N_3140,N_1669,N_586);
and U3141 (N_3141,N_2099,N_931);
or U3142 (N_3142,N_1636,N_675);
or U3143 (N_3143,N_641,N_152);
nand U3144 (N_3144,N_1251,N_742);
nand U3145 (N_3145,N_689,N_584);
and U3146 (N_3146,N_1139,N_817);
nand U3147 (N_3147,N_2200,N_454);
and U3148 (N_3148,N_2398,N_248);
nand U3149 (N_3149,N_1267,N_1745);
or U3150 (N_3150,N_2352,N_1813);
or U3151 (N_3151,N_426,N_1085);
nor U3152 (N_3152,N_774,N_1104);
xnor U3153 (N_3153,N_2222,N_209);
nand U3154 (N_3154,N_1688,N_87);
nand U3155 (N_3155,N_2185,N_1397);
nor U3156 (N_3156,N_1260,N_565);
and U3157 (N_3157,N_1451,N_802);
and U3158 (N_3158,N_1515,N_1610);
or U3159 (N_3159,N_1959,N_1344);
or U3160 (N_3160,N_2184,N_1529);
or U3161 (N_3161,N_105,N_228);
xnor U3162 (N_3162,N_1252,N_1755);
and U3163 (N_3163,N_397,N_1277);
and U3164 (N_3164,N_1766,N_1189);
or U3165 (N_3165,N_338,N_1799);
nor U3166 (N_3166,N_2064,N_897);
and U3167 (N_3167,N_1654,N_423);
nand U3168 (N_3168,N_492,N_832);
and U3169 (N_3169,N_1025,N_582);
and U3170 (N_3170,N_570,N_2334);
nand U3171 (N_3171,N_70,N_2347);
nor U3172 (N_3172,N_1041,N_1742);
and U3173 (N_3173,N_2213,N_1837);
nor U3174 (N_3174,N_2270,N_999);
and U3175 (N_3175,N_1010,N_1828);
and U3176 (N_3176,N_432,N_1940);
nor U3177 (N_3177,N_1632,N_2070);
nor U3178 (N_3178,N_1437,N_497);
nor U3179 (N_3179,N_716,N_1777);
and U3180 (N_3180,N_2294,N_1962);
and U3181 (N_3181,N_734,N_1165);
nor U3182 (N_3182,N_102,N_1865);
and U3183 (N_3183,N_151,N_2458);
and U3184 (N_3184,N_1235,N_95);
or U3185 (N_3185,N_1953,N_905);
nor U3186 (N_3186,N_288,N_1826);
nor U3187 (N_3187,N_1858,N_170);
nor U3188 (N_3188,N_2331,N_34);
or U3189 (N_3189,N_1501,N_384);
nor U3190 (N_3190,N_1017,N_1478);
nand U3191 (N_3191,N_2265,N_1811);
nor U3192 (N_3192,N_2080,N_914);
nor U3193 (N_3193,N_1984,N_948);
and U3194 (N_3194,N_1433,N_595);
nand U3195 (N_3195,N_679,N_2436);
and U3196 (N_3196,N_1623,N_1640);
or U3197 (N_3197,N_883,N_1708);
nand U3198 (N_3198,N_2268,N_1310);
and U3199 (N_3199,N_1769,N_773);
and U3200 (N_3200,N_429,N_1914);
and U3201 (N_3201,N_391,N_502);
nor U3202 (N_3202,N_922,N_706);
or U3203 (N_3203,N_1557,N_1530);
or U3204 (N_3204,N_1771,N_2163);
or U3205 (N_3205,N_2291,N_495);
and U3206 (N_3206,N_222,N_2049);
nor U3207 (N_3207,N_745,N_22);
and U3208 (N_3208,N_596,N_1890);
nor U3209 (N_3209,N_441,N_1089);
and U3210 (N_3210,N_1014,N_1699);
and U3211 (N_3211,N_1206,N_223);
nand U3212 (N_3212,N_845,N_1182);
nor U3213 (N_3213,N_1715,N_297);
nand U3214 (N_3214,N_2212,N_1123);
nor U3215 (N_3215,N_790,N_1871);
nor U3216 (N_3216,N_1377,N_272);
nor U3217 (N_3217,N_461,N_988);
and U3218 (N_3218,N_1677,N_146);
nor U3219 (N_3219,N_566,N_924);
nor U3220 (N_3220,N_2180,N_631);
nor U3221 (N_3221,N_550,N_26);
and U3222 (N_3222,N_493,N_2441);
nand U3223 (N_3223,N_1792,N_1420);
or U3224 (N_3224,N_106,N_2029);
and U3225 (N_3225,N_2216,N_1658);
nor U3226 (N_3226,N_1630,N_583);
nor U3227 (N_3227,N_2391,N_119);
or U3228 (N_3228,N_1937,N_1395);
and U3229 (N_3229,N_943,N_763);
and U3230 (N_3230,N_1812,N_559);
nand U3231 (N_3231,N_2077,N_814);
or U3232 (N_3232,N_263,N_2393);
nand U3233 (N_3233,N_443,N_1845);
nor U3234 (N_3234,N_2384,N_110);
nor U3235 (N_3235,N_1459,N_1161);
and U3236 (N_3236,N_1645,N_719);
and U3237 (N_3237,N_1743,N_1908);
and U3238 (N_3238,N_1929,N_506);
and U3239 (N_3239,N_686,N_656);
nor U3240 (N_3240,N_2335,N_6);
nor U3241 (N_3241,N_1948,N_2365);
nand U3242 (N_3242,N_283,N_576);
nor U3243 (N_3243,N_627,N_346);
and U3244 (N_3244,N_371,N_1783);
nor U3245 (N_3245,N_349,N_857);
nand U3246 (N_3246,N_518,N_828);
nand U3247 (N_3247,N_1925,N_369);
and U3248 (N_3248,N_1576,N_2214);
or U3249 (N_3249,N_545,N_1457);
or U3250 (N_3250,N_1930,N_2063);
or U3251 (N_3251,N_1011,N_932);
or U3252 (N_3252,N_1820,N_1120);
nor U3253 (N_3253,N_711,N_1700);
or U3254 (N_3254,N_1563,N_1254);
nor U3255 (N_3255,N_2190,N_242);
and U3256 (N_3256,N_702,N_1887);
nand U3257 (N_3257,N_2041,N_134);
and U3258 (N_3258,N_1440,N_144);
nor U3259 (N_3259,N_1062,N_980);
or U3260 (N_3260,N_30,N_2048);
nor U3261 (N_3261,N_985,N_521);
nor U3262 (N_3262,N_1918,N_1838);
or U3263 (N_3263,N_101,N_2267);
or U3264 (N_3264,N_639,N_2045);
nor U3265 (N_3265,N_1425,N_947);
nor U3266 (N_3266,N_977,N_1083);
nand U3267 (N_3267,N_2468,N_871);
or U3268 (N_3268,N_2246,N_899);
or U3269 (N_3269,N_1750,N_859);
nand U3270 (N_3270,N_1878,N_623);
and U3271 (N_3271,N_691,N_1188);
or U3272 (N_3272,N_2130,N_1581);
or U3273 (N_3273,N_573,N_1361);
and U3274 (N_3274,N_2155,N_833);
nor U3275 (N_3275,N_1558,N_1121);
nor U3276 (N_3276,N_2446,N_2160);
nor U3277 (N_3277,N_2179,N_551);
nand U3278 (N_3278,N_198,N_1801);
nand U3279 (N_3279,N_1290,N_465);
nand U3280 (N_3280,N_1145,N_715);
nand U3281 (N_3281,N_1467,N_2055);
xnor U3282 (N_3282,N_1497,N_798);
and U3283 (N_3283,N_181,N_1775);
and U3284 (N_3284,N_474,N_2011);
or U3285 (N_3285,N_2293,N_324);
nand U3286 (N_3286,N_96,N_1265);
nor U3287 (N_3287,N_2303,N_1683);
and U3288 (N_3288,N_1758,N_1761);
nand U3289 (N_3289,N_2425,N_2083);
nand U3290 (N_3290,N_163,N_314);
or U3291 (N_3291,N_395,N_1869);
nand U3292 (N_3292,N_613,N_1607);
or U3293 (N_3293,N_1366,N_2112);
and U3294 (N_3294,N_392,N_996);
nand U3295 (N_3295,N_1215,N_1108);
and U3296 (N_3296,N_2354,N_1256);
or U3297 (N_3297,N_301,N_1322);
or U3298 (N_3298,N_1849,N_1609);
nand U3299 (N_3299,N_1852,N_1078);
and U3300 (N_3300,N_149,N_1787);
and U3301 (N_3301,N_1788,N_1413);
or U3302 (N_3302,N_348,N_311);
and U3303 (N_3303,N_25,N_1107);
nand U3304 (N_3304,N_2411,N_1873);
and U3305 (N_3305,N_1825,N_1185);
nor U3306 (N_3306,N_1604,N_2497);
or U3307 (N_3307,N_1904,N_2026);
nor U3308 (N_3308,N_1308,N_543);
or U3309 (N_3309,N_1992,N_1257);
and U3310 (N_3310,N_2371,N_2372);
or U3311 (N_3311,N_2124,N_739);
or U3312 (N_3312,N_1779,N_2465);
or U3313 (N_3313,N_1091,N_731);
nor U3314 (N_3314,N_2341,N_331);
nor U3315 (N_3315,N_484,N_1903);
nand U3316 (N_3316,N_1635,N_1143);
and U3317 (N_3317,N_1985,N_360);
nor U3318 (N_3318,N_316,N_2118);
or U3319 (N_3319,N_2219,N_1464);
nor U3320 (N_3320,N_355,N_2459);
or U3321 (N_3321,N_1528,N_1156);
nand U3322 (N_3322,N_1600,N_487);
nor U3323 (N_3323,N_2369,N_1);
nand U3324 (N_3324,N_2024,N_1416);
and U3325 (N_3325,N_2100,N_1512);
and U3326 (N_3326,N_1652,N_1180);
nor U3327 (N_3327,N_1974,N_2176);
and U3328 (N_3328,N_1084,N_1674);
nor U3329 (N_3329,N_1667,N_500);
or U3330 (N_3330,N_172,N_602);
nand U3331 (N_3331,N_77,N_1884);
nand U3332 (N_3332,N_1407,N_471);
nor U3333 (N_3333,N_1327,N_585);
nor U3334 (N_3334,N_1318,N_2068);
or U3335 (N_3335,N_727,N_2113);
and U3336 (N_3336,N_756,N_1719);
or U3337 (N_3337,N_2457,N_2136);
nor U3338 (N_3338,N_449,N_1717);
or U3339 (N_3339,N_1532,N_1227);
nor U3340 (N_3340,N_1237,N_129);
and U3341 (N_3341,N_2,N_903);
or U3342 (N_3342,N_818,N_2445);
nor U3343 (N_3343,N_1707,N_321);
nand U3344 (N_3344,N_1131,N_2111);
and U3345 (N_3345,N_2452,N_1687);
nor U3346 (N_3346,N_1264,N_713);
nor U3347 (N_3347,N_207,N_1880);
or U3348 (N_3348,N_2296,N_1330);
or U3349 (N_3349,N_1966,N_2107);
nand U3350 (N_3350,N_399,N_530);
nor U3351 (N_3351,N_663,N_1289);
or U3352 (N_3352,N_1483,N_249);
and U3353 (N_3353,N_1448,N_2165);
nor U3354 (N_3354,N_950,N_721);
and U3355 (N_3355,N_1642,N_11);
nand U3356 (N_3356,N_1059,N_2087);
and U3357 (N_3357,N_761,N_937);
nor U3358 (N_3358,N_768,N_80);
nand U3359 (N_3359,N_83,N_781);
and U3360 (N_3360,N_1391,N_376);
or U3361 (N_3361,N_901,N_946);
nor U3362 (N_3362,N_659,N_787);
or U3363 (N_3363,N_69,N_722);
nor U3364 (N_3364,N_1739,N_2178);
nor U3365 (N_3365,N_797,N_1627);
nand U3366 (N_3366,N_1043,N_408);
or U3367 (N_3367,N_1193,N_1831);
nand U3368 (N_3368,N_1651,N_1539);
or U3369 (N_3369,N_1617,N_1740);
and U3370 (N_3370,N_2340,N_1733);
or U3371 (N_3371,N_2115,N_666);
nor U3372 (N_3372,N_1401,N_912);
or U3373 (N_3373,N_2474,N_1234);
nor U3374 (N_3374,N_1292,N_562);
nand U3375 (N_3375,N_1932,N_264);
nand U3376 (N_3376,N_846,N_104);
or U3377 (N_3377,N_1798,N_2007);
or U3378 (N_3378,N_1230,N_2290);
nand U3379 (N_3379,N_1455,N_2253);
nand U3380 (N_3380,N_1994,N_2170);
or U3381 (N_3381,N_1746,N_1248);
or U3382 (N_3382,N_2251,N_485);
or U3383 (N_3383,N_1389,N_2448);
and U3384 (N_3384,N_626,N_2328);
xnor U3385 (N_3385,N_2390,N_19);
and U3386 (N_3386,N_478,N_219);
nand U3387 (N_3387,N_1936,N_1533);
nor U3388 (N_3388,N_2009,N_2203);
nor U3389 (N_3389,N_1855,N_1655);
nor U3390 (N_3390,N_730,N_2434);
or U3391 (N_3391,N_1223,N_2363);
or U3392 (N_3392,N_1201,N_1454);
or U3393 (N_3393,N_971,N_1196);
nor U3394 (N_3394,N_1137,N_1067);
nor U3395 (N_3395,N_2196,N_455);
nand U3396 (N_3396,N_1449,N_289);
and U3397 (N_3397,N_86,N_383);
nand U3398 (N_3398,N_1663,N_668);
xnor U3399 (N_3399,N_1696,N_258);
and U3400 (N_3400,N_771,N_877);
or U3401 (N_3401,N_1470,N_1913);
nand U3402 (N_3402,N_1020,N_1657);
nand U3403 (N_3403,N_377,N_1447);
and U3404 (N_3404,N_608,N_2467);
and U3405 (N_3405,N_1000,N_1220);
nor U3406 (N_3406,N_1815,N_958);
nand U3407 (N_3407,N_231,N_2056);
and U3408 (N_3408,N_53,N_902);
nor U3409 (N_3409,N_359,N_2275);
nor U3410 (N_3410,N_1099,N_2420);
nor U3411 (N_3411,N_1814,N_1428);
or U3412 (N_3412,N_1886,N_837);
nand U3413 (N_3413,N_1776,N_801);
or U3414 (N_3414,N_760,N_2271);
or U3415 (N_3415,N_1414,N_2289);
nand U3416 (N_3416,N_1543,N_2478);
nand U3417 (N_3417,N_438,N_1889);
or U3418 (N_3418,N_1704,N_2336);
or U3419 (N_3419,N_1819,N_199);
or U3420 (N_3420,N_476,N_387);
nand U3421 (N_3421,N_202,N_563);
nand U3422 (N_3422,N_1566,N_2416);
or U3423 (N_3423,N_2194,N_1571);
and U3424 (N_3424,N_67,N_1462);
or U3425 (N_3425,N_707,N_2226);
or U3426 (N_3426,N_479,N_1823);
and U3427 (N_3427,N_593,N_524);
or U3428 (N_3428,N_2428,N_269);
nor U3429 (N_3429,N_2315,N_622);
and U3430 (N_3430,N_32,N_2320);
nor U3431 (N_3431,N_412,N_1709);
nor U3432 (N_3432,N_1081,N_1026);
and U3433 (N_3433,N_1784,N_1598);
nor U3434 (N_3434,N_1549,N_824);
and U3435 (N_3435,N_1396,N_1909);
or U3436 (N_3436,N_1229,N_1280);
nor U3437 (N_3437,N_1741,N_1661);
nor U3438 (N_3438,N_1118,N_1096);
or U3439 (N_3439,N_2211,N_1299);
nand U3440 (N_3440,N_2151,N_1970);
xor U3441 (N_3441,N_2231,N_1098);
or U3442 (N_3442,N_1504,N_1309);
xnor U3443 (N_3443,N_1287,N_1379);
and U3444 (N_3444,N_2021,N_328);
nand U3445 (N_3445,N_1232,N_417);
nor U3446 (N_3446,N_48,N_2259);
and U3447 (N_3447,N_1042,N_2311);
nand U3448 (N_3448,N_488,N_490);
and U3449 (N_3449,N_507,N_1142);
and U3450 (N_3450,N_1757,N_1013);
xor U3451 (N_3451,N_2057,N_2027);
or U3452 (N_3452,N_2366,N_575);
and U3453 (N_3453,N_1579,N_1603);
nor U3454 (N_3454,N_1698,N_1731);
nand U3455 (N_3455,N_1112,N_720);
or U3456 (N_3456,N_373,N_1593);
and U3457 (N_3457,N_78,N_789);
or U3458 (N_3458,N_776,N_591);
nor U3459 (N_3459,N_365,N_607);
nand U3460 (N_3460,N_1691,N_1935);
and U3461 (N_3461,N_1403,N_2069);
nand U3462 (N_3462,N_2364,N_915);
and U3463 (N_3463,N_2280,N_805);
nor U3464 (N_3464,N_411,N_1333);
and U3465 (N_3465,N_2031,N_9);
and U3466 (N_3466,N_2003,N_1653);
nand U3467 (N_3467,N_2144,N_862);
nor U3468 (N_3468,N_2260,N_1342);
nor U3469 (N_3469,N_1445,N_1738);
and U3470 (N_3470,N_891,N_1286);
nor U3471 (N_3471,N_1360,N_910);
nor U3472 (N_3472,N_220,N_1614);
nor U3473 (N_3473,N_1618,N_239);
nor U3474 (N_3474,N_1376,N_1187);
nand U3475 (N_3475,N_1927,N_938);
or U3476 (N_3476,N_2088,N_403);
and U3477 (N_3477,N_1130,N_1240);
nor U3478 (N_3478,N_749,N_1587);
and U3479 (N_3479,N_179,N_352);
and U3480 (N_3480,N_1153,N_804);
and U3481 (N_3481,N_416,N_1018);
and U3482 (N_3482,N_519,N_71);
or U3483 (N_3483,N_2332,N_1991);
nand U3484 (N_3484,N_1058,N_98);
nand U3485 (N_3485,N_1117,N_989);
and U3486 (N_3486,N_480,N_1810);
and U3487 (N_3487,N_927,N_122);
or U3488 (N_3488,N_2232,N_92);
or U3489 (N_3489,N_1981,N_2464);
nand U3490 (N_3490,N_599,N_2090);
and U3491 (N_3491,N_558,N_1822);
nor U3492 (N_3492,N_860,N_447);
or U3493 (N_3493,N_2421,N_868);
and U3494 (N_3494,N_2101,N_1957);
or U3495 (N_3495,N_1679,N_1127);
or U3496 (N_3496,N_885,N_350);
nand U3497 (N_3497,N_887,N_2488);
nor U3498 (N_3498,N_677,N_757);
nand U3499 (N_3499,N_2432,N_1648);
nand U3500 (N_3500,N_777,N_450);
and U3501 (N_3501,N_453,N_1197);
and U3502 (N_3502,N_410,N_85);
nor U3503 (N_3503,N_954,N_2181);
or U3504 (N_3504,N_695,N_692);
or U3505 (N_3505,N_93,N_1782);
or U3506 (N_3506,N_114,N_2277);
nand U3507 (N_3507,N_884,N_1056);
nor U3508 (N_3508,N_1211,N_693);
and U3509 (N_3509,N_1381,N_266);
or U3510 (N_3510,N_185,N_676);
nor U3511 (N_3511,N_1987,N_634);
nand U3512 (N_3512,N_1354,N_256);
and U3513 (N_3513,N_1727,N_1178);
or U3514 (N_3514,N_1275,N_1601);
nor U3515 (N_3515,N_414,N_1481);
or U3516 (N_3516,N_167,N_1789);
and U3517 (N_3517,N_1106,N_1208);
or U3518 (N_3518,N_970,N_1382);
and U3519 (N_3519,N_1115,N_567);
and U3520 (N_3520,N_2447,N_993);
or U3521 (N_3521,N_2091,N_2481);
nand U3522 (N_3522,N_1244,N_337);
nand U3523 (N_3523,N_1002,N_1751);
or U3524 (N_3524,N_813,N_1562);
xor U3525 (N_3525,N_250,N_1685);
nand U3526 (N_3526,N_2295,N_2134);
or U3527 (N_3527,N_632,N_647);
nor U3528 (N_3528,N_609,N_1803);
nor U3529 (N_3529,N_212,N_468);
nand U3530 (N_3530,N_1778,N_1129);
or U3531 (N_3531,N_1923,N_697);
and U3532 (N_3532,N_1093,N_525);
nand U3533 (N_3533,N_1666,N_1910);
and U3534 (N_3534,N_285,N_1647);
nand U3535 (N_3535,N_1436,N_2135);
nand U3536 (N_3536,N_1716,N_1148);
and U3537 (N_3537,N_3,N_246);
and U3538 (N_3538,N_1270,N_1399);
xor U3539 (N_3539,N_120,N_1721);
or U3540 (N_3540,N_1963,N_974);
nor U3541 (N_3541,N_1911,N_203);
or U3542 (N_3542,N_617,N_99);
nand U3543 (N_3543,N_746,N_1261);
nor U3544 (N_3544,N_1644,N_354);
nor U3545 (N_3545,N_590,N_2266);
or U3546 (N_3546,N_783,N_15);
and U3547 (N_3547,N_2456,N_1356);
or U3548 (N_3548,N_216,N_243);
nand U3549 (N_3549,N_292,N_799);
and U3550 (N_3550,N_1253,N_1976);
nand U3551 (N_3551,N_2382,N_1134);
and U3552 (N_3552,N_2106,N_1435);
or U3553 (N_3553,N_1489,N_2220);
or U3554 (N_3554,N_1417,N_2262);
nor U3555 (N_3555,N_2065,N_1116);
and U3556 (N_3556,N_1791,N_2473);
nor U3557 (N_3557,N_1737,N_1037);
and U3558 (N_3558,N_139,N_1747);
nor U3559 (N_3559,N_2356,N_1284);
and U3560 (N_3560,N_82,N_494);
or U3561 (N_3561,N_548,N_1170);
and U3562 (N_3562,N_724,N_1154);
or U3563 (N_3563,N_2158,N_1800);
and U3564 (N_3564,N_133,N_1125);
and U3565 (N_3565,N_208,N_1527);
nor U3566 (N_3566,N_1752,N_189);
or U3567 (N_3567,N_1754,N_1519);
and U3568 (N_3568,N_1961,N_1163);
and U3569 (N_3569,N_2370,N_1028);
or U3570 (N_3570,N_1331,N_1538);
nand U3571 (N_3571,N_192,N_1714);
nand U3572 (N_3572,N_2209,N_27);
nor U3573 (N_3573,N_2238,N_1639);
nand U3574 (N_3574,N_1998,N_1352);
nor U3575 (N_3575,N_1242,N_1660);
nor U3576 (N_3576,N_1198,N_458);
and U3577 (N_3577,N_79,N_712);
nor U3578 (N_3578,N_2159,N_620);
or U3579 (N_3579,N_1173,N_2307);
xor U3580 (N_3580,N_2157,N_1646);
nor U3581 (N_3581,N_1582,N_1785);
nor U3582 (N_3582,N_1680,N_1216);
nor U3583 (N_3583,N_362,N_2258);
nand U3584 (N_3584,N_2193,N_2141);
nor U3585 (N_3585,N_1893,N_1368);
nand U3586 (N_3586,N_51,N_2255);
nor U3587 (N_3587,N_579,N_1359);
and U3588 (N_3588,N_1075,N_1348);
nand U3589 (N_3589,N_2431,N_1412);
nor U3590 (N_3590,N_1996,N_317);
or U3591 (N_3591,N_2278,N_72);
nor U3592 (N_3592,N_2052,N_2281);
or U3593 (N_3593,N_2429,N_467);
and U3594 (N_3594,N_1031,N_2476);
nor U3595 (N_3595,N_255,N_2073);
and U3596 (N_3596,N_2454,N_888);
nor U3597 (N_3597,N_895,N_1297);
nor U3598 (N_3598,N_2019,N_1830);
nor U3599 (N_3599,N_2287,N_1077);
nand U3600 (N_3600,N_2108,N_1105);
nor U3601 (N_3601,N_1518,N_265);
or U3602 (N_3602,N_1463,N_1281);
xor U3603 (N_3603,N_498,N_1213);
nor U3604 (N_3604,N_1853,N_113);
nor U3605 (N_3605,N_2081,N_14);
nor U3606 (N_3606,N_323,N_2415);
and U3607 (N_3607,N_1824,N_1924);
and U3608 (N_3608,N_457,N_834);
nand U3609 (N_3609,N_2053,N_234);
or U3610 (N_3610,N_2453,N_1842);
nand U3611 (N_3611,N_2326,N_736);
nor U3612 (N_3612,N_2066,N_2116);
or U3613 (N_3613,N_315,N_470);
or U3614 (N_3614,N_2221,N_1082);
and U3615 (N_3615,N_1616,N_2397);
nand U3616 (N_3616,N_848,N_2120);
or U3617 (N_3617,N_574,N_1901);
and U3618 (N_3618,N_158,N_1585);
nor U3619 (N_3619,N_1508,N_1053);
and U3620 (N_3620,N_890,N_1466);
and U3621 (N_3621,N_238,N_1032);
nor U3622 (N_3622,N_1355,N_1094);
and U3623 (N_3623,N_1502,N_21);
and U3624 (N_3624,N_913,N_227);
nor U3625 (N_3625,N_865,N_1833);
and U3626 (N_3626,N_235,N_1279);
nor U3627 (N_3627,N_125,N_1781);
and U3628 (N_3628,N_270,N_578);
nor U3629 (N_3629,N_764,N_442);
and U3630 (N_3630,N_1526,N_1442);
and U3631 (N_3631,N_1393,N_1875);
or U3632 (N_3632,N_645,N_928);
and U3633 (N_3633,N_18,N_555);
or U3634 (N_3634,N_1706,N_368);
nor U3635 (N_3635,N_705,N_844);
nand U3636 (N_3636,N_2274,N_1323);
nor U3637 (N_3637,N_672,N_1194);
and U3638 (N_3638,N_2161,N_2187);
or U3639 (N_3639,N_1605,N_2095);
nand U3640 (N_3640,N_1954,N_2206);
nand U3641 (N_3641,N_1695,N_594);
nand U3642 (N_3642,N_2349,N_1866);
nand U3643 (N_3643,N_1113,N_1722);
nand U3644 (N_3644,N_1378,N_2337);
or U3645 (N_3645,N_737,N_1574);
nand U3646 (N_3646,N_1898,N_960);
and U3647 (N_3647,N_109,N_221);
nand U3648 (N_3648,N_1864,N_580);
nor U3649 (N_3649,N_2062,N_2383);
and U3650 (N_3650,N_2207,N_1334);
or U3651 (N_3651,N_1262,N_2204);
and U3652 (N_3652,N_2350,N_1338);
or U3653 (N_3653,N_143,N_2305);
nand U3654 (N_3654,N_1128,N_1282);
or U3655 (N_3655,N_322,N_1726);
or U3656 (N_3656,N_1591,N_2042);
and U3657 (N_3657,N_190,N_1863);
or U3658 (N_3658,N_1631,N_908);
nor U3659 (N_3659,N_505,N_334);
nand U3660 (N_3660,N_1087,N_1946);
nand U3661 (N_3661,N_1054,N_1203);
nor U3662 (N_3662,N_698,N_522);
or U3663 (N_3663,N_1971,N_2321);
and U3664 (N_3664,N_1892,N_998);
or U3665 (N_3665,N_1503,N_2319);
or U3666 (N_3666,N_180,N_1022);
nor U3667 (N_3667,N_1958,N_184);
or U3668 (N_3668,N_1577,N_1405);
and U3669 (N_3669,N_1385,N_38);
nor U3670 (N_3670,N_427,N_1487);
nand U3671 (N_3671,N_1559,N_778);
and U3672 (N_3672,N_939,N_1684);
nor U3673 (N_3673,N_343,N_956);
nor U3674 (N_3674,N_1753,N_1857);
nor U3675 (N_3675,N_917,N_1986);
and U3676 (N_3676,N_446,N_581);
nor U3677 (N_3677,N_1305,N_1656);
and U3678 (N_3678,N_2012,N_2498);
nand U3679 (N_3679,N_1384,N_197);
nand U3680 (N_3680,N_874,N_259);
or U3681 (N_3681,N_916,N_1846);
or U3682 (N_3682,N_275,N_942);
or U3683 (N_3683,N_1494,N_2169);
nand U3684 (N_3684,N_1136,N_62);
or U3685 (N_3685,N_130,N_2075);
nor U3686 (N_3686,N_0,N_1228);
nor U3687 (N_3687,N_1029,N_2050);
and U3688 (N_3688,N_1226,N_386);
nor U3689 (N_3689,N_690,N_633);
nor U3690 (N_3690,N_1780,N_1964);
nand U3691 (N_3691,N_1272,N_957);
nand U3692 (N_3692,N_1545,N_400);
or U3693 (N_3693,N_743,N_552);
nand U3694 (N_3694,N_826,N_2496);
or U3695 (N_3695,N_823,N_1968);
or U3696 (N_3696,N_187,N_1770);
and U3697 (N_3697,N_1380,N_1443);
nand U3698 (N_3698,N_951,N_2233);
nor U3699 (N_3699,N_997,N_2044);
xnor U3700 (N_3700,N_2469,N_1409);
and U3701 (N_3701,N_2224,N_491);
or U3702 (N_3702,N_1854,N_1150);
nand U3703 (N_3703,N_850,N_280);
nor U3704 (N_3704,N_1912,N_1169);
or U3705 (N_3705,N_188,N_1877);
nand U3706 (N_3706,N_687,N_1482);
nor U3707 (N_3707,N_2006,N_815);
and U3708 (N_3708,N_547,N_2338);
nor U3709 (N_3709,N_2149,N_431);
and U3710 (N_3710,N_2430,N_1621);
and U3711 (N_3711,N_1659,N_514);
nand U3712 (N_3712,N_1829,N_1588);
or U3713 (N_3713,N_1951,N_516);
nand U3714 (N_3714,N_1146,N_1460);
nor U3715 (N_3715,N_2079,N_984);
nand U3716 (N_3716,N_544,N_2061);
or U3717 (N_3717,N_1217,N_1608);
nor U3718 (N_3718,N_1119,N_1086);
and U3719 (N_3719,N_2493,N_1345);
and U3720 (N_3720,N_28,N_1006);
or U3721 (N_3721,N_1469,N_1786);
and U3722 (N_3722,N_1458,N_49);
and U3723 (N_3723,N_886,N_2210);
and U3724 (N_3724,N_240,N_336);
nor U3725 (N_3725,N_1565,N_841);
nand U3726 (N_3726,N_1628,N_123);
and U3727 (N_3727,N_2375,N_1702);
and U3728 (N_3728,N_261,N_2360);
nor U3729 (N_3729,N_820,N_196);
nand U3730 (N_3730,N_1326,N_1597);
nand U3731 (N_3731,N_1307,N_254);
nor U3732 (N_3732,N_277,N_2318);
and U3733 (N_3733,N_821,N_2156);
nor U3734 (N_3734,N_800,N_308);
or U3735 (N_3735,N_1847,N_229);
nand U3736 (N_3736,N_1862,N_1192);
and U3737 (N_3737,N_2230,N_2435);
and U3738 (N_3738,N_1586,N_893);
or U3739 (N_3739,N_589,N_655);
nor U3740 (N_3740,N_600,N_335);
nand U3741 (N_3741,N_1584,N_2244);
nand U3742 (N_3742,N_772,N_1367);
and U3743 (N_3743,N_1554,N_433);
and U3744 (N_3744,N_1160,N_2123);
nand U3745 (N_3745,N_175,N_132);
or U3746 (N_3746,N_236,N_836);
nor U3747 (N_3747,N_791,N_531);
nand U3748 (N_3748,N_385,N_1513);
nand U3749 (N_3749,N_405,N_2138);
and U3750 (N_3750,N_2418,N_2307);
nor U3751 (N_3751,N_1559,N_1637);
nor U3752 (N_3752,N_569,N_207);
nand U3753 (N_3753,N_779,N_2277);
nor U3754 (N_3754,N_2046,N_1568);
or U3755 (N_3755,N_1927,N_708);
and U3756 (N_3756,N_1718,N_1297);
nand U3757 (N_3757,N_293,N_145);
nand U3758 (N_3758,N_1449,N_1557);
and U3759 (N_3759,N_1619,N_176);
nand U3760 (N_3760,N_175,N_1200);
nand U3761 (N_3761,N_851,N_897);
nand U3762 (N_3762,N_358,N_1281);
and U3763 (N_3763,N_2160,N_668);
nor U3764 (N_3764,N_378,N_1060);
and U3765 (N_3765,N_997,N_2392);
or U3766 (N_3766,N_2023,N_2155);
or U3767 (N_3767,N_618,N_1238);
and U3768 (N_3768,N_1502,N_661);
nor U3769 (N_3769,N_487,N_1062);
nor U3770 (N_3770,N_2433,N_1419);
nand U3771 (N_3771,N_1939,N_1932);
or U3772 (N_3772,N_1833,N_1297);
and U3773 (N_3773,N_382,N_940);
nor U3774 (N_3774,N_283,N_2363);
and U3775 (N_3775,N_21,N_580);
and U3776 (N_3776,N_2315,N_1497);
and U3777 (N_3777,N_1454,N_586);
and U3778 (N_3778,N_901,N_802);
or U3779 (N_3779,N_1138,N_1487);
nand U3780 (N_3780,N_1374,N_1674);
nor U3781 (N_3781,N_905,N_1155);
or U3782 (N_3782,N_1758,N_2208);
nor U3783 (N_3783,N_1730,N_852);
or U3784 (N_3784,N_130,N_426);
or U3785 (N_3785,N_1443,N_2382);
or U3786 (N_3786,N_1891,N_662);
nand U3787 (N_3787,N_1238,N_1940);
nand U3788 (N_3788,N_1056,N_260);
xnor U3789 (N_3789,N_2186,N_2220);
and U3790 (N_3790,N_2450,N_297);
nand U3791 (N_3791,N_680,N_1061);
nand U3792 (N_3792,N_1408,N_2492);
nand U3793 (N_3793,N_217,N_2130);
nor U3794 (N_3794,N_380,N_129);
nor U3795 (N_3795,N_656,N_1045);
nor U3796 (N_3796,N_1615,N_1094);
or U3797 (N_3797,N_1380,N_2398);
nor U3798 (N_3798,N_1421,N_1614);
or U3799 (N_3799,N_772,N_561);
nand U3800 (N_3800,N_1405,N_1478);
nor U3801 (N_3801,N_920,N_1415);
nor U3802 (N_3802,N_1607,N_229);
and U3803 (N_3803,N_2348,N_379);
or U3804 (N_3804,N_2280,N_1757);
nand U3805 (N_3805,N_924,N_1596);
and U3806 (N_3806,N_2441,N_579);
nand U3807 (N_3807,N_2476,N_1287);
nor U3808 (N_3808,N_398,N_1838);
nand U3809 (N_3809,N_1279,N_368);
nor U3810 (N_3810,N_1089,N_2369);
xor U3811 (N_3811,N_1313,N_348);
and U3812 (N_3812,N_550,N_9);
nor U3813 (N_3813,N_886,N_2451);
or U3814 (N_3814,N_2052,N_445);
or U3815 (N_3815,N_1766,N_56);
nand U3816 (N_3816,N_1910,N_553);
and U3817 (N_3817,N_300,N_516);
or U3818 (N_3818,N_391,N_1363);
nor U3819 (N_3819,N_2464,N_2079);
nand U3820 (N_3820,N_592,N_1938);
nor U3821 (N_3821,N_1298,N_1809);
nand U3822 (N_3822,N_1293,N_2215);
nor U3823 (N_3823,N_1791,N_1172);
and U3824 (N_3824,N_1616,N_229);
or U3825 (N_3825,N_2440,N_2053);
nand U3826 (N_3826,N_22,N_2305);
or U3827 (N_3827,N_1064,N_667);
nor U3828 (N_3828,N_1578,N_1774);
nor U3829 (N_3829,N_585,N_2113);
and U3830 (N_3830,N_458,N_1518);
nand U3831 (N_3831,N_493,N_697);
or U3832 (N_3832,N_2140,N_620);
nor U3833 (N_3833,N_1124,N_525);
and U3834 (N_3834,N_1666,N_1226);
and U3835 (N_3835,N_2415,N_92);
nor U3836 (N_3836,N_1500,N_1521);
nand U3837 (N_3837,N_2241,N_1810);
nor U3838 (N_3838,N_2329,N_2153);
nand U3839 (N_3839,N_621,N_734);
and U3840 (N_3840,N_951,N_1656);
and U3841 (N_3841,N_859,N_1188);
and U3842 (N_3842,N_2026,N_1467);
nand U3843 (N_3843,N_1173,N_764);
or U3844 (N_3844,N_1016,N_1235);
and U3845 (N_3845,N_1801,N_708);
nand U3846 (N_3846,N_1831,N_2105);
nor U3847 (N_3847,N_2433,N_566);
nand U3848 (N_3848,N_1318,N_1009);
nand U3849 (N_3849,N_1855,N_2345);
and U3850 (N_3850,N_169,N_1954);
xor U3851 (N_3851,N_36,N_754);
or U3852 (N_3852,N_2392,N_455);
nand U3853 (N_3853,N_2074,N_2220);
nand U3854 (N_3854,N_2040,N_1134);
or U3855 (N_3855,N_911,N_1601);
nor U3856 (N_3856,N_571,N_101);
and U3857 (N_3857,N_591,N_1906);
nand U3858 (N_3858,N_240,N_210);
and U3859 (N_3859,N_2070,N_1546);
nor U3860 (N_3860,N_1659,N_827);
nor U3861 (N_3861,N_1398,N_1438);
and U3862 (N_3862,N_93,N_509);
or U3863 (N_3863,N_2466,N_1946);
nor U3864 (N_3864,N_2330,N_2177);
nand U3865 (N_3865,N_1808,N_2015);
or U3866 (N_3866,N_92,N_1378);
and U3867 (N_3867,N_128,N_910);
nand U3868 (N_3868,N_1128,N_1433);
or U3869 (N_3869,N_266,N_683);
nor U3870 (N_3870,N_1083,N_721);
or U3871 (N_3871,N_800,N_581);
nor U3872 (N_3872,N_1488,N_1806);
or U3873 (N_3873,N_298,N_1155);
nand U3874 (N_3874,N_1316,N_556);
nor U3875 (N_3875,N_1443,N_635);
or U3876 (N_3876,N_277,N_1613);
nor U3877 (N_3877,N_2139,N_57);
and U3878 (N_3878,N_2267,N_1729);
and U3879 (N_3879,N_1788,N_1497);
or U3880 (N_3880,N_2032,N_231);
nand U3881 (N_3881,N_774,N_2097);
nor U3882 (N_3882,N_520,N_545);
nand U3883 (N_3883,N_1152,N_407);
nor U3884 (N_3884,N_2235,N_1138);
or U3885 (N_3885,N_2140,N_1009);
nor U3886 (N_3886,N_1186,N_1148);
nand U3887 (N_3887,N_1709,N_1003);
or U3888 (N_3888,N_2350,N_2377);
nand U3889 (N_3889,N_1833,N_2107);
nor U3890 (N_3890,N_1294,N_773);
and U3891 (N_3891,N_2363,N_329);
and U3892 (N_3892,N_1226,N_148);
nand U3893 (N_3893,N_353,N_2052);
or U3894 (N_3894,N_430,N_1139);
nor U3895 (N_3895,N_193,N_1539);
or U3896 (N_3896,N_1313,N_199);
or U3897 (N_3897,N_457,N_1022);
nand U3898 (N_3898,N_1733,N_2228);
nor U3899 (N_3899,N_1933,N_2249);
and U3900 (N_3900,N_1596,N_1149);
or U3901 (N_3901,N_832,N_1288);
and U3902 (N_3902,N_1994,N_928);
or U3903 (N_3903,N_1836,N_1678);
and U3904 (N_3904,N_1617,N_1220);
or U3905 (N_3905,N_1675,N_1568);
or U3906 (N_3906,N_582,N_430);
nor U3907 (N_3907,N_1440,N_845);
or U3908 (N_3908,N_1464,N_1941);
nand U3909 (N_3909,N_450,N_2312);
or U3910 (N_3910,N_663,N_170);
nand U3911 (N_3911,N_740,N_1962);
nand U3912 (N_3912,N_2363,N_1507);
xor U3913 (N_3913,N_2306,N_2475);
or U3914 (N_3914,N_1771,N_2164);
nor U3915 (N_3915,N_2292,N_1783);
nand U3916 (N_3916,N_998,N_2080);
nor U3917 (N_3917,N_50,N_855);
or U3918 (N_3918,N_1678,N_1112);
nand U3919 (N_3919,N_1212,N_689);
nor U3920 (N_3920,N_1228,N_1729);
or U3921 (N_3921,N_1883,N_93);
and U3922 (N_3922,N_454,N_1814);
and U3923 (N_3923,N_1610,N_62);
nand U3924 (N_3924,N_4,N_220);
and U3925 (N_3925,N_2114,N_962);
or U3926 (N_3926,N_2473,N_1549);
nand U3927 (N_3927,N_1638,N_1166);
xor U3928 (N_3928,N_0,N_1272);
nor U3929 (N_3929,N_1035,N_1252);
nand U3930 (N_3930,N_306,N_1367);
or U3931 (N_3931,N_715,N_2357);
and U3932 (N_3932,N_1676,N_2000);
and U3933 (N_3933,N_919,N_1774);
nor U3934 (N_3934,N_1029,N_2282);
nor U3935 (N_3935,N_381,N_1371);
nor U3936 (N_3936,N_203,N_254);
and U3937 (N_3937,N_1986,N_1656);
nor U3938 (N_3938,N_2439,N_1346);
xor U3939 (N_3939,N_899,N_901);
or U3940 (N_3940,N_471,N_1060);
or U3941 (N_3941,N_280,N_2402);
or U3942 (N_3942,N_614,N_2451);
nand U3943 (N_3943,N_128,N_958);
nand U3944 (N_3944,N_2310,N_91);
and U3945 (N_3945,N_1024,N_1119);
nor U3946 (N_3946,N_2423,N_904);
nand U3947 (N_3947,N_2294,N_1258);
nor U3948 (N_3948,N_1921,N_110);
and U3949 (N_3949,N_1068,N_283);
and U3950 (N_3950,N_77,N_1660);
nand U3951 (N_3951,N_2250,N_981);
or U3952 (N_3952,N_1605,N_1959);
and U3953 (N_3953,N_1513,N_2414);
nor U3954 (N_3954,N_521,N_2081);
nor U3955 (N_3955,N_1903,N_1837);
or U3956 (N_3956,N_297,N_1952);
nand U3957 (N_3957,N_336,N_124);
or U3958 (N_3958,N_1091,N_649);
and U3959 (N_3959,N_511,N_1808);
and U3960 (N_3960,N_277,N_610);
or U3961 (N_3961,N_2474,N_1494);
or U3962 (N_3962,N_1773,N_1921);
and U3963 (N_3963,N_1777,N_1127);
nand U3964 (N_3964,N_781,N_1567);
nor U3965 (N_3965,N_2384,N_2349);
nand U3966 (N_3966,N_2384,N_437);
nor U3967 (N_3967,N_2320,N_116);
and U3968 (N_3968,N_336,N_1381);
nor U3969 (N_3969,N_391,N_2253);
nand U3970 (N_3970,N_1411,N_797);
nand U3971 (N_3971,N_1467,N_651);
or U3972 (N_3972,N_930,N_1348);
nand U3973 (N_3973,N_601,N_1230);
nand U3974 (N_3974,N_620,N_1894);
and U3975 (N_3975,N_447,N_1155);
or U3976 (N_3976,N_180,N_22);
and U3977 (N_3977,N_191,N_402);
and U3978 (N_3978,N_2479,N_194);
and U3979 (N_3979,N_839,N_1875);
nand U3980 (N_3980,N_1284,N_1253);
and U3981 (N_3981,N_2102,N_2168);
and U3982 (N_3982,N_1580,N_1980);
nand U3983 (N_3983,N_548,N_495);
and U3984 (N_3984,N_2163,N_1222);
nor U3985 (N_3985,N_605,N_1000);
or U3986 (N_3986,N_1587,N_1801);
and U3987 (N_3987,N_60,N_1327);
nor U3988 (N_3988,N_1893,N_1332);
nand U3989 (N_3989,N_33,N_1752);
or U3990 (N_3990,N_1541,N_972);
nand U3991 (N_3991,N_104,N_2070);
nand U3992 (N_3992,N_984,N_1031);
xnor U3993 (N_3993,N_1216,N_132);
and U3994 (N_3994,N_171,N_1638);
or U3995 (N_3995,N_427,N_943);
nand U3996 (N_3996,N_1098,N_10);
or U3997 (N_3997,N_888,N_809);
or U3998 (N_3998,N_260,N_2338);
and U3999 (N_3999,N_1853,N_972);
nor U4000 (N_4000,N_526,N_1102);
and U4001 (N_4001,N_691,N_1524);
nand U4002 (N_4002,N_1627,N_1338);
or U4003 (N_4003,N_374,N_632);
and U4004 (N_4004,N_399,N_1337);
nor U4005 (N_4005,N_1332,N_1646);
or U4006 (N_4006,N_265,N_1628);
or U4007 (N_4007,N_344,N_340);
and U4008 (N_4008,N_323,N_1679);
or U4009 (N_4009,N_571,N_1141);
or U4010 (N_4010,N_1812,N_1838);
or U4011 (N_4011,N_1226,N_477);
nor U4012 (N_4012,N_1623,N_2387);
or U4013 (N_4013,N_1460,N_1262);
nor U4014 (N_4014,N_357,N_393);
nor U4015 (N_4015,N_946,N_704);
or U4016 (N_4016,N_790,N_408);
nor U4017 (N_4017,N_356,N_199);
nand U4018 (N_4018,N_219,N_842);
nor U4019 (N_4019,N_1279,N_2238);
nand U4020 (N_4020,N_161,N_2278);
and U4021 (N_4021,N_1232,N_247);
or U4022 (N_4022,N_1133,N_1642);
xnor U4023 (N_4023,N_300,N_2042);
or U4024 (N_4024,N_2263,N_786);
or U4025 (N_4025,N_147,N_319);
xnor U4026 (N_4026,N_818,N_203);
nand U4027 (N_4027,N_1553,N_899);
nand U4028 (N_4028,N_2273,N_2183);
and U4029 (N_4029,N_218,N_1184);
nor U4030 (N_4030,N_150,N_1430);
and U4031 (N_4031,N_660,N_301);
or U4032 (N_4032,N_620,N_1942);
or U4033 (N_4033,N_873,N_1139);
nand U4034 (N_4034,N_1669,N_825);
nand U4035 (N_4035,N_2100,N_2216);
or U4036 (N_4036,N_943,N_1285);
and U4037 (N_4037,N_1859,N_1707);
nand U4038 (N_4038,N_1094,N_2049);
nor U4039 (N_4039,N_1803,N_2335);
and U4040 (N_4040,N_1584,N_2400);
nand U4041 (N_4041,N_27,N_511);
nand U4042 (N_4042,N_712,N_706);
or U4043 (N_4043,N_33,N_1904);
or U4044 (N_4044,N_2184,N_1005);
nor U4045 (N_4045,N_535,N_296);
nor U4046 (N_4046,N_2423,N_1575);
or U4047 (N_4047,N_1643,N_1068);
and U4048 (N_4048,N_2470,N_1050);
nor U4049 (N_4049,N_1659,N_596);
nand U4050 (N_4050,N_1789,N_855);
nor U4051 (N_4051,N_2053,N_2100);
or U4052 (N_4052,N_1007,N_356);
nor U4053 (N_4053,N_672,N_161);
or U4054 (N_4054,N_814,N_853);
nand U4055 (N_4055,N_184,N_1744);
and U4056 (N_4056,N_2402,N_312);
nor U4057 (N_4057,N_218,N_2455);
and U4058 (N_4058,N_591,N_572);
nand U4059 (N_4059,N_2034,N_1961);
or U4060 (N_4060,N_977,N_1739);
and U4061 (N_4061,N_39,N_582);
nor U4062 (N_4062,N_2122,N_401);
or U4063 (N_4063,N_470,N_2087);
nor U4064 (N_4064,N_1903,N_1508);
or U4065 (N_4065,N_1191,N_1290);
and U4066 (N_4066,N_1857,N_1500);
and U4067 (N_4067,N_2331,N_2409);
nor U4068 (N_4068,N_249,N_1614);
and U4069 (N_4069,N_1713,N_1913);
nor U4070 (N_4070,N_1662,N_85);
and U4071 (N_4071,N_1733,N_453);
and U4072 (N_4072,N_1784,N_1611);
nand U4073 (N_4073,N_2186,N_2069);
nand U4074 (N_4074,N_2038,N_2102);
and U4075 (N_4075,N_1501,N_181);
nor U4076 (N_4076,N_817,N_1763);
or U4077 (N_4077,N_2413,N_965);
nor U4078 (N_4078,N_2292,N_26);
and U4079 (N_4079,N_1649,N_668);
and U4080 (N_4080,N_563,N_441);
and U4081 (N_4081,N_2137,N_2470);
and U4082 (N_4082,N_852,N_2145);
nand U4083 (N_4083,N_966,N_800);
or U4084 (N_4084,N_2440,N_2105);
nor U4085 (N_4085,N_1632,N_641);
nand U4086 (N_4086,N_2329,N_2003);
or U4087 (N_4087,N_2213,N_1782);
nor U4088 (N_4088,N_1852,N_1554);
or U4089 (N_4089,N_118,N_1370);
nand U4090 (N_4090,N_2199,N_1729);
or U4091 (N_4091,N_1189,N_705);
and U4092 (N_4092,N_2490,N_2039);
or U4093 (N_4093,N_250,N_885);
nor U4094 (N_4094,N_2464,N_756);
nand U4095 (N_4095,N_2284,N_134);
and U4096 (N_4096,N_1543,N_753);
and U4097 (N_4097,N_985,N_2405);
or U4098 (N_4098,N_1436,N_513);
nor U4099 (N_4099,N_2326,N_693);
nor U4100 (N_4100,N_2288,N_179);
nand U4101 (N_4101,N_2028,N_93);
or U4102 (N_4102,N_322,N_1817);
and U4103 (N_4103,N_743,N_618);
nor U4104 (N_4104,N_1447,N_367);
or U4105 (N_4105,N_238,N_2462);
nor U4106 (N_4106,N_267,N_673);
and U4107 (N_4107,N_1,N_1919);
nor U4108 (N_4108,N_1149,N_1032);
or U4109 (N_4109,N_521,N_44);
nor U4110 (N_4110,N_1834,N_1924);
or U4111 (N_4111,N_1754,N_2216);
or U4112 (N_4112,N_1382,N_528);
and U4113 (N_4113,N_1728,N_522);
nor U4114 (N_4114,N_136,N_1810);
and U4115 (N_4115,N_1157,N_1911);
xnor U4116 (N_4116,N_2198,N_1919);
or U4117 (N_4117,N_2044,N_2420);
or U4118 (N_4118,N_345,N_2086);
or U4119 (N_4119,N_250,N_2128);
nor U4120 (N_4120,N_73,N_1247);
and U4121 (N_4121,N_1084,N_445);
nand U4122 (N_4122,N_2403,N_2316);
nand U4123 (N_4123,N_24,N_327);
or U4124 (N_4124,N_641,N_1907);
and U4125 (N_4125,N_497,N_513);
nor U4126 (N_4126,N_2024,N_151);
or U4127 (N_4127,N_1404,N_912);
and U4128 (N_4128,N_1250,N_855);
nand U4129 (N_4129,N_95,N_27);
and U4130 (N_4130,N_2065,N_1798);
nand U4131 (N_4131,N_1119,N_818);
and U4132 (N_4132,N_454,N_1279);
or U4133 (N_4133,N_2486,N_582);
and U4134 (N_4134,N_2209,N_712);
and U4135 (N_4135,N_2067,N_1105);
and U4136 (N_4136,N_1651,N_1331);
nand U4137 (N_4137,N_1162,N_2279);
or U4138 (N_4138,N_2253,N_927);
nor U4139 (N_4139,N_1388,N_816);
nor U4140 (N_4140,N_553,N_2430);
and U4141 (N_4141,N_540,N_2292);
and U4142 (N_4142,N_1370,N_2398);
nand U4143 (N_4143,N_2332,N_1596);
or U4144 (N_4144,N_102,N_1395);
nor U4145 (N_4145,N_1024,N_410);
and U4146 (N_4146,N_1043,N_574);
and U4147 (N_4147,N_1069,N_1972);
nor U4148 (N_4148,N_2050,N_1459);
nor U4149 (N_4149,N_2478,N_973);
or U4150 (N_4150,N_762,N_507);
and U4151 (N_4151,N_1673,N_1144);
nor U4152 (N_4152,N_1738,N_219);
nor U4153 (N_4153,N_1276,N_500);
nor U4154 (N_4154,N_1318,N_2055);
nand U4155 (N_4155,N_1345,N_1488);
nor U4156 (N_4156,N_2152,N_492);
and U4157 (N_4157,N_1572,N_13);
nand U4158 (N_4158,N_1408,N_1519);
nor U4159 (N_4159,N_1812,N_2268);
nor U4160 (N_4160,N_894,N_2488);
and U4161 (N_4161,N_1663,N_260);
nor U4162 (N_4162,N_1413,N_1116);
nand U4163 (N_4163,N_1990,N_1374);
nor U4164 (N_4164,N_1903,N_1151);
nor U4165 (N_4165,N_597,N_1510);
nor U4166 (N_4166,N_777,N_1401);
nand U4167 (N_4167,N_518,N_812);
xor U4168 (N_4168,N_2211,N_2168);
and U4169 (N_4169,N_957,N_1792);
and U4170 (N_4170,N_1675,N_689);
nand U4171 (N_4171,N_1788,N_2164);
nor U4172 (N_4172,N_227,N_1291);
nor U4173 (N_4173,N_1004,N_933);
nand U4174 (N_4174,N_786,N_1808);
nor U4175 (N_4175,N_947,N_983);
and U4176 (N_4176,N_2017,N_1554);
nand U4177 (N_4177,N_1170,N_1148);
and U4178 (N_4178,N_936,N_2484);
nor U4179 (N_4179,N_874,N_191);
or U4180 (N_4180,N_1827,N_1388);
nor U4181 (N_4181,N_878,N_448);
and U4182 (N_4182,N_1997,N_1129);
and U4183 (N_4183,N_855,N_212);
and U4184 (N_4184,N_476,N_37);
and U4185 (N_4185,N_1408,N_1610);
or U4186 (N_4186,N_881,N_944);
and U4187 (N_4187,N_2115,N_155);
nand U4188 (N_4188,N_365,N_1999);
or U4189 (N_4189,N_2297,N_143);
and U4190 (N_4190,N_2493,N_625);
and U4191 (N_4191,N_2462,N_477);
nor U4192 (N_4192,N_2387,N_1241);
or U4193 (N_4193,N_1340,N_491);
or U4194 (N_4194,N_362,N_484);
or U4195 (N_4195,N_1242,N_2124);
nor U4196 (N_4196,N_1569,N_1373);
or U4197 (N_4197,N_904,N_1190);
nand U4198 (N_4198,N_370,N_1273);
nor U4199 (N_4199,N_887,N_1393);
nand U4200 (N_4200,N_451,N_1548);
and U4201 (N_4201,N_1492,N_2471);
or U4202 (N_4202,N_1506,N_2183);
and U4203 (N_4203,N_56,N_2142);
and U4204 (N_4204,N_770,N_1491);
nor U4205 (N_4205,N_609,N_526);
and U4206 (N_4206,N_1884,N_781);
or U4207 (N_4207,N_437,N_1115);
nand U4208 (N_4208,N_1659,N_1203);
nor U4209 (N_4209,N_1492,N_794);
nor U4210 (N_4210,N_1171,N_694);
nor U4211 (N_4211,N_291,N_259);
nand U4212 (N_4212,N_605,N_2459);
nand U4213 (N_4213,N_1132,N_2374);
nand U4214 (N_4214,N_856,N_1608);
or U4215 (N_4215,N_1350,N_843);
or U4216 (N_4216,N_1401,N_470);
or U4217 (N_4217,N_1451,N_2183);
or U4218 (N_4218,N_717,N_1467);
and U4219 (N_4219,N_1767,N_15);
nor U4220 (N_4220,N_873,N_416);
or U4221 (N_4221,N_1915,N_2311);
and U4222 (N_4222,N_540,N_184);
nor U4223 (N_4223,N_1508,N_1407);
xnor U4224 (N_4224,N_1947,N_587);
or U4225 (N_4225,N_1089,N_1321);
nor U4226 (N_4226,N_901,N_1117);
nor U4227 (N_4227,N_1932,N_162);
nor U4228 (N_4228,N_1506,N_149);
and U4229 (N_4229,N_311,N_1056);
or U4230 (N_4230,N_2395,N_2068);
nand U4231 (N_4231,N_276,N_1132);
and U4232 (N_4232,N_1332,N_350);
nand U4233 (N_4233,N_1440,N_457);
and U4234 (N_4234,N_73,N_949);
nor U4235 (N_4235,N_860,N_780);
nor U4236 (N_4236,N_34,N_1735);
xnor U4237 (N_4237,N_1878,N_1478);
and U4238 (N_4238,N_584,N_1884);
nand U4239 (N_4239,N_854,N_222);
nand U4240 (N_4240,N_561,N_1448);
and U4241 (N_4241,N_510,N_1346);
nor U4242 (N_4242,N_1686,N_1517);
and U4243 (N_4243,N_566,N_1208);
nor U4244 (N_4244,N_1367,N_777);
nor U4245 (N_4245,N_32,N_698);
nor U4246 (N_4246,N_2281,N_573);
nand U4247 (N_4247,N_54,N_250);
nor U4248 (N_4248,N_1848,N_924);
and U4249 (N_4249,N_1258,N_1869);
nor U4250 (N_4250,N_1397,N_296);
and U4251 (N_4251,N_1321,N_1343);
and U4252 (N_4252,N_637,N_1783);
and U4253 (N_4253,N_319,N_1284);
nor U4254 (N_4254,N_835,N_141);
nor U4255 (N_4255,N_313,N_1126);
or U4256 (N_4256,N_2391,N_1190);
nor U4257 (N_4257,N_2320,N_55);
and U4258 (N_4258,N_184,N_2209);
nor U4259 (N_4259,N_1917,N_819);
nand U4260 (N_4260,N_583,N_2415);
nor U4261 (N_4261,N_2344,N_1675);
nand U4262 (N_4262,N_2363,N_694);
and U4263 (N_4263,N_816,N_1765);
and U4264 (N_4264,N_1484,N_865);
xnor U4265 (N_4265,N_452,N_1137);
and U4266 (N_4266,N_835,N_1784);
and U4267 (N_4267,N_1755,N_1433);
or U4268 (N_4268,N_19,N_2007);
xor U4269 (N_4269,N_2448,N_1799);
nand U4270 (N_4270,N_226,N_367);
nand U4271 (N_4271,N_152,N_2416);
nand U4272 (N_4272,N_2486,N_559);
or U4273 (N_4273,N_1837,N_97);
nand U4274 (N_4274,N_2080,N_2442);
or U4275 (N_4275,N_319,N_2100);
or U4276 (N_4276,N_1705,N_145);
and U4277 (N_4277,N_1577,N_160);
nor U4278 (N_4278,N_164,N_1043);
or U4279 (N_4279,N_2035,N_100);
nor U4280 (N_4280,N_2481,N_2369);
or U4281 (N_4281,N_1277,N_745);
nor U4282 (N_4282,N_362,N_80);
and U4283 (N_4283,N_2185,N_779);
and U4284 (N_4284,N_1059,N_2496);
nor U4285 (N_4285,N_1008,N_2275);
nor U4286 (N_4286,N_1775,N_102);
nand U4287 (N_4287,N_2393,N_445);
nor U4288 (N_4288,N_1260,N_1521);
nor U4289 (N_4289,N_2228,N_2031);
or U4290 (N_4290,N_2497,N_1110);
and U4291 (N_4291,N_1879,N_136);
or U4292 (N_4292,N_1161,N_1136);
nor U4293 (N_4293,N_2287,N_169);
nor U4294 (N_4294,N_204,N_1364);
or U4295 (N_4295,N_1197,N_1305);
nor U4296 (N_4296,N_412,N_1908);
and U4297 (N_4297,N_2437,N_1723);
or U4298 (N_4298,N_1077,N_2042);
or U4299 (N_4299,N_2119,N_1201);
nor U4300 (N_4300,N_1502,N_483);
and U4301 (N_4301,N_1001,N_201);
and U4302 (N_4302,N_681,N_1917);
or U4303 (N_4303,N_1818,N_1066);
nand U4304 (N_4304,N_1677,N_826);
or U4305 (N_4305,N_1214,N_2251);
nand U4306 (N_4306,N_1321,N_1965);
nand U4307 (N_4307,N_63,N_121);
and U4308 (N_4308,N_1742,N_410);
nand U4309 (N_4309,N_677,N_472);
or U4310 (N_4310,N_40,N_2248);
and U4311 (N_4311,N_1334,N_1961);
or U4312 (N_4312,N_2110,N_744);
nand U4313 (N_4313,N_1314,N_2263);
or U4314 (N_4314,N_1921,N_1437);
or U4315 (N_4315,N_2374,N_2041);
and U4316 (N_4316,N_1066,N_1876);
and U4317 (N_4317,N_1921,N_403);
or U4318 (N_4318,N_248,N_2326);
nor U4319 (N_4319,N_1518,N_2226);
nand U4320 (N_4320,N_267,N_2055);
or U4321 (N_4321,N_2202,N_1404);
or U4322 (N_4322,N_2409,N_2255);
nand U4323 (N_4323,N_2160,N_1640);
and U4324 (N_4324,N_2300,N_316);
nor U4325 (N_4325,N_848,N_1258);
nor U4326 (N_4326,N_999,N_1588);
xnor U4327 (N_4327,N_1537,N_1377);
or U4328 (N_4328,N_1570,N_1027);
nor U4329 (N_4329,N_1407,N_1959);
and U4330 (N_4330,N_763,N_1931);
or U4331 (N_4331,N_2022,N_1926);
nand U4332 (N_4332,N_1789,N_1587);
or U4333 (N_4333,N_1208,N_1216);
or U4334 (N_4334,N_1069,N_2449);
and U4335 (N_4335,N_1797,N_88);
or U4336 (N_4336,N_238,N_988);
nor U4337 (N_4337,N_2436,N_905);
nor U4338 (N_4338,N_1321,N_512);
and U4339 (N_4339,N_1786,N_2240);
nor U4340 (N_4340,N_890,N_958);
and U4341 (N_4341,N_332,N_1560);
nor U4342 (N_4342,N_1147,N_1406);
nor U4343 (N_4343,N_2100,N_1022);
nor U4344 (N_4344,N_2333,N_453);
and U4345 (N_4345,N_1811,N_1311);
nor U4346 (N_4346,N_2194,N_728);
or U4347 (N_4347,N_1232,N_2170);
nor U4348 (N_4348,N_962,N_1769);
and U4349 (N_4349,N_2123,N_2290);
and U4350 (N_4350,N_1903,N_886);
and U4351 (N_4351,N_1265,N_98);
and U4352 (N_4352,N_629,N_1449);
and U4353 (N_4353,N_1231,N_2376);
and U4354 (N_4354,N_1135,N_397);
and U4355 (N_4355,N_1855,N_1221);
nor U4356 (N_4356,N_2450,N_1248);
and U4357 (N_4357,N_1946,N_798);
or U4358 (N_4358,N_2161,N_1426);
nand U4359 (N_4359,N_1906,N_383);
and U4360 (N_4360,N_1282,N_2204);
and U4361 (N_4361,N_1027,N_1290);
and U4362 (N_4362,N_496,N_1401);
or U4363 (N_4363,N_2265,N_2469);
nand U4364 (N_4364,N_838,N_2308);
nand U4365 (N_4365,N_1937,N_735);
and U4366 (N_4366,N_2009,N_1918);
and U4367 (N_4367,N_227,N_963);
and U4368 (N_4368,N_1697,N_1268);
nor U4369 (N_4369,N_1945,N_1546);
nor U4370 (N_4370,N_1526,N_1114);
nor U4371 (N_4371,N_850,N_910);
nor U4372 (N_4372,N_925,N_1953);
or U4373 (N_4373,N_2493,N_475);
or U4374 (N_4374,N_1413,N_2303);
nor U4375 (N_4375,N_1989,N_440);
nand U4376 (N_4376,N_1423,N_2202);
or U4377 (N_4377,N_2044,N_156);
or U4378 (N_4378,N_1899,N_1444);
nor U4379 (N_4379,N_2310,N_1227);
nand U4380 (N_4380,N_1795,N_1239);
and U4381 (N_4381,N_445,N_1935);
nand U4382 (N_4382,N_1505,N_2149);
nand U4383 (N_4383,N_1097,N_1131);
nand U4384 (N_4384,N_1161,N_1029);
nor U4385 (N_4385,N_1266,N_992);
or U4386 (N_4386,N_1441,N_1148);
nor U4387 (N_4387,N_2309,N_875);
nor U4388 (N_4388,N_1730,N_2250);
nand U4389 (N_4389,N_1897,N_175);
or U4390 (N_4390,N_1208,N_2054);
and U4391 (N_4391,N_2411,N_1407);
and U4392 (N_4392,N_975,N_2332);
nor U4393 (N_4393,N_1701,N_1531);
and U4394 (N_4394,N_575,N_2132);
and U4395 (N_4395,N_2381,N_2439);
nand U4396 (N_4396,N_1409,N_1844);
and U4397 (N_4397,N_1971,N_2014);
and U4398 (N_4398,N_549,N_1557);
and U4399 (N_4399,N_486,N_2152);
nor U4400 (N_4400,N_56,N_664);
or U4401 (N_4401,N_1376,N_1535);
or U4402 (N_4402,N_183,N_84);
nand U4403 (N_4403,N_1545,N_2310);
nand U4404 (N_4404,N_248,N_2150);
nor U4405 (N_4405,N_1871,N_2329);
or U4406 (N_4406,N_1686,N_983);
nand U4407 (N_4407,N_678,N_764);
or U4408 (N_4408,N_2005,N_2232);
xor U4409 (N_4409,N_1743,N_2030);
nor U4410 (N_4410,N_2089,N_1622);
or U4411 (N_4411,N_898,N_814);
or U4412 (N_4412,N_2439,N_1405);
nor U4413 (N_4413,N_3,N_2081);
nor U4414 (N_4414,N_920,N_1009);
nor U4415 (N_4415,N_1294,N_194);
nand U4416 (N_4416,N_1895,N_2333);
nand U4417 (N_4417,N_2351,N_1686);
nor U4418 (N_4418,N_2034,N_2157);
nor U4419 (N_4419,N_421,N_389);
nand U4420 (N_4420,N_934,N_1044);
or U4421 (N_4421,N_558,N_411);
nand U4422 (N_4422,N_2284,N_960);
nand U4423 (N_4423,N_2102,N_177);
or U4424 (N_4424,N_1220,N_1866);
nor U4425 (N_4425,N_1929,N_521);
and U4426 (N_4426,N_1088,N_39);
nor U4427 (N_4427,N_1894,N_1317);
nor U4428 (N_4428,N_1723,N_787);
nor U4429 (N_4429,N_1364,N_2075);
nand U4430 (N_4430,N_1127,N_2385);
or U4431 (N_4431,N_1834,N_490);
and U4432 (N_4432,N_232,N_1595);
xor U4433 (N_4433,N_2247,N_583);
and U4434 (N_4434,N_1224,N_1352);
and U4435 (N_4435,N_536,N_484);
and U4436 (N_4436,N_478,N_1363);
nor U4437 (N_4437,N_959,N_1567);
nand U4438 (N_4438,N_2388,N_422);
nand U4439 (N_4439,N_1752,N_2197);
nor U4440 (N_4440,N_562,N_641);
nand U4441 (N_4441,N_819,N_2056);
or U4442 (N_4442,N_1147,N_515);
nand U4443 (N_4443,N_455,N_199);
or U4444 (N_4444,N_708,N_2038);
and U4445 (N_4445,N_451,N_999);
nor U4446 (N_4446,N_1493,N_1128);
nand U4447 (N_4447,N_1596,N_151);
and U4448 (N_4448,N_576,N_128);
or U4449 (N_4449,N_1746,N_2285);
and U4450 (N_4450,N_873,N_1418);
nand U4451 (N_4451,N_125,N_1096);
nor U4452 (N_4452,N_1761,N_187);
nor U4453 (N_4453,N_2333,N_2278);
or U4454 (N_4454,N_529,N_1034);
or U4455 (N_4455,N_1525,N_2417);
xnor U4456 (N_4456,N_2156,N_1706);
or U4457 (N_4457,N_1526,N_509);
xor U4458 (N_4458,N_197,N_1210);
nor U4459 (N_4459,N_36,N_784);
nand U4460 (N_4460,N_2360,N_318);
nand U4461 (N_4461,N_2304,N_473);
nor U4462 (N_4462,N_994,N_1585);
nand U4463 (N_4463,N_2429,N_1236);
nor U4464 (N_4464,N_1222,N_1440);
nand U4465 (N_4465,N_1129,N_1489);
and U4466 (N_4466,N_2031,N_1064);
nor U4467 (N_4467,N_2491,N_461);
or U4468 (N_4468,N_443,N_1114);
nand U4469 (N_4469,N_195,N_2224);
nand U4470 (N_4470,N_102,N_1002);
or U4471 (N_4471,N_1940,N_1868);
and U4472 (N_4472,N_82,N_1930);
nand U4473 (N_4473,N_2098,N_2430);
and U4474 (N_4474,N_1908,N_296);
nand U4475 (N_4475,N_1787,N_390);
and U4476 (N_4476,N_569,N_2487);
and U4477 (N_4477,N_1480,N_1409);
and U4478 (N_4478,N_2112,N_1682);
nor U4479 (N_4479,N_192,N_1907);
nor U4480 (N_4480,N_2312,N_1041);
or U4481 (N_4481,N_1675,N_723);
nor U4482 (N_4482,N_1793,N_1680);
nor U4483 (N_4483,N_2406,N_1511);
or U4484 (N_4484,N_662,N_468);
nand U4485 (N_4485,N_1380,N_31);
and U4486 (N_4486,N_694,N_1131);
nand U4487 (N_4487,N_799,N_502);
nand U4488 (N_4488,N_2450,N_1262);
nand U4489 (N_4489,N_1940,N_1876);
or U4490 (N_4490,N_102,N_2310);
or U4491 (N_4491,N_2179,N_621);
nor U4492 (N_4492,N_1528,N_2455);
and U4493 (N_4493,N_182,N_961);
nor U4494 (N_4494,N_1561,N_1889);
or U4495 (N_4495,N_2367,N_1883);
nand U4496 (N_4496,N_754,N_234);
or U4497 (N_4497,N_325,N_2084);
nor U4498 (N_4498,N_364,N_760);
nor U4499 (N_4499,N_764,N_2167);
nor U4500 (N_4500,N_2495,N_843);
nand U4501 (N_4501,N_2207,N_975);
or U4502 (N_4502,N_179,N_374);
and U4503 (N_4503,N_892,N_1342);
nand U4504 (N_4504,N_735,N_2383);
or U4505 (N_4505,N_2310,N_1712);
or U4506 (N_4506,N_634,N_456);
nor U4507 (N_4507,N_1560,N_2132);
nand U4508 (N_4508,N_535,N_307);
nand U4509 (N_4509,N_2290,N_2440);
nor U4510 (N_4510,N_1766,N_1007);
or U4511 (N_4511,N_66,N_502);
and U4512 (N_4512,N_90,N_864);
or U4513 (N_4513,N_967,N_78);
nor U4514 (N_4514,N_1795,N_1153);
or U4515 (N_4515,N_1811,N_156);
nor U4516 (N_4516,N_2194,N_1308);
nor U4517 (N_4517,N_1363,N_1368);
nor U4518 (N_4518,N_684,N_1135);
and U4519 (N_4519,N_1958,N_411);
or U4520 (N_4520,N_1446,N_347);
nand U4521 (N_4521,N_1143,N_1544);
or U4522 (N_4522,N_1105,N_1828);
or U4523 (N_4523,N_731,N_2462);
nor U4524 (N_4524,N_1955,N_2216);
nand U4525 (N_4525,N_1112,N_1896);
nand U4526 (N_4526,N_850,N_721);
nor U4527 (N_4527,N_282,N_896);
nand U4528 (N_4528,N_2045,N_1143);
nor U4529 (N_4529,N_471,N_599);
nand U4530 (N_4530,N_1328,N_1141);
nand U4531 (N_4531,N_654,N_572);
nor U4532 (N_4532,N_655,N_2243);
and U4533 (N_4533,N_1306,N_1145);
and U4534 (N_4534,N_1634,N_2256);
and U4535 (N_4535,N_985,N_1791);
or U4536 (N_4536,N_968,N_495);
or U4537 (N_4537,N_524,N_670);
and U4538 (N_4538,N_2463,N_630);
nor U4539 (N_4539,N_1003,N_2182);
and U4540 (N_4540,N_1504,N_1267);
or U4541 (N_4541,N_1777,N_1327);
nor U4542 (N_4542,N_1071,N_1056);
and U4543 (N_4543,N_2033,N_18);
nand U4544 (N_4544,N_1128,N_1155);
and U4545 (N_4545,N_643,N_1110);
or U4546 (N_4546,N_506,N_27);
or U4547 (N_4547,N_1875,N_802);
nand U4548 (N_4548,N_476,N_973);
and U4549 (N_4549,N_829,N_2027);
xor U4550 (N_4550,N_1923,N_1099);
and U4551 (N_4551,N_179,N_2397);
nor U4552 (N_4552,N_1179,N_1229);
nor U4553 (N_4553,N_1154,N_1773);
or U4554 (N_4554,N_1301,N_299);
or U4555 (N_4555,N_134,N_2390);
and U4556 (N_4556,N_853,N_1593);
and U4557 (N_4557,N_992,N_2317);
and U4558 (N_4558,N_2243,N_1500);
nand U4559 (N_4559,N_74,N_2424);
nand U4560 (N_4560,N_2481,N_1918);
nor U4561 (N_4561,N_790,N_2330);
and U4562 (N_4562,N_2408,N_661);
nor U4563 (N_4563,N_1498,N_1134);
nor U4564 (N_4564,N_2450,N_233);
nor U4565 (N_4565,N_42,N_2023);
or U4566 (N_4566,N_546,N_1168);
nor U4567 (N_4567,N_2437,N_1838);
nor U4568 (N_4568,N_1749,N_141);
nand U4569 (N_4569,N_142,N_38);
or U4570 (N_4570,N_2191,N_1086);
and U4571 (N_4571,N_499,N_182);
nor U4572 (N_4572,N_1619,N_186);
nand U4573 (N_4573,N_56,N_1904);
or U4574 (N_4574,N_2110,N_712);
or U4575 (N_4575,N_1809,N_2116);
and U4576 (N_4576,N_2368,N_1432);
or U4577 (N_4577,N_871,N_180);
nor U4578 (N_4578,N_1447,N_175);
nand U4579 (N_4579,N_394,N_939);
and U4580 (N_4580,N_1106,N_1065);
or U4581 (N_4581,N_1617,N_1661);
nor U4582 (N_4582,N_401,N_51);
and U4583 (N_4583,N_330,N_2241);
and U4584 (N_4584,N_378,N_1746);
and U4585 (N_4585,N_1447,N_1086);
nand U4586 (N_4586,N_1631,N_2455);
and U4587 (N_4587,N_1627,N_626);
nor U4588 (N_4588,N_931,N_1749);
or U4589 (N_4589,N_912,N_1595);
nor U4590 (N_4590,N_2131,N_1551);
nor U4591 (N_4591,N_2209,N_110);
xor U4592 (N_4592,N_1535,N_1894);
or U4593 (N_4593,N_2178,N_2208);
nand U4594 (N_4594,N_2366,N_737);
or U4595 (N_4595,N_521,N_1724);
nor U4596 (N_4596,N_1300,N_138);
and U4597 (N_4597,N_1350,N_913);
or U4598 (N_4598,N_1751,N_1204);
or U4599 (N_4599,N_1871,N_1111);
or U4600 (N_4600,N_1547,N_2405);
nor U4601 (N_4601,N_2154,N_700);
nand U4602 (N_4602,N_2017,N_826);
nand U4603 (N_4603,N_317,N_464);
and U4604 (N_4604,N_739,N_993);
nand U4605 (N_4605,N_1779,N_379);
and U4606 (N_4606,N_1405,N_2372);
nor U4607 (N_4607,N_1139,N_189);
nor U4608 (N_4608,N_879,N_2173);
or U4609 (N_4609,N_857,N_554);
and U4610 (N_4610,N_2224,N_564);
nand U4611 (N_4611,N_2418,N_2155);
nor U4612 (N_4612,N_2106,N_400);
or U4613 (N_4613,N_1295,N_586);
nor U4614 (N_4614,N_1058,N_424);
and U4615 (N_4615,N_25,N_2284);
or U4616 (N_4616,N_2002,N_1779);
nand U4617 (N_4617,N_1330,N_1823);
nand U4618 (N_4618,N_495,N_2360);
nor U4619 (N_4619,N_540,N_718);
or U4620 (N_4620,N_2201,N_2427);
or U4621 (N_4621,N_857,N_1831);
nor U4622 (N_4622,N_2446,N_1064);
and U4623 (N_4623,N_1581,N_1584);
nand U4624 (N_4624,N_2320,N_1737);
and U4625 (N_4625,N_1033,N_1672);
or U4626 (N_4626,N_1927,N_2189);
or U4627 (N_4627,N_2431,N_1921);
nand U4628 (N_4628,N_2447,N_2084);
or U4629 (N_4629,N_670,N_335);
nor U4630 (N_4630,N_1263,N_1480);
nor U4631 (N_4631,N_1247,N_211);
and U4632 (N_4632,N_1970,N_1639);
and U4633 (N_4633,N_2364,N_1960);
nor U4634 (N_4634,N_1461,N_2159);
nor U4635 (N_4635,N_1726,N_1806);
nand U4636 (N_4636,N_654,N_679);
nand U4637 (N_4637,N_1928,N_2115);
and U4638 (N_4638,N_2196,N_2138);
and U4639 (N_4639,N_1817,N_153);
or U4640 (N_4640,N_1886,N_507);
and U4641 (N_4641,N_483,N_1878);
and U4642 (N_4642,N_408,N_909);
nand U4643 (N_4643,N_1156,N_2359);
nor U4644 (N_4644,N_1361,N_1281);
or U4645 (N_4645,N_49,N_1906);
nand U4646 (N_4646,N_858,N_1664);
or U4647 (N_4647,N_277,N_2205);
nand U4648 (N_4648,N_1570,N_1643);
xnor U4649 (N_4649,N_589,N_217);
nor U4650 (N_4650,N_1517,N_485);
nor U4651 (N_4651,N_1139,N_2461);
nor U4652 (N_4652,N_468,N_295);
and U4653 (N_4653,N_29,N_2314);
nand U4654 (N_4654,N_165,N_630);
or U4655 (N_4655,N_17,N_2039);
nor U4656 (N_4656,N_2284,N_454);
nor U4657 (N_4657,N_1235,N_1317);
nor U4658 (N_4658,N_2053,N_1195);
or U4659 (N_4659,N_526,N_1880);
nand U4660 (N_4660,N_730,N_1186);
xnor U4661 (N_4661,N_1650,N_364);
or U4662 (N_4662,N_1494,N_1090);
or U4663 (N_4663,N_389,N_2107);
nor U4664 (N_4664,N_1087,N_1361);
and U4665 (N_4665,N_1250,N_2314);
nand U4666 (N_4666,N_79,N_1244);
and U4667 (N_4667,N_694,N_1501);
nand U4668 (N_4668,N_1900,N_885);
nor U4669 (N_4669,N_1883,N_2059);
and U4670 (N_4670,N_265,N_438);
nor U4671 (N_4671,N_2034,N_1591);
or U4672 (N_4672,N_1489,N_1340);
nor U4673 (N_4673,N_686,N_1551);
or U4674 (N_4674,N_474,N_226);
and U4675 (N_4675,N_1262,N_910);
nand U4676 (N_4676,N_432,N_1376);
nand U4677 (N_4677,N_1904,N_437);
nor U4678 (N_4678,N_1382,N_2121);
nand U4679 (N_4679,N_1408,N_542);
nand U4680 (N_4680,N_1055,N_1483);
and U4681 (N_4681,N_741,N_2064);
nor U4682 (N_4682,N_2108,N_998);
nand U4683 (N_4683,N_2089,N_2407);
or U4684 (N_4684,N_672,N_245);
nor U4685 (N_4685,N_238,N_1486);
and U4686 (N_4686,N_2111,N_416);
or U4687 (N_4687,N_75,N_1038);
nand U4688 (N_4688,N_952,N_1639);
xor U4689 (N_4689,N_1713,N_232);
and U4690 (N_4690,N_761,N_1194);
and U4691 (N_4691,N_316,N_1976);
and U4692 (N_4692,N_1294,N_132);
and U4693 (N_4693,N_2167,N_1893);
nand U4694 (N_4694,N_868,N_464);
or U4695 (N_4695,N_2346,N_1426);
and U4696 (N_4696,N_2126,N_2002);
nor U4697 (N_4697,N_2348,N_113);
and U4698 (N_4698,N_2402,N_2049);
or U4699 (N_4699,N_1835,N_2170);
nor U4700 (N_4700,N_183,N_621);
or U4701 (N_4701,N_1654,N_141);
nand U4702 (N_4702,N_1406,N_1719);
or U4703 (N_4703,N_1779,N_1984);
or U4704 (N_4704,N_1273,N_357);
or U4705 (N_4705,N_1898,N_109);
and U4706 (N_4706,N_503,N_122);
and U4707 (N_4707,N_87,N_1179);
or U4708 (N_4708,N_2070,N_1272);
nand U4709 (N_4709,N_1529,N_888);
and U4710 (N_4710,N_2325,N_1478);
and U4711 (N_4711,N_1564,N_545);
nor U4712 (N_4712,N_2163,N_283);
and U4713 (N_4713,N_1140,N_1772);
nor U4714 (N_4714,N_380,N_2184);
and U4715 (N_4715,N_592,N_1756);
and U4716 (N_4716,N_977,N_773);
nand U4717 (N_4717,N_573,N_2420);
or U4718 (N_4718,N_1851,N_639);
or U4719 (N_4719,N_306,N_1223);
nor U4720 (N_4720,N_2024,N_683);
or U4721 (N_4721,N_591,N_1455);
and U4722 (N_4722,N_89,N_2009);
and U4723 (N_4723,N_1219,N_907);
or U4724 (N_4724,N_65,N_1922);
or U4725 (N_4725,N_1696,N_26);
or U4726 (N_4726,N_720,N_734);
and U4727 (N_4727,N_396,N_1173);
nand U4728 (N_4728,N_2288,N_1001);
or U4729 (N_4729,N_2408,N_183);
nand U4730 (N_4730,N_1702,N_1989);
or U4731 (N_4731,N_2032,N_1352);
nand U4732 (N_4732,N_1704,N_312);
or U4733 (N_4733,N_109,N_1500);
or U4734 (N_4734,N_1158,N_227);
nand U4735 (N_4735,N_1111,N_964);
nor U4736 (N_4736,N_459,N_1324);
or U4737 (N_4737,N_241,N_1796);
nand U4738 (N_4738,N_2218,N_581);
nor U4739 (N_4739,N_802,N_957);
and U4740 (N_4740,N_2073,N_1669);
nand U4741 (N_4741,N_1593,N_237);
or U4742 (N_4742,N_1775,N_2433);
nand U4743 (N_4743,N_855,N_1159);
and U4744 (N_4744,N_200,N_2314);
or U4745 (N_4745,N_2337,N_2181);
or U4746 (N_4746,N_1384,N_692);
or U4747 (N_4747,N_1548,N_1134);
and U4748 (N_4748,N_1671,N_1594);
or U4749 (N_4749,N_2301,N_1331);
or U4750 (N_4750,N_1978,N_2485);
or U4751 (N_4751,N_2280,N_2322);
nor U4752 (N_4752,N_1823,N_2284);
or U4753 (N_4753,N_2364,N_2330);
or U4754 (N_4754,N_1551,N_1692);
and U4755 (N_4755,N_2051,N_782);
nand U4756 (N_4756,N_502,N_2380);
nand U4757 (N_4757,N_888,N_2407);
nor U4758 (N_4758,N_2179,N_2176);
nand U4759 (N_4759,N_381,N_1256);
nand U4760 (N_4760,N_947,N_407);
nand U4761 (N_4761,N_1279,N_952);
and U4762 (N_4762,N_1852,N_1343);
nand U4763 (N_4763,N_1617,N_1161);
or U4764 (N_4764,N_570,N_1528);
nand U4765 (N_4765,N_237,N_2274);
or U4766 (N_4766,N_2055,N_544);
nand U4767 (N_4767,N_1353,N_296);
nand U4768 (N_4768,N_2014,N_872);
and U4769 (N_4769,N_1806,N_679);
nand U4770 (N_4770,N_540,N_1302);
and U4771 (N_4771,N_287,N_1179);
and U4772 (N_4772,N_1008,N_7);
nor U4773 (N_4773,N_980,N_1213);
nand U4774 (N_4774,N_383,N_1819);
nor U4775 (N_4775,N_58,N_1274);
and U4776 (N_4776,N_250,N_1457);
nor U4777 (N_4777,N_810,N_202);
or U4778 (N_4778,N_199,N_1343);
and U4779 (N_4779,N_927,N_1736);
and U4780 (N_4780,N_505,N_2);
nand U4781 (N_4781,N_784,N_1271);
xor U4782 (N_4782,N_103,N_718);
nor U4783 (N_4783,N_1859,N_1063);
and U4784 (N_4784,N_1260,N_1224);
and U4785 (N_4785,N_1486,N_934);
nor U4786 (N_4786,N_2490,N_1041);
and U4787 (N_4787,N_642,N_1915);
nand U4788 (N_4788,N_208,N_1347);
nor U4789 (N_4789,N_2079,N_1011);
nand U4790 (N_4790,N_736,N_1189);
or U4791 (N_4791,N_1887,N_762);
nand U4792 (N_4792,N_1759,N_64);
or U4793 (N_4793,N_1001,N_139);
or U4794 (N_4794,N_924,N_617);
or U4795 (N_4795,N_2009,N_1305);
nor U4796 (N_4796,N_958,N_1280);
and U4797 (N_4797,N_1993,N_2181);
or U4798 (N_4798,N_10,N_2256);
or U4799 (N_4799,N_1873,N_1740);
nor U4800 (N_4800,N_619,N_2108);
or U4801 (N_4801,N_1057,N_417);
or U4802 (N_4802,N_1221,N_974);
nand U4803 (N_4803,N_790,N_2259);
nor U4804 (N_4804,N_2298,N_529);
nor U4805 (N_4805,N_453,N_514);
or U4806 (N_4806,N_578,N_1967);
nor U4807 (N_4807,N_1076,N_1672);
nand U4808 (N_4808,N_2173,N_443);
nor U4809 (N_4809,N_1499,N_1974);
nand U4810 (N_4810,N_718,N_48);
xor U4811 (N_4811,N_1524,N_578);
and U4812 (N_4812,N_1467,N_1391);
and U4813 (N_4813,N_166,N_955);
nand U4814 (N_4814,N_226,N_1912);
nand U4815 (N_4815,N_2278,N_1612);
and U4816 (N_4816,N_1453,N_1609);
and U4817 (N_4817,N_1858,N_2172);
nand U4818 (N_4818,N_917,N_1057);
nor U4819 (N_4819,N_229,N_2060);
nor U4820 (N_4820,N_252,N_208);
nor U4821 (N_4821,N_1322,N_713);
and U4822 (N_4822,N_898,N_1454);
nand U4823 (N_4823,N_758,N_186);
or U4824 (N_4824,N_2496,N_268);
nand U4825 (N_4825,N_1355,N_1855);
nor U4826 (N_4826,N_1771,N_2119);
or U4827 (N_4827,N_1654,N_1511);
nor U4828 (N_4828,N_74,N_436);
nand U4829 (N_4829,N_1683,N_2092);
or U4830 (N_4830,N_622,N_1041);
nor U4831 (N_4831,N_2055,N_908);
or U4832 (N_4832,N_2179,N_1198);
nor U4833 (N_4833,N_301,N_131);
and U4834 (N_4834,N_2101,N_992);
or U4835 (N_4835,N_269,N_1622);
nor U4836 (N_4836,N_878,N_1456);
and U4837 (N_4837,N_326,N_965);
nand U4838 (N_4838,N_1536,N_568);
nand U4839 (N_4839,N_1533,N_1913);
nand U4840 (N_4840,N_2313,N_2494);
nand U4841 (N_4841,N_375,N_1591);
nor U4842 (N_4842,N_2119,N_2442);
nor U4843 (N_4843,N_1070,N_2094);
nand U4844 (N_4844,N_1765,N_788);
nor U4845 (N_4845,N_182,N_1632);
and U4846 (N_4846,N_1970,N_1986);
or U4847 (N_4847,N_799,N_2249);
nand U4848 (N_4848,N_1712,N_2034);
nor U4849 (N_4849,N_1015,N_521);
and U4850 (N_4850,N_1469,N_259);
nand U4851 (N_4851,N_7,N_1625);
nor U4852 (N_4852,N_1997,N_1386);
nand U4853 (N_4853,N_1825,N_251);
or U4854 (N_4854,N_1025,N_741);
xor U4855 (N_4855,N_2406,N_791);
and U4856 (N_4856,N_174,N_535);
nand U4857 (N_4857,N_165,N_493);
nand U4858 (N_4858,N_1339,N_183);
or U4859 (N_4859,N_282,N_154);
nand U4860 (N_4860,N_1212,N_2159);
or U4861 (N_4861,N_2070,N_2482);
nand U4862 (N_4862,N_1540,N_557);
nor U4863 (N_4863,N_1028,N_125);
nand U4864 (N_4864,N_2097,N_1593);
nand U4865 (N_4865,N_1722,N_2298);
and U4866 (N_4866,N_1227,N_1083);
nor U4867 (N_4867,N_277,N_2024);
nand U4868 (N_4868,N_973,N_1714);
nand U4869 (N_4869,N_1097,N_48);
nor U4870 (N_4870,N_2050,N_641);
nand U4871 (N_4871,N_1789,N_1052);
nand U4872 (N_4872,N_263,N_1065);
nor U4873 (N_4873,N_2402,N_422);
or U4874 (N_4874,N_1007,N_1262);
nand U4875 (N_4875,N_2074,N_808);
nor U4876 (N_4876,N_2039,N_919);
nand U4877 (N_4877,N_1885,N_404);
and U4878 (N_4878,N_1810,N_1501);
or U4879 (N_4879,N_2250,N_781);
nand U4880 (N_4880,N_1272,N_1921);
nand U4881 (N_4881,N_1115,N_303);
xor U4882 (N_4882,N_1434,N_378);
nor U4883 (N_4883,N_198,N_369);
nand U4884 (N_4884,N_422,N_1477);
or U4885 (N_4885,N_1223,N_1438);
and U4886 (N_4886,N_385,N_1252);
or U4887 (N_4887,N_86,N_537);
and U4888 (N_4888,N_425,N_1681);
nand U4889 (N_4889,N_1350,N_123);
or U4890 (N_4890,N_1729,N_2425);
nor U4891 (N_4891,N_51,N_1500);
and U4892 (N_4892,N_478,N_2222);
or U4893 (N_4893,N_98,N_836);
nor U4894 (N_4894,N_806,N_1461);
nor U4895 (N_4895,N_2297,N_1614);
nand U4896 (N_4896,N_1483,N_1796);
xnor U4897 (N_4897,N_813,N_554);
nor U4898 (N_4898,N_1539,N_512);
or U4899 (N_4899,N_1180,N_1513);
and U4900 (N_4900,N_2404,N_2180);
nor U4901 (N_4901,N_2141,N_1060);
and U4902 (N_4902,N_823,N_2157);
nand U4903 (N_4903,N_2391,N_1182);
or U4904 (N_4904,N_103,N_1541);
or U4905 (N_4905,N_2272,N_2190);
and U4906 (N_4906,N_2072,N_1239);
nor U4907 (N_4907,N_776,N_1503);
or U4908 (N_4908,N_146,N_1307);
or U4909 (N_4909,N_386,N_205);
or U4910 (N_4910,N_1353,N_891);
nor U4911 (N_4911,N_1015,N_813);
and U4912 (N_4912,N_624,N_2268);
and U4913 (N_4913,N_19,N_438);
nor U4914 (N_4914,N_1110,N_1320);
and U4915 (N_4915,N_844,N_2450);
nor U4916 (N_4916,N_2415,N_1447);
nor U4917 (N_4917,N_361,N_141);
or U4918 (N_4918,N_536,N_596);
or U4919 (N_4919,N_1306,N_254);
nor U4920 (N_4920,N_1869,N_291);
and U4921 (N_4921,N_1925,N_1196);
or U4922 (N_4922,N_404,N_1404);
nand U4923 (N_4923,N_1141,N_2058);
xnor U4924 (N_4924,N_708,N_2404);
nand U4925 (N_4925,N_1602,N_284);
and U4926 (N_4926,N_377,N_395);
and U4927 (N_4927,N_2496,N_439);
nor U4928 (N_4928,N_1522,N_64);
or U4929 (N_4929,N_511,N_2047);
nor U4930 (N_4930,N_674,N_879);
and U4931 (N_4931,N_455,N_1952);
or U4932 (N_4932,N_737,N_16);
nor U4933 (N_4933,N_2390,N_160);
or U4934 (N_4934,N_881,N_1287);
nor U4935 (N_4935,N_982,N_192);
nand U4936 (N_4936,N_1213,N_1266);
nand U4937 (N_4937,N_540,N_840);
nand U4938 (N_4938,N_88,N_1648);
or U4939 (N_4939,N_315,N_177);
and U4940 (N_4940,N_641,N_475);
nand U4941 (N_4941,N_1054,N_1177);
and U4942 (N_4942,N_1054,N_525);
or U4943 (N_4943,N_1815,N_109);
nand U4944 (N_4944,N_157,N_1778);
nand U4945 (N_4945,N_683,N_875);
nor U4946 (N_4946,N_53,N_977);
or U4947 (N_4947,N_1777,N_189);
nor U4948 (N_4948,N_1614,N_283);
nor U4949 (N_4949,N_2131,N_77);
nor U4950 (N_4950,N_2196,N_2405);
nand U4951 (N_4951,N_495,N_378);
and U4952 (N_4952,N_2,N_15);
or U4953 (N_4953,N_280,N_1649);
and U4954 (N_4954,N_104,N_2244);
or U4955 (N_4955,N_17,N_1928);
nand U4956 (N_4956,N_2434,N_1484);
nand U4957 (N_4957,N_420,N_106);
nor U4958 (N_4958,N_2267,N_714);
nand U4959 (N_4959,N_2211,N_895);
and U4960 (N_4960,N_789,N_2372);
nand U4961 (N_4961,N_1129,N_2202);
and U4962 (N_4962,N_1063,N_1765);
and U4963 (N_4963,N_865,N_1078);
nor U4964 (N_4964,N_1832,N_127);
or U4965 (N_4965,N_396,N_285);
and U4966 (N_4966,N_640,N_2205);
nor U4967 (N_4967,N_750,N_2175);
nand U4968 (N_4968,N_1625,N_282);
or U4969 (N_4969,N_1443,N_1183);
nand U4970 (N_4970,N_1319,N_2034);
and U4971 (N_4971,N_2206,N_14);
or U4972 (N_4972,N_2254,N_987);
and U4973 (N_4973,N_1309,N_2198);
nand U4974 (N_4974,N_1292,N_1294);
and U4975 (N_4975,N_801,N_1493);
nor U4976 (N_4976,N_1694,N_2332);
and U4977 (N_4977,N_289,N_694);
nand U4978 (N_4978,N_2358,N_289);
xnor U4979 (N_4979,N_1082,N_1844);
nand U4980 (N_4980,N_1498,N_207);
and U4981 (N_4981,N_694,N_1226);
nor U4982 (N_4982,N_1406,N_1342);
nor U4983 (N_4983,N_470,N_439);
and U4984 (N_4984,N_915,N_1129);
nand U4985 (N_4985,N_642,N_1128);
nor U4986 (N_4986,N_903,N_2472);
nand U4987 (N_4987,N_1044,N_1427);
nand U4988 (N_4988,N_2026,N_881);
nand U4989 (N_4989,N_1849,N_811);
nor U4990 (N_4990,N_1073,N_1397);
and U4991 (N_4991,N_1181,N_2242);
nand U4992 (N_4992,N_2107,N_768);
nor U4993 (N_4993,N_373,N_691);
nor U4994 (N_4994,N_1211,N_690);
and U4995 (N_4995,N_2098,N_1600);
nand U4996 (N_4996,N_121,N_1399);
or U4997 (N_4997,N_2266,N_1156);
nor U4998 (N_4998,N_345,N_1057);
and U4999 (N_4999,N_1357,N_1002);
and U5000 (N_5000,N_4147,N_3182);
nor U5001 (N_5001,N_2628,N_2937);
nor U5002 (N_5002,N_4353,N_3920);
nand U5003 (N_5003,N_4197,N_3946);
nand U5004 (N_5004,N_2824,N_4131);
nor U5005 (N_5005,N_4372,N_3836);
and U5006 (N_5006,N_4616,N_3556);
and U5007 (N_5007,N_3979,N_3413);
or U5008 (N_5008,N_3116,N_3329);
or U5009 (N_5009,N_4395,N_3720);
or U5010 (N_5010,N_3553,N_4941);
and U5011 (N_5011,N_3433,N_3305);
nor U5012 (N_5012,N_2781,N_3658);
nand U5013 (N_5013,N_3013,N_2998);
and U5014 (N_5014,N_2896,N_4640);
and U5015 (N_5015,N_3762,N_2785);
or U5016 (N_5016,N_4290,N_4219);
nand U5017 (N_5017,N_2554,N_3494);
or U5018 (N_5018,N_2738,N_4889);
nor U5019 (N_5019,N_2873,N_3291);
and U5020 (N_5020,N_4875,N_3848);
nand U5021 (N_5021,N_3825,N_3301);
nand U5022 (N_5022,N_2877,N_3648);
or U5023 (N_5023,N_2548,N_2701);
or U5024 (N_5024,N_4924,N_4442);
or U5025 (N_5025,N_3128,N_2776);
or U5026 (N_5026,N_4095,N_3109);
nor U5027 (N_5027,N_3850,N_4417);
nand U5028 (N_5028,N_4970,N_3893);
or U5029 (N_5029,N_2968,N_4311);
and U5030 (N_5030,N_4898,N_2811);
nand U5031 (N_5031,N_2804,N_4802);
and U5032 (N_5032,N_3371,N_4226);
nand U5033 (N_5033,N_2726,N_3726);
and U5034 (N_5034,N_2592,N_4482);
or U5035 (N_5035,N_2611,N_3035);
nand U5036 (N_5036,N_3197,N_3717);
nor U5037 (N_5037,N_4656,N_2580);
and U5038 (N_5038,N_3174,N_4388);
or U5039 (N_5039,N_4159,N_3385);
or U5040 (N_5040,N_2661,N_3328);
nand U5041 (N_5041,N_3936,N_4491);
nor U5042 (N_5042,N_2624,N_3377);
xnor U5043 (N_5043,N_3210,N_4668);
nor U5044 (N_5044,N_3804,N_3111);
nor U5045 (N_5045,N_4922,N_4546);
nand U5046 (N_5046,N_3749,N_4454);
or U5047 (N_5047,N_3906,N_4060);
nand U5048 (N_5048,N_4416,N_4078);
nand U5049 (N_5049,N_3084,N_3925);
nor U5050 (N_5050,N_4637,N_3297);
and U5051 (N_5051,N_4854,N_4620);
and U5052 (N_5052,N_4070,N_4991);
nor U5053 (N_5053,N_3712,N_3792);
nand U5054 (N_5054,N_3916,N_3045);
nor U5055 (N_5055,N_4660,N_4731);
nor U5056 (N_5056,N_4526,N_3962);
nand U5057 (N_5057,N_4608,N_3959);
and U5058 (N_5058,N_3880,N_4917);
nor U5059 (N_5059,N_4590,N_3968);
or U5060 (N_5060,N_3955,N_4088);
or U5061 (N_5061,N_2986,N_2637);
and U5062 (N_5062,N_3805,N_3540);
nand U5063 (N_5063,N_2994,N_3692);
nor U5064 (N_5064,N_4401,N_3872);
nor U5065 (N_5065,N_3330,N_3349);
nor U5066 (N_5066,N_4659,N_3633);
nor U5067 (N_5067,N_4649,N_2865);
or U5068 (N_5068,N_2575,N_2569);
nor U5069 (N_5069,N_3500,N_3740);
nand U5070 (N_5070,N_4465,N_3732);
or U5071 (N_5071,N_2845,N_3405);
nand U5072 (N_5072,N_3632,N_4164);
and U5073 (N_5073,N_3316,N_3739);
nand U5074 (N_5074,N_3711,N_4581);
and U5075 (N_5075,N_4457,N_3076);
nor U5076 (N_5076,N_4537,N_4004);
and U5077 (N_5077,N_4080,N_4053);
and U5078 (N_5078,N_3905,N_4574);
and U5079 (N_5079,N_2979,N_4771);
or U5080 (N_5080,N_4866,N_4634);
or U5081 (N_5081,N_3978,N_3830);
nor U5082 (N_5082,N_2832,N_4143);
nand U5083 (N_5083,N_4202,N_4342);
nand U5084 (N_5084,N_3320,N_3376);
or U5085 (N_5085,N_2692,N_3131);
and U5086 (N_5086,N_3409,N_4486);
or U5087 (N_5087,N_3422,N_4603);
nor U5088 (N_5088,N_4007,N_3323);
and U5089 (N_5089,N_3048,N_4560);
and U5090 (N_5090,N_4030,N_3317);
nor U5091 (N_5091,N_4303,N_2674);
nor U5092 (N_5092,N_2601,N_3187);
or U5093 (N_5093,N_4554,N_3009);
or U5094 (N_5094,N_2576,N_3492);
nor U5095 (N_5095,N_4119,N_4717);
and U5096 (N_5096,N_2612,N_4886);
nand U5097 (N_5097,N_4447,N_4831);
nor U5098 (N_5098,N_2943,N_3488);
and U5099 (N_5099,N_2634,N_4432);
nand U5100 (N_5100,N_3304,N_4425);
and U5101 (N_5101,N_2844,N_3584);
and U5102 (N_5102,N_4163,N_4065);
nand U5103 (N_5103,N_2836,N_4724);
nand U5104 (N_5104,N_4497,N_3497);
or U5105 (N_5105,N_4024,N_3443);
or U5106 (N_5106,N_2679,N_3350);
nand U5107 (N_5107,N_3403,N_3242);
nand U5108 (N_5108,N_4257,N_4777);
and U5109 (N_5109,N_3458,N_3679);
nor U5110 (N_5110,N_2620,N_4414);
and U5111 (N_5111,N_4788,N_4208);
nor U5112 (N_5112,N_4250,N_4180);
xnor U5113 (N_5113,N_3032,N_4796);
and U5114 (N_5114,N_4074,N_3236);
nand U5115 (N_5115,N_3384,N_2740);
and U5116 (N_5116,N_3460,N_3463);
and U5117 (N_5117,N_3469,N_3826);
nand U5118 (N_5118,N_2952,N_4089);
nor U5119 (N_5119,N_3431,N_4259);
nor U5120 (N_5120,N_4453,N_2660);
nor U5121 (N_5121,N_3815,N_3481);
and U5122 (N_5122,N_4273,N_3410);
and U5123 (N_5123,N_2543,N_4234);
nand U5124 (N_5124,N_3067,N_3266);
nor U5125 (N_5125,N_3787,N_4549);
nor U5126 (N_5126,N_4309,N_2887);
nor U5127 (N_5127,N_2848,N_3573);
nor U5128 (N_5128,N_3104,N_2756);
nand U5129 (N_5129,N_4919,N_3364);
nand U5130 (N_5130,N_3402,N_3490);
or U5131 (N_5131,N_4185,N_2523);
nand U5132 (N_5132,N_4888,N_3202);
nor U5133 (N_5133,N_2571,N_4695);
and U5134 (N_5134,N_2745,N_3241);
nor U5135 (N_5135,N_3406,N_4179);
nand U5136 (N_5136,N_3583,N_3884);
or U5137 (N_5137,N_4278,N_3341);
xnor U5138 (N_5138,N_4043,N_4613);
and U5139 (N_5139,N_3506,N_3185);
nor U5140 (N_5140,N_3258,N_2878);
nand U5141 (N_5141,N_2656,N_2531);
nand U5142 (N_5142,N_4751,N_4930);
and U5143 (N_5143,N_2578,N_4572);
or U5144 (N_5144,N_2525,N_4085);
xor U5145 (N_5145,N_4477,N_3821);
nand U5146 (N_5146,N_4003,N_3235);
and U5147 (N_5147,N_4748,N_3782);
or U5148 (N_5148,N_2838,N_3829);
or U5149 (N_5149,N_2515,N_3641);
nor U5150 (N_5150,N_4161,N_3003);
or U5151 (N_5151,N_3219,N_3252);
and U5152 (N_5152,N_4284,N_2553);
nor U5153 (N_5153,N_4139,N_3140);
or U5154 (N_5154,N_3943,N_3719);
or U5155 (N_5155,N_4026,N_4718);
or U5156 (N_5156,N_3548,N_3681);
nor U5157 (N_5157,N_4481,N_3630);
or U5158 (N_5158,N_3387,N_2524);
nor U5159 (N_5159,N_4441,N_4715);
nand U5160 (N_5160,N_4364,N_3485);
or U5161 (N_5161,N_2860,N_4765);
nand U5162 (N_5162,N_4320,N_3614);
xor U5163 (N_5163,N_3576,N_4628);
or U5164 (N_5164,N_4846,N_3809);
or U5165 (N_5165,N_4845,N_4907);
and U5166 (N_5166,N_3984,N_2762);
or U5167 (N_5167,N_4368,N_3703);
nand U5168 (N_5168,N_3521,N_4969);
nand U5169 (N_5169,N_4791,N_3053);
nand U5170 (N_5170,N_3563,N_4515);
or U5171 (N_5171,N_4992,N_3801);
nor U5172 (N_5172,N_3810,N_3066);
and U5173 (N_5173,N_3878,N_4399);
and U5174 (N_5174,N_4101,N_4582);
nor U5175 (N_5175,N_4727,N_2849);
nor U5176 (N_5176,N_3147,N_3747);
nor U5177 (N_5177,N_3216,N_3399);
and U5178 (N_5178,N_4997,N_3026);
or U5179 (N_5179,N_4794,N_3750);
nand U5180 (N_5180,N_3107,N_3730);
nand U5181 (N_5181,N_4487,N_4822);
nand U5182 (N_5182,N_3274,N_2978);
nor U5183 (N_5183,N_4901,N_3496);
or U5184 (N_5184,N_4485,N_3394);
nand U5185 (N_5185,N_4819,N_3081);
and U5186 (N_5186,N_2803,N_2714);
nor U5187 (N_5187,N_4955,N_4697);
and U5188 (N_5188,N_4870,N_4657);
and U5189 (N_5189,N_3106,N_3899);
or U5190 (N_5190,N_2667,N_4867);
and U5191 (N_5191,N_4172,N_3868);
or U5192 (N_5192,N_2972,N_3518);
or U5193 (N_5193,N_4424,N_3987);
nor U5194 (N_5194,N_2830,N_4156);
nand U5195 (N_5195,N_2895,N_4860);
nand U5196 (N_5196,N_4701,N_4929);
nor U5197 (N_5197,N_3549,N_3155);
or U5198 (N_5198,N_4123,N_4224);
or U5199 (N_5199,N_2893,N_2642);
and U5200 (N_5200,N_3926,N_4528);
and U5201 (N_5201,N_4036,N_2862);
nor U5202 (N_5202,N_4382,N_3493);
or U5203 (N_5203,N_3339,N_3603);
nor U5204 (N_5204,N_2517,N_4979);
nand U5205 (N_5205,N_3306,N_3284);
nand U5206 (N_5206,N_4687,N_2572);
or U5207 (N_5207,N_3434,N_3575);
and U5208 (N_5208,N_4102,N_4877);
nor U5209 (N_5209,N_2884,N_2956);
nor U5210 (N_5210,N_2589,N_4367);
and U5211 (N_5211,N_4496,N_4317);
nand U5212 (N_5212,N_3662,N_3487);
nor U5213 (N_5213,N_4621,N_4797);
nor U5214 (N_5214,N_4965,N_3578);
and U5215 (N_5215,N_2566,N_3322);
nor U5216 (N_5216,N_3914,N_3784);
nand U5217 (N_5217,N_3967,N_2669);
and U5218 (N_5218,N_3158,N_4712);
nor U5219 (N_5219,N_2919,N_4210);
nand U5220 (N_5220,N_3283,N_4335);
nor U5221 (N_5221,N_4019,N_2530);
nor U5222 (N_5222,N_2960,N_2795);
nor U5223 (N_5223,N_4981,N_4840);
nand U5224 (N_5224,N_3949,N_3938);
nor U5225 (N_5225,N_4493,N_3522);
nor U5226 (N_5226,N_3861,N_3999);
nand U5227 (N_5227,N_3708,N_3800);
nor U5228 (N_5228,N_2903,N_2724);
nand U5229 (N_5229,N_4162,N_3990);
nor U5230 (N_5230,N_3470,N_3477);
or U5231 (N_5231,N_2899,N_3022);
nand U5232 (N_5232,N_4610,N_3611);
or U5233 (N_5233,N_2987,N_4990);
and U5234 (N_5234,N_4556,N_3819);
xnor U5235 (N_5235,N_4461,N_2666);
nand U5236 (N_5236,N_2552,N_4968);
and U5237 (N_5237,N_2562,N_3977);
or U5238 (N_5238,N_4206,N_3562);
or U5239 (N_5239,N_4787,N_2703);
and U5240 (N_5240,N_3253,N_3550);
nor U5241 (N_5241,N_2573,N_4033);
nor U5242 (N_5242,N_4938,N_4275);
nand U5243 (N_5243,N_4961,N_4196);
or U5244 (N_5244,N_4121,N_3054);
nor U5245 (N_5245,N_4440,N_2625);
and U5246 (N_5246,N_3774,N_3234);
and U5247 (N_5247,N_3876,N_4918);
nand U5248 (N_5248,N_4389,N_4795);
or U5249 (N_5249,N_3031,N_4527);
nor U5250 (N_5250,N_3450,N_4125);
nand U5251 (N_5251,N_3890,N_4566);
or U5252 (N_5252,N_2509,N_3199);
and U5253 (N_5253,N_4562,N_4002);
nand U5254 (N_5254,N_4669,N_3640);
nor U5255 (N_5255,N_2591,N_3451);
nand U5256 (N_5256,N_4696,N_3859);
or U5257 (N_5257,N_4861,N_4512);
nor U5258 (N_5258,N_2755,N_3741);
nand U5259 (N_5259,N_4508,N_4267);
nand U5260 (N_5260,N_4058,N_4283);
or U5261 (N_5261,N_2834,N_4577);
or U5262 (N_5262,N_2505,N_4248);
nand U5263 (N_5263,N_3933,N_2963);
or U5264 (N_5264,N_4611,N_3411);
nor U5265 (N_5265,N_3367,N_4298);
nand U5266 (N_5266,N_4381,N_2742);
nor U5267 (N_5267,N_3318,N_3154);
or U5268 (N_5268,N_4539,N_3621);
and U5269 (N_5269,N_4808,N_4218);
and U5270 (N_5270,N_4827,N_4271);
nor U5271 (N_5271,N_3997,N_2833);
or U5272 (N_5272,N_3204,N_3319);
and U5273 (N_5273,N_3922,N_4948);
or U5274 (N_5274,N_3516,N_3218);
and U5275 (N_5275,N_4587,N_4347);
or U5276 (N_5276,N_2704,N_3724);
nand U5277 (N_5277,N_4413,N_4510);
or U5278 (N_5278,N_2827,N_3645);
and U5279 (N_5279,N_3668,N_4314);
nand U5280 (N_5280,N_3574,N_3822);
and U5281 (N_5281,N_2971,N_3956);
nand U5282 (N_5282,N_2613,N_3754);
or U5283 (N_5283,N_3159,N_3526);
nand U5284 (N_5284,N_4722,N_3760);
nor U5285 (N_5285,N_3709,N_3300);
nand U5286 (N_5286,N_2922,N_4470);
and U5287 (N_5287,N_4571,N_3119);
or U5288 (N_5288,N_3271,N_4914);
or U5289 (N_5289,N_3127,N_4263);
or U5290 (N_5290,N_3927,N_2521);
and U5291 (N_5291,N_3126,N_4768);
nand U5292 (N_5292,N_3646,N_3386);
nor U5293 (N_5293,N_4650,N_4490);
nor U5294 (N_5294,N_4268,N_4944);
nor U5295 (N_5295,N_3517,N_4895);
and U5296 (N_5296,N_4471,N_3163);
or U5297 (N_5297,N_4132,N_4770);
nand U5298 (N_5298,N_4458,N_3857);
nand U5299 (N_5299,N_3459,N_3964);
nand U5300 (N_5300,N_4985,N_3923);
nand U5301 (N_5301,N_4792,N_2938);
or U5302 (N_5302,N_3802,N_3581);
and U5303 (N_5303,N_4176,N_2850);
and U5304 (N_5304,N_2821,N_3655);
nand U5305 (N_5305,N_3838,N_4468);
and U5306 (N_5306,N_3212,N_2748);
or U5307 (N_5307,N_3535,N_2853);
and U5308 (N_5308,N_4667,N_4800);
or U5309 (N_5309,N_4115,N_4324);
nand U5310 (N_5310,N_4127,N_4699);
and U5311 (N_5311,N_2977,N_3078);
or U5312 (N_5312,N_4373,N_4077);
or U5313 (N_5313,N_4051,N_2761);
or U5314 (N_5314,N_4448,N_4811);
and U5315 (N_5315,N_2528,N_4570);
and U5316 (N_5316,N_3853,N_4021);
and U5317 (N_5317,N_2790,N_4048);
nor U5318 (N_5318,N_4292,N_4285);
or U5319 (N_5319,N_4222,N_3285);
nor U5320 (N_5320,N_3156,N_3312);
and U5321 (N_5321,N_3102,N_2542);
nor U5322 (N_5322,N_2607,N_2951);
and U5323 (N_5323,N_3108,N_3206);
and U5324 (N_5324,N_3452,N_4144);
or U5325 (N_5325,N_3074,N_3783);
or U5326 (N_5326,N_3120,N_4553);
nand U5327 (N_5327,N_2915,N_4069);
or U5328 (N_5328,N_4034,N_3577);
nor U5329 (N_5329,N_2680,N_3846);
nand U5330 (N_5330,N_3125,N_3524);
nand U5331 (N_5331,N_2683,N_3737);
nor U5332 (N_5332,N_3609,N_3834);
and U5333 (N_5333,N_3296,N_4439);
and U5334 (N_5334,N_3093,N_4774);
and U5335 (N_5335,N_3671,N_4396);
nor U5336 (N_5336,N_4277,N_4322);
nor U5337 (N_5337,N_2947,N_4641);
nand U5338 (N_5338,N_2995,N_3813);
nor U5339 (N_5339,N_2647,N_4685);
and U5340 (N_5340,N_4246,N_2638);
nand U5341 (N_5341,N_4551,N_4882);
nor U5342 (N_5342,N_3921,N_2969);
nand U5343 (N_5343,N_3634,N_4092);
nor U5344 (N_5344,N_3864,N_3795);
nand U5345 (N_5345,N_3250,N_2710);
nand U5346 (N_5346,N_3798,N_4357);
nor U5347 (N_5347,N_4518,N_3596);
or U5348 (N_5348,N_3725,N_4460);
nand U5349 (N_5349,N_3699,N_4530);
and U5350 (N_5350,N_4906,N_3908);
and U5351 (N_5351,N_2962,N_4823);
and U5352 (N_5352,N_3992,N_3336);
nand U5353 (N_5353,N_3309,N_3653);
and U5354 (N_5354,N_2501,N_4511);
and U5355 (N_5355,N_3618,N_3198);
and U5356 (N_5356,N_4564,N_3298);
or U5357 (N_5357,N_4578,N_2691);
and U5358 (N_5358,N_3950,N_4192);
or U5359 (N_5359,N_4343,N_4844);
or U5360 (N_5360,N_3259,N_3001);
and U5361 (N_5361,N_4595,N_2746);
nor U5362 (N_5362,N_3767,N_4896);
nand U5363 (N_5363,N_4666,N_2633);
or U5364 (N_5364,N_4923,N_4466);
nor U5365 (N_5365,N_3040,N_2693);
and U5366 (N_5366,N_4837,N_4557);
nor U5367 (N_5367,N_3696,N_3270);
nand U5368 (N_5368,N_4730,N_3844);
or U5369 (N_5369,N_4747,N_4903);
nor U5370 (N_5370,N_3347,N_2813);
or U5371 (N_5371,N_4175,N_3482);
nor U5372 (N_5372,N_2942,N_3333);
nor U5373 (N_5373,N_3568,N_4384);
nand U5374 (N_5374,N_2739,N_4063);
or U5375 (N_5375,N_2786,N_2897);
or U5376 (N_5376,N_4850,N_3221);
and U5377 (N_5377,N_2920,N_3590);
nor U5378 (N_5378,N_4203,N_4756);
nor U5379 (N_5379,N_2914,N_4517);
and U5380 (N_5380,N_4585,N_3510);
and U5381 (N_5381,N_4690,N_4568);
nor U5382 (N_5382,N_3569,N_4920);
or U5383 (N_5383,N_4719,N_3215);
nand U5384 (N_5384,N_2711,N_2876);
nor U5385 (N_5385,N_3372,N_2616);
or U5386 (N_5386,N_2825,N_2551);
and U5387 (N_5387,N_4565,N_4062);
nand U5388 (N_5388,N_3080,N_3501);
and U5389 (N_5389,N_3513,N_2940);
nor U5390 (N_5390,N_4893,N_3303);
nor U5391 (N_5391,N_4182,N_2772);
nor U5392 (N_5392,N_4394,N_3847);
nand U5393 (N_5393,N_3095,N_3690);
nor U5394 (N_5394,N_4812,N_4438);
nor U5395 (N_5395,N_3585,N_4251);
and U5396 (N_5396,N_4056,N_3171);
or U5397 (N_5397,N_3995,N_3960);
nand U5398 (N_5398,N_3167,N_4201);
nand U5399 (N_5399,N_4632,N_4044);
and U5400 (N_5400,N_4232,N_4535);
nor U5401 (N_5401,N_3564,N_4931);
or U5402 (N_5402,N_3014,N_4529);
and U5403 (N_5403,N_2904,N_3512);
nand U5404 (N_5404,N_3797,N_4307);
nor U5405 (N_5405,N_4361,N_2584);
or U5406 (N_5406,N_2730,N_4684);
nand U5407 (N_5407,N_4910,N_3896);
nor U5408 (N_5408,N_4057,N_3058);
nand U5409 (N_5409,N_4655,N_4714);
nor U5410 (N_5410,N_3932,N_4223);
and U5411 (N_5411,N_4761,N_2950);
nand U5412 (N_5412,N_4514,N_4694);
nand U5413 (N_5413,N_2864,N_2949);
and U5414 (N_5414,N_3788,N_3390);
and U5415 (N_5415,N_2600,N_3000);
nor U5416 (N_5416,N_4341,N_4593);
nor U5417 (N_5417,N_4241,N_4779);
and U5418 (N_5418,N_4966,N_4061);
nor U5419 (N_5419,N_3909,N_3466);
nand U5420 (N_5420,N_4674,N_2538);
nor U5421 (N_5421,N_4445,N_3486);
and U5422 (N_5422,N_4291,N_4187);
nand U5423 (N_5423,N_4780,N_3263);
nand U5424 (N_5424,N_4816,N_3144);
nor U5425 (N_5425,N_2908,N_3059);
or U5426 (N_5426,N_4400,N_3771);
nand U5427 (N_5427,N_3184,N_4405);
or U5428 (N_5428,N_4456,N_4702);
and U5429 (N_5429,N_3276,N_3177);
and U5430 (N_5430,N_3358,N_3162);
nand U5431 (N_5431,N_4337,N_3700);
and U5432 (N_5432,N_3072,N_2640);
or U5433 (N_5433,N_2874,N_2526);
nand U5434 (N_5434,N_4964,N_4707);
nor U5435 (N_5435,N_3183,N_4113);
nand U5436 (N_5436,N_4793,N_3227);
nor U5437 (N_5437,N_4592,N_4782);
nand U5438 (N_5438,N_4605,N_4630);
or U5439 (N_5439,N_4000,N_4737);
nand U5440 (N_5440,N_4018,N_4946);
and U5441 (N_5441,N_2970,N_3468);
or U5442 (N_5442,N_4473,N_3015);
or U5443 (N_5443,N_4740,N_3380);
and U5444 (N_5444,N_3094,N_2775);
nor U5445 (N_5445,N_2644,N_3669);
or U5446 (N_5446,N_2750,N_4244);
nor U5447 (N_5447,N_4863,N_3768);
nor U5448 (N_5448,N_2597,N_2565);
nor U5449 (N_5449,N_3515,N_3400);
and U5450 (N_5450,N_2506,N_2799);
nor U5451 (N_5451,N_4576,N_2665);
or U5452 (N_5452,N_3345,N_4437);
nand U5453 (N_5453,N_3389,N_3855);
or U5454 (N_5454,N_3718,N_4746);
or U5455 (N_5455,N_3554,N_2757);
nor U5456 (N_5456,N_3793,N_3392);
and U5457 (N_5457,N_3430,N_4479);
nor U5458 (N_5458,N_4928,N_3680);
and U5459 (N_5459,N_3523,N_3145);
or U5460 (N_5460,N_3536,N_4904);
nand U5461 (N_5461,N_3153,N_3370);
or U5462 (N_5462,N_3244,N_4409);
nand U5463 (N_5463,N_3361,N_4339);
and U5464 (N_5464,N_4544,N_3401);
and U5465 (N_5465,N_4688,N_3617);
nor U5466 (N_5466,N_4327,N_3441);
nand U5467 (N_5467,N_2751,N_4894);
or U5468 (N_5468,N_4279,N_4094);
or U5469 (N_5469,N_2858,N_4936);
and U5470 (N_5470,N_4921,N_3817);
nor U5471 (N_5471,N_4661,N_2507);
and U5472 (N_5472,N_4871,N_3862);
nand U5473 (N_5473,N_2892,N_3693);
and U5474 (N_5474,N_3912,N_4723);
or U5475 (N_5475,N_4153,N_4642);
nand U5476 (N_5476,N_4807,N_3044);
nand U5477 (N_5477,N_4207,N_4186);
or U5478 (N_5478,N_3539,N_3944);
nand U5479 (N_5479,N_3148,N_4813);
nor U5480 (N_5480,N_3917,N_2901);
nand U5481 (N_5481,N_4825,N_2841);
or U5482 (N_5482,N_4954,N_2609);
nor U5483 (N_5483,N_3706,N_3592);
and U5484 (N_5484,N_3417,N_3308);
or U5485 (N_5485,N_2654,N_3663);
nand U5486 (N_5486,N_4776,N_4494);
nor U5487 (N_5487,N_4803,N_3610);
nand U5488 (N_5488,N_3464,N_2585);
nor U5489 (N_5489,N_4146,N_4829);
and U5490 (N_5490,N_3324,N_3427);
or U5491 (N_5491,N_4989,N_2539);
nor U5492 (N_5492,N_4167,N_4652);
or U5493 (N_5493,N_4011,N_3544);
nand U5494 (N_5494,N_3025,N_2659);
xnor U5495 (N_5495,N_4138,N_4711);
or U5496 (N_5496,N_2555,N_4504);
or U5497 (N_5497,N_4488,N_4880);
and U5498 (N_5498,N_3672,N_2645);
nand U5499 (N_5499,N_2626,N_3674);
and U5500 (N_5500,N_4194,N_4169);
and U5501 (N_5501,N_4272,N_3791);
nor U5502 (N_5502,N_2812,N_3315);
nor U5503 (N_5503,N_2558,N_3005);
or U5504 (N_5504,N_4261,N_4228);
nand U5505 (N_5505,N_2514,N_2948);
and U5506 (N_5506,N_3715,N_3937);
nor U5507 (N_5507,N_3019,N_4166);
and U5508 (N_5508,N_4155,N_3256);
and U5509 (N_5509,N_4635,N_2537);
nand U5510 (N_5510,N_2753,N_2723);
nand U5511 (N_5511,N_4407,N_4449);
nor U5512 (N_5512,N_3842,N_3265);
and U5513 (N_5513,N_2777,N_4977);
and U5514 (N_5514,N_3412,N_2955);
or U5515 (N_5515,N_4658,N_2867);
and U5516 (N_5516,N_3082,N_2907);
nand U5517 (N_5517,N_3223,N_2744);
xor U5518 (N_5518,N_4258,N_3873);
and U5519 (N_5519,N_3975,N_3453);
nor U5520 (N_5520,N_4205,N_4963);
and U5521 (N_5521,N_3713,N_3337);
or U5522 (N_5522,N_4325,N_4227);
nand U5523 (N_5523,N_3351,N_3207);
and U5524 (N_5524,N_4444,N_4098);
or U5525 (N_5525,N_3279,N_4856);
and U5526 (N_5526,N_3063,N_3247);
and U5527 (N_5527,N_3591,N_2502);
or U5528 (N_5528,N_4899,N_4858);
or U5529 (N_5529,N_2682,N_2641);
and U5530 (N_5530,N_3710,N_4545);
xnor U5531 (N_5531,N_2976,N_3904);
nor U5532 (N_5532,N_4391,N_3537);
and U5533 (N_5533,N_2635,N_3444);
or U5534 (N_5534,N_3894,N_4112);
and U5535 (N_5535,N_2518,N_4975);
nor U5536 (N_5536,N_4665,N_3192);
and U5537 (N_5537,N_4902,N_4874);
nand U5538 (N_5538,N_2854,N_2694);
and U5539 (N_5539,N_3666,N_2778);
or U5540 (N_5540,N_3624,N_2513);
nand U5541 (N_5541,N_4911,N_3302);
nor U5542 (N_5542,N_2699,N_3545);
or U5543 (N_5543,N_4499,N_2686);
and U5544 (N_5544,N_4096,N_3061);
nor U5545 (N_5545,N_3143,N_2925);
and U5546 (N_5546,N_3664,N_3856);
nor U5547 (N_5547,N_4001,N_4785);
nor U5548 (N_5548,N_3363,N_3294);
and U5549 (N_5549,N_3166,N_2747);
and U5550 (N_5550,N_4841,N_3678);
or U5551 (N_5551,N_4951,N_3100);
and U5552 (N_5552,N_3877,N_2946);
nand U5553 (N_5553,N_3114,N_3606);
or U5554 (N_5554,N_4976,N_3688);
or U5555 (N_5555,N_3449,N_2820);
or U5556 (N_5556,N_2535,N_3334);
nor U5557 (N_5557,N_4626,N_3023);
or U5558 (N_5558,N_3445,N_4828);
and U5559 (N_5559,N_3502,N_4081);
and U5560 (N_5560,N_4900,N_3806);
or U5561 (N_5561,N_3869,N_4643);
and U5562 (N_5562,N_2767,N_4726);
or U5563 (N_5563,N_2934,N_4297);
and U5564 (N_5564,N_2717,N_4580);
nand U5565 (N_5565,N_2696,N_4725);
and U5566 (N_5566,N_4170,N_4887);
or U5567 (N_5567,N_4378,N_2957);
and U5568 (N_5568,N_4198,N_3299);
and U5569 (N_5569,N_2603,N_4301);
or U5570 (N_5570,N_4212,N_3214);
and U5571 (N_5571,N_4358,N_4713);
nand U5572 (N_5572,N_3911,N_2818);
nand U5573 (N_5573,N_3635,N_4183);
nand U5574 (N_5574,N_4505,N_3652);
or U5575 (N_5575,N_3735,N_3897);
or U5576 (N_5576,N_3701,N_3335);
or U5577 (N_5577,N_4385,N_2540);
nand U5578 (N_5578,N_4993,N_3528);
and U5579 (N_5579,N_4862,N_4996);
nor U5580 (N_5580,N_4883,N_3728);
nand U5581 (N_5581,N_3803,N_3758);
and U5582 (N_5582,N_3217,N_2973);
nor U5583 (N_5583,N_4853,N_4306);
nor U5584 (N_5584,N_2754,N_3068);
or U5585 (N_5585,N_3928,N_4028);
or U5586 (N_5586,N_3599,N_4559);
and U5587 (N_5587,N_4348,N_3340);
nor U5588 (N_5588,N_4766,N_3673);
or U5589 (N_5589,N_2930,N_4937);
nand U5590 (N_5590,N_2814,N_4084);
nor U5591 (N_5591,N_4451,N_2549);
or U5592 (N_5592,N_2577,N_3073);
and U5593 (N_5593,N_4809,N_4738);
or U5594 (N_5594,N_3642,N_4949);
nand U5595 (N_5595,N_4878,N_2615);
nor U5596 (N_5596,N_3050,N_3112);
or U5597 (N_5597,N_3729,N_4463);
or U5598 (N_5598,N_4017,N_4624);
nand U5599 (N_5599,N_2636,N_3232);
nor U5600 (N_5600,N_2911,N_2852);
and U5601 (N_5601,N_3644,N_3004);
nor U5602 (N_5602,N_4220,N_3110);
or U5603 (N_5603,N_3360,N_3261);
nand U5604 (N_5604,N_3619,N_4542);
nor U5605 (N_5605,N_4604,N_4398);
nor U5606 (N_5606,N_4126,N_3559);
nand U5607 (N_5607,N_4371,N_3439);
and U5608 (N_5608,N_4848,N_4558);
nor U5609 (N_5609,N_4673,N_4633);
nor U5610 (N_5610,N_3251,N_4052);
and U5611 (N_5611,N_3142,N_4591);
and U5612 (N_5612,N_4607,N_2961);
nand U5613 (N_5613,N_4299,N_4599);
and U5614 (N_5614,N_3098,N_3875);
or U5615 (N_5615,N_4913,N_3533);
nand U5616 (N_5616,N_2861,N_3356);
and U5617 (N_5617,N_4075,N_4789);
nor U5618 (N_5618,N_2851,N_2631);
nand U5619 (N_5619,N_4264,N_3396);
or U5620 (N_5620,N_2671,N_3665);
or U5621 (N_5621,N_3414,N_4045);
nand U5622 (N_5622,N_3620,N_4638);
nor U5623 (N_5623,N_3379,N_2974);
nand U5624 (N_5624,N_2735,N_4947);
nor U5625 (N_5625,N_4124,N_3047);
nand U5626 (N_5626,N_2604,N_2520);
and U5627 (N_5627,N_4213,N_2688);
or U5628 (N_5628,N_4171,N_4269);
or U5629 (N_5629,N_4188,N_4749);
nand U5630 (N_5630,N_4849,N_4211);
or U5631 (N_5631,N_2632,N_4943);
nor U5632 (N_5632,N_4427,N_4059);
nor U5633 (N_5633,N_4178,N_4190);
and U5634 (N_5634,N_3970,N_3991);
nand U5635 (N_5635,N_2924,N_3461);
and U5636 (N_5636,N_4023,N_2872);
nor U5637 (N_5637,N_4274,N_3507);
nand U5638 (N_5638,N_3357,N_4799);
nand U5639 (N_5639,N_3814,N_2716);
or U5640 (N_5640,N_4729,N_3230);
nand U5641 (N_5641,N_4152,N_3772);
nor U5642 (N_5642,N_2536,N_2796);
and U5643 (N_5643,N_3423,N_3831);
or U5644 (N_5644,N_3687,N_3030);
nand U5645 (N_5645,N_4597,N_4333);
nand U5646 (N_5646,N_4393,N_3429);
and U5647 (N_5647,N_4265,N_3551);
or U5648 (N_5648,N_4679,N_4573);
nor U5649 (N_5649,N_2843,N_3179);
nor U5650 (N_5650,N_4010,N_4217);
or U5651 (N_5651,N_3716,N_2596);
or U5652 (N_5652,N_2828,N_3613);
and U5653 (N_5653,N_4455,N_2610);
nor U5654 (N_5654,N_4934,N_2568);
or U5655 (N_5655,N_3369,N_2719);
and U5656 (N_5656,N_3934,N_3704);
or U5657 (N_5657,N_4925,N_2689);
nand U5658 (N_5658,N_4588,N_4589);
or U5659 (N_5659,N_3683,N_4959);
nand U5660 (N_5660,N_4778,N_3193);
and U5661 (N_5661,N_3752,N_2605);
and U5662 (N_5662,N_3832,N_3029);
nand U5663 (N_5663,N_4513,N_4355);
nor U5664 (N_5664,N_3627,N_4872);
and U5665 (N_5665,N_3837,N_4230);
nor U5666 (N_5666,N_2508,N_4110);
nand U5667 (N_5667,N_4728,N_3761);
or U5668 (N_5668,N_2881,N_3541);
and U5669 (N_5669,N_2988,N_2886);
nor U5670 (N_5670,N_4374,N_4209);
nor U5671 (N_5671,N_3368,N_3115);
nor U5672 (N_5672,N_3457,N_4994);
nand U5673 (N_5673,N_4280,N_3373);
nor U5674 (N_5674,N_2787,N_3565);
nor U5675 (N_5675,N_3751,N_3608);
nand U5676 (N_5676,N_3677,N_3086);
nand U5677 (N_5677,N_4352,N_4752);
nand U5678 (N_5678,N_3191,N_3845);
and U5679 (N_5679,N_4134,N_4647);
or U5680 (N_5680,N_2765,N_2681);
or U5681 (N_5681,N_2687,N_3172);
nand U5682 (N_5682,N_3420,N_2743);
and U5683 (N_5683,N_2588,N_2700);
and U5684 (N_5684,N_4950,N_3508);
xor U5685 (N_5685,N_2650,N_4705);
nor U5686 (N_5686,N_3612,N_4104);
and U5687 (N_5687,N_4140,N_2939);
or U5688 (N_5688,N_3248,N_2856);
or U5689 (N_5689,N_3840,N_2593);
nand U5690 (N_5690,N_4181,N_4359);
and U5691 (N_5691,N_4945,N_2932);
and U5692 (N_5692,N_3675,N_4041);
and U5693 (N_5693,N_3989,N_2857);
nand U5694 (N_5694,N_2527,N_3343);
nand U5695 (N_5695,N_3604,N_4349);
or U5696 (N_5696,N_4027,N_3649);
and U5697 (N_5697,N_4067,N_4814);
nor U5698 (N_5698,N_2898,N_4998);
or U5699 (N_5699,N_4586,N_4820);
nor U5700 (N_5700,N_4760,N_2997);
and U5701 (N_5701,N_3480,N_4255);
nor U5702 (N_5702,N_3647,N_2918);
and U5703 (N_5703,N_4410,N_3629);
or U5704 (N_5704,N_4328,N_2889);
or U5705 (N_5705,N_2668,N_2882);
or U5706 (N_5706,N_4826,N_3395);
and U5707 (N_5707,N_2871,N_4967);
nand U5708 (N_5708,N_3656,N_3293);
nand U5709 (N_5709,N_3176,N_2729);
nor U5710 (N_5710,N_3188,N_3254);
nor U5711 (N_5711,N_4857,N_2880);
and U5712 (N_5712,N_3388,N_4149);
nor U5713 (N_5713,N_4313,N_4214);
nor U5714 (N_5714,N_2670,N_4254);
or U5715 (N_5715,N_4739,N_4029);
and U5716 (N_5716,N_3639,N_4974);
and U5717 (N_5717,N_4236,N_3954);
or U5718 (N_5718,N_4329,N_3201);
and U5719 (N_5719,N_3939,N_4009);
or U5720 (N_5720,N_2759,N_4832);
and U5721 (N_5721,N_4015,N_4534);
and U5722 (N_5722,N_4631,N_4693);
and U5723 (N_5723,N_3542,N_3682);
or U5724 (N_5724,N_3983,N_4336);
or U5725 (N_5725,N_3132,N_2733);
and U5726 (N_5726,N_2999,N_4524);
nand U5727 (N_5727,N_4247,N_3571);
nor U5728 (N_5728,N_4704,N_2639);
and U5729 (N_5729,N_3824,N_4645);
nand U5730 (N_5730,N_3615,N_2953);
and U5731 (N_5731,N_4908,N_4204);
and U5732 (N_5732,N_4020,N_3262);
or U5733 (N_5733,N_3287,N_4567);
or U5734 (N_5734,N_3462,N_2697);
nand U5735 (N_5735,N_4653,N_4680);
nor U5736 (N_5736,N_4745,N_3961);
or U5737 (N_5737,N_2805,N_3245);
or U5738 (N_5738,N_2840,N_3883);
nor U5739 (N_5739,N_2563,N_4318);
nor U5740 (N_5740,N_4376,N_2728);
nor U5741 (N_5741,N_4117,N_2771);
nand U5742 (N_5742,N_2912,N_4536);
or U5743 (N_5743,N_3200,N_2764);
or U5744 (N_5744,N_3657,N_3915);
or U5745 (N_5745,N_3736,N_3616);
nand U5746 (N_5746,N_3173,N_4602);
and U5747 (N_5747,N_4703,N_4689);
or U5748 (N_5748,N_4375,N_4054);
or U5749 (N_5749,N_4775,N_4569);
and U5750 (N_5750,N_3907,N_2931);
or U5751 (N_5751,N_3375,N_3090);
nor U5752 (N_5752,N_4338,N_3779);
or U5753 (N_5753,N_4216,N_4145);
and U5754 (N_5754,N_4129,N_4249);
or U5755 (N_5755,N_3882,N_4363);
and U5756 (N_5756,N_2594,N_3667);
nand U5757 (N_5757,N_3381,N_3888);
and U5758 (N_5758,N_4366,N_4988);
and U5759 (N_5759,N_3440,N_4135);
nand U5760 (N_5760,N_3566,N_2809);
nor U5761 (N_5761,N_4282,N_4881);
nand U5762 (N_5762,N_4885,N_3504);
and U5763 (N_5763,N_4459,N_4781);
nand U5764 (N_5764,N_4351,N_3532);
nor U5765 (N_5765,N_4193,N_3272);
nor U5766 (N_5766,N_3165,N_3233);
nor U5767 (N_5767,N_4741,N_2590);
nor U5768 (N_5768,N_2890,N_2866);
nor U5769 (N_5769,N_2883,N_2807);
or U5770 (N_5770,N_3070,N_3117);
nand U5771 (N_5771,N_4618,N_4744);
and U5772 (N_5772,N_3587,N_3391);
nor U5773 (N_5773,N_4855,N_2855);
nand U5774 (N_5774,N_4916,N_3495);
nand U5775 (N_5775,N_3124,N_4538);
and U5776 (N_5776,N_3756,N_3060);
and U5777 (N_5777,N_3691,N_4288);
or U5778 (N_5778,N_4326,N_2965);
or U5779 (N_5779,N_3697,N_4006);
nor U5780 (N_5780,N_2532,N_4681);
and U5781 (N_5781,N_3966,N_4253);
nor U5782 (N_5782,N_3024,N_4055);
nand U5783 (N_5783,N_3478,N_3881);
nand U5784 (N_5784,N_4046,N_2676);
and U5785 (N_5785,N_3123,N_3538);
or U5786 (N_5786,N_4676,N_3676);
or U5787 (N_5787,N_3224,N_4675);
and U5788 (N_5788,N_2816,N_3727);
nand U5789 (N_5789,N_3940,N_4522);
nor U5790 (N_5790,N_2651,N_3757);
and U5791 (N_5791,N_3973,N_4651);
and U5792 (N_5792,N_3139,N_2606);
nand U5793 (N_5793,N_2663,N_4397);
nor U5794 (N_5794,N_4952,N_4472);
nand U5795 (N_5795,N_2579,N_4281);
nand U5796 (N_5796,N_4215,N_4402);
or U5797 (N_5797,N_3404,N_3455);
nor U5798 (N_5798,N_4999,N_3901);
nand U5799 (N_5799,N_3134,N_3953);
or U5800 (N_5800,N_2736,N_3588);
xor U5801 (N_5801,N_3046,N_3910);
or U5802 (N_5802,N_3010,N_3092);
or U5803 (N_5803,N_3865,N_4252);
nand U5804 (N_5804,N_4435,N_3189);
or U5805 (N_5805,N_4677,N_2608);
nor U5806 (N_5806,N_2831,N_3190);
and U5807 (N_5807,N_3527,N_3879);
or U5808 (N_5808,N_2980,N_2910);
nor U5809 (N_5809,N_2783,N_3998);
nor U5810 (N_5810,N_4256,N_3733);
nor U5811 (N_5811,N_3101,N_4221);
nand U5812 (N_5812,N_4733,N_2715);
or U5813 (N_5813,N_3582,N_4106);
and U5814 (N_5814,N_3467,N_4130);
and U5815 (N_5815,N_3919,N_4810);
or U5816 (N_5816,N_4783,N_2928);
and U5817 (N_5817,N_4245,N_4897);
or U5818 (N_5818,N_4662,N_3625);
nor U5819 (N_5819,N_4184,N_3570);
nand U5820 (N_5820,N_3083,N_3240);
nand U5821 (N_5821,N_4073,N_4103);
nand U5822 (N_5822,N_3454,N_3354);
nand U5823 (N_5823,N_2695,N_2649);
nor U5824 (N_5824,N_2819,N_4933);
and U5825 (N_5825,N_4120,N_4354);
nor U5826 (N_5826,N_4710,N_2936);
or U5827 (N_5827,N_3650,N_4200);
or U5828 (N_5828,N_3898,N_4406);
nor U5829 (N_5829,N_4755,N_4289);
nand U5830 (N_5830,N_3530,N_3605);
or U5831 (N_5831,N_2823,N_2766);
nor U5832 (N_5832,N_3670,N_3579);
nand U5833 (N_5833,N_4225,N_4118);
or U5834 (N_5834,N_2826,N_4422);
nor U5835 (N_5835,N_3175,N_3065);
and U5836 (N_5836,N_3062,N_4821);
nor U5837 (N_5837,N_3456,N_4953);
or U5838 (N_5838,N_3208,N_4623);
or U5839 (N_5839,N_2614,N_3794);
and U5840 (N_5840,N_4876,N_2721);
nand U5841 (N_5841,N_2964,N_2529);
and U5842 (N_5842,N_2734,N_3442);
nor U5843 (N_5843,N_3765,N_4467);
nand U5844 (N_5844,N_2720,N_3169);
nand U5845 (N_5845,N_4984,N_4540);
nor U5846 (N_5846,N_4304,N_2586);
nor U5847 (N_5847,N_4072,N_2652);
nand U5848 (N_5848,N_3448,N_3327);
nor U5849 (N_5849,N_4750,N_4843);
or U5850 (N_5850,N_3012,N_3957);
nor U5851 (N_5851,N_4408,N_2557);
nand U5852 (N_5852,N_4801,N_3808);
nor U5853 (N_5853,N_3891,N_3344);
and U5854 (N_5854,N_4109,N_4547);
nand U5855 (N_5855,N_4978,N_4550);
or U5856 (N_5856,N_4958,N_3476);
and U5857 (N_5857,N_3511,N_4066);
or U5858 (N_5858,N_3011,N_3288);
and U5859 (N_5859,N_4474,N_4412);
nor U5860 (N_5860,N_3622,N_4418);
or U5861 (N_5861,N_4362,N_3714);
nor U5862 (N_5862,N_4068,N_2511);
nor U5863 (N_5863,N_4421,N_3498);
nand U5864 (N_5864,N_3534,N_3543);
nand U5865 (N_5865,N_2879,N_4040);
nor U5866 (N_5866,N_4644,N_4709);
or U5867 (N_5867,N_4443,N_4430);
nor U5868 (N_5868,N_3472,N_3295);
or U5869 (N_5869,N_4772,N_3852);
nor U5870 (N_5870,N_3246,N_4686);
nand U5871 (N_5871,N_3702,N_2900);
nand U5872 (N_5872,N_4022,N_2722);
nand U5873 (N_5873,N_3892,N_3332);
nand U5874 (N_5874,N_4583,N_3269);
nand U5875 (N_5875,N_3561,N_3348);
nand U5876 (N_5876,N_4141,N_2602);
and U5877 (N_5877,N_2797,N_3286);
and U5878 (N_5878,N_3008,N_3325);
nor U5879 (N_5879,N_3777,N_4377);
or U5880 (N_5880,N_4960,N_3407);
and U5881 (N_5881,N_3594,N_3870);
nand U5882 (N_5882,N_3763,N_4506);
nand U5883 (N_5883,N_3827,N_3555);
and U5884 (N_5884,N_4833,N_3428);
nor U5885 (N_5885,N_3273,N_4509);
and U5886 (N_5886,N_4229,N_3249);
nand U5887 (N_5887,N_3597,N_2583);
or U5888 (N_5888,N_4636,N_2789);
and U5889 (N_5889,N_4431,N_4757);
or U5890 (N_5890,N_4331,N_4295);
nor U5891 (N_5891,N_4035,N_3243);
nand U5892 (N_5892,N_4767,N_3151);
and U5893 (N_5893,N_2921,N_3426);
and U5894 (N_5894,N_3866,N_3734);
nand U5895 (N_5895,N_2675,N_2837);
and U5896 (N_5896,N_2713,N_4016);
nand U5897 (N_5897,N_4360,N_3871);
and U5898 (N_5898,N_2810,N_4464);
and U5899 (N_5899,N_4158,N_3133);
nand U5900 (N_5900,N_4671,N_2677);
or U5901 (N_5901,N_4076,N_3918);
nor U5902 (N_5902,N_4122,N_4852);
and U5903 (N_5903,N_2684,N_3796);
nand U5904 (N_5904,N_2545,N_3157);
and U5905 (N_5905,N_3651,N_2662);
or U5906 (N_5906,N_3886,N_2547);
nand U5907 (N_5907,N_4450,N_3421);
or U5908 (N_5908,N_3135,N_4716);
and U5909 (N_5909,N_3393,N_3280);
or U5910 (N_5910,N_4315,N_2582);
nand U5911 (N_5911,N_2891,N_2752);
or U5912 (N_5912,N_3557,N_3425);
or U5913 (N_5913,N_4365,N_3121);
or U5914 (N_5914,N_3948,N_2731);
nor U5915 (N_5915,N_4836,N_3220);
or U5916 (N_5916,N_2705,N_2737);
and U5917 (N_5917,N_4627,N_3705);
or U5918 (N_5918,N_4492,N_2885);
nor U5919 (N_5919,N_4957,N_4762);
nor U5920 (N_5920,N_3161,N_4769);
nand U5921 (N_5921,N_3525,N_3362);
and U5922 (N_5922,N_4165,N_2504);
nor U5923 (N_5923,N_3103,N_3986);
and U5924 (N_5924,N_3519,N_4008);
nor U5925 (N_5925,N_4563,N_3816);
nand U5926 (N_5926,N_4873,N_3408);
nand U5927 (N_5927,N_2712,N_3945);
nor U5928 (N_5928,N_4469,N_3985);
nor U5929 (N_5929,N_2560,N_2727);
and U5930 (N_5930,N_4935,N_4090);
nand U5931 (N_5931,N_4543,N_3007);
nand U5932 (N_5932,N_3436,N_4648);
and U5933 (N_5933,N_4191,N_3994);
and U5934 (N_5934,N_2690,N_3860);
and U5935 (N_5935,N_4742,N_2945);
or U5936 (N_5936,N_4345,N_2793);
nor U5937 (N_5937,N_3505,N_2774);
nor U5938 (N_5938,N_4334,N_3924);
or U5939 (N_5939,N_4423,N_4764);
nand U5940 (N_5940,N_4663,N_3203);
nand U5941 (N_5941,N_3503,N_4721);
and U5942 (N_5942,N_3257,N_2619);
or U5943 (N_5943,N_2773,N_3475);
nand U5944 (N_5944,N_3695,N_4370);
nand U5945 (N_5945,N_3146,N_4622);
or U5946 (N_5946,N_4734,N_4150);
and U5947 (N_5947,N_3972,N_2868);
and U5948 (N_5948,N_2519,N_4064);
nand U5949 (N_5949,N_3623,N_4818);
or U5950 (N_5950,N_3835,N_3113);
or U5951 (N_5951,N_3567,N_3180);
and U5952 (N_5952,N_3415,N_3041);
nor U5953 (N_5953,N_4579,N_2503);
nand U5954 (N_5954,N_2941,N_4199);
nand U5955 (N_5955,N_3499,N_4868);
nand U5956 (N_5956,N_3531,N_3785);
nor U5957 (N_5957,N_2906,N_2935);
nor U5958 (N_5958,N_3419,N_3064);
nand U5959 (N_5959,N_4859,N_3996);
nand U5960 (N_5960,N_4507,N_4332);
and U5961 (N_5961,N_3660,N_3952);
nand U5962 (N_5962,N_3310,N_2926);
nor U5963 (N_5963,N_4160,N_3229);
nand U5964 (N_5964,N_4037,N_4743);
nor U5965 (N_5965,N_3085,N_3572);
and U5966 (N_5966,N_2706,N_2966);
or U5967 (N_5967,N_3194,N_3965);
nand U5968 (N_5968,N_3226,N_3775);
or U5969 (N_5969,N_4942,N_3900);
and U5970 (N_5970,N_2875,N_4380);
xnor U5971 (N_5971,N_3479,N_3277);
nand U5972 (N_5972,N_3483,N_3281);
or U5973 (N_5973,N_4100,N_3353);
or U5974 (N_5974,N_3447,N_3839);
nand U5975 (N_5975,N_2958,N_3424);
nand U5976 (N_5976,N_3289,N_3807);
and U5977 (N_5977,N_4133,N_4817);
or U5978 (N_5978,N_4890,N_4426);
and U5979 (N_5979,N_2769,N_4189);
and U5980 (N_5980,N_4615,N_3593);
nand U5981 (N_5981,N_4982,N_4386);
nand U5982 (N_5982,N_4042,N_3546);
nor U5983 (N_5983,N_4625,N_4790);
nor U5984 (N_5984,N_4962,N_2567);
or U5985 (N_5985,N_4940,N_4099);
or U5986 (N_5986,N_2913,N_4047);
nand U5987 (N_5987,N_3398,N_4523);
nand U5988 (N_5988,N_2929,N_3138);
and U5989 (N_5989,N_2655,N_2516);
or U5990 (N_5990,N_2933,N_4005);
or U5991 (N_5991,N_3267,N_4390);
nand U5992 (N_5992,N_3099,N_3790);
nor U5993 (N_5993,N_3746,N_4032);
nor U5994 (N_5994,N_4495,N_3181);
nor U5995 (N_5995,N_4612,N_4682);
or U5996 (N_5996,N_4157,N_4093);
nor U5997 (N_5997,N_3969,N_2863);
nand U5998 (N_5998,N_3707,N_3776);
nand U5999 (N_5999,N_3438,N_4321);
and U6000 (N_6000,N_2990,N_3885);
nor U6001 (N_6001,N_2808,N_3607);
nor U6002 (N_6002,N_4503,N_4865);
nand U6003 (N_6003,N_3027,N_3659);
nand U6004 (N_6004,N_2664,N_4753);
and U6005 (N_6005,N_4700,N_2500);
xnor U6006 (N_6006,N_2788,N_4784);
and U6007 (N_6007,N_3731,N_4082);
or U6008 (N_6008,N_3586,N_3811);
nor U6009 (N_6009,N_3057,N_3043);
nand U6010 (N_6010,N_2780,N_3863);
nand U6011 (N_6011,N_3021,N_3087);
and U6012 (N_6012,N_3874,N_3435);
nor U6013 (N_6013,N_3552,N_3902);
nand U6014 (N_6014,N_4909,N_4927);
nor U6015 (N_6015,N_4452,N_4483);
nand U6016 (N_6016,N_2725,N_3028);
nor U6017 (N_6017,N_3338,N_3841);
or U6018 (N_6018,N_4233,N_2822);
or U6019 (N_6019,N_3164,N_4884);
nand U6020 (N_6020,N_3205,N_3069);
nand U6021 (N_6021,N_2996,N_4995);
nor U6022 (N_6022,N_4419,N_3951);
nor U6023 (N_6023,N_2770,N_3474);
and U6024 (N_6024,N_2981,N_4555);
nor U6025 (N_6025,N_3264,N_3039);
or U6026 (N_6026,N_3770,N_3122);
nor U6027 (N_6027,N_4356,N_2870);
nor U6028 (N_6028,N_4532,N_4237);
and U6029 (N_6029,N_4433,N_4531);
or U6030 (N_6030,N_3331,N_4097);
or U6031 (N_6031,N_4489,N_4014);
nand U6032 (N_6032,N_4294,N_3359);
or U6033 (N_6033,N_2782,N_4415);
nand U6034 (N_6034,N_3958,N_4429);
or U6035 (N_6035,N_2839,N_4305);
and U6036 (N_6036,N_4892,N_2779);
and U6037 (N_6037,N_3346,N_2570);
nor U6038 (N_6038,N_4038,N_4239);
nand U6039 (N_6039,N_3268,N_4136);
nor U6040 (N_6040,N_4980,N_3748);
or U6041 (N_6041,N_3988,N_2984);
and U6042 (N_6042,N_4720,N_3160);
nor U6043 (N_6043,N_2859,N_4732);
nor U6044 (N_6044,N_3843,N_2846);
nand U6045 (N_6045,N_3947,N_3278);
and U6046 (N_6046,N_4260,N_2621);
nor U6047 (N_6047,N_4344,N_4672);
nor U6048 (N_6048,N_3628,N_3780);
and U6049 (N_6049,N_2902,N_4939);
or U6050 (N_6050,N_4151,N_3383);
nor U6051 (N_6051,N_3769,N_3753);
and U6052 (N_6052,N_3196,N_3759);
nor U6053 (N_6053,N_3077,N_2792);
nor U6054 (N_6054,N_4240,N_4293);
nor U6055 (N_6055,N_3723,N_3721);
nor U6056 (N_6056,N_2510,N_4319);
or U6057 (N_6057,N_2574,N_4050);
nor U6058 (N_6058,N_4646,N_4806);
and U6059 (N_6059,N_2623,N_4462);
nor U6060 (N_6060,N_3773,N_4683);
and U6061 (N_6061,N_4266,N_3326);
nor U6062 (N_6062,N_4932,N_2648);
nand U6063 (N_6063,N_4835,N_2643);
and U6064 (N_6064,N_3694,N_3178);
or U6065 (N_6065,N_3211,N_3786);
and U6066 (N_6066,N_4596,N_2617);
or U6067 (N_6067,N_3096,N_3935);
and U6068 (N_6068,N_3152,N_4798);
xnor U6069 (N_6069,N_4891,N_4238);
or U6070 (N_6070,N_3091,N_4670);
and U6071 (N_6071,N_3820,N_4025);
and U6072 (N_6072,N_4619,N_3366);
nor U6073 (N_6073,N_4691,N_4516);
or U6074 (N_6074,N_3799,N_3186);
or U6075 (N_6075,N_4231,N_2794);
or U6076 (N_6076,N_3689,N_4759);
or U6077 (N_6077,N_2993,N_2829);
or U6078 (N_6078,N_3484,N_3854);
nand U6079 (N_6079,N_2708,N_4879);
or U6080 (N_6080,N_3849,N_3397);
nand U6081 (N_6081,N_2847,N_3755);
and U6082 (N_6082,N_4598,N_4013);
nor U6083 (N_6083,N_4520,N_2541);
and U6084 (N_6084,N_2629,N_3222);
nand U6085 (N_6085,N_3255,N_2658);
or U6086 (N_6086,N_4087,N_3365);
and U6087 (N_6087,N_3105,N_2815);
nor U6088 (N_6088,N_2894,N_4168);
xor U6089 (N_6089,N_2709,N_2749);
or U6090 (N_6090,N_2522,N_4369);
or U6091 (N_6091,N_4847,N_4834);
or U6092 (N_6092,N_4404,N_4926);
nor U6093 (N_6093,N_3598,N_4300);
nor U6094 (N_6094,N_4387,N_3321);
nor U6095 (N_6095,N_3446,N_4533);
or U6096 (N_6096,N_3818,N_4107);
nor U6097 (N_6097,N_2758,N_2561);
nand U6098 (N_6098,N_4428,N_2927);
and U6099 (N_6099,N_3867,N_2581);
nor U6100 (N_6100,N_4575,N_4864);
and U6101 (N_6101,N_3823,N_3352);
nor U6102 (N_6102,N_3231,N_4039);
or U6103 (N_6103,N_4654,N_3282);
nand U6104 (N_6104,N_4956,N_3042);
nor U6105 (N_6105,N_4972,N_4987);
and U6106 (N_6106,N_4276,N_4316);
nand U6107 (N_6107,N_3514,N_4310);
and U6108 (N_6108,N_4758,N_4235);
nand U6109 (N_6109,N_4915,N_3743);
or U6110 (N_6110,N_4173,N_4296);
and U6111 (N_6111,N_4154,N_3685);
and U6112 (N_6112,N_2702,N_2989);
or U6113 (N_6113,N_2905,N_3520);
nand U6114 (N_6114,N_4521,N_2784);
nand U6115 (N_6115,N_4323,N_3292);
or U6116 (N_6116,N_4869,N_4839);
nor U6117 (N_6117,N_4434,N_3118);
nand U6118 (N_6118,N_3631,N_3170);
and U6119 (N_6119,N_2835,N_2657);
nand U6120 (N_6120,N_3942,N_4476);
nor U6121 (N_6121,N_2618,N_3016);
or U6122 (N_6122,N_4108,N_2653);
nand U6123 (N_6123,N_4308,N_2630);
and U6124 (N_6124,N_4692,N_3589);
or U6125 (N_6125,N_4137,N_4735);
or U6126 (N_6126,N_4114,N_3416);
nand U6127 (N_6127,N_4971,N_3698);
and U6128 (N_6128,N_4851,N_3260);
nor U6129 (N_6129,N_4436,N_4480);
and U6130 (N_6130,N_3963,N_2798);
or U6131 (N_6131,N_3473,N_3168);
nand U6132 (N_6132,N_4561,N_4446);
nor U6133 (N_6133,N_4012,N_4420);
nand U6134 (N_6134,N_3311,N_2967);
nand U6135 (N_6135,N_3378,N_4824);
or U6136 (N_6136,N_2741,N_3471);
nor U6137 (N_6137,N_3547,N_4031);
nor U6138 (N_6138,N_4142,N_4079);
and U6139 (N_6139,N_4830,N_4049);
nor U6140 (N_6140,N_4177,N_4195);
or U6141 (N_6141,N_4614,N_4500);
nand U6142 (N_6142,N_4912,N_4128);
nor U6143 (N_6143,N_3006,N_3020);
and U6144 (N_6144,N_3228,N_3049);
or U6145 (N_6145,N_3684,N_2944);
or U6146 (N_6146,N_4484,N_3141);
or U6147 (N_6147,N_2544,N_3913);
and U6148 (N_6148,N_2991,N_3560);
and U6149 (N_6149,N_2564,N_3465);
or U6150 (N_6150,N_3781,N_4392);
nand U6151 (N_6151,N_2959,N_4350);
nor U6152 (N_6152,N_3342,N_3738);
nor U6153 (N_6153,N_4736,N_2732);
or U6154 (N_6154,N_4905,N_3887);
nand U6155 (N_6155,N_4706,N_3638);
nor U6156 (N_6156,N_3744,N_3789);
nand U6157 (N_6157,N_3129,N_4708);
or U6158 (N_6158,N_3930,N_2954);
and U6159 (N_6159,N_3833,N_2982);
nor U6160 (N_6160,N_3654,N_2917);
or U6161 (N_6161,N_4270,N_2707);
nor U6162 (N_6162,N_4815,N_4986);
nor U6163 (N_6163,N_3136,N_3602);
and U6164 (N_6164,N_4478,N_4639);
and U6165 (N_6165,N_3149,N_4594);
or U6166 (N_6166,N_3055,N_3071);
or U6167 (N_6167,N_2975,N_4973);
nand U6168 (N_6168,N_3033,N_2923);
or U6169 (N_6169,N_3643,N_3558);
nand U6170 (N_6170,N_3314,N_3971);
nor U6171 (N_6171,N_4600,N_3636);
nor U6172 (N_6172,N_4552,N_3929);
nand U6173 (N_6173,N_4519,N_4243);
nand U6174 (N_6174,N_2763,N_4286);
nor U6175 (N_6175,N_3600,N_4501);
nor U6176 (N_6176,N_2992,N_3075);
nor U6177 (N_6177,N_4174,N_3778);
or U6178 (N_6178,N_3097,N_3509);
or U6179 (N_6179,N_3742,N_4786);
nand U6180 (N_6180,N_3418,N_4116);
nand U6181 (N_6181,N_3974,N_3313);
nand U6182 (N_6182,N_4148,N_4606);
or U6183 (N_6183,N_3150,N_4340);
or U6184 (N_6184,N_3812,N_3038);
nand U6185 (N_6185,N_3766,N_4411);
nand U6186 (N_6186,N_4383,N_3290);
nor U6187 (N_6187,N_3981,N_4086);
nand U6188 (N_6188,N_2768,N_3851);
nand U6189 (N_6189,N_3764,N_3903);
nor U6190 (N_6190,N_3307,N_2698);
nor U6191 (N_6191,N_3491,N_3056);
and U6192 (N_6192,N_4403,N_3993);
and U6193 (N_6193,N_3034,N_3489);
nor U6194 (N_6194,N_4287,N_3355);
and U6195 (N_6195,N_3686,N_4312);
nand U6196 (N_6196,N_2556,N_4111);
nand U6197 (N_6197,N_4242,N_3661);
and U6198 (N_6198,N_3858,N_3275);
or U6199 (N_6199,N_3982,N_4804);
nor U6200 (N_6200,N_3017,N_2598);
or U6201 (N_6201,N_3195,N_4379);
nor U6202 (N_6202,N_4678,N_2599);
nand U6203 (N_6203,N_4105,N_2983);
or U6204 (N_6204,N_2672,N_3052);
and U6205 (N_6205,N_3626,N_2685);
nand U6206 (N_6206,N_2646,N_3432);
nor U6207 (N_6207,N_4664,N_3722);
nand U6208 (N_6208,N_3941,N_4629);
and U6209 (N_6209,N_2791,N_4842);
and U6210 (N_6210,N_3002,N_3595);
nand U6211 (N_6211,N_2985,N_2869);
nand U6212 (N_6212,N_2802,N_2817);
nor U6213 (N_6213,N_2546,N_3980);
and U6214 (N_6214,N_3238,N_4498);
or U6215 (N_6215,N_2533,N_3437);
nand U6216 (N_6216,N_4601,N_4773);
or U6217 (N_6217,N_4502,N_4302);
nor U6218 (N_6218,N_3209,N_3088);
or U6219 (N_6219,N_3828,N_3037);
nand U6220 (N_6220,N_2512,N_2916);
and U6221 (N_6221,N_4584,N_3018);
or U6222 (N_6222,N_4262,N_3079);
nor U6223 (N_6223,N_2800,N_3374);
nor U6224 (N_6224,N_3130,N_3225);
and U6225 (N_6225,N_3239,N_3931);
and U6226 (N_6226,N_2678,N_3529);
nand U6227 (N_6227,N_3976,N_4609);
and U6228 (N_6228,N_2673,N_4071);
and U6229 (N_6229,N_4091,N_3895);
and U6230 (N_6230,N_4083,N_3637);
nand U6231 (N_6231,N_4838,N_3089);
and U6232 (N_6232,N_2909,N_4617);
and U6233 (N_6233,N_2627,N_4541);
and U6234 (N_6234,N_3237,N_2806);
nand U6235 (N_6235,N_2550,N_2559);
nand U6236 (N_6236,N_2801,N_4525);
xnor U6237 (N_6237,N_4754,N_4763);
or U6238 (N_6238,N_4346,N_4548);
nor U6239 (N_6239,N_3601,N_2534);
and U6240 (N_6240,N_4983,N_3745);
nor U6241 (N_6241,N_3051,N_3580);
nand U6242 (N_6242,N_2595,N_2718);
nor U6243 (N_6243,N_3889,N_2760);
nand U6244 (N_6244,N_4805,N_3382);
nand U6245 (N_6245,N_3036,N_4698);
nor U6246 (N_6246,N_3213,N_4330);
xor U6247 (N_6247,N_2842,N_2888);
or U6248 (N_6248,N_2622,N_2587);
nand U6249 (N_6249,N_4475,N_3137);
and U6250 (N_6250,N_4850,N_3502);
or U6251 (N_6251,N_3015,N_4298);
or U6252 (N_6252,N_4539,N_3109);
or U6253 (N_6253,N_3774,N_2889);
nand U6254 (N_6254,N_2584,N_4096);
and U6255 (N_6255,N_4797,N_4757);
or U6256 (N_6256,N_4592,N_4332);
nor U6257 (N_6257,N_3899,N_4508);
nor U6258 (N_6258,N_3855,N_3022);
nand U6259 (N_6259,N_4722,N_3774);
nor U6260 (N_6260,N_2962,N_3992);
nor U6261 (N_6261,N_4720,N_2847);
nand U6262 (N_6262,N_2592,N_4218);
nand U6263 (N_6263,N_3589,N_2722);
nand U6264 (N_6264,N_3102,N_3059);
and U6265 (N_6265,N_4854,N_3981);
and U6266 (N_6266,N_4554,N_4516);
or U6267 (N_6267,N_4375,N_4840);
and U6268 (N_6268,N_2755,N_3654);
and U6269 (N_6269,N_4746,N_2670);
nor U6270 (N_6270,N_3845,N_2599);
and U6271 (N_6271,N_3617,N_3321);
nand U6272 (N_6272,N_4303,N_2719);
nor U6273 (N_6273,N_3447,N_3931);
and U6274 (N_6274,N_3776,N_3119);
nand U6275 (N_6275,N_3469,N_4974);
nand U6276 (N_6276,N_2966,N_4178);
or U6277 (N_6277,N_3435,N_4123);
nor U6278 (N_6278,N_2825,N_4226);
nand U6279 (N_6279,N_3816,N_3594);
nand U6280 (N_6280,N_4208,N_3726);
or U6281 (N_6281,N_4433,N_3476);
and U6282 (N_6282,N_4300,N_4778);
nor U6283 (N_6283,N_4718,N_2689);
or U6284 (N_6284,N_4535,N_3886);
nand U6285 (N_6285,N_4759,N_2832);
nand U6286 (N_6286,N_3706,N_4163);
or U6287 (N_6287,N_4323,N_3969);
or U6288 (N_6288,N_4710,N_2525);
or U6289 (N_6289,N_3164,N_3602);
nor U6290 (N_6290,N_4511,N_3871);
nand U6291 (N_6291,N_3420,N_4822);
nand U6292 (N_6292,N_2824,N_4032);
and U6293 (N_6293,N_2597,N_4751);
nor U6294 (N_6294,N_4866,N_2924);
or U6295 (N_6295,N_3932,N_2513);
nor U6296 (N_6296,N_3349,N_2805);
or U6297 (N_6297,N_2920,N_2654);
or U6298 (N_6298,N_2690,N_2918);
and U6299 (N_6299,N_4504,N_3684);
nor U6300 (N_6300,N_2661,N_3637);
nand U6301 (N_6301,N_3736,N_4099);
nor U6302 (N_6302,N_3235,N_2697);
nand U6303 (N_6303,N_4916,N_2504);
and U6304 (N_6304,N_3512,N_2606);
and U6305 (N_6305,N_4822,N_3746);
nor U6306 (N_6306,N_4455,N_3045);
nor U6307 (N_6307,N_2527,N_4073);
or U6308 (N_6308,N_3470,N_4311);
nand U6309 (N_6309,N_4960,N_3728);
nor U6310 (N_6310,N_4337,N_3580);
or U6311 (N_6311,N_4333,N_3184);
and U6312 (N_6312,N_2597,N_3767);
nand U6313 (N_6313,N_3122,N_4731);
or U6314 (N_6314,N_3086,N_3639);
nand U6315 (N_6315,N_2586,N_3692);
nand U6316 (N_6316,N_3462,N_3461);
and U6317 (N_6317,N_4281,N_3174);
or U6318 (N_6318,N_4708,N_4105);
nand U6319 (N_6319,N_2562,N_4269);
nand U6320 (N_6320,N_4829,N_3728);
and U6321 (N_6321,N_4761,N_2721);
nand U6322 (N_6322,N_4159,N_4944);
nor U6323 (N_6323,N_4011,N_4080);
nand U6324 (N_6324,N_2841,N_3762);
and U6325 (N_6325,N_3698,N_3811);
and U6326 (N_6326,N_4912,N_4224);
nand U6327 (N_6327,N_3682,N_3097);
nor U6328 (N_6328,N_3169,N_4429);
and U6329 (N_6329,N_2747,N_2607);
nand U6330 (N_6330,N_4094,N_3991);
or U6331 (N_6331,N_2847,N_2787);
nor U6332 (N_6332,N_4663,N_3850);
and U6333 (N_6333,N_3058,N_4963);
nor U6334 (N_6334,N_3399,N_4809);
nor U6335 (N_6335,N_4811,N_4531);
nand U6336 (N_6336,N_3532,N_4887);
nor U6337 (N_6337,N_4555,N_3610);
or U6338 (N_6338,N_2546,N_4008);
nor U6339 (N_6339,N_4311,N_3472);
and U6340 (N_6340,N_3666,N_3707);
or U6341 (N_6341,N_2764,N_2862);
nor U6342 (N_6342,N_2833,N_2954);
or U6343 (N_6343,N_3959,N_4829);
nor U6344 (N_6344,N_3617,N_4629);
and U6345 (N_6345,N_2667,N_4320);
or U6346 (N_6346,N_3193,N_3286);
nor U6347 (N_6347,N_4746,N_3363);
or U6348 (N_6348,N_3395,N_2929);
nand U6349 (N_6349,N_3026,N_3824);
nand U6350 (N_6350,N_4698,N_4327);
or U6351 (N_6351,N_3432,N_2930);
and U6352 (N_6352,N_4106,N_3962);
or U6353 (N_6353,N_4777,N_3431);
or U6354 (N_6354,N_4021,N_4777);
nand U6355 (N_6355,N_2580,N_2598);
nor U6356 (N_6356,N_3854,N_2988);
nor U6357 (N_6357,N_2749,N_3998);
nand U6358 (N_6358,N_4963,N_3278);
or U6359 (N_6359,N_3872,N_3279);
or U6360 (N_6360,N_4100,N_4059);
nor U6361 (N_6361,N_3700,N_4074);
or U6362 (N_6362,N_4325,N_3480);
or U6363 (N_6363,N_4773,N_4907);
nor U6364 (N_6364,N_3277,N_3872);
nor U6365 (N_6365,N_2658,N_3099);
or U6366 (N_6366,N_2920,N_3470);
and U6367 (N_6367,N_3057,N_3284);
nor U6368 (N_6368,N_4957,N_4159);
nor U6369 (N_6369,N_2611,N_4887);
nand U6370 (N_6370,N_2775,N_3568);
and U6371 (N_6371,N_4641,N_3642);
and U6372 (N_6372,N_2627,N_4743);
or U6373 (N_6373,N_4154,N_3139);
or U6374 (N_6374,N_4763,N_4303);
and U6375 (N_6375,N_4651,N_3319);
nand U6376 (N_6376,N_3549,N_3563);
or U6377 (N_6377,N_3474,N_4642);
and U6378 (N_6378,N_4086,N_2742);
and U6379 (N_6379,N_3029,N_4874);
nand U6380 (N_6380,N_4645,N_4864);
nor U6381 (N_6381,N_3873,N_4361);
and U6382 (N_6382,N_4626,N_4230);
and U6383 (N_6383,N_3984,N_3410);
or U6384 (N_6384,N_4045,N_4455);
nor U6385 (N_6385,N_2835,N_3455);
nor U6386 (N_6386,N_3140,N_3397);
or U6387 (N_6387,N_4138,N_3025);
nand U6388 (N_6388,N_2545,N_2854);
and U6389 (N_6389,N_2532,N_4864);
or U6390 (N_6390,N_3667,N_2963);
or U6391 (N_6391,N_2534,N_4050);
nor U6392 (N_6392,N_3314,N_2773);
and U6393 (N_6393,N_4768,N_4424);
nand U6394 (N_6394,N_2700,N_3394);
nor U6395 (N_6395,N_4213,N_3789);
or U6396 (N_6396,N_2572,N_3133);
nor U6397 (N_6397,N_3983,N_2686);
and U6398 (N_6398,N_2763,N_3930);
and U6399 (N_6399,N_4468,N_3486);
or U6400 (N_6400,N_4454,N_3127);
or U6401 (N_6401,N_4798,N_2948);
nand U6402 (N_6402,N_4362,N_2623);
or U6403 (N_6403,N_3491,N_4964);
and U6404 (N_6404,N_3166,N_3356);
and U6405 (N_6405,N_3685,N_2934);
or U6406 (N_6406,N_4800,N_4444);
or U6407 (N_6407,N_3982,N_4880);
nand U6408 (N_6408,N_3744,N_4316);
and U6409 (N_6409,N_3252,N_2959);
nand U6410 (N_6410,N_4275,N_4704);
nand U6411 (N_6411,N_3106,N_3466);
nor U6412 (N_6412,N_4291,N_3358);
and U6413 (N_6413,N_4153,N_3222);
nor U6414 (N_6414,N_4768,N_2869);
nor U6415 (N_6415,N_4450,N_2744);
nand U6416 (N_6416,N_4974,N_3173);
nor U6417 (N_6417,N_3159,N_4168);
and U6418 (N_6418,N_4097,N_4765);
or U6419 (N_6419,N_2627,N_3614);
nor U6420 (N_6420,N_3207,N_3902);
nand U6421 (N_6421,N_3037,N_4946);
or U6422 (N_6422,N_3536,N_3746);
and U6423 (N_6423,N_3223,N_3392);
nor U6424 (N_6424,N_4128,N_3030);
nand U6425 (N_6425,N_2957,N_4972);
and U6426 (N_6426,N_4679,N_3004);
and U6427 (N_6427,N_3800,N_4838);
and U6428 (N_6428,N_3558,N_4661);
and U6429 (N_6429,N_3266,N_3881);
and U6430 (N_6430,N_4251,N_4439);
or U6431 (N_6431,N_3486,N_4002);
nor U6432 (N_6432,N_3711,N_3323);
nor U6433 (N_6433,N_4271,N_2672);
or U6434 (N_6434,N_4074,N_2998);
and U6435 (N_6435,N_3469,N_3556);
nor U6436 (N_6436,N_3289,N_2688);
nor U6437 (N_6437,N_4912,N_3847);
nor U6438 (N_6438,N_4409,N_4446);
or U6439 (N_6439,N_3854,N_3714);
and U6440 (N_6440,N_4282,N_3147);
and U6441 (N_6441,N_4225,N_3553);
and U6442 (N_6442,N_4718,N_2643);
and U6443 (N_6443,N_3561,N_3958);
nor U6444 (N_6444,N_2532,N_3003);
and U6445 (N_6445,N_3766,N_2606);
nand U6446 (N_6446,N_3170,N_3835);
xor U6447 (N_6447,N_3019,N_3665);
and U6448 (N_6448,N_4011,N_4320);
or U6449 (N_6449,N_4230,N_3024);
nor U6450 (N_6450,N_4710,N_3981);
nand U6451 (N_6451,N_3338,N_4872);
or U6452 (N_6452,N_4951,N_4643);
nor U6453 (N_6453,N_2996,N_4051);
or U6454 (N_6454,N_4394,N_3851);
and U6455 (N_6455,N_2922,N_3508);
or U6456 (N_6456,N_4449,N_3832);
nor U6457 (N_6457,N_3015,N_3122);
or U6458 (N_6458,N_2605,N_2939);
and U6459 (N_6459,N_2845,N_3030);
and U6460 (N_6460,N_3696,N_3656);
nand U6461 (N_6461,N_3830,N_3995);
nor U6462 (N_6462,N_4955,N_4980);
nor U6463 (N_6463,N_3009,N_4585);
and U6464 (N_6464,N_2656,N_3328);
or U6465 (N_6465,N_2578,N_3711);
and U6466 (N_6466,N_2569,N_4471);
and U6467 (N_6467,N_4022,N_2980);
and U6468 (N_6468,N_2847,N_4649);
and U6469 (N_6469,N_3405,N_3421);
or U6470 (N_6470,N_4829,N_3827);
or U6471 (N_6471,N_4983,N_2821);
nand U6472 (N_6472,N_4589,N_3378);
and U6473 (N_6473,N_3549,N_3849);
nand U6474 (N_6474,N_4124,N_2990);
nor U6475 (N_6475,N_3366,N_4371);
and U6476 (N_6476,N_3175,N_2792);
nor U6477 (N_6477,N_4988,N_3116);
nand U6478 (N_6478,N_4236,N_4525);
nand U6479 (N_6479,N_3524,N_4155);
nand U6480 (N_6480,N_3565,N_3716);
xnor U6481 (N_6481,N_3818,N_4140);
and U6482 (N_6482,N_3290,N_2869);
nand U6483 (N_6483,N_4339,N_3980);
nor U6484 (N_6484,N_4963,N_3527);
nor U6485 (N_6485,N_4091,N_3526);
xor U6486 (N_6486,N_3044,N_3966);
and U6487 (N_6487,N_3761,N_4351);
and U6488 (N_6488,N_4600,N_4870);
nor U6489 (N_6489,N_3054,N_3833);
and U6490 (N_6490,N_4626,N_3165);
or U6491 (N_6491,N_4267,N_4922);
and U6492 (N_6492,N_3791,N_3082);
nor U6493 (N_6493,N_3587,N_2768);
and U6494 (N_6494,N_3921,N_3188);
nand U6495 (N_6495,N_2744,N_3285);
nand U6496 (N_6496,N_3290,N_4114);
or U6497 (N_6497,N_2827,N_2600);
and U6498 (N_6498,N_4484,N_4781);
or U6499 (N_6499,N_4908,N_4907);
or U6500 (N_6500,N_2644,N_3338);
nor U6501 (N_6501,N_4520,N_3863);
or U6502 (N_6502,N_3283,N_3436);
and U6503 (N_6503,N_4625,N_4577);
or U6504 (N_6504,N_3746,N_4133);
nand U6505 (N_6505,N_3503,N_4454);
nor U6506 (N_6506,N_4018,N_3171);
or U6507 (N_6507,N_4348,N_4761);
nand U6508 (N_6508,N_4377,N_3500);
nand U6509 (N_6509,N_4054,N_2997);
nor U6510 (N_6510,N_4732,N_3456);
nand U6511 (N_6511,N_4318,N_4677);
and U6512 (N_6512,N_2981,N_3488);
nor U6513 (N_6513,N_4069,N_4765);
nand U6514 (N_6514,N_2838,N_4931);
or U6515 (N_6515,N_4984,N_4875);
and U6516 (N_6516,N_2521,N_3645);
or U6517 (N_6517,N_3249,N_3648);
and U6518 (N_6518,N_2735,N_2967);
and U6519 (N_6519,N_2864,N_3245);
and U6520 (N_6520,N_3822,N_3313);
nor U6521 (N_6521,N_4531,N_3953);
or U6522 (N_6522,N_2843,N_3719);
nor U6523 (N_6523,N_4108,N_3153);
nand U6524 (N_6524,N_4169,N_2805);
or U6525 (N_6525,N_3394,N_3342);
and U6526 (N_6526,N_4114,N_3444);
nor U6527 (N_6527,N_4155,N_4964);
nor U6528 (N_6528,N_2806,N_4295);
nor U6529 (N_6529,N_4221,N_3853);
or U6530 (N_6530,N_4797,N_4182);
and U6531 (N_6531,N_3098,N_3097);
nor U6532 (N_6532,N_4667,N_3274);
nor U6533 (N_6533,N_4713,N_4614);
and U6534 (N_6534,N_3157,N_3685);
nor U6535 (N_6535,N_4224,N_2938);
and U6536 (N_6536,N_4949,N_4956);
nor U6537 (N_6537,N_4700,N_4654);
or U6538 (N_6538,N_4851,N_3357);
or U6539 (N_6539,N_4970,N_4308);
or U6540 (N_6540,N_2873,N_4713);
nor U6541 (N_6541,N_4882,N_4398);
nor U6542 (N_6542,N_4471,N_3803);
nand U6543 (N_6543,N_2710,N_3292);
nand U6544 (N_6544,N_3370,N_4842);
or U6545 (N_6545,N_4040,N_3458);
nor U6546 (N_6546,N_4593,N_4082);
and U6547 (N_6547,N_2533,N_4639);
nor U6548 (N_6548,N_4285,N_3206);
nor U6549 (N_6549,N_3935,N_3417);
and U6550 (N_6550,N_4764,N_3440);
and U6551 (N_6551,N_4156,N_4244);
nand U6552 (N_6552,N_4899,N_4348);
and U6553 (N_6553,N_4086,N_3242);
or U6554 (N_6554,N_3952,N_4499);
or U6555 (N_6555,N_4629,N_4903);
or U6556 (N_6556,N_4085,N_3974);
nor U6557 (N_6557,N_3952,N_2744);
nor U6558 (N_6558,N_3355,N_2894);
and U6559 (N_6559,N_3907,N_2606);
nor U6560 (N_6560,N_4438,N_4375);
and U6561 (N_6561,N_4361,N_3524);
or U6562 (N_6562,N_4583,N_3988);
nand U6563 (N_6563,N_3543,N_3938);
or U6564 (N_6564,N_3204,N_2976);
nor U6565 (N_6565,N_4250,N_4560);
nand U6566 (N_6566,N_3134,N_4770);
nor U6567 (N_6567,N_4375,N_3343);
nor U6568 (N_6568,N_4982,N_4646);
nor U6569 (N_6569,N_3836,N_2588);
nand U6570 (N_6570,N_3338,N_4179);
nor U6571 (N_6571,N_3878,N_3250);
nor U6572 (N_6572,N_3102,N_4316);
nor U6573 (N_6573,N_3748,N_2824);
nand U6574 (N_6574,N_4850,N_4335);
or U6575 (N_6575,N_3515,N_3237);
and U6576 (N_6576,N_4165,N_4336);
nand U6577 (N_6577,N_4887,N_2910);
nand U6578 (N_6578,N_4645,N_2968);
nand U6579 (N_6579,N_4663,N_2589);
or U6580 (N_6580,N_2826,N_3679);
nor U6581 (N_6581,N_4121,N_3090);
nand U6582 (N_6582,N_3302,N_3005);
and U6583 (N_6583,N_4097,N_3093);
nor U6584 (N_6584,N_3117,N_3594);
and U6585 (N_6585,N_3487,N_4927);
or U6586 (N_6586,N_4509,N_3024);
nor U6587 (N_6587,N_4014,N_4916);
nand U6588 (N_6588,N_2814,N_3877);
and U6589 (N_6589,N_4784,N_4775);
and U6590 (N_6590,N_4241,N_4107);
or U6591 (N_6591,N_3296,N_2995);
nand U6592 (N_6592,N_3488,N_4333);
nand U6593 (N_6593,N_3628,N_3409);
or U6594 (N_6594,N_2710,N_4230);
nor U6595 (N_6595,N_4385,N_3866);
nor U6596 (N_6596,N_3202,N_4894);
and U6597 (N_6597,N_3867,N_2677);
nor U6598 (N_6598,N_3792,N_3802);
nor U6599 (N_6599,N_4926,N_4326);
or U6600 (N_6600,N_2839,N_2584);
or U6601 (N_6601,N_3613,N_4929);
and U6602 (N_6602,N_2781,N_2993);
or U6603 (N_6603,N_4313,N_4847);
and U6604 (N_6604,N_2854,N_2703);
and U6605 (N_6605,N_2505,N_3058);
nor U6606 (N_6606,N_2909,N_3375);
and U6607 (N_6607,N_3873,N_4320);
nand U6608 (N_6608,N_3804,N_3133);
or U6609 (N_6609,N_4427,N_2579);
and U6610 (N_6610,N_4986,N_3211);
and U6611 (N_6611,N_4230,N_3217);
or U6612 (N_6612,N_2671,N_3582);
or U6613 (N_6613,N_2658,N_4825);
and U6614 (N_6614,N_2588,N_3790);
nor U6615 (N_6615,N_4771,N_2864);
nand U6616 (N_6616,N_3844,N_3487);
or U6617 (N_6617,N_4269,N_4089);
or U6618 (N_6618,N_4257,N_3652);
nor U6619 (N_6619,N_2518,N_3296);
or U6620 (N_6620,N_4326,N_4325);
nor U6621 (N_6621,N_2929,N_4377);
nor U6622 (N_6622,N_2655,N_2583);
nor U6623 (N_6623,N_3857,N_2595);
nor U6624 (N_6624,N_4131,N_3695);
and U6625 (N_6625,N_4626,N_3766);
nand U6626 (N_6626,N_4306,N_4204);
or U6627 (N_6627,N_4947,N_2816);
nor U6628 (N_6628,N_3750,N_4743);
or U6629 (N_6629,N_4023,N_3656);
nand U6630 (N_6630,N_3889,N_2853);
or U6631 (N_6631,N_3874,N_3967);
or U6632 (N_6632,N_2818,N_3546);
or U6633 (N_6633,N_4096,N_3998);
and U6634 (N_6634,N_2870,N_4630);
and U6635 (N_6635,N_3975,N_4470);
or U6636 (N_6636,N_3029,N_2798);
nand U6637 (N_6637,N_3759,N_3600);
or U6638 (N_6638,N_4877,N_4798);
nand U6639 (N_6639,N_4763,N_2676);
or U6640 (N_6640,N_4019,N_3846);
and U6641 (N_6641,N_4635,N_3308);
nor U6642 (N_6642,N_3301,N_3240);
nand U6643 (N_6643,N_3177,N_3604);
and U6644 (N_6644,N_3824,N_4335);
nor U6645 (N_6645,N_4494,N_4889);
and U6646 (N_6646,N_2724,N_4804);
nor U6647 (N_6647,N_3516,N_4500);
and U6648 (N_6648,N_3051,N_2557);
nand U6649 (N_6649,N_3120,N_3131);
or U6650 (N_6650,N_3165,N_3351);
and U6651 (N_6651,N_2936,N_2814);
and U6652 (N_6652,N_3340,N_3473);
nor U6653 (N_6653,N_4586,N_4944);
and U6654 (N_6654,N_2561,N_2541);
xnor U6655 (N_6655,N_4159,N_3686);
nor U6656 (N_6656,N_2669,N_2721);
nand U6657 (N_6657,N_4361,N_3364);
nand U6658 (N_6658,N_3958,N_2832);
nand U6659 (N_6659,N_3736,N_3761);
or U6660 (N_6660,N_4434,N_4345);
nor U6661 (N_6661,N_3661,N_3978);
nand U6662 (N_6662,N_2664,N_2578);
nor U6663 (N_6663,N_3301,N_3095);
nand U6664 (N_6664,N_4402,N_2596);
nand U6665 (N_6665,N_4140,N_3007);
or U6666 (N_6666,N_3028,N_3202);
nand U6667 (N_6667,N_3382,N_3279);
and U6668 (N_6668,N_3214,N_3540);
xnor U6669 (N_6669,N_2882,N_3738);
nand U6670 (N_6670,N_3041,N_3629);
or U6671 (N_6671,N_3588,N_3108);
nand U6672 (N_6672,N_4210,N_3672);
and U6673 (N_6673,N_4986,N_3406);
or U6674 (N_6674,N_3416,N_3154);
and U6675 (N_6675,N_3124,N_4028);
and U6676 (N_6676,N_3287,N_3153);
nor U6677 (N_6677,N_3795,N_3000);
nand U6678 (N_6678,N_3325,N_4468);
or U6679 (N_6679,N_4154,N_4906);
and U6680 (N_6680,N_3144,N_4136);
nand U6681 (N_6681,N_4253,N_4392);
or U6682 (N_6682,N_4795,N_2709);
nand U6683 (N_6683,N_4826,N_2969);
or U6684 (N_6684,N_2624,N_3260);
and U6685 (N_6685,N_3158,N_4454);
and U6686 (N_6686,N_2656,N_4778);
and U6687 (N_6687,N_3295,N_4760);
nor U6688 (N_6688,N_2536,N_3670);
nor U6689 (N_6689,N_3655,N_4675);
nor U6690 (N_6690,N_2645,N_4052);
nand U6691 (N_6691,N_3505,N_3802);
or U6692 (N_6692,N_4911,N_4279);
nand U6693 (N_6693,N_3463,N_4111);
and U6694 (N_6694,N_3104,N_3501);
nor U6695 (N_6695,N_3040,N_3166);
or U6696 (N_6696,N_4183,N_3261);
or U6697 (N_6697,N_3883,N_3230);
nor U6698 (N_6698,N_4593,N_4582);
and U6699 (N_6699,N_3584,N_4481);
nor U6700 (N_6700,N_2610,N_3641);
and U6701 (N_6701,N_4264,N_4374);
nand U6702 (N_6702,N_2995,N_3740);
nor U6703 (N_6703,N_3405,N_4584);
nand U6704 (N_6704,N_3657,N_4981);
and U6705 (N_6705,N_3569,N_4987);
nor U6706 (N_6706,N_3355,N_4965);
nor U6707 (N_6707,N_2878,N_3264);
and U6708 (N_6708,N_3999,N_4753);
and U6709 (N_6709,N_3589,N_4151);
or U6710 (N_6710,N_2711,N_2860);
and U6711 (N_6711,N_4359,N_4188);
or U6712 (N_6712,N_4317,N_4840);
or U6713 (N_6713,N_4800,N_4270);
nand U6714 (N_6714,N_3393,N_2787);
nor U6715 (N_6715,N_3324,N_4100);
or U6716 (N_6716,N_4975,N_4023);
nand U6717 (N_6717,N_2706,N_3386);
or U6718 (N_6718,N_2601,N_3559);
nand U6719 (N_6719,N_3405,N_3331);
and U6720 (N_6720,N_4187,N_4536);
or U6721 (N_6721,N_2815,N_3405);
and U6722 (N_6722,N_3234,N_4175);
and U6723 (N_6723,N_4817,N_3592);
or U6724 (N_6724,N_3374,N_2805);
nand U6725 (N_6725,N_2844,N_3909);
nor U6726 (N_6726,N_2536,N_4138);
xnor U6727 (N_6727,N_3320,N_4054);
or U6728 (N_6728,N_3164,N_4294);
and U6729 (N_6729,N_4941,N_4503);
or U6730 (N_6730,N_4295,N_3574);
and U6731 (N_6731,N_3555,N_2925);
nor U6732 (N_6732,N_4054,N_3296);
nor U6733 (N_6733,N_3657,N_3928);
and U6734 (N_6734,N_3998,N_4985);
and U6735 (N_6735,N_4208,N_3697);
or U6736 (N_6736,N_3289,N_4198);
nor U6737 (N_6737,N_4507,N_3208);
nand U6738 (N_6738,N_3297,N_2860);
or U6739 (N_6739,N_3725,N_2695);
or U6740 (N_6740,N_2596,N_2692);
or U6741 (N_6741,N_4368,N_3593);
nor U6742 (N_6742,N_4516,N_4902);
and U6743 (N_6743,N_4973,N_4124);
and U6744 (N_6744,N_3895,N_2997);
nand U6745 (N_6745,N_4781,N_4022);
or U6746 (N_6746,N_2612,N_3889);
or U6747 (N_6747,N_4083,N_3997);
and U6748 (N_6748,N_3963,N_4308);
nor U6749 (N_6749,N_4250,N_4105);
nor U6750 (N_6750,N_3378,N_4058);
nor U6751 (N_6751,N_2529,N_3966);
and U6752 (N_6752,N_4592,N_3754);
or U6753 (N_6753,N_4836,N_3709);
xnor U6754 (N_6754,N_4844,N_3247);
nand U6755 (N_6755,N_3823,N_3242);
nor U6756 (N_6756,N_3864,N_4564);
nand U6757 (N_6757,N_3407,N_3608);
and U6758 (N_6758,N_4608,N_4239);
nand U6759 (N_6759,N_4746,N_4429);
and U6760 (N_6760,N_4189,N_2727);
and U6761 (N_6761,N_3186,N_2607);
or U6762 (N_6762,N_3979,N_4457);
xnor U6763 (N_6763,N_2618,N_4121);
nand U6764 (N_6764,N_4945,N_4009);
or U6765 (N_6765,N_3209,N_4874);
nor U6766 (N_6766,N_3967,N_2762);
nand U6767 (N_6767,N_4106,N_3878);
nor U6768 (N_6768,N_4507,N_3970);
or U6769 (N_6769,N_3542,N_2711);
and U6770 (N_6770,N_4422,N_4536);
and U6771 (N_6771,N_3957,N_2943);
nor U6772 (N_6772,N_4281,N_2832);
or U6773 (N_6773,N_4280,N_4752);
nor U6774 (N_6774,N_4729,N_4286);
and U6775 (N_6775,N_3117,N_2755);
or U6776 (N_6776,N_4534,N_3993);
or U6777 (N_6777,N_3720,N_3596);
nand U6778 (N_6778,N_2748,N_4018);
and U6779 (N_6779,N_2585,N_2594);
or U6780 (N_6780,N_3402,N_4974);
or U6781 (N_6781,N_2539,N_3811);
nand U6782 (N_6782,N_3588,N_2577);
nor U6783 (N_6783,N_3817,N_3318);
nor U6784 (N_6784,N_3835,N_3492);
or U6785 (N_6785,N_3743,N_3898);
xor U6786 (N_6786,N_4006,N_3360);
and U6787 (N_6787,N_2867,N_3022);
and U6788 (N_6788,N_4854,N_4405);
nor U6789 (N_6789,N_2947,N_3853);
nand U6790 (N_6790,N_4153,N_4736);
nand U6791 (N_6791,N_4201,N_3642);
and U6792 (N_6792,N_2612,N_3949);
nand U6793 (N_6793,N_3635,N_4773);
or U6794 (N_6794,N_4686,N_2591);
or U6795 (N_6795,N_3787,N_3538);
or U6796 (N_6796,N_4817,N_3164);
or U6797 (N_6797,N_4961,N_3826);
and U6798 (N_6798,N_3361,N_4781);
and U6799 (N_6799,N_4143,N_2721);
nor U6800 (N_6800,N_3639,N_4262);
and U6801 (N_6801,N_3406,N_4719);
nor U6802 (N_6802,N_3853,N_4090);
or U6803 (N_6803,N_3116,N_3405);
and U6804 (N_6804,N_4770,N_3580);
nor U6805 (N_6805,N_3121,N_3493);
nor U6806 (N_6806,N_2982,N_4600);
and U6807 (N_6807,N_4168,N_3048);
and U6808 (N_6808,N_4650,N_3781);
and U6809 (N_6809,N_4326,N_2872);
and U6810 (N_6810,N_4057,N_4226);
nand U6811 (N_6811,N_3739,N_4991);
nor U6812 (N_6812,N_4729,N_4888);
and U6813 (N_6813,N_4611,N_3484);
nor U6814 (N_6814,N_3731,N_4075);
and U6815 (N_6815,N_3673,N_3505);
or U6816 (N_6816,N_2915,N_4320);
nor U6817 (N_6817,N_4665,N_3540);
nor U6818 (N_6818,N_2968,N_3428);
or U6819 (N_6819,N_4208,N_2888);
nand U6820 (N_6820,N_3169,N_3739);
nand U6821 (N_6821,N_4867,N_4522);
and U6822 (N_6822,N_3547,N_3131);
nor U6823 (N_6823,N_4514,N_3598);
and U6824 (N_6824,N_3410,N_4768);
nor U6825 (N_6825,N_2536,N_3360);
or U6826 (N_6826,N_3755,N_4112);
nand U6827 (N_6827,N_3248,N_4646);
or U6828 (N_6828,N_2617,N_4546);
nor U6829 (N_6829,N_3879,N_3801);
nand U6830 (N_6830,N_3510,N_4803);
or U6831 (N_6831,N_2816,N_3769);
nor U6832 (N_6832,N_3684,N_4813);
and U6833 (N_6833,N_4897,N_3117);
or U6834 (N_6834,N_2840,N_4626);
nand U6835 (N_6835,N_2546,N_2764);
and U6836 (N_6836,N_2529,N_2638);
nor U6837 (N_6837,N_2677,N_3718);
nor U6838 (N_6838,N_3859,N_3927);
nand U6839 (N_6839,N_4368,N_4037);
or U6840 (N_6840,N_2939,N_2640);
or U6841 (N_6841,N_4184,N_3803);
nor U6842 (N_6842,N_2911,N_4685);
nor U6843 (N_6843,N_4438,N_3514);
nor U6844 (N_6844,N_2633,N_4508);
nand U6845 (N_6845,N_3240,N_2973);
or U6846 (N_6846,N_3139,N_3579);
nand U6847 (N_6847,N_2547,N_2928);
nand U6848 (N_6848,N_2713,N_4778);
nor U6849 (N_6849,N_4947,N_3229);
xnor U6850 (N_6850,N_3250,N_4116);
or U6851 (N_6851,N_2956,N_3159);
nand U6852 (N_6852,N_4197,N_4388);
nand U6853 (N_6853,N_4912,N_4635);
nand U6854 (N_6854,N_2682,N_3651);
or U6855 (N_6855,N_3728,N_2795);
nor U6856 (N_6856,N_2998,N_4697);
nor U6857 (N_6857,N_3371,N_3414);
nor U6858 (N_6858,N_4817,N_4057);
and U6859 (N_6859,N_4302,N_3586);
and U6860 (N_6860,N_3307,N_3248);
and U6861 (N_6861,N_3740,N_4517);
nor U6862 (N_6862,N_4836,N_2618);
or U6863 (N_6863,N_4726,N_3215);
and U6864 (N_6864,N_4934,N_2935);
or U6865 (N_6865,N_4611,N_4667);
and U6866 (N_6866,N_3931,N_2624);
nand U6867 (N_6867,N_3293,N_4886);
nand U6868 (N_6868,N_3512,N_3829);
or U6869 (N_6869,N_3199,N_4662);
nand U6870 (N_6870,N_3356,N_2782);
and U6871 (N_6871,N_2653,N_4315);
and U6872 (N_6872,N_2686,N_3987);
nor U6873 (N_6873,N_3914,N_2768);
nor U6874 (N_6874,N_2923,N_3710);
and U6875 (N_6875,N_3442,N_3650);
nor U6876 (N_6876,N_2593,N_3555);
nand U6877 (N_6877,N_4680,N_3309);
nand U6878 (N_6878,N_3179,N_4373);
and U6879 (N_6879,N_4342,N_4041);
xnor U6880 (N_6880,N_2627,N_3454);
and U6881 (N_6881,N_2642,N_4681);
or U6882 (N_6882,N_3552,N_3388);
and U6883 (N_6883,N_3271,N_2928);
and U6884 (N_6884,N_3693,N_4002);
and U6885 (N_6885,N_3546,N_2726);
nor U6886 (N_6886,N_2933,N_4220);
nor U6887 (N_6887,N_2904,N_4090);
and U6888 (N_6888,N_4012,N_2897);
nand U6889 (N_6889,N_4505,N_4414);
nor U6890 (N_6890,N_3903,N_3701);
or U6891 (N_6891,N_4285,N_3642);
nor U6892 (N_6892,N_4647,N_4561);
and U6893 (N_6893,N_3291,N_3203);
or U6894 (N_6894,N_4220,N_3316);
nor U6895 (N_6895,N_4099,N_2880);
or U6896 (N_6896,N_3017,N_2994);
or U6897 (N_6897,N_4249,N_4369);
nor U6898 (N_6898,N_4185,N_4770);
or U6899 (N_6899,N_3663,N_4221);
or U6900 (N_6900,N_3378,N_2637);
and U6901 (N_6901,N_3595,N_2749);
nor U6902 (N_6902,N_3545,N_3238);
nand U6903 (N_6903,N_4182,N_4360);
or U6904 (N_6904,N_4888,N_4429);
and U6905 (N_6905,N_3404,N_4678);
nand U6906 (N_6906,N_3768,N_2942);
nand U6907 (N_6907,N_3687,N_3953);
or U6908 (N_6908,N_3836,N_2863);
nor U6909 (N_6909,N_4590,N_3057);
and U6910 (N_6910,N_4870,N_3176);
nor U6911 (N_6911,N_4939,N_4964);
nand U6912 (N_6912,N_4603,N_2706);
or U6913 (N_6913,N_3500,N_2916);
nor U6914 (N_6914,N_2866,N_3728);
and U6915 (N_6915,N_2527,N_4502);
and U6916 (N_6916,N_3868,N_3856);
nand U6917 (N_6917,N_4087,N_2656);
and U6918 (N_6918,N_2631,N_2719);
or U6919 (N_6919,N_3074,N_4901);
nor U6920 (N_6920,N_3703,N_2789);
and U6921 (N_6921,N_3440,N_3888);
nor U6922 (N_6922,N_4889,N_2573);
and U6923 (N_6923,N_4673,N_4875);
nand U6924 (N_6924,N_2609,N_3715);
and U6925 (N_6925,N_2542,N_2660);
and U6926 (N_6926,N_3411,N_2672);
nand U6927 (N_6927,N_3166,N_4366);
and U6928 (N_6928,N_3559,N_3801);
and U6929 (N_6929,N_4535,N_2531);
nor U6930 (N_6930,N_3863,N_3748);
nand U6931 (N_6931,N_3753,N_3900);
nor U6932 (N_6932,N_4886,N_3252);
and U6933 (N_6933,N_3397,N_4612);
xnor U6934 (N_6934,N_4510,N_4294);
or U6935 (N_6935,N_3152,N_3788);
or U6936 (N_6936,N_2928,N_3531);
nand U6937 (N_6937,N_4280,N_3809);
nor U6938 (N_6938,N_4029,N_3121);
nor U6939 (N_6939,N_4602,N_2936);
or U6940 (N_6940,N_4915,N_4537);
or U6941 (N_6941,N_3640,N_4156);
and U6942 (N_6942,N_4316,N_4270);
nor U6943 (N_6943,N_4791,N_4294);
nor U6944 (N_6944,N_2620,N_4238);
nor U6945 (N_6945,N_3209,N_3293);
nand U6946 (N_6946,N_3252,N_4398);
or U6947 (N_6947,N_4103,N_4886);
nand U6948 (N_6948,N_3593,N_3808);
nand U6949 (N_6949,N_3890,N_4310);
nand U6950 (N_6950,N_4744,N_2502);
or U6951 (N_6951,N_4051,N_4125);
or U6952 (N_6952,N_3598,N_4214);
nand U6953 (N_6953,N_2717,N_4388);
and U6954 (N_6954,N_4480,N_3079);
or U6955 (N_6955,N_4821,N_4353);
nand U6956 (N_6956,N_2786,N_2712);
nor U6957 (N_6957,N_4682,N_3756);
and U6958 (N_6958,N_3928,N_4928);
nand U6959 (N_6959,N_2718,N_4884);
or U6960 (N_6960,N_3767,N_4920);
and U6961 (N_6961,N_4837,N_3859);
and U6962 (N_6962,N_2961,N_4060);
or U6963 (N_6963,N_3565,N_4549);
and U6964 (N_6964,N_4554,N_3426);
or U6965 (N_6965,N_3233,N_4546);
nand U6966 (N_6966,N_2660,N_4490);
nor U6967 (N_6967,N_2564,N_3213);
nand U6968 (N_6968,N_4287,N_4934);
and U6969 (N_6969,N_3529,N_3266);
nand U6970 (N_6970,N_4238,N_4074);
nand U6971 (N_6971,N_3299,N_4656);
and U6972 (N_6972,N_4051,N_4918);
or U6973 (N_6973,N_3711,N_2527);
nand U6974 (N_6974,N_4886,N_4377);
nand U6975 (N_6975,N_3639,N_3178);
and U6976 (N_6976,N_3213,N_3925);
and U6977 (N_6977,N_4825,N_4490);
or U6978 (N_6978,N_4997,N_4571);
and U6979 (N_6979,N_4499,N_4473);
nor U6980 (N_6980,N_2617,N_4451);
nand U6981 (N_6981,N_4405,N_4345);
nor U6982 (N_6982,N_2826,N_3782);
nor U6983 (N_6983,N_4244,N_2681);
or U6984 (N_6984,N_3442,N_3204);
and U6985 (N_6985,N_4072,N_2874);
and U6986 (N_6986,N_2556,N_2662);
or U6987 (N_6987,N_4912,N_3593);
or U6988 (N_6988,N_3494,N_3288);
or U6989 (N_6989,N_4208,N_4381);
and U6990 (N_6990,N_4953,N_4545);
nand U6991 (N_6991,N_4428,N_3701);
nor U6992 (N_6992,N_4025,N_3776);
and U6993 (N_6993,N_4022,N_3026);
nand U6994 (N_6994,N_2906,N_2716);
nand U6995 (N_6995,N_3340,N_3983);
and U6996 (N_6996,N_2806,N_2712);
or U6997 (N_6997,N_2814,N_2668);
or U6998 (N_6998,N_4818,N_4219);
nor U6999 (N_6999,N_3196,N_3657);
nor U7000 (N_7000,N_4483,N_4196);
nor U7001 (N_7001,N_4491,N_4099);
nor U7002 (N_7002,N_3630,N_4995);
nor U7003 (N_7003,N_3951,N_2808);
nor U7004 (N_7004,N_3543,N_3351);
nand U7005 (N_7005,N_2725,N_3744);
nand U7006 (N_7006,N_4392,N_3067);
and U7007 (N_7007,N_4745,N_3547);
nand U7008 (N_7008,N_4404,N_2693);
nor U7009 (N_7009,N_4425,N_3644);
or U7010 (N_7010,N_4023,N_2568);
and U7011 (N_7011,N_4972,N_4188);
nand U7012 (N_7012,N_4363,N_2668);
nor U7013 (N_7013,N_2577,N_3463);
and U7014 (N_7014,N_3401,N_2793);
or U7015 (N_7015,N_4762,N_3086);
or U7016 (N_7016,N_3574,N_4604);
nand U7017 (N_7017,N_3274,N_4437);
or U7018 (N_7018,N_4951,N_3187);
nor U7019 (N_7019,N_4229,N_3881);
and U7020 (N_7020,N_4001,N_3768);
nor U7021 (N_7021,N_3481,N_4234);
nor U7022 (N_7022,N_4027,N_3654);
or U7023 (N_7023,N_2687,N_4781);
and U7024 (N_7024,N_4754,N_4662);
or U7025 (N_7025,N_3727,N_2792);
and U7026 (N_7026,N_3833,N_4472);
nand U7027 (N_7027,N_3650,N_4181);
and U7028 (N_7028,N_3671,N_3314);
or U7029 (N_7029,N_2642,N_3985);
nor U7030 (N_7030,N_3893,N_4287);
or U7031 (N_7031,N_2949,N_2920);
nand U7032 (N_7032,N_2832,N_3076);
nor U7033 (N_7033,N_3258,N_4336);
and U7034 (N_7034,N_3435,N_4463);
and U7035 (N_7035,N_3903,N_4751);
or U7036 (N_7036,N_2648,N_3554);
and U7037 (N_7037,N_2784,N_4678);
or U7038 (N_7038,N_4161,N_4398);
or U7039 (N_7039,N_3056,N_3165);
or U7040 (N_7040,N_3151,N_3827);
nor U7041 (N_7041,N_3917,N_3392);
xor U7042 (N_7042,N_3889,N_3718);
or U7043 (N_7043,N_4099,N_4907);
and U7044 (N_7044,N_4092,N_4109);
nand U7045 (N_7045,N_4515,N_3059);
or U7046 (N_7046,N_2989,N_3402);
nand U7047 (N_7047,N_2789,N_3361);
and U7048 (N_7048,N_3283,N_3370);
nand U7049 (N_7049,N_3092,N_3640);
and U7050 (N_7050,N_3067,N_4442);
or U7051 (N_7051,N_3212,N_4560);
nor U7052 (N_7052,N_4264,N_2524);
nor U7053 (N_7053,N_4207,N_3304);
nor U7054 (N_7054,N_2831,N_2556);
nor U7055 (N_7055,N_4646,N_3924);
or U7056 (N_7056,N_4892,N_4076);
or U7057 (N_7057,N_2709,N_2992);
nand U7058 (N_7058,N_3087,N_4557);
nand U7059 (N_7059,N_4589,N_4152);
nor U7060 (N_7060,N_4978,N_4233);
nor U7061 (N_7061,N_3772,N_2957);
and U7062 (N_7062,N_3916,N_4318);
or U7063 (N_7063,N_3566,N_3499);
or U7064 (N_7064,N_4546,N_3535);
nor U7065 (N_7065,N_4982,N_3161);
nor U7066 (N_7066,N_2874,N_2983);
and U7067 (N_7067,N_3158,N_4677);
and U7068 (N_7068,N_3187,N_3899);
nor U7069 (N_7069,N_3464,N_3780);
and U7070 (N_7070,N_2881,N_3385);
and U7071 (N_7071,N_2549,N_3213);
nand U7072 (N_7072,N_4644,N_2685);
nor U7073 (N_7073,N_3754,N_4820);
nor U7074 (N_7074,N_3839,N_3817);
xnor U7075 (N_7075,N_2575,N_2960);
nand U7076 (N_7076,N_4767,N_3609);
nand U7077 (N_7077,N_3311,N_4521);
or U7078 (N_7078,N_4543,N_3921);
or U7079 (N_7079,N_4406,N_4930);
nor U7080 (N_7080,N_3389,N_3199);
nor U7081 (N_7081,N_2853,N_3752);
or U7082 (N_7082,N_3895,N_4389);
nor U7083 (N_7083,N_2642,N_2994);
nor U7084 (N_7084,N_4207,N_2875);
and U7085 (N_7085,N_4684,N_2981);
nor U7086 (N_7086,N_2897,N_4479);
or U7087 (N_7087,N_3090,N_3795);
and U7088 (N_7088,N_3989,N_4881);
or U7089 (N_7089,N_3729,N_3089);
and U7090 (N_7090,N_2906,N_3628);
or U7091 (N_7091,N_2939,N_4522);
nor U7092 (N_7092,N_2838,N_4044);
or U7093 (N_7093,N_4012,N_4306);
nor U7094 (N_7094,N_4905,N_4121);
or U7095 (N_7095,N_4034,N_4783);
or U7096 (N_7096,N_3180,N_3450);
nor U7097 (N_7097,N_3066,N_3531);
nand U7098 (N_7098,N_3577,N_3443);
and U7099 (N_7099,N_3154,N_3424);
nand U7100 (N_7100,N_3717,N_3058);
nor U7101 (N_7101,N_4824,N_3167);
nand U7102 (N_7102,N_3871,N_3363);
nand U7103 (N_7103,N_4738,N_3963);
or U7104 (N_7104,N_4316,N_4008);
nor U7105 (N_7105,N_4158,N_4355);
and U7106 (N_7106,N_3278,N_3288);
or U7107 (N_7107,N_4596,N_3579);
and U7108 (N_7108,N_3687,N_2596);
nand U7109 (N_7109,N_4557,N_3216);
nand U7110 (N_7110,N_3618,N_2829);
and U7111 (N_7111,N_2840,N_2649);
nor U7112 (N_7112,N_4555,N_2723);
nand U7113 (N_7113,N_2529,N_4274);
or U7114 (N_7114,N_3493,N_2944);
and U7115 (N_7115,N_3487,N_4606);
or U7116 (N_7116,N_3288,N_3141);
and U7117 (N_7117,N_3437,N_3577);
nand U7118 (N_7118,N_2672,N_4766);
or U7119 (N_7119,N_3094,N_3851);
or U7120 (N_7120,N_4430,N_4530);
nand U7121 (N_7121,N_3405,N_3897);
nand U7122 (N_7122,N_4160,N_4759);
nor U7123 (N_7123,N_4634,N_2574);
nor U7124 (N_7124,N_2780,N_2532);
and U7125 (N_7125,N_3466,N_4796);
or U7126 (N_7126,N_3634,N_4982);
nand U7127 (N_7127,N_2934,N_4278);
nor U7128 (N_7128,N_3382,N_4673);
or U7129 (N_7129,N_4572,N_3119);
and U7130 (N_7130,N_3366,N_4941);
or U7131 (N_7131,N_2787,N_2973);
and U7132 (N_7132,N_2840,N_3834);
nor U7133 (N_7133,N_4736,N_2579);
nand U7134 (N_7134,N_4180,N_4036);
nor U7135 (N_7135,N_4284,N_4073);
or U7136 (N_7136,N_3910,N_2886);
nand U7137 (N_7137,N_2615,N_2864);
and U7138 (N_7138,N_4152,N_2970);
nor U7139 (N_7139,N_4528,N_3873);
nor U7140 (N_7140,N_4045,N_4461);
or U7141 (N_7141,N_4576,N_2590);
nand U7142 (N_7142,N_4933,N_4581);
nor U7143 (N_7143,N_3683,N_3438);
and U7144 (N_7144,N_4114,N_4979);
nand U7145 (N_7145,N_4789,N_4228);
and U7146 (N_7146,N_3380,N_3811);
nor U7147 (N_7147,N_3362,N_4553);
nand U7148 (N_7148,N_4077,N_2547);
nor U7149 (N_7149,N_3774,N_3394);
nand U7150 (N_7150,N_4845,N_4807);
nand U7151 (N_7151,N_4008,N_4189);
nand U7152 (N_7152,N_3631,N_4827);
or U7153 (N_7153,N_4053,N_2904);
nand U7154 (N_7154,N_3810,N_4491);
nor U7155 (N_7155,N_4504,N_4431);
nand U7156 (N_7156,N_2616,N_2500);
and U7157 (N_7157,N_3820,N_3423);
or U7158 (N_7158,N_3236,N_4046);
nand U7159 (N_7159,N_4494,N_3332);
or U7160 (N_7160,N_3713,N_3817);
nor U7161 (N_7161,N_4113,N_2528);
or U7162 (N_7162,N_4062,N_3307);
nand U7163 (N_7163,N_4189,N_4281);
nor U7164 (N_7164,N_3826,N_3656);
nor U7165 (N_7165,N_2927,N_4452);
nor U7166 (N_7166,N_3100,N_3566);
and U7167 (N_7167,N_3615,N_4553);
or U7168 (N_7168,N_2738,N_3898);
nand U7169 (N_7169,N_2603,N_3337);
nand U7170 (N_7170,N_4205,N_4925);
nor U7171 (N_7171,N_4619,N_4117);
nand U7172 (N_7172,N_3950,N_4654);
nor U7173 (N_7173,N_3302,N_4234);
nor U7174 (N_7174,N_4207,N_2630);
or U7175 (N_7175,N_3025,N_4444);
or U7176 (N_7176,N_3699,N_4317);
and U7177 (N_7177,N_4440,N_4051);
or U7178 (N_7178,N_3476,N_3027);
and U7179 (N_7179,N_2634,N_3731);
nand U7180 (N_7180,N_4793,N_2577);
or U7181 (N_7181,N_4357,N_3914);
and U7182 (N_7182,N_4218,N_4633);
or U7183 (N_7183,N_4731,N_3906);
and U7184 (N_7184,N_3721,N_3916);
nor U7185 (N_7185,N_3193,N_4143);
or U7186 (N_7186,N_4281,N_3172);
or U7187 (N_7187,N_3320,N_3604);
or U7188 (N_7188,N_2893,N_4229);
and U7189 (N_7189,N_2663,N_2714);
and U7190 (N_7190,N_4796,N_4368);
nor U7191 (N_7191,N_3738,N_2562);
and U7192 (N_7192,N_3136,N_3090);
nor U7193 (N_7193,N_3865,N_3352);
nor U7194 (N_7194,N_3264,N_3985);
or U7195 (N_7195,N_3295,N_4570);
nand U7196 (N_7196,N_4529,N_2790);
nor U7197 (N_7197,N_3122,N_3790);
nand U7198 (N_7198,N_4576,N_4560);
nor U7199 (N_7199,N_2575,N_3337);
nand U7200 (N_7200,N_2901,N_2848);
nand U7201 (N_7201,N_4835,N_4490);
and U7202 (N_7202,N_4897,N_3668);
and U7203 (N_7203,N_4090,N_3303);
nand U7204 (N_7204,N_3189,N_3212);
nand U7205 (N_7205,N_3746,N_4954);
or U7206 (N_7206,N_3816,N_3482);
or U7207 (N_7207,N_4105,N_3584);
or U7208 (N_7208,N_4571,N_2686);
and U7209 (N_7209,N_2737,N_4046);
or U7210 (N_7210,N_2968,N_2673);
and U7211 (N_7211,N_3325,N_3605);
nand U7212 (N_7212,N_4153,N_4321);
nor U7213 (N_7213,N_4221,N_3647);
or U7214 (N_7214,N_4384,N_3134);
nor U7215 (N_7215,N_4343,N_3664);
nor U7216 (N_7216,N_4639,N_2806);
nand U7217 (N_7217,N_3300,N_4692);
nand U7218 (N_7218,N_4566,N_4636);
xor U7219 (N_7219,N_4834,N_4311);
and U7220 (N_7220,N_3014,N_2517);
nand U7221 (N_7221,N_3053,N_4669);
nor U7222 (N_7222,N_4887,N_3428);
nand U7223 (N_7223,N_3534,N_4416);
or U7224 (N_7224,N_3657,N_4190);
or U7225 (N_7225,N_4985,N_4864);
or U7226 (N_7226,N_3708,N_3041);
or U7227 (N_7227,N_3200,N_3431);
and U7228 (N_7228,N_3502,N_4101);
nor U7229 (N_7229,N_3566,N_2753);
nand U7230 (N_7230,N_3979,N_4316);
or U7231 (N_7231,N_2768,N_4127);
nand U7232 (N_7232,N_4607,N_3073);
and U7233 (N_7233,N_4350,N_4761);
nand U7234 (N_7234,N_4051,N_3096);
and U7235 (N_7235,N_3283,N_3012);
or U7236 (N_7236,N_3744,N_4083);
nor U7237 (N_7237,N_3407,N_3870);
or U7238 (N_7238,N_4319,N_3063);
nor U7239 (N_7239,N_2873,N_4629);
and U7240 (N_7240,N_4432,N_2869);
or U7241 (N_7241,N_2511,N_3057);
nor U7242 (N_7242,N_3789,N_4070);
nor U7243 (N_7243,N_2695,N_3501);
or U7244 (N_7244,N_4212,N_3334);
nor U7245 (N_7245,N_2886,N_4250);
nand U7246 (N_7246,N_3110,N_4319);
or U7247 (N_7247,N_3435,N_4263);
and U7248 (N_7248,N_4344,N_2794);
or U7249 (N_7249,N_3302,N_4051);
nor U7250 (N_7250,N_4956,N_2597);
or U7251 (N_7251,N_3954,N_2750);
nor U7252 (N_7252,N_4804,N_4916);
or U7253 (N_7253,N_3992,N_2515);
and U7254 (N_7254,N_4174,N_4810);
nand U7255 (N_7255,N_4603,N_4895);
or U7256 (N_7256,N_2543,N_3890);
and U7257 (N_7257,N_3655,N_3289);
xnor U7258 (N_7258,N_3115,N_3694);
nor U7259 (N_7259,N_4506,N_3550);
or U7260 (N_7260,N_2819,N_4405);
nor U7261 (N_7261,N_4228,N_4648);
nor U7262 (N_7262,N_4352,N_2593);
nor U7263 (N_7263,N_4410,N_4677);
xnor U7264 (N_7264,N_4449,N_4761);
and U7265 (N_7265,N_3059,N_2654);
or U7266 (N_7266,N_2957,N_4941);
nand U7267 (N_7267,N_4933,N_2894);
nor U7268 (N_7268,N_3139,N_4690);
and U7269 (N_7269,N_3901,N_4632);
or U7270 (N_7270,N_4662,N_4148);
nor U7271 (N_7271,N_4065,N_4219);
nand U7272 (N_7272,N_3204,N_2925);
or U7273 (N_7273,N_4835,N_4664);
nand U7274 (N_7274,N_4607,N_4340);
or U7275 (N_7275,N_3551,N_3160);
xor U7276 (N_7276,N_3387,N_3921);
and U7277 (N_7277,N_3964,N_4054);
and U7278 (N_7278,N_4178,N_3879);
and U7279 (N_7279,N_3768,N_4391);
nand U7280 (N_7280,N_4516,N_3711);
xor U7281 (N_7281,N_3993,N_3393);
nor U7282 (N_7282,N_3990,N_4214);
nand U7283 (N_7283,N_4894,N_2805);
and U7284 (N_7284,N_3360,N_2653);
or U7285 (N_7285,N_2558,N_4892);
nand U7286 (N_7286,N_3984,N_3615);
nand U7287 (N_7287,N_4256,N_4849);
nor U7288 (N_7288,N_2657,N_3099);
nor U7289 (N_7289,N_2580,N_3151);
nand U7290 (N_7290,N_3898,N_2521);
and U7291 (N_7291,N_2781,N_3765);
nand U7292 (N_7292,N_4250,N_4777);
and U7293 (N_7293,N_2891,N_4838);
or U7294 (N_7294,N_2637,N_4278);
or U7295 (N_7295,N_3136,N_4282);
nor U7296 (N_7296,N_4238,N_4292);
and U7297 (N_7297,N_3011,N_2523);
or U7298 (N_7298,N_2547,N_3250);
nor U7299 (N_7299,N_4322,N_4458);
nand U7300 (N_7300,N_3621,N_4300);
or U7301 (N_7301,N_2994,N_4352);
nor U7302 (N_7302,N_4568,N_4231);
nand U7303 (N_7303,N_3973,N_2963);
or U7304 (N_7304,N_2995,N_4992);
or U7305 (N_7305,N_3273,N_2899);
nor U7306 (N_7306,N_4923,N_2535);
nand U7307 (N_7307,N_3131,N_3394);
nand U7308 (N_7308,N_4034,N_3209);
and U7309 (N_7309,N_3141,N_4882);
nor U7310 (N_7310,N_4645,N_3183);
nand U7311 (N_7311,N_3547,N_4071);
or U7312 (N_7312,N_4786,N_2908);
or U7313 (N_7313,N_4317,N_4630);
nor U7314 (N_7314,N_2756,N_4852);
and U7315 (N_7315,N_3779,N_4746);
and U7316 (N_7316,N_3407,N_4818);
nor U7317 (N_7317,N_2582,N_2541);
and U7318 (N_7318,N_2999,N_3839);
or U7319 (N_7319,N_3774,N_3421);
and U7320 (N_7320,N_2742,N_3861);
xnor U7321 (N_7321,N_4842,N_4035);
and U7322 (N_7322,N_4761,N_3567);
or U7323 (N_7323,N_3697,N_2528);
and U7324 (N_7324,N_3411,N_2823);
or U7325 (N_7325,N_3308,N_3268);
nor U7326 (N_7326,N_4271,N_2721);
and U7327 (N_7327,N_4862,N_3395);
nand U7328 (N_7328,N_4029,N_2637);
or U7329 (N_7329,N_3929,N_2773);
and U7330 (N_7330,N_4141,N_2979);
or U7331 (N_7331,N_4436,N_2762);
or U7332 (N_7332,N_3965,N_3169);
or U7333 (N_7333,N_2523,N_3743);
nor U7334 (N_7334,N_3233,N_3900);
or U7335 (N_7335,N_2995,N_3521);
or U7336 (N_7336,N_4633,N_3453);
and U7337 (N_7337,N_2587,N_2754);
or U7338 (N_7338,N_4177,N_3117);
nor U7339 (N_7339,N_4165,N_3100);
and U7340 (N_7340,N_4496,N_2922);
nand U7341 (N_7341,N_3372,N_4466);
nand U7342 (N_7342,N_2893,N_4466);
nand U7343 (N_7343,N_3484,N_3648);
and U7344 (N_7344,N_3475,N_2778);
nor U7345 (N_7345,N_3282,N_3205);
nor U7346 (N_7346,N_4219,N_2774);
and U7347 (N_7347,N_2646,N_3093);
or U7348 (N_7348,N_3424,N_4004);
nor U7349 (N_7349,N_2768,N_4634);
nand U7350 (N_7350,N_3277,N_4814);
nand U7351 (N_7351,N_3796,N_4184);
or U7352 (N_7352,N_2651,N_3562);
nand U7353 (N_7353,N_3686,N_3542);
and U7354 (N_7354,N_4043,N_3502);
nor U7355 (N_7355,N_4965,N_4619);
nor U7356 (N_7356,N_3685,N_4511);
or U7357 (N_7357,N_3999,N_4024);
and U7358 (N_7358,N_3298,N_4817);
nor U7359 (N_7359,N_3672,N_3892);
nor U7360 (N_7360,N_2573,N_2735);
nor U7361 (N_7361,N_2522,N_4987);
and U7362 (N_7362,N_3794,N_4064);
or U7363 (N_7363,N_4624,N_3004);
nor U7364 (N_7364,N_4601,N_3144);
and U7365 (N_7365,N_2572,N_2651);
nor U7366 (N_7366,N_3621,N_3827);
and U7367 (N_7367,N_2701,N_4408);
nand U7368 (N_7368,N_4423,N_3589);
nand U7369 (N_7369,N_3342,N_2812);
nand U7370 (N_7370,N_3529,N_3085);
and U7371 (N_7371,N_3593,N_3048);
nor U7372 (N_7372,N_3074,N_4968);
nor U7373 (N_7373,N_3400,N_3431);
xnor U7374 (N_7374,N_3641,N_2885);
and U7375 (N_7375,N_3278,N_4995);
nor U7376 (N_7376,N_3064,N_3937);
nor U7377 (N_7377,N_4620,N_2978);
nor U7378 (N_7378,N_2628,N_3680);
or U7379 (N_7379,N_3456,N_2649);
nand U7380 (N_7380,N_3526,N_4020);
nand U7381 (N_7381,N_3135,N_3656);
nand U7382 (N_7382,N_3749,N_4573);
or U7383 (N_7383,N_4069,N_4809);
and U7384 (N_7384,N_3997,N_3459);
nand U7385 (N_7385,N_4215,N_3118);
or U7386 (N_7386,N_4531,N_3213);
nand U7387 (N_7387,N_3910,N_2971);
and U7388 (N_7388,N_4761,N_3557);
or U7389 (N_7389,N_3338,N_4670);
and U7390 (N_7390,N_4813,N_3931);
and U7391 (N_7391,N_4004,N_4705);
and U7392 (N_7392,N_4608,N_4741);
nor U7393 (N_7393,N_4620,N_3336);
or U7394 (N_7394,N_2687,N_3223);
and U7395 (N_7395,N_4815,N_4781);
and U7396 (N_7396,N_3327,N_3235);
nor U7397 (N_7397,N_2584,N_4455);
and U7398 (N_7398,N_4052,N_4704);
nor U7399 (N_7399,N_4871,N_4407);
nand U7400 (N_7400,N_4790,N_3232);
and U7401 (N_7401,N_2556,N_4434);
and U7402 (N_7402,N_3687,N_4614);
or U7403 (N_7403,N_4115,N_4926);
and U7404 (N_7404,N_3151,N_4300);
nand U7405 (N_7405,N_4884,N_2979);
and U7406 (N_7406,N_4137,N_4965);
or U7407 (N_7407,N_3840,N_2842);
or U7408 (N_7408,N_4374,N_2591);
or U7409 (N_7409,N_3973,N_4308);
or U7410 (N_7410,N_4879,N_4103);
xor U7411 (N_7411,N_2542,N_4663);
and U7412 (N_7412,N_3983,N_4038);
or U7413 (N_7413,N_4830,N_4321);
nand U7414 (N_7414,N_3547,N_2829);
nand U7415 (N_7415,N_2930,N_3520);
nor U7416 (N_7416,N_4543,N_4633);
nand U7417 (N_7417,N_3993,N_3948);
nand U7418 (N_7418,N_4581,N_2600);
nor U7419 (N_7419,N_4090,N_2553);
or U7420 (N_7420,N_2773,N_3153);
or U7421 (N_7421,N_4599,N_4431);
and U7422 (N_7422,N_3688,N_4208);
or U7423 (N_7423,N_4258,N_4439);
nand U7424 (N_7424,N_2518,N_4449);
nand U7425 (N_7425,N_3130,N_4415);
nor U7426 (N_7426,N_4763,N_4575);
nor U7427 (N_7427,N_3939,N_2802);
and U7428 (N_7428,N_3081,N_3487);
nor U7429 (N_7429,N_4227,N_3073);
nand U7430 (N_7430,N_2986,N_2755);
or U7431 (N_7431,N_3786,N_3438);
or U7432 (N_7432,N_4383,N_3417);
nand U7433 (N_7433,N_3281,N_3127);
and U7434 (N_7434,N_3000,N_3701);
or U7435 (N_7435,N_2667,N_2914);
nor U7436 (N_7436,N_3064,N_4482);
or U7437 (N_7437,N_3616,N_3605);
and U7438 (N_7438,N_3898,N_3472);
or U7439 (N_7439,N_4517,N_2929);
and U7440 (N_7440,N_3381,N_2548);
and U7441 (N_7441,N_4218,N_4434);
nor U7442 (N_7442,N_3276,N_2834);
or U7443 (N_7443,N_4454,N_2916);
or U7444 (N_7444,N_3647,N_4485);
and U7445 (N_7445,N_3184,N_3105);
nand U7446 (N_7446,N_3234,N_3214);
and U7447 (N_7447,N_3575,N_4849);
or U7448 (N_7448,N_3541,N_2754);
and U7449 (N_7449,N_3355,N_3213);
nor U7450 (N_7450,N_4820,N_3036);
nand U7451 (N_7451,N_3005,N_4643);
nor U7452 (N_7452,N_4074,N_4041);
nand U7453 (N_7453,N_2506,N_3899);
nor U7454 (N_7454,N_4750,N_3243);
nand U7455 (N_7455,N_2537,N_4869);
nand U7456 (N_7456,N_3480,N_2627);
or U7457 (N_7457,N_4461,N_4498);
nor U7458 (N_7458,N_4886,N_3960);
or U7459 (N_7459,N_4598,N_2939);
and U7460 (N_7460,N_2959,N_3640);
or U7461 (N_7461,N_2602,N_4827);
and U7462 (N_7462,N_4802,N_4929);
nand U7463 (N_7463,N_3833,N_2579);
nand U7464 (N_7464,N_4146,N_4439);
or U7465 (N_7465,N_4084,N_2936);
or U7466 (N_7466,N_3340,N_4435);
nor U7467 (N_7467,N_3818,N_3676);
or U7468 (N_7468,N_3192,N_4671);
or U7469 (N_7469,N_2623,N_4891);
nand U7470 (N_7470,N_4803,N_4523);
nand U7471 (N_7471,N_3594,N_4260);
nor U7472 (N_7472,N_4245,N_3437);
nor U7473 (N_7473,N_3669,N_4232);
nor U7474 (N_7474,N_4840,N_3172);
or U7475 (N_7475,N_3429,N_2586);
nand U7476 (N_7476,N_3631,N_2540);
and U7477 (N_7477,N_3936,N_4535);
and U7478 (N_7478,N_2710,N_2864);
and U7479 (N_7479,N_3039,N_4486);
nor U7480 (N_7480,N_2774,N_4218);
nand U7481 (N_7481,N_3062,N_2898);
and U7482 (N_7482,N_4543,N_4125);
or U7483 (N_7483,N_4019,N_4147);
nand U7484 (N_7484,N_2778,N_4672);
nand U7485 (N_7485,N_4791,N_4550);
nor U7486 (N_7486,N_2666,N_3269);
or U7487 (N_7487,N_4328,N_4634);
and U7488 (N_7488,N_3546,N_4152);
nor U7489 (N_7489,N_4363,N_2521);
nand U7490 (N_7490,N_4475,N_4774);
nand U7491 (N_7491,N_3442,N_4908);
nand U7492 (N_7492,N_2535,N_4701);
and U7493 (N_7493,N_4318,N_2952);
nand U7494 (N_7494,N_2602,N_4676);
nand U7495 (N_7495,N_2745,N_2743);
or U7496 (N_7496,N_4525,N_4024);
or U7497 (N_7497,N_4037,N_3080);
nor U7498 (N_7498,N_4708,N_3390);
and U7499 (N_7499,N_3391,N_3698);
nor U7500 (N_7500,N_6908,N_7069);
nand U7501 (N_7501,N_6895,N_5346);
nor U7502 (N_7502,N_5932,N_5894);
or U7503 (N_7503,N_6667,N_7100);
or U7504 (N_7504,N_5676,N_5411);
nand U7505 (N_7505,N_5367,N_6362);
nor U7506 (N_7506,N_5500,N_7105);
nor U7507 (N_7507,N_5088,N_6503);
nor U7508 (N_7508,N_7060,N_5529);
and U7509 (N_7509,N_6113,N_7458);
nand U7510 (N_7510,N_6153,N_7264);
and U7511 (N_7511,N_5548,N_6190);
nand U7512 (N_7512,N_5139,N_5574);
or U7513 (N_7513,N_6636,N_5859);
nand U7514 (N_7514,N_6025,N_5908);
nand U7515 (N_7515,N_6757,N_5007);
or U7516 (N_7516,N_6334,N_7297);
and U7517 (N_7517,N_6480,N_6534);
nand U7518 (N_7518,N_6183,N_7445);
xor U7519 (N_7519,N_5535,N_5419);
nor U7520 (N_7520,N_6612,N_6373);
and U7521 (N_7521,N_7462,N_6106);
and U7522 (N_7522,N_5295,N_7189);
nor U7523 (N_7523,N_5552,N_5846);
or U7524 (N_7524,N_6098,N_6846);
nand U7525 (N_7525,N_7490,N_5654);
or U7526 (N_7526,N_5710,N_5178);
nand U7527 (N_7527,N_5871,N_5637);
or U7528 (N_7528,N_5168,N_6316);
and U7529 (N_7529,N_6478,N_6269);
nor U7530 (N_7530,N_5076,N_7292);
and U7531 (N_7531,N_6795,N_5935);
and U7532 (N_7532,N_7349,N_6450);
or U7533 (N_7533,N_7203,N_6767);
nor U7534 (N_7534,N_5200,N_5928);
nor U7535 (N_7535,N_5747,N_6763);
or U7536 (N_7536,N_7233,N_6035);
nand U7537 (N_7537,N_6713,N_5551);
xor U7538 (N_7538,N_6927,N_6909);
nand U7539 (N_7539,N_6651,N_5721);
or U7540 (N_7540,N_5426,N_7312);
and U7541 (N_7541,N_5353,N_6443);
nand U7542 (N_7542,N_5463,N_7088);
or U7543 (N_7543,N_5105,N_6003);
nand U7544 (N_7544,N_5695,N_6185);
nor U7545 (N_7545,N_5015,N_5366);
or U7546 (N_7546,N_5328,N_6387);
or U7547 (N_7547,N_7428,N_6009);
or U7548 (N_7548,N_5153,N_7115);
nand U7549 (N_7549,N_5011,N_6738);
nor U7550 (N_7550,N_5931,N_5691);
nor U7551 (N_7551,N_5503,N_5387);
or U7552 (N_7552,N_7262,N_6735);
and U7553 (N_7553,N_5762,N_7104);
or U7554 (N_7554,N_6550,N_6408);
nor U7555 (N_7555,N_6785,N_5425);
nand U7556 (N_7556,N_6426,N_6622);
and U7557 (N_7557,N_5855,N_6322);
nor U7558 (N_7558,N_5126,N_5711);
nor U7559 (N_7559,N_6123,N_7291);
and U7560 (N_7560,N_5818,N_6541);
and U7561 (N_7561,N_6463,N_7273);
nor U7562 (N_7562,N_6770,N_6119);
nand U7563 (N_7563,N_6732,N_5286);
or U7564 (N_7564,N_5669,N_5285);
nand U7565 (N_7565,N_5980,N_5441);
nand U7566 (N_7566,N_7194,N_6931);
or U7567 (N_7567,N_7110,N_5201);
and U7568 (N_7568,N_5761,N_6028);
nand U7569 (N_7569,N_6089,N_6220);
nand U7570 (N_7570,N_7023,N_7006);
or U7571 (N_7571,N_5939,N_5730);
and U7572 (N_7572,N_6553,N_7496);
nor U7573 (N_7573,N_6414,N_5892);
nor U7574 (N_7574,N_5712,N_6386);
or U7575 (N_7575,N_6876,N_5505);
or U7576 (N_7576,N_7204,N_5331);
nand U7577 (N_7577,N_5584,N_5190);
or U7578 (N_7578,N_7219,N_6068);
nand U7579 (N_7579,N_6234,N_6883);
or U7580 (N_7580,N_6142,N_5432);
or U7581 (N_7581,N_6283,N_7393);
nor U7582 (N_7582,N_5262,N_5434);
nor U7583 (N_7583,N_5448,N_6049);
nor U7584 (N_7584,N_5949,N_6349);
and U7585 (N_7585,N_7282,N_5655);
nand U7586 (N_7586,N_5388,N_5922);
or U7587 (N_7587,N_6700,N_6392);
nand U7588 (N_7588,N_5351,N_7119);
and U7589 (N_7589,N_6706,N_6157);
nor U7590 (N_7590,N_5031,N_5142);
or U7591 (N_7591,N_5720,N_5451);
nand U7592 (N_7592,N_6808,N_7321);
or U7593 (N_7593,N_6370,N_7420);
xnor U7594 (N_7594,N_6340,N_5072);
and U7595 (N_7595,N_6248,N_5945);
nor U7596 (N_7596,N_6102,N_7187);
and U7597 (N_7597,N_7185,N_6921);
or U7598 (N_7598,N_7410,N_5498);
and U7599 (N_7599,N_5148,N_5150);
and U7600 (N_7600,N_5116,N_6026);
nand U7601 (N_7601,N_7146,N_5942);
and U7602 (N_7602,N_5917,N_7357);
nor U7603 (N_7603,N_6029,N_5728);
nand U7604 (N_7604,N_5677,N_5996);
and U7605 (N_7605,N_5336,N_7228);
nor U7606 (N_7606,N_5350,N_7396);
or U7607 (N_7607,N_7113,N_7293);
nor U7608 (N_7608,N_6860,N_6532);
nor U7609 (N_7609,N_6440,N_5363);
and U7610 (N_7610,N_7141,N_5035);
nor U7611 (N_7611,N_7055,N_6189);
or U7612 (N_7612,N_5239,N_7376);
or U7613 (N_7613,N_5110,N_6052);
nor U7614 (N_7614,N_5540,N_5335);
nand U7615 (N_7615,N_6292,N_5061);
and U7616 (N_7616,N_5970,N_7386);
nor U7617 (N_7617,N_6829,N_7181);
nand U7618 (N_7618,N_5471,N_6156);
nor U7619 (N_7619,N_5050,N_5990);
and U7620 (N_7620,N_5074,N_6716);
or U7621 (N_7621,N_6796,N_7003);
and U7622 (N_7622,N_6634,N_6941);
nand U7623 (N_7623,N_5319,N_5330);
nand U7624 (N_7624,N_5054,N_6525);
or U7625 (N_7625,N_6179,N_5971);
and U7626 (N_7626,N_6528,N_5482);
nand U7627 (N_7627,N_5428,N_5863);
nor U7628 (N_7628,N_6261,N_6662);
nand U7629 (N_7629,N_7412,N_6653);
nor U7630 (N_7630,N_6586,N_6849);
or U7631 (N_7631,N_6213,N_7150);
and U7632 (N_7632,N_6658,N_7478);
nor U7633 (N_7633,N_7070,N_5468);
nand U7634 (N_7634,N_6229,N_5296);
or U7635 (N_7635,N_5784,N_5927);
nor U7636 (N_7636,N_5310,N_7295);
nor U7637 (N_7637,N_6843,N_7008);
nand U7638 (N_7638,N_7179,N_5359);
or U7639 (N_7639,N_5872,N_5699);
or U7640 (N_7640,N_6290,N_5660);
nor U7641 (N_7641,N_7311,N_6080);
and U7642 (N_7642,N_6556,N_5853);
or U7643 (N_7643,N_6875,N_6365);
nand U7644 (N_7644,N_7417,N_7419);
nor U7645 (N_7645,N_5952,N_5356);
nand U7646 (N_7646,N_6902,N_5571);
and U7647 (N_7647,N_6639,N_5521);
nor U7648 (N_7648,N_6115,N_6050);
and U7649 (N_7649,N_6991,N_7495);
and U7650 (N_7650,N_6898,N_6524);
nand U7651 (N_7651,N_5983,N_6238);
or U7652 (N_7652,N_6637,N_5948);
nand U7653 (N_7653,N_6583,N_6800);
nor U7654 (N_7654,N_5824,N_5467);
nor U7655 (N_7655,N_7031,N_5206);
or U7656 (N_7656,N_6314,N_6342);
nor U7657 (N_7657,N_5257,N_6014);
nor U7658 (N_7658,N_7235,N_5140);
or U7659 (N_7659,N_7245,N_6221);
nand U7660 (N_7660,N_6228,N_5458);
nor U7661 (N_7661,N_5687,N_6685);
and U7662 (N_7662,N_5003,N_5197);
nand U7663 (N_7663,N_5659,N_5213);
and U7664 (N_7664,N_7036,N_5183);
or U7665 (N_7665,N_5809,N_5134);
and U7666 (N_7666,N_6859,N_5272);
and U7667 (N_7667,N_6212,N_6928);
nor U7668 (N_7668,N_6704,N_5758);
nand U7669 (N_7669,N_7373,N_6818);
nand U7670 (N_7670,N_6660,N_7002);
nand U7671 (N_7671,N_5370,N_6057);
xor U7672 (N_7672,N_6648,N_5533);
nor U7673 (N_7673,N_6776,N_6574);
and U7674 (N_7674,N_6851,N_5947);
and U7675 (N_7675,N_6522,N_6817);
nor U7676 (N_7676,N_7168,N_6451);
and U7677 (N_7677,N_5217,N_5186);
nand U7678 (N_7678,N_7431,N_6870);
or U7679 (N_7679,N_7184,N_5369);
xnor U7680 (N_7680,N_5610,N_5019);
and U7681 (N_7681,N_6599,N_6638);
and U7682 (N_7682,N_6493,N_6078);
nand U7683 (N_7683,N_6861,N_6878);
and U7684 (N_7684,N_5974,N_5967);
nand U7685 (N_7685,N_5819,N_6570);
and U7686 (N_7686,N_5080,N_6620);
or U7687 (N_7687,N_5991,N_5680);
nand U7688 (N_7688,N_7065,N_5430);
and U7689 (N_7689,N_6589,N_5511);
nand U7690 (N_7690,N_5643,N_7337);
nor U7691 (N_7691,N_6232,N_5534);
and U7692 (N_7692,N_5668,N_7134);
nor U7693 (N_7693,N_7378,N_5175);
and U7694 (N_7694,N_5044,N_5266);
or U7695 (N_7695,N_6930,N_7080);
or U7696 (N_7696,N_6202,N_6852);
and U7697 (N_7697,N_5666,N_6762);
and U7698 (N_7698,N_7310,N_5166);
and U7699 (N_7699,N_7379,N_6251);
or U7700 (N_7700,N_5913,N_5856);
nor U7701 (N_7701,N_6975,N_5324);
xnor U7702 (N_7702,N_5544,N_7405);
or U7703 (N_7703,N_7126,N_5864);
nor U7704 (N_7704,N_6823,N_5941);
nand U7705 (N_7705,N_7016,N_6847);
and U7706 (N_7706,N_6429,N_5705);
and U7707 (N_7707,N_6799,N_5321);
or U7708 (N_7708,N_5121,N_5787);
and U7709 (N_7709,N_7047,N_5724);
nand U7710 (N_7710,N_5499,N_6977);
nor U7711 (N_7711,N_5365,N_7129);
or U7712 (N_7712,N_5156,N_6786);
and U7713 (N_7713,N_5953,N_5915);
nor U7714 (N_7714,N_6871,N_6476);
nor U7715 (N_7715,N_6237,N_6358);
or U7716 (N_7716,N_7304,N_6814);
nor U7717 (N_7717,N_5905,N_6730);
nor U7718 (N_7718,N_5027,N_6301);
nor U7719 (N_7719,N_5848,N_7195);
and U7720 (N_7720,N_5263,N_6621);
nand U7721 (N_7721,N_5603,N_6647);
and U7722 (N_7722,N_5767,N_6067);
or U7723 (N_7723,N_6967,N_6798);
nor U7724 (N_7724,N_5601,N_6084);
and U7725 (N_7725,N_5706,N_5563);
and U7726 (N_7726,N_6598,N_7358);
nor U7727 (N_7727,N_5934,N_6545);
or U7728 (N_7728,N_7395,N_6791);
nor U7729 (N_7729,N_5009,N_5043);
nand U7730 (N_7730,N_7025,N_7201);
nor U7731 (N_7731,N_6372,N_5822);
nand U7732 (N_7732,N_5250,N_5636);
or U7733 (N_7733,N_5128,N_7413);
nor U7734 (N_7734,N_5982,N_6579);
nand U7735 (N_7735,N_5984,N_6596);
and U7736 (N_7736,N_5966,N_6766);
nand U7737 (N_7737,N_7452,N_5661);
or U7738 (N_7738,N_5798,N_7045);
and U7739 (N_7739,N_6580,N_5355);
and U7740 (N_7740,N_5412,N_6956);
or U7741 (N_7741,N_5987,N_7300);
nor U7742 (N_7742,N_5943,N_6491);
nor U7743 (N_7743,N_6855,N_6572);
or U7744 (N_7744,N_5879,N_5746);
nor U7745 (N_7745,N_6425,N_6768);
or U7746 (N_7746,N_7248,N_6371);
and U7747 (N_7747,N_6148,N_6402);
nand U7748 (N_7748,N_7352,N_5813);
and U7749 (N_7749,N_5360,N_7165);
nor U7750 (N_7750,N_6311,N_5958);
nor U7751 (N_7751,N_6893,N_7402);
and U7752 (N_7752,N_6465,N_5522);
nand U7753 (N_7753,N_7131,N_5994);
nand U7754 (N_7754,N_6201,N_6203);
and U7755 (N_7755,N_5502,N_5218);
or U7756 (N_7756,N_7019,N_6635);
nand U7757 (N_7757,N_7062,N_6282);
and U7758 (N_7758,N_5821,N_6812);
nand U7759 (N_7759,N_5289,N_6173);
nor U7760 (N_7760,N_5878,N_6448);
nor U7761 (N_7761,N_5543,N_6015);
or U7762 (N_7762,N_6656,N_7385);
nand U7763 (N_7763,N_7064,N_6184);
and U7764 (N_7764,N_7261,N_5777);
or U7765 (N_7765,N_5851,N_7154);
nand U7766 (N_7766,N_5665,N_7294);
nor U7767 (N_7767,N_7192,N_6728);
or U7768 (N_7768,N_7360,N_5438);
and U7769 (N_7769,N_5111,N_5518);
or U7770 (N_7770,N_6108,N_6519);
nand U7771 (N_7771,N_7313,N_6987);
and U7772 (N_7772,N_6864,N_5199);
and U7773 (N_7773,N_6320,N_6219);
and U7774 (N_7774,N_7318,N_7058);
nand U7775 (N_7775,N_7037,N_7281);
and U7776 (N_7776,N_6527,N_5656);
or U7777 (N_7777,N_6710,N_7087);
nand U7778 (N_7778,N_7017,N_5163);
or U7779 (N_7779,N_6146,N_5442);
nand U7780 (N_7780,N_5246,N_6200);
and U7781 (N_7781,N_6266,N_6310);
nand U7782 (N_7782,N_5252,N_6935);
or U7783 (N_7783,N_6291,N_5796);
nor U7784 (N_7784,N_5021,N_5023);
nor U7785 (N_7785,N_6894,N_5267);
and U7786 (N_7786,N_5006,N_6518);
nand U7787 (N_7787,N_5307,N_6573);
or U7788 (N_7788,N_6815,N_6912);
nand U7789 (N_7789,N_5688,N_5383);
nand U7790 (N_7790,N_5870,N_5527);
and U7791 (N_7791,N_6077,N_5338);
and U7792 (N_7792,N_7299,N_7483);
or U7793 (N_7793,N_5597,N_6124);
or U7794 (N_7794,N_6794,N_5689);
nor U7795 (N_7795,N_5165,N_6252);
nor U7796 (N_7796,N_6952,N_6787);
nand U7797 (N_7797,N_7265,N_5833);
and U7798 (N_7798,N_6492,N_6711);
nand U7799 (N_7799,N_5089,N_6037);
nor U7800 (N_7800,N_5159,N_6903);
or U7801 (N_7801,N_6222,N_5042);
or U7802 (N_7802,N_5577,N_5647);
nor U7803 (N_7803,N_7053,N_5466);
or U7804 (N_7804,N_5398,N_5567);
and U7805 (N_7805,N_5269,N_6126);
nor U7806 (N_7806,N_5024,N_6976);
and U7807 (N_7807,N_6592,N_5133);
xor U7808 (N_7808,N_5093,N_7473);
or U7809 (N_7809,N_5480,N_5607);
nor U7810 (N_7810,N_5646,N_6646);
and U7811 (N_7811,N_5684,N_5125);
nor U7812 (N_7812,N_5944,N_6147);
nand U7813 (N_7813,N_7137,N_5137);
nor U7814 (N_7814,N_7120,N_7035);
nand U7815 (N_7815,N_5769,N_6932);
nand U7816 (N_7816,N_6990,N_6957);
nand U7817 (N_7817,N_6420,N_6705);
or U7818 (N_7818,N_5611,N_6582);
nand U7819 (N_7819,N_6442,N_6922);
nand U7820 (N_7820,N_6982,N_5802);
or U7821 (N_7821,N_6929,N_6023);
and U7822 (N_7822,N_6074,N_5616);
nor U7823 (N_7823,N_5354,N_5118);
xnor U7824 (N_7824,N_6474,N_5575);
or U7825 (N_7825,N_6198,N_6937);
nor U7826 (N_7826,N_7167,N_6216);
nand U7827 (N_7827,N_6194,N_6994);
and U7828 (N_7828,N_7488,N_5379);
nand U7829 (N_7829,N_7450,N_7421);
or U7830 (N_7830,N_5397,N_5858);
and U7831 (N_7831,N_5337,N_5897);
or U7832 (N_7832,N_6950,N_6407);
and U7833 (N_7833,N_6830,N_6769);
or U7834 (N_7834,N_6666,N_5185);
and U7835 (N_7835,N_5674,N_5946);
and U7836 (N_7836,N_7365,N_7033);
nor U7837 (N_7837,N_7253,N_6970);
or U7838 (N_7838,N_5051,N_5475);
nor U7839 (N_7839,N_5599,N_5733);
nor U7840 (N_7840,N_6630,N_5243);
and U7841 (N_7841,N_7086,N_6267);
nor U7842 (N_7842,N_7277,N_6286);
and U7843 (N_7843,N_5339,N_7072);
nor U7844 (N_7844,N_5248,N_5612);
or U7845 (N_7845,N_7079,N_5632);
nand U7846 (N_7846,N_5719,N_6946);
nor U7847 (N_7847,N_6918,N_5075);
nor U7848 (N_7848,N_7459,N_5176);
nor U7849 (N_7849,N_5594,N_6243);
and U7850 (N_7850,N_6816,N_5002);
or U7851 (N_7851,N_5483,N_5057);
nand U7852 (N_7852,N_7005,N_6192);
xnor U7853 (N_7853,N_6778,N_6703);
nand U7854 (N_7854,N_6784,N_7392);
nor U7855 (N_7855,N_5929,N_6754);
or U7856 (N_7856,N_6717,N_6724);
and U7857 (N_7857,N_5161,N_6743);
and U7858 (N_7858,N_6385,N_7461);
or U7859 (N_7859,N_6539,N_5580);
and U7860 (N_7860,N_5454,N_7007);
or U7861 (N_7861,N_5617,N_5315);
nand U7862 (N_7862,N_6718,N_5032);
and U7863 (N_7863,N_6629,N_5247);
nor U7864 (N_7864,N_7447,N_5470);
nand U7865 (N_7865,N_7470,N_5487);
nand U7866 (N_7866,N_5672,N_5145);
nor U7867 (N_7867,N_7403,N_5226);
or U7868 (N_7868,N_5961,N_5760);
nand U7869 (N_7869,N_5536,N_6974);
and U7870 (N_7870,N_5595,N_5249);
nor U7871 (N_7871,N_5107,N_6240);
nor U7872 (N_7872,N_6775,N_6032);
and U7873 (N_7873,N_5079,N_6178);
nor U7874 (N_7874,N_6661,N_5625);
and U7875 (N_7875,N_5129,N_6566);
nand U7876 (N_7876,N_6693,N_5405);
and U7877 (N_7877,N_5839,N_5293);
nand U7878 (N_7878,N_5083,N_5361);
nor U7879 (N_7879,N_6765,N_7375);
or U7880 (N_7880,N_7389,N_6617);
nand U7881 (N_7881,N_5431,N_5385);
or U7882 (N_7882,N_7116,N_5708);
or U7883 (N_7883,N_7381,N_5357);
nand U7884 (N_7884,N_5343,N_7399);
and U7885 (N_7885,N_6172,N_5332);
or U7886 (N_7886,N_6277,N_5070);
nand U7887 (N_7887,N_6033,N_7001);
nor U7888 (N_7888,N_6678,N_6809);
or U7889 (N_7889,N_6761,N_6403);
nand U7890 (N_7890,N_6208,N_7362);
and U7891 (N_7891,N_6838,N_7238);
nor U7892 (N_7892,N_5576,N_5582);
or U7893 (N_7893,N_5675,N_5488);
nor U7894 (N_7894,N_6038,N_6013);
nand U7895 (N_7895,N_6565,N_6313);
nand U7896 (N_7896,N_6563,N_5790);
nand U7897 (N_7897,N_5236,N_7229);
and U7898 (N_7898,N_6874,N_7174);
or U7899 (N_7899,N_5736,N_6684);
or U7900 (N_7900,N_6427,N_6613);
nor U7901 (N_7901,N_6307,N_6054);
nand U7902 (N_7902,N_6502,N_5960);
and U7903 (N_7903,N_6865,N_7152);
nand U7904 (N_7904,N_7372,N_7114);
nor U7905 (N_7905,N_7054,N_5400);
nor U7906 (N_7906,N_5745,N_5423);
or U7907 (N_7907,N_5566,N_6643);
or U7908 (N_7908,N_6933,N_6345);
nand U7909 (N_7909,N_6008,N_5222);
nand U7910 (N_7910,N_6597,N_6366);
nor U7911 (N_7911,N_6329,N_5472);
nand U7912 (N_7912,N_7198,N_7480);
and U7913 (N_7913,N_6915,N_6432);
nand U7914 (N_7914,N_6979,N_5352);
and U7915 (N_7915,N_7288,N_6083);
or U7916 (N_7916,N_5657,N_5341);
nor U7917 (N_7917,N_5390,N_5969);
and U7918 (N_7918,N_6632,N_7040);
and U7919 (N_7919,N_6352,N_6674);
nand U7920 (N_7920,N_5086,N_6961);
and U7921 (N_7921,N_6332,N_7454);
and U7922 (N_7922,N_6231,N_5826);
nand U7923 (N_7923,N_6577,N_7332);
nor U7924 (N_7924,N_5903,N_5744);
or U7925 (N_7925,N_7316,N_6835);
or U7926 (N_7926,N_6672,N_6584);
nand U7927 (N_7927,N_6335,N_6531);
or U7928 (N_7928,N_6422,N_7342);
nand U7929 (N_7929,N_6047,N_5737);
nand U7930 (N_7930,N_5055,N_6164);
or U7931 (N_7931,N_5810,N_7096);
and U7932 (N_7932,N_6547,N_6694);
nand U7933 (N_7933,N_6107,N_6917);
and U7934 (N_7934,N_5520,N_6182);
nand U7935 (N_7935,N_5697,N_5664);
nor U7936 (N_7936,N_6368,N_7144);
nand U7937 (N_7937,N_6681,N_5182);
or U7938 (N_7938,N_7051,N_5874);
or U7939 (N_7939,N_6390,N_7092);
nand U7940 (N_7940,N_5800,N_5038);
or U7941 (N_7941,N_6910,N_5381);
nor U7942 (N_7942,N_6697,N_5840);
nand U7943 (N_7943,N_5375,N_5590);
or U7944 (N_7944,N_7394,N_6030);
and U7945 (N_7945,N_6832,N_5741);
nand U7946 (N_7946,N_5732,N_5493);
nand U7947 (N_7947,N_6789,N_5513);
or U7948 (N_7948,N_5170,N_5081);
nor U7949 (N_7949,N_5241,N_5399);
nand U7950 (N_7950,N_7117,N_6866);
nor U7951 (N_7951,N_7247,N_5022);
nand U7952 (N_7952,N_5312,N_5010);
nor U7953 (N_7953,N_5287,N_5937);
or U7954 (N_7954,N_5530,N_6328);
nand U7955 (N_7955,N_7441,N_7382);
nor U7956 (N_7956,N_6459,N_6309);
nor U7957 (N_7957,N_6317,N_7324);
nand U7958 (N_7958,N_5000,N_6304);
nand U7959 (N_7959,N_6343,N_5804);
or U7960 (N_7960,N_6842,N_6544);
nand U7961 (N_7961,N_5144,N_6399);
and U7962 (N_7962,N_6051,N_6092);
nand U7963 (N_7963,N_5933,N_6130);
and U7964 (N_7964,N_6170,N_5198);
nor U7965 (N_7965,N_6455,N_6125);
or U7966 (N_7966,N_7391,N_6230);
or U7967 (N_7967,N_6073,N_7400);
nor U7968 (N_7968,N_7259,N_5794);
and U7969 (N_7969,N_5301,N_5273);
and U7970 (N_7970,N_6751,N_7455);
nand U7971 (N_7971,N_7449,N_6306);
and U7972 (N_7972,N_5828,N_5701);
and U7973 (N_7973,N_7415,N_7170);
nor U7974 (N_7974,N_5427,N_7061);
nand U7975 (N_7975,N_7308,N_6276);
nor U7976 (N_7976,N_6939,N_5275);
and U7977 (N_7977,N_5538,N_5885);
and U7978 (N_7978,N_5342,N_6535);
and U7979 (N_7979,N_5756,N_7084);
nor U7980 (N_7980,N_6076,N_7212);
and U7981 (N_7981,N_6065,N_6246);
nand U7982 (N_7982,N_5334,N_7498);
and U7983 (N_7983,N_7186,N_5151);
and U7984 (N_7984,N_5694,N_6516);
and U7985 (N_7985,N_6430,N_5436);
nand U7986 (N_7986,N_7401,N_6406);
and U7987 (N_7987,N_7284,N_6682);
nor U7988 (N_7988,N_5208,N_6241);
or U7989 (N_7989,N_7029,N_6161);
nand U7990 (N_7990,N_7028,N_5344);
or U7991 (N_7991,N_5755,N_6802);
nor U7992 (N_7992,N_5773,N_5670);
nand U7993 (N_7993,N_6327,N_7135);
or U7994 (N_7994,N_6564,N_5205);
or U7995 (N_7995,N_7098,N_7239);
nand U7996 (N_7996,N_5896,N_5146);
or U7997 (N_7997,N_6159,N_5384);
or U7998 (N_7998,N_6141,N_7083);
nor U7999 (N_7999,N_5995,N_6374);
and U8000 (N_8000,N_6548,N_5469);
nand U8001 (N_8001,N_5781,N_6217);
and U8002 (N_8002,N_5378,N_5834);
and U8003 (N_8003,N_5591,N_6677);
nor U8004 (N_8004,N_7177,N_6578);
or U8005 (N_8005,N_5377,N_5526);
and U8006 (N_8006,N_5555,N_6945);
nor U8007 (N_8007,N_5805,N_5512);
nor U8008 (N_8008,N_5622,N_5709);
nor U8009 (N_8009,N_5882,N_5026);
and U8010 (N_8010,N_6249,N_7370);
and U8011 (N_8011,N_5866,N_7090);
nor U8012 (N_8012,N_5649,N_6034);
or U8013 (N_8013,N_7099,N_5320);
nor U8014 (N_8014,N_6591,N_6740);
nor U8015 (N_8015,N_7387,N_5553);
or U8016 (N_8016,N_6568,N_5508);
nor U8017 (N_8017,N_6360,N_6278);
nand U8018 (N_8018,N_6122,N_5037);
or U8019 (N_8019,N_7207,N_5765);
nand U8020 (N_8020,N_5778,N_5314);
nand U8021 (N_8021,N_6603,N_6485);
nor U8022 (N_8022,N_6642,N_5223);
nand U8023 (N_8023,N_7094,N_5465);
or U8024 (N_8024,N_5306,N_6773);
and U8025 (N_8025,N_5406,N_6947);
nand U8026 (N_8026,N_7298,N_6060);
nor U8027 (N_8027,N_7444,N_5417);
or U8028 (N_8028,N_5780,N_6687);
or U8029 (N_8029,N_5396,N_6176);
nor U8030 (N_8030,N_5829,N_5507);
nor U8031 (N_8031,N_6268,N_5349);
nor U8032 (N_8032,N_6040,N_6383);
or U8033 (N_8033,N_6120,N_7091);
or U8034 (N_8034,N_6722,N_7232);
or U8035 (N_8035,N_6379,N_5638);
and U8036 (N_8036,N_6749,N_6145);
and U8037 (N_8037,N_5847,N_6714);
or U8038 (N_8038,N_5259,N_5868);
nor U8039 (N_8039,N_5380,N_7442);
nand U8040 (N_8040,N_6689,N_5416);
or U8041 (N_8041,N_7075,N_5046);
nand U8042 (N_8042,N_6433,N_7034);
and U8043 (N_8043,N_5734,N_6719);
nor U8044 (N_8044,N_7202,N_6691);
nor U8045 (N_8045,N_7303,N_5726);
or U8046 (N_8046,N_6562,N_6044);
nand U8047 (N_8047,N_7024,N_7271);
nor U8048 (N_8048,N_6271,N_7089);
or U8049 (N_8049,N_5421,N_5963);
nor U8050 (N_8050,N_6488,N_5449);
nand U8051 (N_8051,N_5005,N_6273);
and U8052 (N_8052,N_6560,N_6610);
nand U8053 (N_8053,N_7260,N_6367);
nor U8054 (N_8054,N_6224,N_7275);
nand U8055 (N_8055,N_5564,N_7171);
nand U8056 (N_8056,N_6558,N_6100);
or U8057 (N_8057,N_7082,N_5158);
and U8058 (N_8058,N_6364,N_5578);
or U8059 (N_8059,N_5298,N_5231);
and U8060 (N_8060,N_5883,N_6211);
or U8061 (N_8061,N_6165,N_7436);
nor U8062 (N_8062,N_7145,N_7249);
or U8063 (N_8063,N_5092,N_5254);
nor U8064 (N_8064,N_6513,N_6275);
nand U8065 (N_8065,N_7237,N_5194);
nand U8066 (N_8066,N_6081,N_5753);
or U8067 (N_8067,N_6435,N_5880);
nor U8068 (N_8068,N_6116,N_6020);
and U8069 (N_8069,N_5340,N_7158);
nor U8070 (N_8070,N_6167,N_5886);
or U8071 (N_8071,N_6663,N_6836);
nand U8072 (N_8072,N_6103,N_6188);
and U8073 (N_8073,N_6397,N_5914);
nand U8074 (N_8074,N_5841,N_6742);
and U8075 (N_8075,N_6175,N_5364);
nor U8076 (N_8076,N_6131,N_5525);
or U8077 (N_8077,N_6062,N_5069);
nand U8078 (N_8078,N_5270,N_6668);
or U8079 (N_8079,N_6325,N_6308);
or U8080 (N_8080,N_5783,N_6105);
nand U8081 (N_8081,N_5362,N_7157);
or U8082 (N_8082,N_5562,N_6396);
nor U8083 (N_8083,N_5509,N_6777);
nor U8084 (N_8084,N_6348,N_5347);
nand U8085 (N_8085,N_6441,N_6361);
and U8086 (N_8086,N_6012,N_6300);
and U8087 (N_8087,N_5018,N_5811);
or U8088 (N_8088,N_5799,N_5925);
nor U8089 (N_8089,N_6760,N_7283);
or U8090 (N_8090,N_6482,N_7435);
nor U8091 (N_8091,N_5389,N_5221);
nor U8092 (N_8092,N_6294,N_6059);
xor U8093 (N_8093,N_6319,N_7346);
nand U8094 (N_8094,N_7314,N_7102);
and U8095 (N_8095,N_6394,N_6581);
or U8096 (N_8096,N_5234,N_5951);
or U8097 (N_8097,N_5113,N_6953);
and U8098 (N_8098,N_6096,N_5678);
and U8099 (N_8099,N_6288,N_5714);
nand U8100 (N_8100,N_7408,N_5311);
and U8101 (N_8101,N_5975,N_5986);
or U8102 (N_8102,N_5593,N_6293);
and U8103 (N_8103,N_5748,N_6355);
or U8104 (N_8104,N_6608,N_6111);
and U8105 (N_8105,N_6168,N_5496);
and U8106 (N_8106,N_5401,N_6456);
nand U8107 (N_8107,N_6747,N_5481);
nand U8108 (N_8108,N_7121,N_5830);
and U8109 (N_8109,N_6091,N_6315);
or U8110 (N_8110,N_6436,N_6439);
nand U8111 (N_8111,N_6058,N_7209);
nor U8112 (N_8112,N_5279,N_6899);
and U8113 (N_8113,N_6772,N_5094);
nor U8114 (N_8114,N_7039,N_6413);
or U8115 (N_8115,N_5460,N_6454);
and U8116 (N_8116,N_7411,N_6152);
or U8117 (N_8117,N_5624,N_5752);
xnor U8118 (N_8118,N_5294,N_5180);
nand U8119 (N_8119,N_5317,N_5997);
nand U8120 (N_8120,N_6764,N_5253);
nand U8121 (N_8121,N_5028,N_6468);
and U8122 (N_8122,N_6460,N_6954);
nor U8123 (N_8123,N_6803,N_6771);
nand U8124 (N_8124,N_5309,N_5358);
nand U8125 (N_8125,N_5123,N_5230);
or U8126 (N_8126,N_5959,N_6353);
nor U8127 (N_8127,N_7156,N_6127);
or U8128 (N_8128,N_5912,N_6494);
nand U8129 (N_8129,N_6886,N_6998);
or U8130 (N_8130,N_6813,N_6887);
or U8131 (N_8131,N_5673,N_5924);
or U8132 (N_8132,N_6913,N_6417);
and U8133 (N_8133,N_6257,N_6758);
and U8134 (N_8134,N_7343,N_6053);
or U8135 (N_8135,N_6186,N_6896);
nand U8136 (N_8136,N_6983,N_7492);
nand U8137 (N_8137,N_6699,N_6393);
or U8138 (N_8138,N_6279,N_5523);
or U8139 (N_8139,N_5573,N_6128);
and U8140 (N_8140,N_6326,N_5102);
and U8141 (N_8141,N_5095,N_7221);
and U8142 (N_8142,N_6960,N_5962);
and U8143 (N_8143,N_6330,N_7359);
or U8144 (N_8144,N_6036,N_6723);
and U8145 (N_8145,N_6181,N_6788);
and U8146 (N_8146,N_5245,N_6986);
and U8147 (N_8147,N_5702,N_5053);
or U8148 (N_8148,N_6605,N_6966);
nand U8149 (N_8149,N_5082,N_6604);
or U8150 (N_8150,N_6099,N_5119);
nand U8151 (N_8151,N_5743,N_7467);
and U8152 (N_8152,N_7268,N_6418);
and U8153 (N_8153,N_5909,N_6272);
nand U8154 (N_8154,N_6690,N_6398);
nor U8155 (N_8155,N_6748,N_6000);
nand U8156 (N_8156,N_6239,N_7018);
and U8157 (N_8157,N_5403,N_5172);
or U8158 (N_8158,N_5435,N_5001);
nand U8159 (N_8159,N_5288,N_6024);
nor U8160 (N_8160,N_6999,N_6972);
and U8161 (N_8161,N_6404,N_5550);
or U8162 (N_8162,N_6045,N_5147);
nor U8163 (N_8163,N_7466,N_6701);
nand U8164 (N_8164,N_5938,N_6464);
nor U8165 (N_8165,N_7361,N_5189);
and U8166 (N_8166,N_7164,N_7424);
nand U8167 (N_8167,N_7009,N_5067);
nand U8168 (N_8168,N_5973,N_6759);
or U8169 (N_8169,N_5130,N_6569);
nand U8170 (N_8170,N_5029,N_7351);
nand U8171 (N_8171,N_7050,N_6965);
and U8172 (N_8172,N_6538,N_7038);
nor U8173 (N_8173,N_7108,N_5763);
nor U8174 (N_8174,N_7356,N_5779);
nand U8175 (N_8175,N_6191,N_6948);
nor U8176 (N_8176,N_6811,N_6477);
and U8177 (N_8177,N_5774,N_6741);
nor U8178 (N_8178,N_7138,N_5203);
or U8179 (N_8179,N_5652,N_5628);
and U8180 (N_8180,N_7042,N_7468);
nor U8181 (N_8181,N_5060,N_7149);
and U8182 (N_8182,N_6138,N_7364);
or U8183 (N_8183,N_7166,N_5570);
or U8184 (N_8184,N_6197,N_5989);
and U8185 (N_8185,N_5725,N_6698);
nor U8186 (N_8186,N_7255,N_5136);
and U8187 (N_8187,N_6114,N_6043);
nand U8188 (N_8188,N_6039,N_6779);
or U8189 (N_8189,N_6624,N_6302);
or U8190 (N_8190,N_6223,N_6409);
nand U8191 (N_8191,N_5477,N_5402);
or U8192 (N_8192,N_5844,N_6263);
nand U8193 (N_8193,N_5237,N_6782);
nor U8194 (N_8194,N_6207,N_7012);
or U8195 (N_8195,N_6139,N_6318);
and U8196 (N_8196,N_6136,N_5141);
or U8197 (N_8197,N_5227,N_6424);
or U8198 (N_8198,N_7407,N_6495);
nor U8199 (N_8199,N_6828,N_5907);
nand U8200 (N_8200,N_5440,N_5849);
and U8201 (N_8201,N_7326,N_6466);
nand U8202 (N_8202,N_7437,N_5073);
nor U8203 (N_8203,N_5167,N_7251);
nor U8204 (N_8204,N_6007,N_5683);
or U8205 (N_8205,N_7074,N_5860);
nor U8206 (N_8206,N_6774,N_5519);
nor U8207 (N_8207,N_5348,N_6906);
and U8208 (N_8208,N_6801,N_5554);
nand U8209 (N_8209,N_7477,N_6844);
nor U8210 (N_8210,N_7339,N_7497);
nor U8211 (N_8211,N_6911,N_6657);
xor U8212 (N_8212,N_7476,N_5209);
nand U8213 (N_8213,N_7112,N_5501);
nand U8214 (N_8214,N_6920,N_6696);
nand U8215 (N_8215,N_7127,N_7254);
or U8216 (N_8216,N_5751,N_6428);
nand U8217 (N_8217,N_6312,N_5211);
nand U8218 (N_8218,N_5174,N_5988);
nor U8219 (N_8219,N_7429,N_5572);
or U8220 (N_8220,N_5817,N_7124);
nand U8221 (N_8221,N_6727,N_5723);
or U8222 (N_8222,N_7015,N_6962);
and U8223 (N_8223,N_6631,N_6733);
nor U8224 (N_8224,N_6063,N_6853);
and U8225 (N_8225,N_7451,N_5302);
nor U8226 (N_8226,N_5921,N_7366);
or U8227 (N_8227,N_5604,N_7482);
or U8228 (N_8228,N_6521,N_6093);
xnor U8229 (N_8229,N_6337,N_7128);
nor U8230 (N_8230,N_5479,N_5539);
nand U8231 (N_8231,N_6590,N_6472);
nand U8232 (N_8232,N_5662,N_6686);
and U8233 (N_8233,N_6154,N_6625);
nor U8234 (N_8234,N_5485,N_6321);
or U8235 (N_8235,N_5106,N_7418);
or U8236 (N_8236,N_6511,N_5663);
nor U8237 (N_8237,N_7246,N_5492);
nand U8238 (N_8238,N_6171,N_7236);
or U8239 (N_8239,N_6822,N_5154);
or U8240 (N_8240,N_6226,N_6992);
or U8241 (N_8241,N_7081,N_6546);
nand U8242 (N_8242,N_6845,N_6255);
nand U8243 (N_8243,N_5443,N_5559);
and U8244 (N_8244,N_6016,N_5558);
or U8245 (N_8245,N_6551,N_6375);
nand U8246 (N_8246,N_6438,N_5993);
or U8247 (N_8247,N_7026,N_6297);
and U8248 (N_8248,N_7010,N_6163);
or U8249 (N_8249,N_5979,N_6410);
nor U8250 (N_8250,N_5631,N_7188);
or U8251 (N_8251,N_6389,N_6341);
nand U8252 (N_8252,N_6680,N_5606);
nand U8253 (N_8253,N_7469,N_7279);
and U8254 (N_8254,N_6529,N_5160);
nor U8255 (N_8255,N_5097,N_6021);
nor U8256 (N_8256,N_5735,N_5803);
or U8257 (N_8257,N_5965,N_7223);
nor U8258 (N_8258,N_5926,N_5825);
nor U8259 (N_8259,N_5936,N_5056);
nand U8260 (N_8260,N_5613,N_6489);
nand U8261 (N_8261,N_6506,N_7208);
or U8262 (N_8262,N_7301,N_6055);
or U8263 (N_8263,N_5700,N_5329);
xor U8264 (N_8264,N_5517,N_6151);
and U8265 (N_8265,N_7206,N_5045);
nor U8266 (N_8266,N_6287,N_7471);
nor U8267 (N_8267,N_5495,N_6810);
or U8268 (N_8268,N_6869,N_5464);
or U8269 (N_8269,N_6242,N_5282);
and U8270 (N_8270,N_7434,N_7041);
nor U8271 (N_8271,N_5409,N_5462);
nand U8272 (N_8272,N_5889,N_7344);
nor U8273 (N_8273,N_5797,N_7175);
nand U8274 (N_8274,N_6160,N_6180);
or U8275 (N_8275,N_7153,N_5256);
nand U8276 (N_8276,N_6737,N_7052);
or U8277 (N_8277,N_5108,N_5100);
nor U8278 (N_8278,N_7190,N_5524);
nor U8279 (N_8279,N_7250,N_5157);
or U8280 (N_8280,N_5327,N_7220);
nor U8281 (N_8281,N_5169,N_5025);
or U8282 (N_8282,N_5515,N_7196);
or U8283 (N_8283,N_5586,N_6709);
or U8284 (N_8284,N_6260,N_6174);
or U8285 (N_8285,N_5473,N_6351);
nand U8286 (N_8286,N_6989,N_5233);
nor U8287 (N_8287,N_6006,N_6623);
or U8288 (N_8288,N_5704,N_5770);
and U8289 (N_8289,N_5392,N_7147);
nor U8290 (N_8290,N_6499,N_7280);
or U8291 (N_8291,N_5992,N_7290);
or U8292 (N_8292,N_5474,N_7390);
nand U8293 (N_8293,N_7139,N_6218);
nor U8294 (N_8294,N_6780,N_5771);
or U8295 (N_8295,N_5195,N_6447);
nand U8296 (N_8296,N_5077,N_7085);
nor U8297 (N_8297,N_6940,N_6042);
xor U8298 (N_8298,N_6400,N_5598);
and U8299 (N_8299,N_6133,N_5382);
and U8300 (N_8300,N_7377,N_5651);
or U8301 (N_8301,N_7244,N_6072);
nor U8302 (N_8302,N_5906,N_7464);
and U8303 (N_8303,N_7241,N_6981);
and U8304 (N_8304,N_5801,N_6675);
nor U8305 (N_8305,N_6419,N_7243);
or U8306 (N_8306,N_5857,N_7032);
or U8307 (N_8307,N_5602,N_6395);
nor U8308 (N_8308,N_7021,N_5549);
or U8309 (N_8309,N_5012,N_5059);
or U8310 (N_8310,N_5875,N_5395);
nor U8311 (N_8311,N_6452,N_5193);
nand U8312 (N_8312,N_7263,N_7491);
or U8313 (N_8313,N_7136,N_6688);
nor U8314 (N_8314,N_7432,N_6926);
or U8315 (N_8315,N_6885,N_6633);
nor U8316 (N_8316,N_5835,N_6137);
or U8317 (N_8317,N_6745,N_6336);
nor U8318 (N_8318,N_5972,N_5615);
nor U8319 (N_8319,N_5215,N_6889);
nor U8320 (N_8320,N_7214,N_5418);
or U8321 (N_8321,N_5455,N_6143);
nand U8322 (N_8322,N_5977,N_5703);
nor U8323 (N_8323,N_5827,N_5484);
nand U8324 (N_8324,N_7148,N_6381);
and U8325 (N_8325,N_6101,N_5569);
or U8326 (N_8326,N_7354,N_6019);
nand U8327 (N_8327,N_6487,N_6753);
nand U8328 (N_8328,N_5033,N_6097);
nand U8329 (N_8329,N_6296,N_6199);
and U8330 (N_8330,N_6069,N_6654);
nand U8331 (N_8331,N_5066,N_6619);
nor U8332 (N_8332,N_6888,N_5609);
or U8333 (N_8333,N_6444,N_6245);
nor U8334 (N_8334,N_6356,N_6606);
nor U8335 (N_8335,N_6149,N_6095);
nand U8336 (N_8336,N_5394,N_7142);
nor U8337 (N_8337,N_7140,N_6509);
nand U8338 (N_8338,N_5323,N_5098);
nand U8339 (N_8339,N_7011,N_7191);
or U8340 (N_8340,N_6649,N_5838);
nand U8341 (N_8341,N_6378,N_5556);
nand U8342 (N_8342,N_7274,N_6980);
nor U8343 (N_8343,N_5785,N_6504);
nor U8344 (N_8344,N_5731,N_7077);
nor U8345 (N_8345,N_7494,N_6734);
xor U8346 (N_8346,N_5087,N_6496);
nand U8347 (N_8347,N_6274,N_6821);
and U8348 (N_8348,N_5117,N_5162);
and U8349 (N_8349,N_7071,N_7384);
xor U8350 (N_8350,N_5281,N_6559);
nand U8351 (N_8351,N_6209,N_7216);
or U8352 (N_8352,N_7151,N_5837);
and U8353 (N_8353,N_6567,N_6609);
nor U8354 (N_8354,N_5634,N_5476);
nand U8355 (N_8355,N_6295,N_5910);
nor U8356 (N_8356,N_6576,N_6520);
nor U8357 (N_8357,N_5642,N_5084);
nor U8358 (N_8358,N_7414,N_6434);
nor U8359 (N_8359,N_6508,N_6254);
nand U8360 (N_8360,N_5196,N_5681);
nand U8361 (N_8361,N_5715,N_6473);
nor U8362 (N_8362,N_5698,N_6963);
or U8363 (N_8363,N_5143,N_5177);
nand U8364 (N_8364,N_6324,N_5985);
nand U8365 (N_8365,N_7252,N_6923);
nor U8366 (N_8366,N_7287,N_5920);
and U8367 (N_8367,N_7169,N_6018);
and U8368 (N_8368,N_5494,N_5999);
and U8369 (N_8369,N_5276,N_5904);
nand U8370 (N_8370,N_6500,N_6721);
or U8371 (N_8371,N_5489,N_7161);
nor U8372 (N_8372,N_5738,N_6575);
xnor U8373 (N_8373,N_6155,N_5453);
xor U8374 (N_8374,N_5188,N_7327);
and U8375 (N_8375,N_6215,N_6840);
nand U8376 (N_8376,N_6514,N_7240);
nor U8377 (N_8377,N_7227,N_7296);
or U8378 (N_8378,N_6897,N_6346);
nor U8379 (N_8379,N_5039,N_6259);
or U8380 (N_8380,N_7388,N_6523);
nor U8381 (N_8381,N_5300,N_5291);
nand U8382 (N_8382,N_6914,N_6150);
nor U8383 (N_8383,N_6475,N_6530);
or U8384 (N_8384,N_6391,N_5930);
nand U8385 (N_8385,N_7183,N_6262);
or U8386 (N_8386,N_6736,N_5976);
nand U8387 (N_8387,N_5852,N_5957);
or U8388 (N_8388,N_6571,N_6616);
nand U8389 (N_8389,N_6793,N_7132);
nor U8390 (N_8390,N_6664,N_5408);
nand U8391 (N_8391,N_6880,N_5096);
or U8392 (N_8392,N_5303,N_5568);
nor U8393 (N_8393,N_5124,N_7347);
nor U8394 (N_8394,N_7374,N_5202);
and U8395 (N_8395,N_6117,N_5016);
and U8396 (N_8396,N_6628,N_6542);
or U8397 (N_8397,N_6431,N_6498);
or U8398 (N_8398,N_5545,N_7159);
nor U8399 (N_8399,N_5542,N_5255);
or U8400 (N_8400,N_7286,N_6792);
nand U8401 (N_8401,N_7307,N_7371);
nor U8402 (N_8402,N_7162,N_7440);
nand U8403 (N_8403,N_5374,N_5583);
nor U8404 (N_8404,N_5414,N_5184);
and U8405 (N_8405,N_7160,N_5807);
or U8406 (N_8406,N_7457,N_7200);
or U8407 (N_8407,N_6618,N_6862);
or U8408 (N_8408,N_5173,N_5793);
or U8409 (N_8409,N_5008,N_7397);
nand U8410 (N_8410,N_6086,N_6943);
nand U8411 (N_8411,N_5954,N_6892);
nor U8412 (N_8412,N_7348,N_5235);
or U8413 (N_8413,N_5047,N_6884);
nor U8414 (N_8414,N_5068,N_5322);
nor U8415 (N_8415,N_6641,N_7317);
and U8416 (N_8416,N_6993,N_7472);
and U8417 (N_8417,N_5393,N_5890);
nor U8418 (N_8418,N_5630,N_6985);
or U8419 (N_8419,N_6934,N_6350);
and U8420 (N_8420,N_6453,N_5528);
nor U8421 (N_8421,N_6824,N_5614);
nand U8422 (N_8422,N_6484,N_7234);
nor U8423 (N_8423,N_5696,N_6955);
nor U8424 (N_8424,N_5820,N_7199);
and U8425 (N_8425,N_6225,N_6357);
and U8426 (N_8426,N_5138,N_5629);
or U8427 (N_8427,N_5099,N_5621);
nor U8428 (N_8428,N_5090,N_7330);
nor U8429 (N_8429,N_5017,N_6075);
nand U8430 (N_8430,N_5112,N_6193);
nand U8431 (N_8431,N_7328,N_5478);
nand U8432 (N_8432,N_6627,N_6462);
nor U8433 (N_8433,N_6247,N_5103);
and U8434 (N_8434,N_6919,N_5816);
and U8435 (N_8435,N_5115,N_7049);
nand U8436 (N_8436,N_5041,N_5297);
nor U8437 (N_8437,N_6916,N_7460);
nand U8438 (N_8438,N_7059,N_5547);
nor U8439 (N_8439,N_6405,N_5459);
nor U8440 (N_8440,N_6907,N_6968);
and U8441 (N_8441,N_6118,N_5444);
nand U8442 (N_8442,N_6449,N_6665);
and U8443 (N_8443,N_7380,N_6347);
and U8444 (N_8444,N_6299,N_7122);
and U8445 (N_8445,N_6087,N_5653);
nor U8446 (N_8446,N_6333,N_6607);
nand U8447 (N_8447,N_6041,N_7231);
nor U8448 (N_8448,N_5212,N_6936);
nor U8449 (N_8449,N_6601,N_7197);
and U8450 (N_8450,N_6995,N_7499);
or U8451 (N_8451,N_6858,N_5058);
nor U8452 (N_8452,N_6692,N_6984);
nand U8453 (N_8453,N_6210,N_6715);
and U8454 (N_8454,N_6094,N_5600);
or U8455 (N_8455,N_5795,N_5750);
and U8456 (N_8456,N_5486,N_5919);
nand U8457 (N_8457,N_6650,N_6423);
and U8458 (N_8458,N_5713,N_6958);
and U8459 (N_8459,N_5313,N_5633);
nand U8460 (N_8460,N_5065,N_6557);
nor U8461 (N_8461,N_6594,N_5537);
nand U8462 (N_8462,N_6206,N_6533);
nor U8463 (N_8463,N_7363,N_5120);
and U8464 (N_8464,N_5034,N_5504);
nor U8465 (N_8465,N_5333,N_5439);
and U8466 (N_8466,N_6951,N_5749);
nand U8467 (N_8467,N_5596,N_5998);
and U8468 (N_8468,N_6265,N_7325);
nand U8469 (N_8469,N_5085,N_5955);
xnor U8470 (N_8470,N_5843,N_7107);
and U8471 (N_8471,N_6856,N_6805);
or U8472 (N_8472,N_5114,N_5179);
nand U8473 (N_8473,N_6515,N_6505);
nand U8474 (N_8474,N_6833,N_6807);
nor U8475 (N_8475,N_6820,N_6826);
nor U8476 (N_8476,N_5876,N_5579);
and U8477 (N_8477,N_6781,N_5639);
and U8478 (N_8478,N_6614,N_5901);
nand U8479 (N_8479,N_7270,N_5278);
and U8480 (N_8480,N_5740,N_5588);
nor U8481 (N_8481,N_5832,N_6806);
and U8482 (N_8482,N_6790,N_5923);
nand U8483 (N_8483,N_6540,N_7320);
or U8484 (N_8484,N_6825,N_6804);
or U8485 (N_8485,N_5881,N_6380);
nand U8486 (N_8486,N_6323,N_7485);
or U8487 (N_8487,N_7266,N_6944);
nand U8488 (N_8488,N_6001,N_6959);
nand U8489 (N_8489,N_6725,N_5260);
and U8490 (N_8490,N_5325,N_6305);
nand U8491 (N_8491,N_5030,N_5623);
nor U8492 (N_8492,N_6890,N_5373);
or U8493 (N_8493,N_5891,N_5238);
and U8494 (N_8494,N_6264,N_6082);
and U8495 (N_8495,N_5902,N_6289);
or U8496 (N_8496,N_6863,N_5242);
nor U8497 (N_8497,N_7425,N_6344);
and U8498 (N_8498,N_5831,N_7106);
nor U8499 (N_8499,N_5229,N_6924);
nand U8500 (N_8500,N_5277,N_6048);
nor U8501 (N_8501,N_6595,N_5693);
nor U8502 (N_8502,N_7355,N_5895);
nand U8503 (N_8503,N_6831,N_6109);
nor U8504 (N_8504,N_5978,N_7125);
nand U8505 (N_8505,N_6281,N_7044);
nor U8506 (N_8506,N_6090,N_5204);
nand U8507 (N_8507,N_5316,N_6669);
xnor U8508 (N_8508,N_5240,N_6708);
nand U8509 (N_8509,N_6158,N_6258);
nor U8510 (N_8510,N_5812,N_7073);
nor U8511 (N_8511,N_5754,N_5326);
nand U8512 (N_8512,N_7111,N_6022);
or U8513 (N_8513,N_5707,N_5063);
or U8514 (N_8514,N_5532,N_7067);
or U8515 (N_8515,N_7426,N_6978);
and U8516 (N_8516,N_5557,N_5433);
nor U8517 (N_8517,N_5561,N_6512);
or U8518 (N_8518,N_5768,N_6561);
or U8519 (N_8519,N_7453,N_6002);
nand U8520 (N_8520,N_6483,N_5514);
or U8521 (N_8521,N_5127,N_7109);
or U8522 (N_8522,N_7256,N_6611);
nand U8523 (N_8523,N_5516,N_7481);
and U8524 (N_8524,N_7057,N_6486);
nor U8525 (N_8525,N_5013,N_5048);
or U8526 (N_8526,N_6552,N_5268);
and U8527 (N_8527,N_5759,N_7463);
nand U8528 (N_8528,N_6079,N_7123);
nor U8529 (N_8529,N_6384,N_6490);
nor U8530 (N_8530,N_7013,N_6270);
nand U8531 (N_8531,N_5424,N_7048);
nand U8532 (N_8532,N_5718,N_7143);
and U8533 (N_8533,N_7258,N_5372);
nand U8534 (N_8534,N_6250,N_7319);
and U8535 (N_8535,N_6437,N_6676);
nor U8536 (N_8536,N_6536,N_6244);
or U8537 (N_8537,N_6416,N_6469);
and U8538 (N_8538,N_7336,N_6005);
nor U8539 (N_8539,N_5191,N_6872);
nor U8540 (N_8540,N_6027,N_5132);
or U8541 (N_8541,N_7331,N_6848);
nor U8542 (N_8542,N_6411,N_7224);
nand U8543 (N_8543,N_7215,N_6731);
or U8544 (N_8544,N_7433,N_6881);
or U8545 (N_8545,N_7334,N_5592);
nor U8546 (N_8546,N_7172,N_6507);
and U8547 (N_8547,N_5109,N_5456);
xnor U8548 (N_8548,N_6104,N_5786);
nor U8549 (N_8549,N_5682,N_7341);
and U8550 (N_8550,N_7333,N_6501);
or U8551 (N_8551,N_5626,N_5152);
or U8552 (N_8552,N_6827,N_5589);
and U8553 (N_8553,N_6354,N_6602);
nand U8554 (N_8554,N_7213,N_5224);
nand U8555 (N_8555,N_5232,N_6298);
and U8556 (N_8556,N_5171,N_5836);
nor U8557 (N_8557,N_5766,N_6587);
nand U8558 (N_8558,N_6555,N_6112);
or U8559 (N_8559,N_5271,N_6461);
or U8560 (N_8560,N_6303,N_6510);
nand U8561 (N_8561,N_6064,N_6671);
or U8562 (N_8562,N_6783,N_5415);
nand U8563 (N_8563,N_5404,N_7474);
xor U8564 (N_8564,N_6739,N_6481);
or U8565 (N_8565,N_6988,N_5679);
and U8566 (N_8566,N_6549,N_5968);
and U8567 (N_8567,N_6205,N_5071);
nor U8568 (N_8568,N_5292,N_7222);
and U8569 (N_8569,N_5608,N_5581);
nor U8570 (N_8570,N_5950,N_7272);
nand U8571 (N_8571,N_5187,N_6061);
nand U8572 (N_8572,N_6712,N_6363);
or U8573 (N_8573,N_5648,N_7210);
xor U8574 (N_8574,N_5956,N_5207);
or U8575 (N_8575,N_6331,N_6683);
nor U8576 (N_8576,N_5620,N_6695);
nand U8577 (N_8577,N_6949,N_7020);
and U8578 (N_8578,N_5104,N_5155);
nor U8579 (N_8579,N_5437,N_6129);
nor U8580 (N_8580,N_7218,N_7267);
nand U8581 (N_8581,N_6195,N_7486);
and U8582 (N_8582,N_7438,N_5192);
or U8583 (N_8583,N_7022,N_7302);
and U8584 (N_8584,N_7306,N_6882);
and U8585 (N_8585,N_5014,N_5772);
nor U8586 (N_8586,N_5911,N_6233);
nand U8587 (N_8587,N_6729,N_5587);
nand U8588 (N_8588,N_5605,N_5635);
nand U8589 (N_8589,N_6750,N_6744);
nand U8590 (N_8590,N_6971,N_5862);
or U8591 (N_8591,N_7030,N_6746);
nand U8592 (N_8592,N_5280,N_7479);
or U8593 (N_8593,N_7368,N_6997);
and U8594 (N_8594,N_5727,N_7309);
nand U8595 (N_8595,N_6707,N_7097);
and U8596 (N_8596,N_5510,N_6467);
nand U8597 (N_8597,N_6011,N_6236);
or U8598 (N_8598,N_7487,N_7173);
nor U8599 (N_8599,N_6615,N_5877);
or U8600 (N_8600,N_5101,N_5490);
or U8601 (N_8601,N_5447,N_5214);
xor U8602 (N_8602,N_7046,N_6187);
and U8603 (N_8603,N_5806,N_7118);
nor U8604 (N_8604,N_5887,N_7226);
nand U8605 (N_8605,N_5228,N_5420);
and U8606 (N_8606,N_6938,N_5842);
nor U8607 (N_8607,N_6285,N_5808);
and U8608 (N_8608,N_5641,N_5265);
or U8609 (N_8609,N_6640,N_6359);
and U8610 (N_8610,N_7367,N_7066);
or U8611 (N_8611,N_5645,N_5219);
nor U8612 (N_8612,N_5004,N_5290);
nand U8613 (N_8613,N_6479,N_6854);
or U8614 (N_8614,N_5814,N_7257);
or U8615 (N_8615,N_5618,N_7014);
nor U8616 (N_8616,N_5422,N_7205);
nand U8617 (N_8617,N_6526,N_6537);
or U8618 (N_8618,N_5220,N_5251);
and U8619 (N_8619,N_7335,N_5722);
or U8620 (N_8620,N_5918,N_7350);
and U8621 (N_8621,N_5052,N_7211);
nor U8622 (N_8622,N_7278,N_6867);
or U8623 (N_8623,N_5900,N_7093);
or U8624 (N_8624,N_6543,N_7383);
nand U8625 (N_8625,N_5413,N_5531);
nor U8626 (N_8626,N_6850,N_5888);
and U8627 (N_8627,N_7484,N_7409);
nand U8628 (N_8628,N_6121,N_7475);
and U8629 (N_8629,N_6891,N_5457);
nor U8630 (N_8630,N_6670,N_7217);
nand U8631 (N_8631,N_5898,N_5658);
or U8632 (N_8632,N_7276,N_7068);
or U8633 (N_8633,N_6857,N_7176);
nor U8634 (N_8634,N_5640,N_6470);
nand U8635 (N_8635,N_5446,N_5216);
nor U8636 (N_8636,N_5850,N_5899);
nand U8637 (N_8637,N_5506,N_7329);
nor U8638 (N_8638,N_7063,N_6196);
nor U8639 (N_8639,N_6756,N_7056);
and U8640 (N_8640,N_7225,N_6905);
nor U8641 (N_8641,N_5869,N_6284);
and U8642 (N_8642,N_6726,N_7163);
nor U8643 (N_8643,N_6162,N_5078);
and U8644 (N_8644,N_7230,N_7289);
nand U8645 (N_8645,N_6659,N_5452);
and U8646 (N_8646,N_6004,N_5845);
nor U8647 (N_8647,N_5261,N_6445);
nor U8648 (N_8648,N_5667,N_7493);
or U8649 (N_8649,N_6376,N_6837);
or U8650 (N_8650,N_6702,N_6056);
or U8651 (N_8651,N_6227,N_5776);
nand U8652 (N_8652,N_5873,N_5823);
and U8653 (N_8653,N_5345,N_7448);
or U8654 (N_8654,N_7369,N_5020);
nand U8655 (N_8655,N_6720,N_5585);
nand U8656 (N_8656,N_6177,N_7338);
and U8657 (N_8657,N_5717,N_6879);
or U8658 (N_8658,N_6140,N_6655);
nand U8659 (N_8659,N_7340,N_6214);
or U8660 (N_8660,N_6925,N_5884);
nand U8661 (N_8661,N_7422,N_6382);
and U8662 (N_8662,N_6070,N_6169);
or U8663 (N_8663,N_7076,N_6797);
or U8664 (N_8664,N_5775,N_7353);
nand U8665 (N_8665,N_6877,N_5305);
or U8666 (N_8666,N_5686,N_7430);
and U8667 (N_8667,N_7182,N_5764);
nor U8668 (N_8668,N_5036,N_6973);
or U8669 (N_8669,N_5546,N_7095);
nand U8670 (N_8670,N_5491,N_6868);
nand U8671 (N_8671,N_5135,N_5122);
or U8672 (N_8672,N_5964,N_6401);
nand U8673 (N_8673,N_5854,N_6046);
nor U8674 (N_8674,N_7178,N_6645);
nand U8675 (N_8675,N_7404,N_5541);
or U8676 (N_8676,N_7193,N_7242);
and U8677 (N_8677,N_6942,N_7465);
nor U8678 (N_8678,N_5916,N_6588);
nand U8679 (N_8679,N_5210,N_5739);
nor U8680 (N_8680,N_6204,N_7027);
nor U8681 (N_8681,N_6017,N_6600);
nand U8682 (N_8682,N_5304,N_6673);
and U8683 (N_8683,N_5565,N_7323);
or U8684 (N_8684,N_7439,N_5560);
or U8685 (N_8685,N_5644,N_5497);
or U8686 (N_8686,N_5692,N_6144);
nor U8687 (N_8687,N_6446,N_5792);
nand U8688 (N_8688,N_6593,N_6755);
or U8689 (N_8689,N_7000,N_7416);
nand U8690 (N_8690,N_5283,N_6134);
nand U8691 (N_8691,N_5690,N_7180);
and U8692 (N_8692,N_7305,N_5264);
or U8693 (N_8693,N_6626,N_7423);
nor U8694 (N_8694,N_5685,N_5429);
or U8695 (N_8695,N_5742,N_7103);
or U8696 (N_8696,N_5258,N_6457);
and U8697 (N_8697,N_6841,N_5064);
xor U8698 (N_8698,N_6458,N_5782);
nand U8699 (N_8699,N_6644,N_5308);
xnor U8700 (N_8700,N_6873,N_5225);
or U8701 (N_8701,N_6819,N_5371);
nand U8702 (N_8702,N_5149,N_6132);
or U8703 (N_8703,N_6253,N_5091);
nor U8704 (N_8704,N_6652,N_6031);
nor U8705 (N_8705,N_7406,N_6388);
nor U8706 (N_8706,N_7322,N_5244);
nor U8707 (N_8707,N_5791,N_7043);
nand U8708 (N_8708,N_6085,N_5376);
or U8709 (N_8709,N_7133,N_5789);
and U8710 (N_8710,N_6517,N_5450);
nand U8711 (N_8711,N_5788,N_6339);
and U8712 (N_8712,N_6901,N_6071);
nand U8713 (N_8713,N_6679,N_5040);
and U8714 (N_8714,N_5729,N_5619);
or U8715 (N_8715,N_5627,N_5391);
xor U8716 (N_8716,N_5716,N_7398);
nor U8717 (N_8717,N_5299,N_6088);
nand U8718 (N_8718,N_5049,N_5410);
and U8719 (N_8719,N_5671,N_5940);
nor U8720 (N_8720,N_7130,N_7489);
and U8721 (N_8721,N_5650,N_7446);
nor U8722 (N_8722,N_5062,N_6066);
nand U8723 (N_8723,N_6369,N_7443);
or U8724 (N_8724,N_7285,N_6256);
and U8725 (N_8725,N_6554,N_6969);
or U8726 (N_8726,N_6377,N_6235);
nand U8727 (N_8727,N_7004,N_6421);
nand U8728 (N_8728,N_6135,N_6996);
nand U8729 (N_8729,N_5386,N_5181);
nor U8730 (N_8730,N_6415,N_6280);
and U8731 (N_8731,N_5815,N_5861);
and U8732 (N_8732,N_6497,N_7456);
nor U8733 (N_8733,N_6166,N_7101);
or U8734 (N_8734,N_6338,N_7078);
nand U8735 (N_8735,N_5865,N_5164);
or U8736 (N_8736,N_5407,N_5757);
or U8737 (N_8737,N_5274,N_6010);
or U8738 (N_8738,N_6904,N_6900);
or U8739 (N_8739,N_5284,N_6839);
and U8740 (N_8740,N_6110,N_7315);
nor U8741 (N_8741,N_6834,N_6585);
nor U8742 (N_8742,N_5368,N_5981);
nor U8743 (N_8743,N_5318,N_5867);
or U8744 (N_8744,N_5131,N_5461);
or U8745 (N_8745,N_7427,N_6412);
nor U8746 (N_8746,N_7345,N_6964);
nand U8747 (N_8747,N_6752,N_6471);
and U8748 (N_8748,N_5893,N_7269);
or U8749 (N_8749,N_7155,N_5445);
nor U8750 (N_8750,N_5697,N_7102);
and U8751 (N_8751,N_6172,N_7196);
nand U8752 (N_8752,N_5524,N_5065);
nand U8753 (N_8753,N_7263,N_7039);
nand U8754 (N_8754,N_7160,N_6674);
nor U8755 (N_8755,N_5585,N_6519);
nor U8756 (N_8756,N_7474,N_5344);
and U8757 (N_8757,N_5264,N_5949);
xnor U8758 (N_8758,N_5524,N_5151);
nand U8759 (N_8759,N_7495,N_7449);
or U8760 (N_8760,N_6223,N_6894);
or U8761 (N_8761,N_7203,N_6881);
nand U8762 (N_8762,N_6345,N_5355);
nand U8763 (N_8763,N_5648,N_7489);
nand U8764 (N_8764,N_7382,N_6853);
or U8765 (N_8765,N_7048,N_7350);
or U8766 (N_8766,N_6804,N_5938);
or U8767 (N_8767,N_5604,N_7172);
nor U8768 (N_8768,N_6094,N_5019);
and U8769 (N_8769,N_5178,N_6913);
or U8770 (N_8770,N_5776,N_5924);
nor U8771 (N_8771,N_5375,N_5224);
and U8772 (N_8772,N_5041,N_5147);
nor U8773 (N_8773,N_5919,N_5242);
nand U8774 (N_8774,N_7156,N_7206);
xnor U8775 (N_8775,N_6647,N_5570);
and U8776 (N_8776,N_6580,N_6807);
nor U8777 (N_8777,N_6691,N_7024);
nand U8778 (N_8778,N_5521,N_5075);
or U8779 (N_8779,N_6109,N_5349);
nand U8780 (N_8780,N_7048,N_7303);
nor U8781 (N_8781,N_5227,N_7281);
and U8782 (N_8782,N_6339,N_6844);
and U8783 (N_8783,N_5175,N_7355);
xnor U8784 (N_8784,N_5612,N_5011);
nor U8785 (N_8785,N_7384,N_6751);
or U8786 (N_8786,N_5415,N_7242);
nor U8787 (N_8787,N_6336,N_6296);
or U8788 (N_8788,N_6632,N_5055);
or U8789 (N_8789,N_7354,N_5123);
nand U8790 (N_8790,N_5220,N_7345);
and U8791 (N_8791,N_6528,N_6471);
nand U8792 (N_8792,N_5220,N_5431);
nor U8793 (N_8793,N_5896,N_5652);
or U8794 (N_8794,N_7054,N_5097);
or U8795 (N_8795,N_6967,N_5292);
nand U8796 (N_8796,N_5460,N_7245);
and U8797 (N_8797,N_7463,N_7484);
or U8798 (N_8798,N_6658,N_5969);
nor U8799 (N_8799,N_7252,N_5543);
and U8800 (N_8800,N_6698,N_5061);
or U8801 (N_8801,N_6436,N_5327);
nor U8802 (N_8802,N_6223,N_6723);
nor U8803 (N_8803,N_6114,N_6570);
nor U8804 (N_8804,N_5998,N_5002);
or U8805 (N_8805,N_5581,N_7261);
nand U8806 (N_8806,N_6723,N_7288);
or U8807 (N_8807,N_6210,N_7419);
or U8808 (N_8808,N_5065,N_5715);
or U8809 (N_8809,N_5234,N_6281);
or U8810 (N_8810,N_7377,N_6747);
and U8811 (N_8811,N_6976,N_5158);
nor U8812 (N_8812,N_6192,N_6386);
nor U8813 (N_8813,N_6895,N_5714);
nand U8814 (N_8814,N_6748,N_5275);
or U8815 (N_8815,N_6427,N_7392);
and U8816 (N_8816,N_7285,N_5500);
and U8817 (N_8817,N_7165,N_6694);
or U8818 (N_8818,N_5054,N_5372);
or U8819 (N_8819,N_5474,N_6703);
or U8820 (N_8820,N_5098,N_6766);
or U8821 (N_8821,N_6617,N_5926);
or U8822 (N_8822,N_5959,N_5302);
or U8823 (N_8823,N_5129,N_5191);
and U8824 (N_8824,N_5819,N_6402);
and U8825 (N_8825,N_6962,N_5981);
and U8826 (N_8826,N_7016,N_6511);
nor U8827 (N_8827,N_5618,N_6612);
or U8828 (N_8828,N_5579,N_7268);
nand U8829 (N_8829,N_7487,N_7064);
nor U8830 (N_8830,N_6026,N_5932);
or U8831 (N_8831,N_5668,N_7285);
or U8832 (N_8832,N_6866,N_6700);
nor U8833 (N_8833,N_5153,N_7087);
or U8834 (N_8834,N_6576,N_5346);
nand U8835 (N_8835,N_5544,N_6230);
or U8836 (N_8836,N_5299,N_6247);
nor U8837 (N_8837,N_6190,N_5648);
nand U8838 (N_8838,N_7407,N_5882);
nor U8839 (N_8839,N_7259,N_5410);
and U8840 (N_8840,N_5170,N_7128);
nor U8841 (N_8841,N_5893,N_5332);
and U8842 (N_8842,N_5142,N_6776);
nand U8843 (N_8843,N_5207,N_7405);
and U8844 (N_8844,N_6097,N_6019);
nor U8845 (N_8845,N_5492,N_5795);
nor U8846 (N_8846,N_5137,N_7095);
and U8847 (N_8847,N_6458,N_5062);
or U8848 (N_8848,N_5861,N_7153);
or U8849 (N_8849,N_6673,N_7167);
nand U8850 (N_8850,N_6027,N_5881);
nor U8851 (N_8851,N_6156,N_5275);
or U8852 (N_8852,N_5070,N_6507);
nor U8853 (N_8853,N_5866,N_7149);
or U8854 (N_8854,N_6602,N_7051);
and U8855 (N_8855,N_6770,N_5693);
or U8856 (N_8856,N_7232,N_5193);
nand U8857 (N_8857,N_6223,N_6060);
or U8858 (N_8858,N_7180,N_7019);
or U8859 (N_8859,N_6107,N_5489);
nand U8860 (N_8860,N_5236,N_6677);
nand U8861 (N_8861,N_5507,N_5980);
nor U8862 (N_8862,N_5523,N_5255);
and U8863 (N_8863,N_5626,N_6126);
and U8864 (N_8864,N_7467,N_6604);
or U8865 (N_8865,N_7270,N_5735);
nor U8866 (N_8866,N_5717,N_5042);
nand U8867 (N_8867,N_6857,N_7430);
nand U8868 (N_8868,N_6327,N_6724);
nor U8869 (N_8869,N_5897,N_6044);
or U8870 (N_8870,N_6220,N_6848);
and U8871 (N_8871,N_6525,N_5938);
or U8872 (N_8872,N_5389,N_7377);
nor U8873 (N_8873,N_5883,N_5948);
nand U8874 (N_8874,N_5054,N_6763);
nor U8875 (N_8875,N_5472,N_5379);
and U8876 (N_8876,N_6376,N_5092);
and U8877 (N_8877,N_6118,N_6604);
nor U8878 (N_8878,N_6458,N_5582);
nor U8879 (N_8879,N_6793,N_5114);
nand U8880 (N_8880,N_5554,N_7475);
nand U8881 (N_8881,N_5765,N_5253);
and U8882 (N_8882,N_6384,N_6420);
nor U8883 (N_8883,N_6938,N_5250);
nor U8884 (N_8884,N_6527,N_5189);
nand U8885 (N_8885,N_5782,N_5445);
or U8886 (N_8886,N_5453,N_6209);
xor U8887 (N_8887,N_5234,N_6102);
nand U8888 (N_8888,N_5495,N_6722);
or U8889 (N_8889,N_5460,N_6878);
or U8890 (N_8890,N_6720,N_6959);
nor U8891 (N_8891,N_6187,N_7132);
and U8892 (N_8892,N_7264,N_5488);
nor U8893 (N_8893,N_5858,N_7111);
nor U8894 (N_8894,N_5954,N_6278);
and U8895 (N_8895,N_5830,N_5840);
nand U8896 (N_8896,N_7037,N_6301);
nand U8897 (N_8897,N_6335,N_5120);
nor U8898 (N_8898,N_6331,N_5811);
and U8899 (N_8899,N_5745,N_5366);
nand U8900 (N_8900,N_5210,N_5383);
and U8901 (N_8901,N_5604,N_6512);
or U8902 (N_8902,N_6181,N_6638);
nor U8903 (N_8903,N_5959,N_7418);
and U8904 (N_8904,N_6861,N_5798);
and U8905 (N_8905,N_6859,N_7031);
and U8906 (N_8906,N_5754,N_5197);
or U8907 (N_8907,N_7379,N_5152);
nor U8908 (N_8908,N_5541,N_7311);
nand U8909 (N_8909,N_5691,N_6866);
nor U8910 (N_8910,N_6164,N_5750);
and U8911 (N_8911,N_6703,N_6742);
nand U8912 (N_8912,N_6258,N_6014);
nand U8913 (N_8913,N_6494,N_6580);
and U8914 (N_8914,N_5895,N_5994);
or U8915 (N_8915,N_7483,N_6219);
and U8916 (N_8916,N_7043,N_6710);
nor U8917 (N_8917,N_7337,N_6122);
nand U8918 (N_8918,N_7236,N_7316);
xor U8919 (N_8919,N_6387,N_5585);
nand U8920 (N_8920,N_6157,N_6252);
nor U8921 (N_8921,N_6808,N_5232);
or U8922 (N_8922,N_6317,N_6443);
nand U8923 (N_8923,N_7165,N_6801);
or U8924 (N_8924,N_6249,N_5341);
and U8925 (N_8925,N_6406,N_6350);
or U8926 (N_8926,N_5611,N_6824);
nand U8927 (N_8927,N_5271,N_7470);
or U8928 (N_8928,N_5918,N_5357);
and U8929 (N_8929,N_7437,N_7080);
nor U8930 (N_8930,N_5057,N_6157);
nand U8931 (N_8931,N_5833,N_7209);
nand U8932 (N_8932,N_6227,N_5683);
and U8933 (N_8933,N_6666,N_6346);
nand U8934 (N_8934,N_6235,N_7398);
and U8935 (N_8935,N_6388,N_6981);
or U8936 (N_8936,N_6562,N_7010);
nor U8937 (N_8937,N_6053,N_5136);
nor U8938 (N_8938,N_6337,N_5829);
or U8939 (N_8939,N_6180,N_6984);
nand U8940 (N_8940,N_5174,N_7494);
or U8941 (N_8941,N_5606,N_6440);
and U8942 (N_8942,N_5258,N_6487);
or U8943 (N_8943,N_6313,N_7304);
and U8944 (N_8944,N_7377,N_6852);
nor U8945 (N_8945,N_5561,N_6469);
and U8946 (N_8946,N_6506,N_5722);
nand U8947 (N_8947,N_7079,N_6871);
and U8948 (N_8948,N_5898,N_5544);
or U8949 (N_8949,N_5738,N_5134);
or U8950 (N_8950,N_5823,N_6905);
nand U8951 (N_8951,N_6556,N_7081);
nand U8952 (N_8952,N_5269,N_5156);
and U8953 (N_8953,N_7241,N_5357);
nand U8954 (N_8954,N_6304,N_6729);
nand U8955 (N_8955,N_5584,N_6768);
nor U8956 (N_8956,N_6940,N_7246);
nor U8957 (N_8957,N_5145,N_7262);
or U8958 (N_8958,N_7166,N_7042);
nand U8959 (N_8959,N_5294,N_5592);
xnor U8960 (N_8960,N_5733,N_5890);
and U8961 (N_8961,N_6818,N_5440);
or U8962 (N_8962,N_5069,N_6036);
nor U8963 (N_8963,N_5871,N_5729);
nand U8964 (N_8964,N_5356,N_5879);
nand U8965 (N_8965,N_7368,N_6485);
nor U8966 (N_8966,N_7362,N_6328);
nor U8967 (N_8967,N_5216,N_7029);
nor U8968 (N_8968,N_5535,N_5275);
or U8969 (N_8969,N_5063,N_6417);
nor U8970 (N_8970,N_7087,N_7192);
or U8971 (N_8971,N_7167,N_6117);
nor U8972 (N_8972,N_5404,N_7047);
nand U8973 (N_8973,N_6110,N_7430);
nor U8974 (N_8974,N_6941,N_7481);
or U8975 (N_8975,N_5556,N_5788);
nand U8976 (N_8976,N_6610,N_6907);
or U8977 (N_8977,N_6640,N_6681);
nand U8978 (N_8978,N_6202,N_5841);
nor U8979 (N_8979,N_5806,N_7230);
and U8980 (N_8980,N_5638,N_7153);
or U8981 (N_8981,N_6846,N_6234);
or U8982 (N_8982,N_7195,N_7276);
and U8983 (N_8983,N_6064,N_6378);
nor U8984 (N_8984,N_6065,N_5214);
nor U8985 (N_8985,N_7102,N_5340);
nor U8986 (N_8986,N_7180,N_7376);
or U8987 (N_8987,N_5534,N_6991);
nand U8988 (N_8988,N_6540,N_6375);
nand U8989 (N_8989,N_5429,N_7165);
nor U8990 (N_8990,N_7267,N_7098);
nand U8991 (N_8991,N_5716,N_5883);
nand U8992 (N_8992,N_5251,N_6931);
nand U8993 (N_8993,N_6649,N_5163);
or U8994 (N_8994,N_5796,N_6822);
nor U8995 (N_8995,N_5372,N_7318);
nand U8996 (N_8996,N_5691,N_5280);
xor U8997 (N_8997,N_5256,N_7409);
or U8998 (N_8998,N_5559,N_6868);
or U8999 (N_8999,N_5829,N_6149);
nand U9000 (N_9000,N_5372,N_6092);
or U9001 (N_9001,N_6437,N_5537);
nor U9002 (N_9002,N_6698,N_7123);
and U9003 (N_9003,N_5717,N_7395);
nor U9004 (N_9004,N_7385,N_7491);
nand U9005 (N_9005,N_5785,N_5218);
or U9006 (N_9006,N_7125,N_5510);
or U9007 (N_9007,N_6563,N_5089);
nand U9008 (N_9008,N_6346,N_5603);
or U9009 (N_9009,N_6831,N_6059);
and U9010 (N_9010,N_5181,N_6417);
and U9011 (N_9011,N_6278,N_6900);
or U9012 (N_9012,N_5952,N_6791);
nand U9013 (N_9013,N_5784,N_7473);
nand U9014 (N_9014,N_7047,N_5742);
and U9015 (N_9015,N_7406,N_6671);
nor U9016 (N_9016,N_6456,N_6292);
and U9017 (N_9017,N_5151,N_5436);
nor U9018 (N_9018,N_7116,N_5660);
or U9019 (N_9019,N_6136,N_5765);
nand U9020 (N_9020,N_6176,N_5970);
or U9021 (N_9021,N_5682,N_6721);
or U9022 (N_9022,N_5318,N_5880);
and U9023 (N_9023,N_7047,N_7149);
nand U9024 (N_9024,N_6744,N_5196);
and U9025 (N_9025,N_5532,N_7199);
nand U9026 (N_9026,N_6256,N_5903);
nand U9027 (N_9027,N_6496,N_5851);
nand U9028 (N_9028,N_5293,N_5345);
or U9029 (N_9029,N_6386,N_5836);
and U9030 (N_9030,N_5971,N_6118);
nor U9031 (N_9031,N_5928,N_5128);
nor U9032 (N_9032,N_7360,N_6921);
nand U9033 (N_9033,N_6562,N_5067);
nand U9034 (N_9034,N_6521,N_7221);
nand U9035 (N_9035,N_5963,N_7099);
and U9036 (N_9036,N_5527,N_6307);
and U9037 (N_9037,N_5994,N_5397);
nand U9038 (N_9038,N_5273,N_6705);
or U9039 (N_9039,N_6034,N_5709);
or U9040 (N_9040,N_6898,N_5392);
nor U9041 (N_9041,N_5441,N_7499);
and U9042 (N_9042,N_5066,N_5550);
or U9043 (N_9043,N_7134,N_6498);
nor U9044 (N_9044,N_6673,N_5912);
or U9045 (N_9045,N_5755,N_6980);
nand U9046 (N_9046,N_5058,N_7075);
nor U9047 (N_9047,N_5255,N_5649);
nand U9048 (N_9048,N_5037,N_7453);
nand U9049 (N_9049,N_5690,N_5765);
nor U9050 (N_9050,N_5068,N_6116);
or U9051 (N_9051,N_6557,N_7345);
and U9052 (N_9052,N_5967,N_5505);
nor U9053 (N_9053,N_5540,N_5401);
nand U9054 (N_9054,N_5601,N_5305);
nor U9055 (N_9055,N_5938,N_6374);
or U9056 (N_9056,N_7446,N_7374);
and U9057 (N_9057,N_5278,N_5309);
nand U9058 (N_9058,N_5615,N_7056);
nor U9059 (N_9059,N_6620,N_5483);
and U9060 (N_9060,N_7272,N_7009);
or U9061 (N_9061,N_5848,N_6131);
nand U9062 (N_9062,N_5444,N_5713);
nor U9063 (N_9063,N_6929,N_5373);
nor U9064 (N_9064,N_5481,N_5258);
or U9065 (N_9065,N_5554,N_5345);
or U9066 (N_9066,N_6448,N_6248);
and U9067 (N_9067,N_6186,N_5480);
nor U9068 (N_9068,N_7212,N_6686);
and U9069 (N_9069,N_6520,N_7194);
and U9070 (N_9070,N_6483,N_5595);
or U9071 (N_9071,N_5581,N_5353);
nand U9072 (N_9072,N_5042,N_5845);
or U9073 (N_9073,N_5536,N_6071);
nor U9074 (N_9074,N_5749,N_7448);
nor U9075 (N_9075,N_5661,N_7247);
nand U9076 (N_9076,N_6086,N_5825);
and U9077 (N_9077,N_5011,N_6980);
or U9078 (N_9078,N_7420,N_5232);
or U9079 (N_9079,N_5332,N_5275);
nand U9080 (N_9080,N_7277,N_5642);
and U9081 (N_9081,N_5499,N_7476);
nor U9082 (N_9082,N_6802,N_6355);
and U9083 (N_9083,N_5257,N_5556);
nand U9084 (N_9084,N_5336,N_7064);
nor U9085 (N_9085,N_5561,N_7319);
and U9086 (N_9086,N_5198,N_5829);
and U9087 (N_9087,N_6231,N_6119);
nand U9088 (N_9088,N_7247,N_7025);
nor U9089 (N_9089,N_5789,N_7135);
nor U9090 (N_9090,N_5764,N_7138);
xnor U9091 (N_9091,N_7184,N_7001);
nor U9092 (N_9092,N_6334,N_6276);
nand U9093 (N_9093,N_7477,N_6965);
nand U9094 (N_9094,N_5810,N_5947);
nor U9095 (N_9095,N_6036,N_5186);
nor U9096 (N_9096,N_5202,N_5477);
and U9097 (N_9097,N_5449,N_5434);
nand U9098 (N_9098,N_6172,N_5707);
or U9099 (N_9099,N_6426,N_5808);
and U9100 (N_9100,N_5924,N_6978);
nor U9101 (N_9101,N_5592,N_5880);
nand U9102 (N_9102,N_5597,N_6732);
and U9103 (N_9103,N_5283,N_6864);
nor U9104 (N_9104,N_6423,N_6735);
and U9105 (N_9105,N_5704,N_5235);
nor U9106 (N_9106,N_7413,N_6122);
nand U9107 (N_9107,N_7259,N_7336);
nor U9108 (N_9108,N_5554,N_6315);
nor U9109 (N_9109,N_7402,N_6471);
and U9110 (N_9110,N_5416,N_5638);
and U9111 (N_9111,N_7002,N_5274);
nand U9112 (N_9112,N_7087,N_7057);
or U9113 (N_9113,N_6625,N_6854);
and U9114 (N_9114,N_5083,N_5470);
and U9115 (N_9115,N_7343,N_6748);
and U9116 (N_9116,N_6211,N_6377);
and U9117 (N_9117,N_6292,N_6391);
and U9118 (N_9118,N_6092,N_5804);
or U9119 (N_9119,N_6567,N_5117);
nand U9120 (N_9120,N_5879,N_5643);
nand U9121 (N_9121,N_6912,N_7032);
nor U9122 (N_9122,N_5719,N_7018);
and U9123 (N_9123,N_7274,N_6956);
and U9124 (N_9124,N_6390,N_5493);
or U9125 (N_9125,N_5721,N_5671);
nor U9126 (N_9126,N_7182,N_6040);
and U9127 (N_9127,N_6983,N_6455);
nand U9128 (N_9128,N_6189,N_6064);
or U9129 (N_9129,N_7387,N_5103);
nand U9130 (N_9130,N_5026,N_5120);
and U9131 (N_9131,N_6200,N_6066);
nor U9132 (N_9132,N_6442,N_5357);
and U9133 (N_9133,N_7273,N_7481);
nor U9134 (N_9134,N_7465,N_6289);
nand U9135 (N_9135,N_6669,N_6529);
and U9136 (N_9136,N_6096,N_5779);
nor U9137 (N_9137,N_5537,N_5221);
and U9138 (N_9138,N_5812,N_5544);
and U9139 (N_9139,N_6147,N_5865);
nor U9140 (N_9140,N_6756,N_6603);
nand U9141 (N_9141,N_7043,N_5688);
or U9142 (N_9142,N_6630,N_6539);
and U9143 (N_9143,N_5335,N_6252);
and U9144 (N_9144,N_5980,N_7442);
nand U9145 (N_9145,N_6296,N_5889);
nand U9146 (N_9146,N_5695,N_6190);
or U9147 (N_9147,N_5079,N_5572);
or U9148 (N_9148,N_5918,N_5944);
and U9149 (N_9149,N_7235,N_5895);
and U9150 (N_9150,N_5376,N_6119);
nand U9151 (N_9151,N_5777,N_6327);
or U9152 (N_9152,N_6441,N_5109);
nand U9153 (N_9153,N_5719,N_5061);
or U9154 (N_9154,N_7237,N_6141);
or U9155 (N_9155,N_5505,N_5630);
and U9156 (N_9156,N_6274,N_5154);
or U9157 (N_9157,N_6197,N_7385);
and U9158 (N_9158,N_6641,N_7051);
nand U9159 (N_9159,N_6040,N_5125);
nand U9160 (N_9160,N_7109,N_6259);
nor U9161 (N_9161,N_5675,N_5368);
and U9162 (N_9162,N_5593,N_6987);
and U9163 (N_9163,N_6704,N_5091);
or U9164 (N_9164,N_7305,N_5555);
nor U9165 (N_9165,N_6980,N_5428);
nand U9166 (N_9166,N_5643,N_7230);
nand U9167 (N_9167,N_5794,N_5065);
nand U9168 (N_9168,N_6039,N_7137);
and U9169 (N_9169,N_7325,N_5133);
nor U9170 (N_9170,N_6763,N_6753);
nand U9171 (N_9171,N_5691,N_7276);
nor U9172 (N_9172,N_6379,N_6499);
nor U9173 (N_9173,N_6469,N_5765);
and U9174 (N_9174,N_6570,N_7221);
or U9175 (N_9175,N_6931,N_5512);
nor U9176 (N_9176,N_5798,N_6382);
or U9177 (N_9177,N_5386,N_5099);
and U9178 (N_9178,N_5135,N_6075);
or U9179 (N_9179,N_5610,N_5078);
and U9180 (N_9180,N_6846,N_6254);
and U9181 (N_9181,N_7326,N_5262);
or U9182 (N_9182,N_6528,N_6779);
and U9183 (N_9183,N_6695,N_5338);
nor U9184 (N_9184,N_5242,N_7301);
or U9185 (N_9185,N_6903,N_5865);
or U9186 (N_9186,N_7240,N_7056);
nor U9187 (N_9187,N_6086,N_6720);
nand U9188 (N_9188,N_7328,N_7157);
or U9189 (N_9189,N_6186,N_6233);
and U9190 (N_9190,N_6884,N_7127);
nand U9191 (N_9191,N_6407,N_7311);
and U9192 (N_9192,N_5981,N_5051);
nand U9193 (N_9193,N_7162,N_7407);
nor U9194 (N_9194,N_5486,N_6491);
and U9195 (N_9195,N_7355,N_5845);
or U9196 (N_9196,N_6798,N_7078);
nand U9197 (N_9197,N_5285,N_5095);
xnor U9198 (N_9198,N_5354,N_5934);
and U9199 (N_9199,N_6087,N_5969);
nor U9200 (N_9200,N_6426,N_5466);
nand U9201 (N_9201,N_7420,N_5063);
nand U9202 (N_9202,N_5495,N_5509);
and U9203 (N_9203,N_7324,N_6342);
or U9204 (N_9204,N_6457,N_6707);
nand U9205 (N_9205,N_7064,N_6940);
and U9206 (N_9206,N_6354,N_7412);
nand U9207 (N_9207,N_6782,N_5564);
and U9208 (N_9208,N_6822,N_6725);
or U9209 (N_9209,N_5039,N_7370);
and U9210 (N_9210,N_5084,N_6977);
and U9211 (N_9211,N_7006,N_5381);
nor U9212 (N_9212,N_5374,N_7233);
or U9213 (N_9213,N_6601,N_6549);
nor U9214 (N_9214,N_6882,N_7005);
or U9215 (N_9215,N_5710,N_5303);
or U9216 (N_9216,N_6508,N_6354);
and U9217 (N_9217,N_5016,N_6542);
nor U9218 (N_9218,N_7358,N_5266);
and U9219 (N_9219,N_6664,N_6860);
or U9220 (N_9220,N_7439,N_6542);
or U9221 (N_9221,N_5221,N_7018);
nand U9222 (N_9222,N_6101,N_7166);
nor U9223 (N_9223,N_6967,N_7116);
and U9224 (N_9224,N_6359,N_7140);
nand U9225 (N_9225,N_5078,N_5761);
and U9226 (N_9226,N_6278,N_5463);
nand U9227 (N_9227,N_7028,N_5666);
or U9228 (N_9228,N_7155,N_5506);
or U9229 (N_9229,N_5092,N_5913);
or U9230 (N_9230,N_5139,N_6966);
or U9231 (N_9231,N_6090,N_5158);
nand U9232 (N_9232,N_5667,N_5821);
or U9233 (N_9233,N_7116,N_7460);
nor U9234 (N_9234,N_6615,N_7287);
xnor U9235 (N_9235,N_5358,N_6445);
or U9236 (N_9236,N_6785,N_7371);
nand U9237 (N_9237,N_5013,N_6167);
nand U9238 (N_9238,N_7244,N_6795);
and U9239 (N_9239,N_7384,N_6814);
nor U9240 (N_9240,N_5141,N_6164);
and U9241 (N_9241,N_6458,N_6762);
or U9242 (N_9242,N_7454,N_5723);
nor U9243 (N_9243,N_6885,N_5483);
or U9244 (N_9244,N_6615,N_5442);
xor U9245 (N_9245,N_5240,N_6889);
nor U9246 (N_9246,N_7418,N_6897);
and U9247 (N_9247,N_5820,N_5637);
nor U9248 (N_9248,N_6941,N_7100);
or U9249 (N_9249,N_6387,N_5090);
or U9250 (N_9250,N_5182,N_6559);
or U9251 (N_9251,N_7303,N_5273);
nand U9252 (N_9252,N_6362,N_6690);
nor U9253 (N_9253,N_5411,N_7480);
or U9254 (N_9254,N_6821,N_6898);
and U9255 (N_9255,N_5688,N_7446);
and U9256 (N_9256,N_5470,N_7181);
and U9257 (N_9257,N_6844,N_6854);
and U9258 (N_9258,N_6068,N_6063);
or U9259 (N_9259,N_6762,N_5530);
nand U9260 (N_9260,N_6673,N_6801);
or U9261 (N_9261,N_5446,N_6197);
nand U9262 (N_9262,N_5469,N_5094);
or U9263 (N_9263,N_6962,N_6281);
nor U9264 (N_9264,N_6286,N_6563);
nand U9265 (N_9265,N_7462,N_6692);
or U9266 (N_9266,N_5898,N_6467);
and U9267 (N_9267,N_5645,N_5686);
nor U9268 (N_9268,N_6171,N_5313);
nand U9269 (N_9269,N_6514,N_5661);
and U9270 (N_9270,N_5966,N_7266);
or U9271 (N_9271,N_7400,N_6545);
or U9272 (N_9272,N_6475,N_5614);
nor U9273 (N_9273,N_5584,N_7427);
nor U9274 (N_9274,N_7371,N_7090);
nand U9275 (N_9275,N_6745,N_5923);
nand U9276 (N_9276,N_5232,N_7319);
nand U9277 (N_9277,N_6153,N_5805);
or U9278 (N_9278,N_5924,N_5562);
or U9279 (N_9279,N_5182,N_6745);
xor U9280 (N_9280,N_5069,N_6155);
or U9281 (N_9281,N_6975,N_5099);
nand U9282 (N_9282,N_6912,N_7293);
or U9283 (N_9283,N_7145,N_7451);
or U9284 (N_9284,N_6530,N_6612);
nor U9285 (N_9285,N_5019,N_5225);
or U9286 (N_9286,N_6861,N_7429);
nand U9287 (N_9287,N_7431,N_7197);
and U9288 (N_9288,N_6260,N_5089);
and U9289 (N_9289,N_5861,N_5158);
nand U9290 (N_9290,N_5083,N_6341);
and U9291 (N_9291,N_5033,N_5472);
and U9292 (N_9292,N_5093,N_6746);
and U9293 (N_9293,N_5558,N_6830);
or U9294 (N_9294,N_5210,N_6846);
nor U9295 (N_9295,N_5196,N_5297);
and U9296 (N_9296,N_6801,N_5036);
nor U9297 (N_9297,N_7464,N_5926);
or U9298 (N_9298,N_6729,N_5316);
or U9299 (N_9299,N_6719,N_7105);
and U9300 (N_9300,N_6871,N_6218);
nand U9301 (N_9301,N_6229,N_6275);
nor U9302 (N_9302,N_6002,N_7242);
nor U9303 (N_9303,N_7439,N_6076);
nor U9304 (N_9304,N_5930,N_5450);
nand U9305 (N_9305,N_6721,N_6958);
or U9306 (N_9306,N_6459,N_5199);
nor U9307 (N_9307,N_6955,N_6922);
or U9308 (N_9308,N_5043,N_5008);
and U9309 (N_9309,N_5973,N_6175);
nand U9310 (N_9310,N_5972,N_5961);
and U9311 (N_9311,N_5457,N_5518);
or U9312 (N_9312,N_7480,N_6503);
or U9313 (N_9313,N_7130,N_6143);
nor U9314 (N_9314,N_6027,N_6479);
nand U9315 (N_9315,N_5096,N_7277);
or U9316 (N_9316,N_6895,N_6080);
nor U9317 (N_9317,N_6002,N_6086);
nor U9318 (N_9318,N_6939,N_5510);
and U9319 (N_9319,N_5947,N_5305);
nor U9320 (N_9320,N_7497,N_5490);
and U9321 (N_9321,N_5826,N_6332);
or U9322 (N_9322,N_6448,N_5662);
and U9323 (N_9323,N_5339,N_5603);
or U9324 (N_9324,N_7361,N_5832);
nand U9325 (N_9325,N_5318,N_7307);
or U9326 (N_9326,N_6336,N_7278);
nor U9327 (N_9327,N_6250,N_6659);
or U9328 (N_9328,N_5171,N_6518);
nand U9329 (N_9329,N_7016,N_6041);
nand U9330 (N_9330,N_7286,N_5532);
nor U9331 (N_9331,N_5788,N_6385);
nor U9332 (N_9332,N_5062,N_6233);
nor U9333 (N_9333,N_6646,N_6702);
nand U9334 (N_9334,N_6542,N_6685);
or U9335 (N_9335,N_5799,N_5603);
nand U9336 (N_9336,N_6749,N_6854);
nor U9337 (N_9337,N_5561,N_6397);
nand U9338 (N_9338,N_6198,N_5968);
nand U9339 (N_9339,N_5154,N_6910);
nand U9340 (N_9340,N_5886,N_5336);
nand U9341 (N_9341,N_6714,N_5345);
nand U9342 (N_9342,N_7103,N_6040);
nand U9343 (N_9343,N_5613,N_6169);
nand U9344 (N_9344,N_5982,N_5379);
nand U9345 (N_9345,N_6757,N_6916);
or U9346 (N_9346,N_6911,N_6433);
nor U9347 (N_9347,N_6481,N_7401);
or U9348 (N_9348,N_7200,N_6075);
nor U9349 (N_9349,N_6381,N_5130);
and U9350 (N_9350,N_6957,N_6010);
and U9351 (N_9351,N_6218,N_6913);
or U9352 (N_9352,N_6686,N_6797);
nor U9353 (N_9353,N_7280,N_7282);
nor U9354 (N_9354,N_5283,N_7244);
nand U9355 (N_9355,N_5780,N_7490);
or U9356 (N_9356,N_5267,N_5520);
and U9357 (N_9357,N_5163,N_6024);
and U9358 (N_9358,N_5960,N_5691);
xnor U9359 (N_9359,N_5951,N_5131);
and U9360 (N_9360,N_6298,N_5602);
nor U9361 (N_9361,N_5582,N_7492);
nor U9362 (N_9362,N_5273,N_5581);
nor U9363 (N_9363,N_5917,N_6498);
or U9364 (N_9364,N_7116,N_6897);
or U9365 (N_9365,N_6420,N_6049);
or U9366 (N_9366,N_5090,N_5213);
or U9367 (N_9367,N_5660,N_6504);
or U9368 (N_9368,N_6303,N_7383);
nand U9369 (N_9369,N_5965,N_7050);
and U9370 (N_9370,N_6794,N_5642);
nor U9371 (N_9371,N_6837,N_5320);
and U9372 (N_9372,N_7462,N_6176);
nor U9373 (N_9373,N_5918,N_5793);
or U9374 (N_9374,N_5629,N_6419);
nand U9375 (N_9375,N_6137,N_7361);
nor U9376 (N_9376,N_5109,N_6576);
nor U9377 (N_9377,N_5534,N_5441);
nand U9378 (N_9378,N_5349,N_5320);
or U9379 (N_9379,N_6591,N_5167);
nand U9380 (N_9380,N_7111,N_7408);
nor U9381 (N_9381,N_5581,N_5434);
nand U9382 (N_9382,N_5296,N_7174);
nand U9383 (N_9383,N_5122,N_6706);
or U9384 (N_9384,N_5966,N_7402);
xnor U9385 (N_9385,N_7066,N_5141);
nand U9386 (N_9386,N_7360,N_5477);
nor U9387 (N_9387,N_6164,N_6868);
nand U9388 (N_9388,N_5061,N_5553);
nor U9389 (N_9389,N_6089,N_5330);
nor U9390 (N_9390,N_6568,N_6116);
nor U9391 (N_9391,N_7275,N_7036);
nor U9392 (N_9392,N_5912,N_5778);
and U9393 (N_9393,N_5523,N_5039);
and U9394 (N_9394,N_6059,N_7264);
nor U9395 (N_9395,N_6215,N_5297);
nor U9396 (N_9396,N_5931,N_6212);
or U9397 (N_9397,N_7183,N_6281);
nand U9398 (N_9398,N_7026,N_5659);
and U9399 (N_9399,N_6969,N_5341);
and U9400 (N_9400,N_6779,N_5327);
nor U9401 (N_9401,N_5109,N_6442);
nor U9402 (N_9402,N_5971,N_6667);
nor U9403 (N_9403,N_5144,N_6594);
nand U9404 (N_9404,N_7469,N_5280);
and U9405 (N_9405,N_5070,N_7027);
nand U9406 (N_9406,N_6319,N_7351);
and U9407 (N_9407,N_6112,N_5539);
nand U9408 (N_9408,N_7306,N_7163);
nand U9409 (N_9409,N_5591,N_5323);
nor U9410 (N_9410,N_5166,N_6438);
nor U9411 (N_9411,N_6836,N_7218);
and U9412 (N_9412,N_5300,N_6964);
nor U9413 (N_9413,N_6286,N_6172);
and U9414 (N_9414,N_6211,N_6574);
or U9415 (N_9415,N_6079,N_5415);
nand U9416 (N_9416,N_6611,N_5836);
nor U9417 (N_9417,N_6886,N_7087);
nand U9418 (N_9418,N_6842,N_5480);
nand U9419 (N_9419,N_6768,N_5432);
nor U9420 (N_9420,N_6006,N_5543);
nor U9421 (N_9421,N_6144,N_6429);
and U9422 (N_9422,N_7318,N_5534);
or U9423 (N_9423,N_7097,N_5406);
or U9424 (N_9424,N_6366,N_5995);
or U9425 (N_9425,N_7443,N_6508);
or U9426 (N_9426,N_5951,N_6870);
or U9427 (N_9427,N_5938,N_6526);
nor U9428 (N_9428,N_6965,N_6388);
and U9429 (N_9429,N_5562,N_5075);
and U9430 (N_9430,N_6169,N_5460);
and U9431 (N_9431,N_6960,N_7217);
nor U9432 (N_9432,N_5764,N_5835);
and U9433 (N_9433,N_5327,N_6010);
nand U9434 (N_9434,N_6228,N_5364);
nand U9435 (N_9435,N_5414,N_6839);
nand U9436 (N_9436,N_7193,N_7278);
nand U9437 (N_9437,N_6980,N_5961);
and U9438 (N_9438,N_7477,N_5353);
nand U9439 (N_9439,N_6423,N_6951);
nand U9440 (N_9440,N_6839,N_5589);
and U9441 (N_9441,N_5342,N_6517);
or U9442 (N_9442,N_6546,N_5766);
or U9443 (N_9443,N_5355,N_6697);
nand U9444 (N_9444,N_7319,N_5295);
nor U9445 (N_9445,N_5358,N_6137);
or U9446 (N_9446,N_6263,N_6802);
nor U9447 (N_9447,N_7161,N_7271);
or U9448 (N_9448,N_6853,N_6292);
nor U9449 (N_9449,N_7489,N_6071);
nor U9450 (N_9450,N_7195,N_5889);
nor U9451 (N_9451,N_6034,N_7401);
nor U9452 (N_9452,N_5192,N_6477);
nor U9453 (N_9453,N_6210,N_6262);
or U9454 (N_9454,N_7374,N_5731);
or U9455 (N_9455,N_5870,N_6234);
nor U9456 (N_9456,N_7144,N_5662);
and U9457 (N_9457,N_5661,N_6215);
nor U9458 (N_9458,N_7141,N_6896);
nand U9459 (N_9459,N_5967,N_6807);
or U9460 (N_9460,N_5254,N_5068);
nor U9461 (N_9461,N_6945,N_6715);
or U9462 (N_9462,N_6005,N_5957);
and U9463 (N_9463,N_7086,N_5401);
and U9464 (N_9464,N_5167,N_5908);
or U9465 (N_9465,N_5735,N_6507);
nor U9466 (N_9466,N_6556,N_7415);
or U9467 (N_9467,N_5341,N_6928);
or U9468 (N_9468,N_5493,N_6350);
or U9469 (N_9469,N_6071,N_5930);
and U9470 (N_9470,N_5278,N_5820);
and U9471 (N_9471,N_6135,N_6155);
or U9472 (N_9472,N_6300,N_6154);
nor U9473 (N_9473,N_5077,N_7320);
nand U9474 (N_9474,N_5910,N_5204);
and U9475 (N_9475,N_7299,N_5964);
nor U9476 (N_9476,N_6360,N_7243);
xor U9477 (N_9477,N_5747,N_7083);
nor U9478 (N_9478,N_7375,N_6931);
nand U9479 (N_9479,N_5134,N_5463);
and U9480 (N_9480,N_5664,N_5625);
nand U9481 (N_9481,N_7410,N_7257);
or U9482 (N_9482,N_7225,N_5735);
or U9483 (N_9483,N_6987,N_5701);
or U9484 (N_9484,N_5067,N_5177);
nand U9485 (N_9485,N_6863,N_5417);
and U9486 (N_9486,N_6290,N_7136);
nand U9487 (N_9487,N_5472,N_5523);
nor U9488 (N_9488,N_6665,N_6203);
and U9489 (N_9489,N_5249,N_5531);
nor U9490 (N_9490,N_7126,N_6670);
or U9491 (N_9491,N_7001,N_5087);
nand U9492 (N_9492,N_6794,N_7447);
nor U9493 (N_9493,N_6903,N_7222);
and U9494 (N_9494,N_5391,N_5176);
nor U9495 (N_9495,N_6312,N_6453);
nand U9496 (N_9496,N_6078,N_6253);
nand U9497 (N_9497,N_7265,N_5203);
nor U9498 (N_9498,N_5643,N_5746);
nand U9499 (N_9499,N_5008,N_5417);
nor U9500 (N_9500,N_5982,N_6559);
and U9501 (N_9501,N_5621,N_5986);
and U9502 (N_9502,N_5748,N_6537);
nand U9503 (N_9503,N_6812,N_5142);
and U9504 (N_9504,N_7256,N_5930);
nand U9505 (N_9505,N_6307,N_6230);
and U9506 (N_9506,N_6909,N_5240);
or U9507 (N_9507,N_7206,N_7154);
nand U9508 (N_9508,N_5872,N_5993);
and U9509 (N_9509,N_6547,N_5896);
nand U9510 (N_9510,N_6614,N_5643);
or U9511 (N_9511,N_6056,N_6787);
and U9512 (N_9512,N_6349,N_7367);
and U9513 (N_9513,N_6340,N_5557);
and U9514 (N_9514,N_6316,N_5959);
nor U9515 (N_9515,N_6878,N_7317);
or U9516 (N_9516,N_6309,N_6315);
xor U9517 (N_9517,N_7067,N_6976);
nor U9518 (N_9518,N_6564,N_5696);
and U9519 (N_9519,N_7396,N_6176);
nand U9520 (N_9520,N_5098,N_7192);
nand U9521 (N_9521,N_5036,N_5785);
nand U9522 (N_9522,N_5544,N_5636);
nand U9523 (N_9523,N_5377,N_7280);
or U9524 (N_9524,N_6260,N_6870);
nor U9525 (N_9525,N_5906,N_6465);
or U9526 (N_9526,N_5863,N_5662);
or U9527 (N_9527,N_6295,N_6448);
nor U9528 (N_9528,N_5890,N_5106);
nand U9529 (N_9529,N_5502,N_5120);
and U9530 (N_9530,N_5144,N_5446);
nand U9531 (N_9531,N_6288,N_5600);
nor U9532 (N_9532,N_5444,N_7441);
xor U9533 (N_9533,N_5039,N_5205);
or U9534 (N_9534,N_5253,N_6617);
and U9535 (N_9535,N_5300,N_7381);
nor U9536 (N_9536,N_5724,N_6648);
nand U9537 (N_9537,N_5850,N_6529);
nor U9538 (N_9538,N_5456,N_6492);
and U9539 (N_9539,N_5936,N_6821);
and U9540 (N_9540,N_7268,N_6147);
or U9541 (N_9541,N_5617,N_7400);
and U9542 (N_9542,N_6094,N_6840);
or U9543 (N_9543,N_7295,N_5453);
and U9544 (N_9544,N_5337,N_5299);
and U9545 (N_9545,N_5813,N_6950);
or U9546 (N_9546,N_7295,N_6677);
nand U9547 (N_9547,N_6740,N_6446);
nand U9548 (N_9548,N_5864,N_6542);
nor U9549 (N_9549,N_5562,N_6618);
and U9550 (N_9550,N_6324,N_6477);
or U9551 (N_9551,N_7122,N_6495);
and U9552 (N_9552,N_5488,N_5350);
nand U9553 (N_9553,N_5286,N_5839);
xor U9554 (N_9554,N_7481,N_5269);
nor U9555 (N_9555,N_6139,N_5052);
or U9556 (N_9556,N_5818,N_6950);
or U9557 (N_9557,N_5641,N_5754);
nand U9558 (N_9558,N_6574,N_7268);
nor U9559 (N_9559,N_7256,N_5987);
nand U9560 (N_9560,N_5888,N_5241);
or U9561 (N_9561,N_7284,N_6901);
nor U9562 (N_9562,N_6762,N_6298);
or U9563 (N_9563,N_6355,N_6440);
nor U9564 (N_9564,N_5478,N_6228);
nor U9565 (N_9565,N_6998,N_5992);
and U9566 (N_9566,N_5893,N_5615);
nor U9567 (N_9567,N_7213,N_5425);
nor U9568 (N_9568,N_5281,N_5280);
xnor U9569 (N_9569,N_5536,N_6654);
or U9570 (N_9570,N_5830,N_7093);
or U9571 (N_9571,N_6435,N_6786);
nor U9572 (N_9572,N_5833,N_6290);
nand U9573 (N_9573,N_6939,N_5483);
and U9574 (N_9574,N_7071,N_6190);
nor U9575 (N_9575,N_5004,N_5271);
or U9576 (N_9576,N_6659,N_6571);
or U9577 (N_9577,N_5285,N_6442);
nand U9578 (N_9578,N_5744,N_5998);
or U9579 (N_9579,N_5890,N_6731);
and U9580 (N_9580,N_7044,N_6837);
and U9581 (N_9581,N_7250,N_6109);
or U9582 (N_9582,N_7179,N_5631);
and U9583 (N_9583,N_5293,N_5559);
or U9584 (N_9584,N_5342,N_7032);
nor U9585 (N_9585,N_5720,N_7089);
or U9586 (N_9586,N_7220,N_5243);
and U9587 (N_9587,N_5698,N_6371);
nor U9588 (N_9588,N_6249,N_7091);
and U9589 (N_9589,N_5216,N_5245);
and U9590 (N_9590,N_6112,N_7398);
nand U9591 (N_9591,N_5526,N_5437);
or U9592 (N_9592,N_7392,N_5012);
or U9593 (N_9593,N_5278,N_7203);
or U9594 (N_9594,N_5775,N_5509);
and U9595 (N_9595,N_6463,N_5205);
nand U9596 (N_9596,N_6070,N_7276);
nand U9597 (N_9597,N_5127,N_7472);
nand U9598 (N_9598,N_5641,N_5475);
nand U9599 (N_9599,N_6298,N_5542);
nor U9600 (N_9600,N_6168,N_6302);
or U9601 (N_9601,N_7041,N_6822);
nor U9602 (N_9602,N_5916,N_5236);
nand U9603 (N_9603,N_6214,N_6796);
nand U9604 (N_9604,N_6160,N_6424);
nand U9605 (N_9605,N_7417,N_7470);
nor U9606 (N_9606,N_6697,N_6338);
or U9607 (N_9607,N_6431,N_6454);
and U9608 (N_9608,N_5492,N_5316);
nor U9609 (N_9609,N_5434,N_5049);
or U9610 (N_9610,N_7012,N_5291);
and U9611 (N_9611,N_5945,N_5249);
or U9612 (N_9612,N_5416,N_6262);
nor U9613 (N_9613,N_5464,N_5654);
nor U9614 (N_9614,N_7029,N_6041);
nor U9615 (N_9615,N_5737,N_6729);
xor U9616 (N_9616,N_6667,N_7375);
and U9617 (N_9617,N_5202,N_7260);
xnor U9618 (N_9618,N_6410,N_5725);
or U9619 (N_9619,N_7053,N_5325);
or U9620 (N_9620,N_6407,N_7060);
nand U9621 (N_9621,N_5193,N_5204);
or U9622 (N_9622,N_5773,N_6119);
nor U9623 (N_9623,N_5918,N_5323);
and U9624 (N_9624,N_6938,N_7333);
or U9625 (N_9625,N_5042,N_7102);
or U9626 (N_9626,N_5584,N_5939);
nand U9627 (N_9627,N_6941,N_5174);
or U9628 (N_9628,N_6409,N_5222);
nand U9629 (N_9629,N_5691,N_5549);
and U9630 (N_9630,N_5044,N_5744);
or U9631 (N_9631,N_6109,N_7281);
and U9632 (N_9632,N_6909,N_5692);
nor U9633 (N_9633,N_6314,N_6501);
nor U9634 (N_9634,N_6960,N_6332);
and U9635 (N_9635,N_5490,N_5273);
nor U9636 (N_9636,N_6969,N_6971);
nor U9637 (N_9637,N_6161,N_6826);
or U9638 (N_9638,N_6611,N_7103);
or U9639 (N_9639,N_6566,N_6556);
nand U9640 (N_9640,N_6654,N_7045);
nand U9641 (N_9641,N_6973,N_6576);
nand U9642 (N_9642,N_6759,N_5995);
nor U9643 (N_9643,N_6941,N_5573);
and U9644 (N_9644,N_5770,N_6856);
nand U9645 (N_9645,N_5517,N_5188);
and U9646 (N_9646,N_5025,N_6491);
nor U9647 (N_9647,N_5775,N_6347);
nor U9648 (N_9648,N_5186,N_6913);
or U9649 (N_9649,N_6993,N_7016);
or U9650 (N_9650,N_5603,N_5123);
nand U9651 (N_9651,N_7267,N_6969);
and U9652 (N_9652,N_6143,N_5567);
nand U9653 (N_9653,N_5214,N_5638);
nor U9654 (N_9654,N_5202,N_6784);
nand U9655 (N_9655,N_6300,N_6523);
nand U9656 (N_9656,N_6112,N_7373);
nand U9657 (N_9657,N_6808,N_7115);
and U9658 (N_9658,N_7361,N_7346);
nand U9659 (N_9659,N_7423,N_6988);
and U9660 (N_9660,N_6426,N_5238);
nand U9661 (N_9661,N_6776,N_5627);
nor U9662 (N_9662,N_5044,N_6255);
nand U9663 (N_9663,N_6238,N_5209);
and U9664 (N_9664,N_6099,N_5721);
nor U9665 (N_9665,N_6576,N_5222);
or U9666 (N_9666,N_5961,N_6982);
or U9667 (N_9667,N_5950,N_6908);
nor U9668 (N_9668,N_7082,N_7432);
and U9669 (N_9669,N_5818,N_7140);
nor U9670 (N_9670,N_7286,N_5242);
nor U9671 (N_9671,N_6300,N_5569);
nand U9672 (N_9672,N_7349,N_6235);
and U9673 (N_9673,N_5590,N_5072);
and U9674 (N_9674,N_5257,N_6525);
nor U9675 (N_9675,N_5114,N_7202);
nand U9676 (N_9676,N_5519,N_5748);
nor U9677 (N_9677,N_5465,N_6957);
nand U9678 (N_9678,N_5013,N_6224);
nor U9679 (N_9679,N_5883,N_6476);
nor U9680 (N_9680,N_5915,N_7261);
or U9681 (N_9681,N_5927,N_6110);
or U9682 (N_9682,N_5431,N_5128);
nand U9683 (N_9683,N_6286,N_6511);
nor U9684 (N_9684,N_6444,N_6588);
and U9685 (N_9685,N_5359,N_6441);
nor U9686 (N_9686,N_6727,N_6386);
or U9687 (N_9687,N_5940,N_7438);
or U9688 (N_9688,N_5339,N_5193);
nand U9689 (N_9689,N_6671,N_7478);
and U9690 (N_9690,N_5668,N_5552);
or U9691 (N_9691,N_7463,N_6466);
and U9692 (N_9692,N_6937,N_6376);
nor U9693 (N_9693,N_7390,N_5891);
and U9694 (N_9694,N_5767,N_5265);
and U9695 (N_9695,N_6330,N_5102);
nand U9696 (N_9696,N_6430,N_6216);
or U9697 (N_9697,N_7410,N_7330);
or U9698 (N_9698,N_7083,N_5560);
and U9699 (N_9699,N_5995,N_6923);
nand U9700 (N_9700,N_6006,N_6462);
nor U9701 (N_9701,N_6142,N_6601);
and U9702 (N_9702,N_5127,N_6208);
or U9703 (N_9703,N_7420,N_7170);
and U9704 (N_9704,N_6569,N_6341);
nor U9705 (N_9705,N_7114,N_7417);
nand U9706 (N_9706,N_6933,N_5567);
nor U9707 (N_9707,N_5324,N_5984);
nand U9708 (N_9708,N_5777,N_7059);
nor U9709 (N_9709,N_5352,N_7149);
nor U9710 (N_9710,N_5413,N_7014);
and U9711 (N_9711,N_7289,N_7085);
or U9712 (N_9712,N_5418,N_5646);
and U9713 (N_9713,N_5756,N_5920);
and U9714 (N_9714,N_6524,N_6299);
and U9715 (N_9715,N_7383,N_6481);
and U9716 (N_9716,N_5583,N_7163);
and U9717 (N_9717,N_5829,N_5374);
nand U9718 (N_9718,N_5777,N_7017);
nor U9719 (N_9719,N_6768,N_5824);
or U9720 (N_9720,N_6476,N_7392);
nand U9721 (N_9721,N_5719,N_5064);
and U9722 (N_9722,N_6502,N_6637);
or U9723 (N_9723,N_6232,N_6326);
nand U9724 (N_9724,N_5417,N_6184);
nand U9725 (N_9725,N_7047,N_6184);
and U9726 (N_9726,N_7254,N_5795);
and U9727 (N_9727,N_5521,N_7105);
xor U9728 (N_9728,N_5831,N_6501);
nand U9729 (N_9729,N_6296,N_6963);
nor U9730 (N_9730,N_6791,N_6190);
nand U9731 (N_9731,N_6828,N_6626);
or U9732 (N_9732,N_5120,N_5418);
nand U9733 (N_9733,N_6529,N_6397);
and U9734 (N_9734,N_6299,N_5822);
and U9735 (N_9735,N_6998,N_5514);
or U9736 (N_9736,N_7147,N_6693);
nand U9737 (N_9737,N_6869,N_5425);
and U9738 (N_9738,N_5889,N_7267);
or U9739 (N_9739,N_5552,N_6591);
or U9740 (N_9740,N_5537,N_5824);
and U9741 (N_9741,N_6921,N_5322);
nor U9742 (N_9742,N_5111,N_6788);
or U9743 (N_9743,N_5986,N_7291);
and U9744 (N_9744,N_5886,N_6776);
nor U9745 (N_9745,N_6476,N_6068);
nor U9746 (N_9746,N_7359,N_6957);
nand U9747 (N_9747,N_7374,N_6121);
and U9748 (N_9748,N_6297,N_5851);
or U9749 (N_9749,N_5671,N_5090);
nor U9750 (N_9750,N_6539,N_7391);
nor U9751 (N_9751,N_6546,N_5204);
nor U9752 (N_9752,N_5720,N_5062);
or U9753 (N_9753,N_5495,N_5925);
and U9754 (N_9754,N_6770,N_6877);
and U9755 (N_9755,N_5764,N_6756);
and U9756 (N_9756,N_6344,N_5673);
and U9757 (N_9757,N_5251,N_5703);
or U9758 (N_9758,N_6495,N_6370);
nand U9759 (N_9759,N_6933,N_7095);
nand U9760 (N_9760,N_5086,N_7129);
or U9761 (N_9761,N_6304,N_6743);
and U9762 (N_9762,N_7156,N_7261);
nand U9763 (N_9763,N_6073,N_6400);
nor U9764 (N_9764,N_5515,N_6194);
nor U9765 (N_9765,N_5579,N_6486);
nor U9766 (N_9766,N_6234,N_7089);
nor U9767 (N_9767,N_5064,N_6504);
nor U9768 (N_9768,N_6951,N_6634);
nor U9769 (N_9769,N_6792,N_7012);
nand U9770 (N_9770,N_5934,N_5058);
nand U9771 (N_9771,N_7136,N_5762);
and U9772 (N_9772,N_7452,N_5368);
nor U9773 (N_9773,N_7324,N_5547);
nand U9774 (N_9774,N_6320,N_6114);
and U9775 (N_9775,N_5681,N_5116);
nand U9776 (N_9776,N_5114,N_5962);
nand U9777 (N_9777,N_6804,N_7232);
nand U9778 (N_9778,N_5024,N_7220);
and U9779 (N_9779,N_6359,N_7360);
and U9780 (N_9780,N_7413,N_7478);
and U9781 (N_9781,N_6470,N_6637);
or U9782 (N_9782,N_7488,N_5219);
nor U9783 (N_9783,N_5856,N_5131);
and U9784 (N_9784,N_5303,N_5353);
and U9785 (N_9785,N_6097,N_5824);
and U9786 (N_9786,N_5570,N_7277);
nor U9787 (N_9787,N_5974,N_5959);
or U9788 (N_9788,N_5973,N_5780);
nor U9789 (N_9789,N_5391,N_7114);
nor U9790 (N_9790,N_6257,N_5941);
and U9791 (N_9791,N_5248,N_6132);
or U9792 (N_9792,N_5693,N_6206);
or U9793 (N_9793,N_5400,N_7188);
nand U9794 (N_9794,N_5872,N_6166);
nor U9795 (N_9795,N_6373,N_7026);
and U9796 (N_9796,N_7435,N_6219);
nor U9797 (N_9797,N_6787,N_7343);
and U9798 (N_9798,N_5297,N_6361);
nand U9799 (N_9799,N_7032,N_6239);
nand U9800 (N_9800,N_6858,N_5272);
and U9801 (N_9801,N_5820,N_6661);
nand U9802 (N_9802,N_5967,N_7436);
or U9803 (N_9803,N_5607,N_5300);
nand U9804 (N_9804,N_6341,N_6538);
nor U9805 (N_9805,N_7240,N_7480);
nor U9806 (N_9806,N_5855,N_5874);
nand U9807 (N_9807,N_6651,N_5245);
and U9808 (N_9808,N_7416,N_6728);
nand U9809 (N_9809,N_5009,N_7358);
or U9810 (N_9810,N_5427,N_7158);
or U9811 (N_9811,N_6855,N_7441);
or U9812 (N_9812,N_5926,N_6684);
nand U9813 (N_9813,N_5307,N_6015);
and U9814 (N_9814,N_6896,N_6329);
and U9815 (N_9815,N_6891,N_7025);
or U9816 (N_9816,N_5265,N_5591);
and U9817 (N_9817,N_6630,N_6898);
nand U9818 (N_9818,N_6573,N_6103);
nor U9819 (N_9819,N_6910,N_6346);
nand U9820 (N_9820,N_5953,N_6690);
and U9821 (N_9821,N_7222,N_6782);
and U9822 (N_9822,N_6051,N_7011);
nand U9823 (N_9823,N_5737,N_7261);
nand U9824 (N_9824,N_6529,N_7072);
nor U9825 (N_9825,N_5219,N_7361);
nor U9826 (N_9826,N_6852,N_5452);
nor U9827 (N_9827,N_6761,N_7323);
and U9828 (N_9828,N_5811,N_7134);
and U9829 (N_9829,N_5605,N_6049);
and U9830 (N_9830,N_6447,N_6735);
xnor U9831 (N_9831,N_6632,N_6343);
nor U9832 (N_9832,N_5473,N_7213);
and U9833 (N_9833,N_5244,N_5180);
or U9834 (N_9834,N_5662,N_6510);
nand U9835 (N_9835,N_5810,N_7022);
nand U9836 (N_9836,N_6727,N_7479);
nand U9837 (N_9837,N_6780,N_5943);
nor U9838 (N_9838,N_5307,N_5970);
and U9839 (N_9839,N_5807,N_5870);
and U9840 (N_9840,N_7097,N_5907);
and U9841 (N_9841,N_5504,N_6336);
nor U9842 (N_9842,N_6557,N_6291);
and U9843 (N_9843,N_5848,N_5476);
nand U9844 (N_9844,N_5463,N_6402);
and U9845 (N_9845,N_5706,N_6579);
nand U9846 (N_9846,N_7419,N_7176);
and U9847 (N_9847,N_5250,N_6311);
nand U9848 (N_9848,N_7158,N_6621);
nor U9849 (N_9849,N_6157,N_6273);
or U9850 (N_9850,N_6387,N_6229);
or U9851 (N_9851,N_5940,N_5027);
and U9852 (N_9852,N_5074,N_6248);
or U9853 (N_9853,N_6026,N_5421);
nor U9854 (N_9854,N_5447,N_5842);
and U9855 (N_9855,N_6079,N_6148);
or U9856 (N_9856,N_5821,N_5084);
and U9857 (N_9857,N_6151,N_6453);
nor U9858 (N_9858,N_5030,N_6150);
nand U9859 (N_9859,N_5779,N_7008);
nor U9860 (N_9860,N_5190,N_6986);
or U9861 (N_9861,N_5988,N_6838);
nor U9862 (N_9862,N_5220,N_5736);
nor U9863 (N_9863,N_5083,N_6506);
or U9864 (N_9864,N_6458,N_5491);
or U9865 (N_9865,N_7223,N_6488);
nand U9866 (N_9866,N_6430,N_5269);
nand U9867 (N_9867,N_5073,N_5210);
or U9868 (N_9868,N_7018,N_5187);
and U9869 (N_9869,N_5800,N_6982);
and U9870 (N_9870,N_5424,N_5196);
and U9871 (N_9871,N_5007,N_5061);
or U9872 (N_9872,N_6127,N_5818);
nor U9873 (N_9873,N_6413,N_6460);
nand U9874 (N_9874,N_5811,N_6665);
or U9875 (N_9875,N_5296,N_6916);
nand U9876 (N_9876,N_5670,N_6674);
and U9877 (N_9877,N_5920,N_6944);
nor U9878 (N_9878,N_6543,N_6706);
and U9879 (N_9879,N_6025,N_6419);
or U9880 (N_9880,N_5583,N_7037);
nand U9881 (N_9881,N_5193,N_6199);
or U9882 (N_9882,N_6579,N_5133);
or U9883 (N_9883,N_6403,N_6496);
and U9884 (N_9884,N_6287,N_7366);
nor U9885 (N_9885,N_5535,N_6929);
xnor U9886 (N_9886,N_5660,N_6971);
nand U9887 (N_9887,N_6328,N_7332);
or U9888 (N_9888,N_7252,N_7287);
nand U9889 (N_9889,N_7221,N_6698);
nor U9890 (N_9890,N_6357,N_5493);
nand U9891 (N_9891,N_5475,N_6029);
or U9892 (N_9892,N_7452,N_7267);
or U9893 (N_9893,N_6115,N_6815);
nor U9894 (N_9894,N_6134,N_5175);
nand U9895 (N_9895,N_6756,N_6901);
or U9896 (N_9896,N_6005,N_6471);
and U9897 (N_9897,N_5828,N_6571);
nand U9898 (N_9898,N_5770,N_5071);
or U9899 (N_9899,N_7263,N_5653);
xnor U9900 (N_9900,N_5358,N_6547);
nand U9901 (N_9901,N_5546,N_5114);
and U9902 (N_9902,N_6083,N_6604);
and U9903 (N_9903,N_6471,N_5358);
nor U9904 (N_9904,N_6584,N_6692);
and U9905 (N_9905,N_6875,N_7383);
or U9906 (N_9906,N_5344,N_6174);
nor U9907 (N_9907,N_6850,N_6054);
nand U9908 (N_9908,N_6884,N_7134);
nor U9909 (N_9909,N_7103,N_6716);
nand U9910 (N_9910,N_6980,N_5237);
nor U9911 (N_9911,N_6397,N_5030);
nand U9912 (N_9912,N_5836,N_7491);
or U9913 (N_9913,N_7487,N_6521);
nand U9914 (N_9914,N_6864,N_7379);
nand U9915 (N_9915,N_7307,N_6254);
nand U9916 (N_9916,N_7196,N_6529);
or U9917 (N_9917,N_7322,N_6193);
and U9918 (N_9918,N_5910,N_7371);
nand U9919 (N_9919,N_6024,N_6412);
or U9920 (N_9920,N_5286,N_7157);
or U9921 (N_9921,N_7422,N_5903);
nor U9922 (N_9922,N_6798,N_7263);
or U9923 (N_9923,N_6510,N_7348);
or U9924 (N_9924,N_6435,N_6022);
nand U9925 (N_9925,N_5725,N_5754);
nand U9926 (N_9926,N_6045,N_5305);
and U9927 (N_9927,N_6716,N_7221);
nor U9928 (N_9928,N_5898,N_5325);
or U9929 (N_9929,N_6853,N_5104);
and U9930 (N_9930,N_6851,N_5024);
nor U9931 (N_9931,N_6673,N_6702);
and U9932 (N_9932,N_5739,N_6364);
and U9933 (N_9933,N_7375,N_7160);
and U9934 (N_9934,N_6093,N_7025);
nand U9935 (N_9935,N_6301,N_6955);
nand U9936 (N_9936,N_7218,N_5048);
or U9937 (N_9937,N_7272,N_6269);
nand U9938 (N_9938,N_7043,N_5728);
or U9939 (N_9939,N_5256,N_6941);
nand U9940 (N_9940,N_5831,N_7198);
or U9941 (N_9941,N_5094,N_7135);
or U9942 (N_9942,N_6466,N_5256);
nand U9943 (N_9943,N_5402,N_5310);
or U9944 (N_9944,N_6913,N_6161);
or U9945 (N_9945,N_5866,N_5703);
or U9946 (N_9946,N_7163,N_5804);
or U9947 (N_9947,N_5786,N_6914);
or U9948 (N_9948,N_7273,N_7442);
and U9949 (N_9949,N_5846,N_5557);
nand U9950 (N_9950,N_5132,N_5064);
and U9951 (N_9951,N_5718,N_7302);
xnor U9952 (N_9952,N_5639,N_7278);
or U9953 (N_9953,N_5636,N_7497);
and U9954 (N_9954,N_6148,N_7002);
or U9955 (N_9955,N_5616,N_5209);
nand U9956 (N_9956,N_7262,N_6466);
nand U9957 (N_9957,N_7043,N_6188);
and U9958 (N_9958,N_7390,N_5347);
or U9959 (N_9959,N_6591,N_7228);
nor U9960 (N_9960,N_5515,N_6741);
or U9961 (N_9961,N_5751,N_5577);
nand U9962 (N_9962,N_5585,N_6001);
nor U9963 (N_9963,N_5873,N_5915);
or U9964 (N_9964,N_6112,N_5073);
nand U9965 (N_9965,N_7445,N_5686);
and U9966 (N_9966,N_6772,N_5451);
and U9967 (N_9967,N_7033,N_5237);
or U9968 (N_9968,N_6834,N_5288);
and U9969 (N_9969,N_6574,N_5959);
nor U9970 (N_9970,N_5319,N_7077);
and U9971 (N_9971,N_5900,N_6082);
and U9972 (N_9972,N_6786,N_5331);
nand U9973 (N_9973,N_7234,N_6446);
and U9974 (N_9974,N_5770,N_6035);
nand U9975 (N_9975,N_6926,N_6142);
nand U9976 (N_9976,N_5120,N_6563);
or U9977 (N_9977,N_6299,N_6422);
nand U9978 (N_9978,N_6570,N_5681);
nand U9979 (N_9979,N_7255,N_6231);
or U9980 (N_9980,N_7236,N_5267);
and U9981 (N_9981,N_5858,N_6403);
nor U9982 (N_9982,N_5266,N_5445);
and U9983 (N_9983,N_5864,N_5661);
nor U9984 (N_9984,N_6648,N_7001);
nor U9985 (N_9985,N_6964,N_5247);
nand U9986 (N_9986,N_6783,N_6512);
nand U9987 (N_9987,N_6834,N_5699);
nand U9988 (N_9988,N_6032,N_5601);
and U9989 (N_9989,N_6263,N_6632);
nor U9990 (N_9990,N_6439,N_5056);
nand U9991 (N_9991,N_5179,N_7135);
nand U9992 (N_9992,N_6559,N_5129);
and U9993 (N_9993,N_6401,N_5579);
nor U9994 (N_9994,N_6177,N_5853);
and U9995 (N_9995,N_7480,N_5345);
nand U9996 (N_9996,N_5815,N_6150);
nand U9997 (N_9997,N_5926,N_6874);
xor U9998 (N_9998,N_5861,N_5615);
and U9999 (N_9999,N_5385,N_7416);
and UO_0 (O_0,N_9256,N_7957);
and UO_1 (O_1,N_7591,N_8993);
nor UO_2 (O_2,N_9170,N_8901);
nor UO_3 (O_3,N_9777,N_8027);
and UO_4 (O_4,N_9944,N_7815);
nand UO_5 (O_5,N_8018,N_7817);
nand UO_6 (O_6,N_9375,N_8302);
nand UO_7 (O_7,N_8968,N_9175);
or UO_8 (O_8,N_8982,N_8924);
or UO_9 (O_9,N_9756,N_8391);
nand UO_10 (O_10,N_9366,N_8477);
nand UO_11 (O_11,N_8701,N_7663);
and UO_12 (O_12,N_8271,N_9925);
nor UO_13 (O_13,N_8972,N_9966);
or UO_14 (O_14,N_8078,N_7735);
or UO_15 (O_15,N_8292,N_9161);
or UO_16 (O_16,N_9315,N_9746);
nor UO_17 (O_17,N_8570,N_7910);
nand UO_18 (O_18,N_8408,N_8463);
or UO_19 (O_19,N_8455,N_8547);
or UO_20 (O_20,N_9960,N_8709);
or UO_21 (O_21,N_8697,N_8638);
and UO_22 (O_22,N_7792,N_9783);
or UO_23 (O_23,N_7725,N_8702);
nor UO_24 (O_24,N_7516,N_9159);
and UO_25 (O_25,N_9360,N_8413);
nand UO_26 (O_26,N_8025,N_7846);
nor UO_27 (O_27,N_9294,N_7612);
and UO_28 (O_28,N_9290,N_9677);
and UO_29 (O_29,N_8526,N_7970);
nor UO_30 (O_30,N_8171,N_9518);
and UO_31 (O_31,N_7597,N_9621);
nor UO_32 (O_32,N_9338,N_9964);
and UO_33 (O_33,N_9370,N_9114);
and UO_34 (O_34,N_8161,N_7893);
or UO_35 (O_35,N_9619,N_8269);
nand UO_36 (O_36,N_7934,N_9562);
and UO_37 (O_37,N_8783,N_9324);
or UO_38 (O_38,N_7992,N_7944);
or UO_39 (O_39,N_8437,N_8444);
or UO_40 (O_40,N_8263,N_7829);
or UO_41 (O_41,N_8754,N_9646);
or UO_42 (O_42,N_8022,N_8943);
nor UO_43 (O_43,N_8604,N_9647);
nor UO_44 (O_44,N_9005,N_7985);
nand UO_45 (O_45,N_8154,N_9818);
and UO_46 (O_46,N_8106,N_9982);
or UO_47 (O_47,N_8453,N_9631);
nand UO_48 (O_48,N_9716,N_8726);
and UO_49 (O_49,N_9356,N_9786);
nand UO_50 (O_50,N_9549,N_9962);
nand UO_51 (O_51,N_9392,N_8124);
nor UO_52 (O_52,N_9204,N_9140);
nand UO_53 (O_53,N_9916,N_7736);
and UO_54 (O_54,N_9792,N_8258);
or UO_55 (O_55,N_9595,N_7621);
or UO_56 (O_56,N_9116,N_8228);
nor UO_57 (O_57,N_7716,N_9842);
nor UO_58 (O_58,N_9468,N_8693);
or UO_59 (O_59,N_8670,N_7564);
and UO_60 (O_60,N_8435,N_9115);
or UO_61 (O_61,N_8385,N_9267);
or UO_62 (O_62,N_9227,N_7654);
nor UO_63 (O_63,N_8575,N_8946);
nand UO_64 (O_64,N_9914,N_8746);
nand UO_65 (O_65,N_7857,N_9233);
nor UO_66 (O_66,N_8801,N_7835);
nand UO_67 (O_67,N_7898,N_8328);
xnor UO_68 (O_68,N_7974,N_9053);
or UO_69 (O_69,N_9876,N_9734);
nor UO_70 (O_70,N_8997,N_7997);
or UO_71 (O_71,N_9197,N_9093);
nand UO_72 (O_72,N_9440,N_7603);
and UO_73 (O_73,N_7524,N_8777);
or UO_74 (O_74,N_8190,N_8093);
or UO_75 (O_75,N_7780,N_8865);
or UO_76 (O_76,N_9453,N_8793);
nor UO_77 (O_77,N_7783,N_7720);
and UO_78 (O_78,N_7634,N_9515);
and UO_79 (O_79,N_7924,N_9067);
and UO_80 (O_80,N_9046,N_9735);
and UO_81 (O_81,N_8928,N_9903);
and UO_82 (O_82,N_8878,N_7662);
nand UO_83 (O_83,N_9832,N_9456);
and UO_84 (O_84,N_8465,N_9146);
nor UO_85 (O_85,N_7952,N_8316);
nand UO_86 (O_86,N_7682,N_8525);
nor UO_87 (O_87,N_8276,N_8070);
nor UO_88 (O_88,N_9107,N_9537);
and UO_89 (O_89,N_9901,N_8551);
or UO_90 (O_90,N_8239,N_8436);
and UO_91 (O_91,N_9153,N_9286);
and UO_92 (O_92,N_8019,N_9494);
nor UO_93 (O_93,N_8415,N_8198);
or UO_94 (O_94,N_8137,N_8768);
and UO_95 (O_95,N_9345,N_8874);
nor UO_96 (O_96,N_9166,N_8553);
nand UO_97 (O_97,N_9834,N_9889);
nor UO_98 (O_98,N_8935,N_9464);
and UO_99 (O_99,N_7620,N_9433);
xnor UO_100 (O_100,N_7703,N_7672);
and UO_101 (O_101,N_8488,N_8255);
nor UO_102 (O_102,N_7980,N_7750);
nor UO_103 (O_103,N_8936,N_9314);
nor UO_104 (O_104,N_8808,N_9711);
and UO_105 (O_105,N_9241,N_8917);
nand UO_106 (O_106,N_7752,N_8026);
or UO_107 (O_107,N_8744,N_8877);
and UO_108 (O_108,N_8075,N_8049);
nand UO_109 (O_109,N_8994,N_9047);
and UO_110 (O_110,N_8885,N_8405);
or UO_111 (O_111,N_9303,N_8097);
nand UO_112 (O_112,N_9181,N_7978);
nor UO_113 (O_113,N_8466,N_9346);
nor UO_114 (O_114,N_8535,N_9608);
nand UO_115 (O_115,N_9905,N_8967);
nand UO_116 (O_116,N_7791,N_8760);
nand UO_117 (O_117,N_8521,N_8434);
nor UO_118 (O_118,N_7686,N_9763);
nand UO_119 (O_119,N_9132,N_9061);
and UO_120 (O_120,N_8441,N_9831);
nor UO_121 (O_121,N_7950,N_8774);
and UO_122 (O_122,N_9733,N_9576);
and UO_123 (O_123,N_7511,N_9878);
and UO_124 (O_124,N_9369,N_9555);
nand UO_125 (O_125,N_9376,N_8305);
nor UO_126 (O_126,N_9695,N_8473);
nand UO_127 (O_127,N_9623,N_8470);
and UO_128 (O_128,N_7513,N_9069);
nor UO_129 (O_129,N_9134,N_9675);
or UO_130 (O_130,N_7825,N_9242);
or UO_131 (O_131,N_7954,N_7856);
and UO_132 (O_132,N_8146,N_9997);
nand UO_133 (O_133,N_9393,N_7656);
or UO_134 (O_134,N_9498,N_9023);
or UO_135 (O_135,N_7589,N_8445);
nand UO_136 (O_136,N_9796,N_8129);
and UO_137 (O_137,N_9096,N_8736);
and UO_138 (O_138,N_8134,N_8661);
nand UO_139 (O_139,N_9372,N_9450);
nor UO_140 (O_140,N_9015,N_8595);
and UO_141 (O_141,N_8919,N_7531);
and UO_142 (O_142,N_9932,N_7529);
and UO_143 (O_143,N_8794,N_8597);
and UO_144 (O_144,N_8400,N_7776);
nand UO_145 (O_145,N_8791,N_8688);
or UO_146 (O_146,N_8557,N_9036);
nor UO_147 (O_147,N_7623,N_8028);
xor UO_148 (O_148,N_9615,N_8071);
or UO_149 (O_149,N_8867,N_8851);
nor UO_150 (O_150,N_9434,N_9686);
or UO_151 (O_151,N_8663,N_9122);
or UO_152 (O_152,N_8607,N_9682);
nand UO_153 (O_153,N_9766,N_9496);
or UO_154 (O_154,N_9341,N_8576);
nand UO_155 (O_155,N_9165,N_9899);
or UO_156 (O_156,N_9702,N_7811);
and UO_157 (O_157,N_9177,N_9040);
nand UO_158 (O_158,N_7868,N_9416);
or UO_159 (O_159,N_7520,N_7973);
and UO_160 (O_160,N_8889,N_8217);
or UO_161 (O_161,N_9262,N_9541);
nor UO_162 (O_162,N_8428,N_9467);
nor UO_163 (O_163,N_8191,N_7535);
or UO_164 (O_164,N_8962,N_7998);
nor UO_165 (O_165,N_8662,N_8964);
and UO_166 (O_166,N_8121,N_9910);
nor UO_167 (O_167,N_7818,N_8064);
nor UO_168 (O_168,N_9331,N_9632);
nand UO_169 (O_169,N_7912,N_9124);
xnor UO_170 (O_170,N_9748,N_7572);
nand UO_171 (O_171,N_8287,N_8092);
or UO_172 (O_172,N_8817,N_8800);
nand UO_173 (O_173,N_9073,N_9694);
nor UO_174 (O_174,N_8298,N_9004);
or UO_175 (O_175,N_9861,N_9846);
nor UO_176 (O_176,N_7855,N_9239);
nand UO_177 (O_177,N_9034,N_9415);
nand UO_178 (O_178,N_7981,N_8756);
nor UO_179 (O_179,N_9998,N_7707);
or UO_180 (O_180,N_9979,N_9712);
and UO_181 (O_181,N_8925,N_9397);
or UO_182 (O_182,N_8512,N_7645);
or UO_183 (O_183,N_8763,N_9614);
nand UO_184 (O_184,N_7743,N_8762);
or UO_185 (O_185,N_8420,N_8222);
and UO_186 (O_186,N_8723,N_9493);
or UO_187 (O_187,N_9249,N_7918);
and UO_188 (O_188,N_9190,N_8614);
and UO_189 (O_189,N_9176,N_8003);
nand UO_190 (O_190,N_7769,N_9228);
and UO_191 (O_191,N_9143,N_8494);
nor UO_192 (O_192,N_9969,N_9913);
or UO_193 (O_193,N_8355,N_9026);
and UO_194 (O_194,N_9542,N_9007);
or UO_195 (O_195,N_7800,N_7805);
or UO_196 (O_196,N_7674,N_9109);
nor UO_197 (O_197,N_7886,N_8956);
nand UO_198 (O_198,N_8695,N_9984);
nand UO_199 (O_199,N_9081,N_9781);
or UO_200 (O_200,N_8552,N_8087);
nand UO_201 (O_201,N_7861,N_8920);
and UO_202 (O_202,N_7537,N_7779);
and UO_203 (O_203,N_8244,N_9907);
or UO_204 (O_204,N_8755,N_7586);
or UO_205 (O_205,N_9002,N_7814);
and UO_206 (O_206,N_8619,N_7732);
nor UO_207 (O_207,N_9957,N_9798);
nand UO_208 (O_208,N_9250,N_8529);
and UO_209 (O_209,N_9483,N_8496);
or UO_210 (O_210,N_8324,N_8327);
and UO_211 (O_211,N_9764,N_9288);
nor UO_212 (O_212,N_8632,N_8440);
nor UO_213 (O_213,N_7504,N_9856);
nor UO_214 (O_214,N_9025,N_9282);
nor UO_215 (O_215,N_8211,N_9474);
or UO_216 (O_216,N_9429,N_8912);
or UO_217 (O_217,N_9826,N_8480);
or UO_218 (O_218,N_8241,N_8834);
or UO_219 (O_219,N_7566,N_8144);
nor UO_220 (O_220,N_8119,N_8761);
nor UO_221 (O_221,N_9441,N_8074);
nor UO_222 (O_222,N_9355,N_7718);
or UO_223 (O_223,N_8771,N_9155);
or UO_224 (O_224,N_8299,N_8537);
nor UO_225 (O_225,N_8034,N_8242);
nor UO_226 (O_226,N_9509,N_8598);
nand UO_227 (O_227,N_8206,N_8212);
nand UO_228 (O_228,N_8174,N_7554);
nand UO_229 (O_229,N_8564,N_8591);
nor UO_230 (O_230,N_9714,N_9887);
nand UO_231 (O_231,N_9626,N_7657);
nor UO_232 (O_232,N_7770,N_9451);
and UO_233 (O_233,N_8718,N_8665);
nand UO_234 (O_234,N_8220,N_9519);
nand UO_235 (O_235,N_8542,N_9362);
and UO_236 (O_236,N_7648,N_9954);
nand UO_237 (O_237,N_8035,N_9285);
or UO_238 (O_238,N_9755,N_8176);
nor UO_239 (O_239,N_9212,N_9524);
nand UO_240 (O_240,N_9521,N_8293);
and UO_241 (O_241,N_8231,N_9062);
or UO_242 (O_242,N_8296,N_8630);
nor UO_243 (O_243,N_8417,N_9545);
nand UO_244 (O_244,N_9209,N_9996);
or UO_245 (O_245,N_8959,N_8030);
nor UO_246 (O_246,N_8281,N_7570);
nor UO_247 (O_247,N_8448,N_7806);
or UO_248 (O_248,N_9784,N_9948);
and UO_249 (O_249,N_8843,N_8085);
or UO_250 (O_250,N_9084,N_8876);
or UO_251 (O_251,N_7804,N_8310);
and UO_252 (O_252,N_7842,N_8905);
and UO_253 (O_253,N_8479,N_9971);
nand UO_254 (O_254,N_9191,N_8080);
nand UO_255 (O_255,N_8061,N_7667);
nor UO_256 (O_256,N_9071,N_8921);
and UO_257 (O_257,N_7911,N_8010);
nand UO_258 (O_258,N_9550,N_8402);
nor UO_259 (O_259,N_8548,N_9037);
nor UO_260 (O_260,N_7797,N_9789);
nand UO_261 (O_261,N_8066,N_8857);
nor UO_262 (O_262,N_9157,N_7712);
nor UO_263 (O_263,N_7534,N_9877);
nand UO_264 (O_264,N_7896,N_9504);
and UO_265 (O_265,N_8374,N_9928);
and UO_266 (O_266,N_8950,N_9131);
nand UO_267 (O_267,N_9339,N_7757);
nand UO_268 (O_268,N_8045,N_8043);
nor UO_269 (O_269,N_8472,N_8165);
or UO_270 (O_270,N_9724,N_8218);
nor UO_271 (O_271,N_8179,N_8397);
nand UO_272 (O_272,N_9893,N_9237);
nor UO_273 (O_273,N_9946,N_9909);
nor UO_274 (O_274,N_9231,N_8699);
and UO_275 (O_275,N_8136,N_9216);
and UO_276 (O_276,N_8563,N_8724);
nor UO_277 (O_277,N_7899,N_8303);
and UO_278 (O_278,N_9730,N_9649);
and UO_279 (O_279,N_8544,N_9323);
and UO_280 (O_280,N_9029,N_9731);
nand UO_281 (O_281,N_8795,N_9880);
or UO_282 (O_282,N_8871,N_9717);
nand UO_283 (O_283,N_8516,N_9357);
nor UO_284 (O_284,N_8691,N_8007);
and UO_285 (O_285,N_9300,N_8185);
or UO_286 (O_286,N_8960,N_9317);
nor UO_287 (O_287,N_9548,N_8647);
nand UO_288 (O_288,N_9321,N_7668);
xnor UO_289 (O_289,N_9863,N_8603);
and UO_290 (O_290,N_9021,N_8425);
nor UO_291 (O_291,N_9050,N_9757);
nor UO_292 (O_292,N_7517,N_9651);
nand UO_293 (O_293,N_9059,N_9726);
nand UO_294 (O_294,N_9455,N_8536);
nor UO_295 (O_295,N_8325,N_9691);
or UO_296 (O_296,N_8990,N_7598);
or UO_297 (O_297,N_7945,N_9754);
nor UO_298 (O_298,N_9701,N_7552);
nor UO_299 (O_299,N_8958,N_7715);
or UO_300 (O_300,N_8684,N_7688);
xor UO_301 (O_301,N_8349,N_9927);
nand UO_302 (O_302,N_7580,N_8804);
or UO_303 (O_303,N_7755,N_8622);
and UO_304 (O_304,N_7894,N_9382);
nand UO_305 (O_305,N_9201,N_7664);
or UO_306 (O_306,N_7587,N_7926);
or UO_307 (O_307,N_8615,N_8459);
and UO_308 (O_308,N_8854,N_9475);
nor UO_309 (O_309,N_9703,N_7721);
or UO_310 (O_310,N_7556,N_9874);
or UO_311 (O_311,N_9297,N_8780);
or UO_312 (O_312,N_7938,N_9171);
nand UO_313 (O_313,N_8369,N_7958);
and UO_314 (O_314,N_9400,N_7533);
or UO_315 (O_315,N_9981,N_8449);
nand UO_316 (O_316,N_8214,N_7638);
nand UO_317 (O_317,N_8451,N_7819);
nor UO_318 (O_318,N_7644,N_9813);
or UO_319 (O_319,N_8054,N_7871);
nor UO_320 (O_320,N_8913,N_8083);
or UO_321 (O_321,N_9095,N_8730);
or UO_322 (O_322,N_9926,N_7676);
and UO_323 (O_323,N_7613,N_7508);
nand UO_324 (O_324,N_7710,N_7576);
nand UO_325 (O_325,N_9513,N_8384);
or UO_326 (O_326,N_9525,N_7632);
nand UO_327 (O_327,N_7538,N_8481);
and UO_328 (O_328,N_7851,N_8235);
or UO_329 (O_329,N_8898,N_8133);
nor UO_330 (O_330,N_8099,N_8065);
and UO_331 (O_331,N_9895,N_8351);
nor UO_332 (O_332,N_8584,N_8819);
nand UO_333 (O_333,N_9459,N_8100);
nand UO_334 (O_334,N_8013,N_8923);
or UO_335 (O_335,N_7543,N_8502);
or UO_336 (O_336,N_8633,N_9224);
and UO_337 (O_337,N_9989,N_9318);
and UO_338 (O_338,N_7813,N_8404);
nand UO_339 (O_339,N_8224,N_7585);
and UO_340 (O_340,N_8856,N_9384);
nand UO_341 (O_341,N_9210,N_8954);
xor UO_342 (O_342,N_8585,N_9961);
nor UO_343 (O_343,N_9090,N_9890);
and UO_344 (O_344,N_9501,N_8234);
nor UO_345 (O_345,N_9172,N_8433);
nand UO_346 (O_346,N_7913,N_7775);
nor UO_347 (O_347,N_8862,N_7904);
and UO_348 (O_348,N_9698,N_8411);
nand UO_349 (O_349,N_8414,N_8170);
and UO_350 (O_350,N_9918,N_8478);
or UO_351 (O_351,N_8505,N_9472);
nand UO_352 (O_352,N_9873,N_7975);
and UO_353 (O_353,N_8352,N_9943);
nand UO_354 (O_354,N_7946,N_8860);
nor UO_355 (O_355,N_8875,N_8558);
and UO_356 (O_356,N_7873,N_8519);
or UO_357 (O_357,N_9829,N_9640);
nand UO_358 (O_358,N_8141,N_7820);
or UO_359 (O_359,N_8992,N_8152);
or UO_360 (O_360,N_8458,N_8897);
or UO_361 (O_361,N_8908,N_8456);
and UO_362 (O_362,N_7614,N_7840);
nor UO_363 (O_363,N_8069,N_7879);
and UO_364 (O_364,N_9184,N_8401);
xor UO_365 (O_365,N_7728,N_9923);
and UO_366 (O_366,N_9641,N_8318);
or UO_367 (O_367,N_9130,N_8252);
nor UO_368 (O_368,N_9517,N_8050);
xor UO_369 (O_369,N_9394,N_8983);
nand UO_370 (O_370,N_8423,N_8509);
nand UO_371 (O_371,N_9902,N_8256);
or UO_372 (O_372,N_7746,N_9374);
nor UO_373 (O_373,N_9859,N_8902);
nand UO_374 (O_374,N_8758,N_9092);
nand UO_375 (O_375,N_8005,N_8012);
nor UO_376 (O_376,N_9410,N_9436);
or UO_377 (O_377,N_9666,N_9431);
nor UO_378 (O_378,N_8036,N_9495);
and UO_379 (O_379,N_8601,N_9148);
or UO_380 (O_380,N_8764,N_9558);
and UO_381 (O_381,N_7518,N_9693);
or UO_382 (O_382,N_9739,N_9908);
nor UO_383 (O_383,N_8084,N_7907);
nand UO_384 (O_384,N_9316,N_9919);
or UO_385 (O_385,N_9043,N_9688);
or UO_386 (O_386,N_9728,N_9546);
nor UO_387 (O_387,N_8418,N_9458);
nor UO_388 (O_388,N_9779,N_8940);
nand UO_389 (O_389,N_9591,N_7847);
or UO_390 (O_390,N_8814,N_8679);
and UO_391 (O_391,N_8205,N_8264);
nor UO_392 (O_392,N_9349,N_7699);
or UO_393 (O_393,N_9547,N_8965);
nand UO_394 (O_394,N_8766,N_8787);
nand UO_395 (O_395,N_8500,N_7802);
nor UO_396 (O_396,N_8782,N_8461);
nor UO_397 (O_397,N_7767,N_7774);
nor UO_398 (O_398,N_7906,N_9083);
nand UO_399 (O_399,N_9138,N_7558);
nor UO_400 (O_400,N_8914,N_9729);
nor UO_401 (O_401,N_8107,N_8095);
and UO_402 (O_402,N_7512,N_8979);
nand UO_403 (O_403,N_8356,N_8790);
or UO_404 (O_404,N_9295,N_7850);
nand UO_405 (O_405,N_9635,N_9065);
nor UO_406 (O_406,N_7569,N_8720);
nor UO_407 (O_407,N_9853,N_8491);
nand UO_408 (O_408,N_7714,N_9800);
and UO_409 (O_409,N_9612,N_8117);
and UO_410 (O_410,N_8559,N_8123);
and UO_411 (O_411,N_8254,N_9778);
or UO_412 (O_412,N_7984,N_8672);
and UO_413 (O_413,N_9390,N_8442);
nand UO_414 (O_414,N_7691,N_8202);
or UO_415 (O_415,N_8503,N_8329);
nand UO_416 (O_416,N_7836,N_8499);
nor UO_417 (O_417,N_9139,N_9343);
nor UO_418 (O_418,N_9484,N_8274);
nor UO_419 (O_419,N_9014,N_9643);
or UO_420 (O_420,N_8606,N_8775);
nor UO_421 (O_421,N_8753,N_9674);
and UO_422 (O_422,N_9113,N_9101);
nand UO_423 (O_423,N_9882,N_9975);
nor UO_424 (O_424,N_8053,N_9992);
nand UO_425 (O_425,N_9560,N_8589);
or UO_426 (O_426,N_9312,N_9031);
or UO_427 (O_427,N_9951,N_9775);
and UO_428 (O_428,N_8151,N_7812);
nor UO_429 (O_429,N_9274,N_9770);
or UO_430 (O_430,N_7737,N_9751);
and UO_431 (O_431,N_9543,N_9743);
nor UO_432 (O_432,N_9788,N_9364);
nor UO_433 (O_433,N_7690,N_7961);
nand UO_434 (O_434,N_8246,N_7740);
nand UO_435 (O_435,N_9683,N_9858);
or UO_436 (O_436,N_9767,N_9602);
nor UO_437 (O_437,N_8520,N_8398);
or UO_438 (O_438,N_8197,N_9719);
or UO_439 (O_439,N_9886,N_8098);
nor UO_440 (O_440,N_7649,N_9535);
nand UO_441 (O_441,N_9888,N_7724);
nor UO_442 (O_442,N_9489,N_8781);
and UO_443 (O_443,N_9179,N_8315);
nand UO_444 (O_444,N_8339,N_9950);
and UO_445 (O_445,N_9298,N_8634);
or UO_446 (O_446,N_7573,N_9596);
and UO_447 (O_447,N_9252,N_8784);
nand UO_448 (O_448,N_7921,N_9803);
nand UO_449 (O_449,N_8184,N_8476);
xnor UO_450 (O_450,N_7567,N_8673);
and UO_451 (O_451,N_9446,N_7647);
and UO_452 (O_452,N_9502,N_9055);
nor UO_453 (O_453,N_9263,N_9306);
nor UO_454 (O_454,N_8360,N_9147);
nor UO_455 (O_455,N_7935,N_8227);
and UO_456 (O_456,N_7990,N_7697);
nor UO_457 (O_457,N_8802,N_9968);
or UO_458 (O_458,N_8855,N_9505);
nor UO_459 (O_459,N_8868,N_8706);
and UO_460 (O_460,N_8278,N_9042);
nand UO_461 (O_461,N_7994,N_9532);
nor UO_462 (O_462,N_9884,N_8249);
nand UO_463 (O_463,N_8290,N_9921);
and UO_464 (O_464,N_8565,N_8534);
or UO_465 (O_465,N_8850,N_9830);
and UO_466 (O_466,N_8248,N_8033);
and UO_467 (O_467,N_8739,N_8969);
xor UO_468 (O_468,N_7604,N_8259);
or UO_469 (O_469,N_9277,N_9287);
nand UO_470 (O_470,N_9665,N_8431);
or UO_471 (O_471,N_9636,N_9010);
nand UO_472 (O_472,N_9658,N_9638);
or UO_473 (O_473,N_8826,N_8167);
or UO_474 (O_474,N_8113,N_8906);
nor UO_475 (O_475,N_8307,N_9942);
nand UO_476 (O_476,N_9673,N_9963);
or UO_477 (O_477,N_8926,N_8268);
xnor UO_478 (O_478,N_9354,N_9432);
nor UO_479 (O_479,N_7677,N_7988);
nor UO_480 (O_480,N_8628,N_8737);
nand UO_481 (O_481,N_8980,N_8941);
or UO_482 (O_482,N_9697,N_9747);
and UO_483 (O_483,N_7547,N_8362);
or UO_484 (O_484,N_9955,N_9327);
nand UO_485 (O_485,N_9854,N_8984);
and UO_486 (O_486,N_9388,N_9938);
or UO_487 (O_487,N_9534,N_8389);
nand UO_488 (O_488,N_9885,N_8785);
or UO_489 (O_489,N_7681,N_9707);
nand UO_490 (O_490,N_7982,N_7949);
nor UO_491 (O_491,N_9144,N_9120);
nand UO_492 (O_492,N_9822,N_9852);
or UO_493 (O_493,N_9685,N_7849);
or UO_494 (O_494,N_7793,N_8769);
or UO_495 (O_495,N_8273,N_9089);
and UO_496 (O_496,N_7930,N_8751);
or UO_497 (O_497,N_8068,N_9452);
or UO_498 (O_498,N_8655,N_7919);
nand UO_499 (O_499,N_9564,N_7966);
and UO_500 (O_500,N_9213,N_8443);
or UO_501 (O_501,N_9760,N_8974);
nor UO_502 (O_502,N_9470,N_7749);
nand UO_503 (O_503,N_9308,N_9567);
and UO_504 (O_504,N_9465,N_9395);
nand UO_505 (O_505,N_9389,N_9597);
nand UO_506 (O_506,N_7758,N_8543);
nor UO_507 (O_507,N_9833,N_9396);
and UO_508 (O_508,N_9387,N_9618);
nand UO_509 (O_509,N_7652,N_8393);
xor UO_510 (O_510,N_9361,N_9278);
xnor UO_511 (O_511,N_8947,N_9839);
and UO_512 (O_512,N_9797,N_9229);
nor UO_513 (O_513,N_8710,N_9438);
nor UO_514 (O_514,N_9523,N_7661);
nand UO_515 (O_515,N_8640,N_7734);
and UO_516 (O_516,N_9772,N_8858);
nand UO_517 (O_517,N_9736,N_7897);
nor UO_518 (O_518,N_9230,N_9710);
or UO_519 (O_519,N_9804,N_8951);
and UO_520 (O_520,N_7659,N_8178);
and UO_521 (O_521,N_9108,N_8289);
nand UO_522 (O_522,N_8829,N_9079);
nand UO_523 (O_523,N_9559,N_9644);
nor UO_524 (O_524,N_9569,N_8999);
and UO_525 (O_525,N_8407,N_8890);
xnor UO_526 (O_526,N_9019,N_7548);
nand UO_527 (O_527,N_7553,N_9817);
or UO_528 (O_528,N_7584,N_8122);
xnor UO_529 (O_529,N_8247,N_9573);
nor UO_530 (O_530,N_8600,N_9953);
and UO_531 (O_531,N_7565,N_7713);
nor UO_532 (O_532,N_9566,N_8531);
and UO_533 (O_533,N_7540,N_9299);
nor UO_534 (O_534,N_7601,N_9648);
and UO_535 (O_535,N_9225,N_9825);
nor UO_536 (O_536,N_9154,N_9363);
or UO_537 (O_537,N_8367,N_7727);
nor UO_538 (O_538,N_9232,N_8574);
nand UO_539 (O_539,N_8143,N_7506);
nand UO_540 (O_540,N_8240,N_7925);
and UO_541 (O_541,N_7942,N_9572);
nand UO_542 (O_542,N_8577,N_8142);
and UO_543 (O_543,N_8060,N_8991);
or UO_544 (O_544,N_7561,N_8166);
or UO_545 (O_545,N_8429,N_9582);
nor UO_546 (O_546,N_9087,N_8955);
or UO_547 (O_547,N_7704,N_8588);
nor UO_548 (O_548,N_8326,N_7678);
or UO_549 (O_549,N_8823,N_7848);
nand UO_550 (O_550,N_8009,N_7941);
nand UO_551 (O_551,N_9974,N_8037);
nand UO_552 (O_552,N_9268,N_9266);
nor UO_553 (O_553,N_7844,N_9684);
nand UO_554 (O_554,N_8409,N_9377);
nand UO_555 (O_555,N_9408,N_8546);
and UO_556 (O_556,N_9607,N_9553);
nand UO_557 (O_557,N_8301,N_9912);
or UO_558 (O_558,N_8284,N_8334);
and UO_559 (O_559,N_9808,N_9407);
and UO_560 (O_560,N_8421,N_7505);
nor UO_561 (O_561,N_7568,N_9304);
nor UO_562 (O_562,N_8815,N_8931);
and UO_563 (O_563,N_9012,N_8394);
and UO_564 (O_564,N_8741,N_9127);
and UO_565 (O_565,N_9855,N_9080);
and UO_566 (O_566,N_9845,N_8841);
or UO_567 (O_567,N_9310,N_7937);
nor UO_568 (O_568,N_8900,N_8610);
or UO_569 (O_569,N_7976,N_9347);
nor UO_570 (O_570,N_9473,N_8798);
or UO_571 (O_571,N_8611,N_7995);
or UO_572 (O_572,N_9149,N_9869);
and UO_573 (O_573,N_7999,N_9482);
and UO_574 (O_574,N_8396,N_8139);
nand UO_575 (O_575,N_9843,N_8708);
nor UO_576 (O_576,N_9900,N_8297);
nand UO_577 (O_577,N_9600,N_9413);
and UO_578 (O_578,N_8957,N_7625);
and UO_579 (O_579,N_8116,N_8338);
nor UO_580 (O_580,N_7539,N_8359);
or UO_581 (O_581,N_9732,N_7762);
nand UO_582 (O_582,N_9871,N_9585);
and UO_583 (O_583,N_9780,N_9592);
or UO_584 (O_584,N_8377,N_7655);
nand UO_585 (O_585,N_9851,N_7521);
and UO_586 (O_586,N_7550,N_8742);
or UO_587 (O_587,N_8942,N_7618);
and UO_588 (O_588,N_7541,N_8583);
nor UO_589 (O_589,N_8430,N_8233);
nand UO_590 (O_590,N_7617,N_7519);
or UO_591 (O_591,N_8637,N_7600);
and UO_592 (O_592,N_8562,N_7642);
nor UO_593 (O_593,N_9082,N_9481);
nor UO_594 (O_594,N_8938,N_9758);
nand UO_595 (O_595,N_8617,N_8593);
or UO_596 (O_596,N_7768,N_7731);
nand UO_597 (O_597,N_9412,N_7694);
nand UO_598 (O_598,N_8788,N_8930);
and UO_599 (O_599,N_9516,N_9454);
and UO_600 (O_600,N_8825,N_8091);
and UO_601 (O_601,N_7687,N_9214);
nor UO_602 (O_602,N_7948,N_8530);
or UO_603 (O_603,N_7546,N_8306);
nor UO_604 (O_604,N_8872,N_8830);
and UO_605 (O_605,N_9409,N_8677);
nor UO_606 (O_606,N_8805,N_7522);
nand UO_607 (O_607,N_7581,N_8966);
or UO_608 (O_608,N_8732,N_8545);
nand UO_609 (O_609,N_8734,N_7876);
xnor UO_610 (O_610,N_7593,N_8948);
nand UO_611 (O_611,N_7765,N_8285);
nand UO_612 (O_612,N_9810,N_7964);
and UO_613 (O_613,N_9654,N_8569);
nor UO_614 (O_614,N_8752,N_8474);
nand UO_615 (O_615,N_7863,N_7588);
or UO_616 (O_616,N_8344,N_8376);
or UO_617 (O_617,N_9028,N_8403);
nor UO_618 (O_618,N_7833,N_8852);
nand UO_619 (O_619,N_8267,N_7599);
nand UO_620 (O_620,N_9531,N_8975);
nand UO_621 (O_621,N_9174,N_9422);
nor UO_622 (O_622,N_7900,N_8952);
and UO_623 (O_623,N_9794,N_9709);
nor UO_624 (O_624,N_7549,N_8020);
and UO_625 (O_625,N_9348,N_8177);
nand UO_626 (O_626,N_7875,N_9194);
and UO_627 (O_627,N_9088,N_8067);
or UO_628 (O_628,N_8842,N_8105);
and UO_629 (O_629,N_8438,N_8213);
nand UO_630 (O_630,N_7760,N_8250);
nor UO_631 (O_631,N_8910,N_9275);
or UO_632 (O_632,N_9583,N_9898);
and UO_633 (O_633,N_9617,N_8038);
and UO_634 (O_634,N_8887,N_9243);
or UO_635 (O_635,N_8566,N_9744);
or UO_636 (O_636,N_9344,N_9167);
or UO_637 (O_637,N_8528,N_9258);
nor UO_638 (O_638,N_8147,N_8131);
nand UO_639 (O_639,N_7932,N_8772);
and UO_640 (O_640,N_8015,N_9245);
and UO_641 (O_641,N_9661,N_9049);
and UO_642 (O_642,N_8533,N_8406);
nor UO_643 (O_643,N_8981,N_9575);
or UO_644 (O_644,N_7684,N_9063);
nor UO_645 (O_645,N_8288,N_8809);
nor UO_646 (O_646,N_8039,N_9106);
or UO_647 (O_647,N_7862,N_8668);
nor UO_648 (O_648,N_8884,N_7890);
or UO_649 (O_649,N_9352,N_8811);
nand UO_650 (O_650,N_8643,N_9935);
or UO_651 (O_651,N_8319,N_9958);
nor UO_652 (O_652,N_9151,N_9325);
or UO_653 (O_653,N_9740,N_9561);
nor UO_654 (O_654,N_7641,N_9064);
or UO_655 (O_655,N_9750,N_9983);
nor UO_656 (O_656,N_9203,N_8322);
nor UO_657 (O_657,N_8594,N_8158);
nand UO_658 (O_658,N_9514,N_8703);
nor UO_659 (O_659,N_9520,N_9508);
nand UO_660 (O_660,N_9060,N_9041);
or UO_661 (O_661,N_9580,N_7895);
nand UO_662 (O_662,N_8767,N_8579);
nor UO_663 (O_663,N_9715,N_9491);
and UO_664 (O_664,N_8332,N_8101);
and UO_665 (O_665,N_9152,N_7920);
and UO_666 (O_666,N_8280,N_9398);
nor UO_667 (O_667,N_9189,N_8682);
and UO_668 (O_668,N_7726,N_8698);
and UO_669 (O_669,N_8381,N_8412);
nand UO_670 (O_670,N_7931,N_8199);
nor UO_671 (O_671,N_9264,N_9336);
nor UO_672 (O_672,N_9795,N_9444);
and UO_673 (O_673,N_7739,N_9721);
or UO_674 (O_674,N_8062,N_9044);
and UO_675 (O_675,N_9259,N_7789);
and UO_676 (O_676,N_7754,N_9637);
or UO_677 (O_677,N_9284,N_7616);
xor UO_678 (O_678,N_8282,N_7653);
and UO_679 (O_679,N_7622,N_9430);
nand UO_680 (O_680,N_9411,N_9185);
or UO_681 (O_681,N_8357,N_7808);
and UO_682 (O_682,N_8773,N_7559);
and UO_683 (O_683,N_7670,N_8765);
or UO_684 (O_684,N_8072,N_8094);
and UO_685 (O_685,N_8261,N_9499);
and UO_686 (O_686,N_7689,N_9426);
and UO_687 (O_687,N_8337,N_9811);
and UO_688 (O_688,N_8778,N_8079);
and UO_689 (O_689,N_9329,N_9442);
or UO_690 (O_690,N_7872,N_8426);
nor UO_691 (O_691,N_9727,N_8138);
or UO_692 (O_692,N_7870,N_8846);
nand UO_693 (O_693,N_7650,N_8104);
nand UO_694 (O_694,N_8873,N_9799);
nand UO_695 (O_695,N_7636,N_7979);
nand UO_696 (O_696,N_9659,N_9223);
nor UO_697 (O_697,N_7685,N_8156);
or UO_698 (O_698,N_7673,N_8939);
nor UO_699 (O_699,N_8922,N_7914);
nand UO_700 (O_700,N_9771,N_9183);
or UO_701 (O_701,N_8343,N_9342);
nor UO_702 (O_702,N_9590,N_9460);
nor UO_703 (O_703,N_8148,N_7956);
or UO_704 (O_704,N_8363,N_8024);
nor UO_705 (O_705,N_9018,N_8410);
xor UO_706 (O_706,N_9078,N_8486);
or UO_707 (O_707,N_8721,N_8824);
and UO_708 (O_708,N_9841,N_9479);
nand UO_709 (O_709,N_8891,N_9812);
or UO_710 (O_710,N_9568,N_8489);
and UO_711 (O_711,N_7542,N_8118);
and UO_712 (O_712,N_9696,N_9690);
or UO_713 (O_713,N_7888,N_9386);
and UO_714 (O_714,N_9391,N_8625);
nand UO_715 (O_715,N_8613,N_9949);
and UO_716 (O_716,N_7729,N_7928);
and UO_717 (O_717,N_9445,N_8649);
or UO_718 (O_718,N_8317,N_8193);
and UO_719 (O_719,N_7764,N_9340);
and UO_720 (O_720,N_8230,N_9599);
and UO_721 (O_721,N_8627,N_9035);
nand UO_722 (O_722,N_9419,N_9222);
or UO_723 (O_723,N_8109,N_8669);
and UO_724 (O_724,N_9773,N_8368);
nor UO_725 (O_725,N_8893,N_8432);
and UO_726 (O_726,N_8916,N_9098);
or UO_727 (O_727,N_8493,N_7582);
nor UO_728 (O_728,N_8294,N_8738);
nor UO_729 (O_729,N_8807,N_8056);
or UO_730 (O_730,N_9313,N_9350);
nand UO_731 (O_731,N_7671,N_7903);
nor UO_732 (O_732,N_9689,N_9443);
and UO_733 (O_733,N_7562,N_9126);
and UO_734 (O_734,N_8620,N_8308);
or UO_735 (O_735,N_7852,N_7891);
and UO_736 (O_736,N_9985,N_8386);
xor UO_737 (O_737,N_8446,N_8243);
nand UO_738 (O_738,N_9009,N_7602);
or UO_739 (O_739,N_8475,N_7882);
nor UO_740 (O_740,N_8115,N_9967);
and UO_741 (O_741,N_9202,N_8399);
or UO_742 (O_742,N_8279,N_8631);
and UO_743 (O_743,N_9401,N_8204);
and UO_744 (O_744,N_8717,N_8194);
or UO_745 (O_745,N_8970,N_7741);
or UO_746 (O_746,N_7838,N_7683);
nor UO_747 (O_747,N_7742,N_9669);
and UO_748 (O_748,N_9253,N_7708);
and UO_749 (O_749,N_8680,N_9931);
nor UO_750 (O_750,N_9248,N_8195);
and UO_751 (O_751,N_8978,N_8153);
nand UO_752 (O_752,N_8330,N_8175);
or UO_753 (O_753,N_7960,N_9768);
and UO_754 (O_754,N_7883,N_8485);
nand UO_755 (O_755,N_7747,N_8513);
or UO_756 (O_756,N_8057,N_7853);
or UO_757 (O_757,N_7693,N_9738);
nor UO_758 (O_758,N_9198,N_8295);
nand UO_759 (O_759,N_9381,N_9506);
nor UO_760 (O_760,N_9200,N_9774);
nand UO_761 (O_761,N_8257,N_8870);
or UO_762 (O_762,N_8590,N_9236);
nand UO_763 (O_763,N_9305,N_8382);
nand UO_764 (O_764,N_8309,N_7763);
and UO_765 (O_765,N_8864,N_9112);
nand UO_766 (O_766,N_7501,N_7615);
nor UO_767 (O_767,N_9218,N_8342);
and UO_768 (O_768,N_8008,N_8618);
or UO_769 (O_769,N_9844,N_9296);
nand UO_770 (O_770,N_8102,N_7608);
nor UO_771 (O_771,N_8853,N_9164);
nand UO_772 (O_772,N_8731,N_8652);
and UO_773 (O_773,N_7936,N_9058);
nand UO_774 (O_774,N_9234,N_9604);
and UO_775 (O_775,N_9332,N_9006);
nand UO_776 (O_776,N_9497,N_9420);
nor UO_777 (O_777,N_8770,N_8827);
nand UO_778 (O_778,N_9672,N_7631);
nand UO_779 (O_779,N_9039,N_9883);
and UO_780 (O_780,N_8483,N_9680);
or UO_781 (O_781,N_9838,N_7916);
nor UO_782 (O_782,N_9463,N_9867);
nand UO_783 (O_783,N_9879,N_9471);
nand UO_784 (O_784,N_7590,N_7834);
or UO_785 (O_785,N_8927,N_8651);
nor UO_786 (O_786,N_7733,N_7830);
nor UO_787 (O_787,N_8266,N_9706);
and UO_788 (O_788,N_9207,N_8882);
nor UO_789 (O_789,N_8722,N_7705);
and UO_790 (O_790,N_8869,N_9894);
or UO_791 (O_791,N_8712,N_9605);
and UO_792 (O_792,N_8096,N_8985);
nor UO_793 (O_793,N_8689,N_8286);
and UO_794 (O_794,N_8540,N_7557);
nor UO_795 (O_795,N_9333,N_9368);
or UO_796 (O_796,N_9142,N_7860);
nor UO_797 (O_797,N_8125,N_8110);
nand UO_798 (O_798,N_8861,N_9085);
nand UO_799 (O_799,N_7700,N_8989);
nand UO_800 (O_800,N_9850,N_9868);
or UO_801 (O_801,N_9309,N_8484);
nor UO_802 (O_802,N_9965,N_7771);
and UO_803 (O_803,N_7807,N_7816);
xor UO_804 (O_804,N_8073,N_8886);
nand UO_805 (O_805,N_7788,N_8725);
nor UO_806 (O_806,N_9616,N_9038);
nor UO_807 (O_807,N_8506,N_9097);
nor UO_808 (O_808,N_7963,N_8321);
xnor UO_809 (O_809,N_7983,N_9123);
and UO_810 (O_810,N_8687,N_9301);
or UO_811 (O_811,N_9681,N_9761);
or UO_812 (O_812,N_8987,N_7709);
and UO_813 (O_813,N_7880,N_8727);
nand UO_814 (O_814,N_7555,N_9156);
or UO_815 (O_815,N_9718,N_8892);
and UO_816 (O_816,N_8354,N_9820);
nor UO_817 (O_817,N_8029,N_9540);
nor UO_818 (O_818,N_9100,N_8644);
and UO_819 (O_819,N_7881,N_8498);
or UO_820 (O_820,N_7646,N_7666);
nand UO_821 (O_821,N_8172,N_8032);
and UO_822 (O_822,N_8812,N_9897);
and UO_823 (O_823,N_7629,N_9787);
nor UO_824 (O_824,N_9920,N_9435);
xnor UO_825 (O_825,N_8283,N_8364);
and UO_826 (O_826,N_9586,N_8135);
or UO_827 (O_827,N_9414,N_7675);
or UO_828 (O_828,N_9246,N_9933);
and UO_829 (O_829,N_8311,N_7843);
or UO_830 (O_830,N_8127,N_8998);
nand UO_831 (O_831,N_9173,N_9215);
nor UO_832 (O_832,N_8532,N_8082);
nand UO_833 (O_833,N_8747,N_7692);
nand UO_834 (O_834,N_9461,N_8348);
or UO_835 (O_835,N_9425,N_9815);
or UO_836 (O_836,N_9319,N_8896);
and UO_837 (O_837,N_9941,N_9337);
nor UO_838 (O_838,N_8017,N_8487);
nand UO_839 (O_839,N_7753,N_8238);
nor UO_840 (O_840,N_9424,N_7943);
or UO_841 (O_841,N_8707,N_8888);
or UO_842 (O_842,N_9801,N_8561);
and UO_843 (O_843,N_8648,N_8799);
nand UO_844 (O_844,N_8323,N_7786);
nand UO_845 (O_845,N_9809,N_7523);
nor UO_846 (O_846,N_9490,N_9522);
or UO_847 (O_847,N_8077,N_8658);
and UO_848 (O_848,N_7575,N_9137);
nor UO_849 (O_849,N_9678,N_9819);
and UO_850 (O_850,N_9529,N_9477);
and UO_851 (O_851,N_9652,N_8749);
and UO_852 (O_852,N_7627,N_8346);
nor UO_853 (O_853,N_8859,N_7854);
nor UO_854 (O_854,N_7730,N_8582);
and UO_855 (O_855,N_9977,N_8666);
nand UO_856 (O_856,N_9598,N_9574);
nand UO_857 (O_857,N_8705,N_9986);
or UO_858 (O_858,N_9270,N_8977);
nand UO_859 (O_859,N_9959,N_7766);
and UO_860 (O_860,N_8508,N_9260);
or UO_861 (O_861,N_9466,N_7571);
nor UO_862 (O_862,N_9503,N_7831);
and UO_863 (O_863,N_8743,N_9406);
nor UO_864 (O_864,N_9462,N_7909);
nand UO_865 (O_865,N_9821,N_8664);
and UO_866 (O_866,N_7821,N_7606);
and UO_867 (O_867,N_7658,N_8714);
nand UO_868 (O_868,N_9922,N_9291);
nand UO_869 (O_869,N_9627,N_8656);
nand UO_870 (O_870,N_7971,N_7706);
and UO_871 (O_871,N_8353,N_8729);
and UO_872 (O_872,N_8929,N_8314);
or UO_873 (O_873,N_9128,N_8903);
and UO_874 (O_874,N_9956,N_8149);
nand UO_875 (O_875,N_9423,N_8592);
nor UO_876 (O_876,N_8646,N_7722);
nand UO_877 (O_877,N_9168,N_9528);
nor UO_878 (O_878,N_8208,N_7528);
nor UO_879 (O_879,N_8051,N_7594);
nand UO_880 (O_880,N_9000,N_9358);
nor UO_881 (O_881,N_9917,N_7514);
or UO_882 (O_882,N_7560,N_8055);
and UO_883 (O_883,N_8621,N_7502);
nor UO_884 (O_884,N_8572,N_9995);
or UO_885 (O_885,N_9273,N_8365);
nand UO_886 (O_886,N_8216,N_9102);
and UO_887 (O_887,N_8145,N_9970);
or UO_888 (O_888,N_8011,N_7951);
or UO_889 (O_889,N_9539,N_9380);
nor UO_890 (O_890,N_8126,N_9105);
nor UO_891 (O_891,N_7977,N_8424);
nand UO_892 (O_892,N_9993,N_9526);
nor UO_893 (O_893,N_9133,N_8789);
or UO_894 (O_894,N_8757,N_7832);
nand UO_895 (O_895,N_7643,N_8047);
nor UO_896 (O_896,N_8963,N_9807);
and UO_897 (O_897,N_9280,N_8567);
or UO_898 (O_898,N_8909,N_9713);
nor UO_899 (O_899,N_9662,N_9269);
nand UO_900 (O_900,N_8245,N_9837);
nor UO_901 (O_901,N_8392,N_8629);
and UO_902 (O_902,N_8510,N_8821);
nor UO_903 (O_903,N_7917,N_8378);
nand UO_904 (O_904,N_9244,N_8160);
nor UO_905 (O_905,N_8642,N_7778);
and UO_906 (O_906,N_8945,N_9762);
or UO_907 (O_907,N_8675,N_7665);
nand UO_908 (O_908,N_8608,N_8186);
nor UO_909 (O_909,N_9469,N_7723);
nor UO_910 (O_910,N_7962,N_8223);
or UO_911 (O_911,N_8182,N_9024);
nor UO_912 (O_912,N_7939,N_8659);
and UO_913 (O_913,N_8996,N_9593);
or UO_914 (O_914,N_8275,N_7991);
nand UO_915 (O_915,N_9664,N_7826);
and UO_916 (O_916,N_9782,N_9251);
nand UO_917 (O_917,N_8635,N_7969);
nor UO_918 (O_918,N_8340,N_8626);
nor UO_919 (O_919,N_9074,N_7790);
nand UO_920 (O_920,N_8609,N_7711);
nand UO_921 (O_921,N_9150,N_9973);
nor UO_922 (O_922,N_8336,N_8155);
nor UO_923 (O_923,N_9554,N_8300);
or UO_924 (O_924,N_7507,N_9577);
and UO_925 (O_925,N_8023,N_8740);
and UO_926 (O_926,N_9980,N_9749);
nor UO_927 (O_927,N_9642,N_9988);
or UO_928 (O_928,N_9320,N_8112);
nor UO_929 (O_929,N_8696,N_9584);
nand UO_930 (O_930,N_9011,N_9033);
and UO_931 (O_931,N_9556,N_9500);
or UO_932 (O_932,N_8745,N_8671);
and UO_933 (O_933,N_9565,N_9571);
nand UO_934 (O_934,N_7884,N_9056);
nand UO_935 (O_935,N_9195,N_8000);
nand UO_936 (O_936,N_9952,N_8040);
nor UO_937 (O_937,N_8650,N_9848);
and UO_938 (O_938,N_8568,N_8422);
nand UO_939 (O_939,N_9929,N_8539);
nand UO_940 (O_940,N_8894,N_7837);
or UO_941 (O_941,N_9939,N_8847);
nand UO_942 (O_942,N_9379,N_8210);
and UO_943 (O_943,N_9991,N_8462);
or UO_944 (O_944,N_9220,N_8495);
nor UO_945 (O_945,N_9335,N_9563);
or UO_946 (O_946,N_9418,N_7965);
and UO_947 (O_947,N_9987,N_8232);
and UO_948 (O_948,N_9178,N_9557);
nor UO_949 (O_949,N_9052,N_9639);
nor UO_950 (O_950,N_9570,N_7509);
or UO_951 (O_951,N_8373,N_9551);
nand UO_952 (O_952,N_9492,N_8103);
and UO_953 (O_953,N_8120,N_8716);
or UO_954 (O_954,N_8490,N_8835);
nor UO_955 (O_955,N_8832,N_9129);
nor UO_956 (O_956,N_8918,N_9103);
nand UO_957 (O_957,N_8641,N_7525);
nand UO_958 (O_958,N_8460,N_8719);
or UO_959 (O_959,N_8866,N_8653);
xor UO_960 (O_960,N_8586,N_8953);
nand UO_961 (O_961,N_7609,N_8236);
nand UO_962 (O_962,N_9182,N_9199);
and UO_963 (O_963,N_7719,N_8692);
nand UO_964 (O_964,N_9937,N_8140);
nor UO_965 (O_965,N_8237,N_8587);
or UO_966 (O_966,N_8820,N_9657);
and UO_967 (O_967,N_9704,N_8159);
or UO_968 (O_968,N_9307,N_8674);
or UO_969 (O_969,N_9099,N_8181);
or UO_970 (O_970,N_9587,N_8961);
nand UO_971 (O_971,N_9723,N_8046);
or UO_972 (O_972,N_7596,N_9692);
xor UO_973 (O_973,N_9145,N_8678);
nor UO_974 (O_974,N_9741,N_8380);
nand UO_975 (O_975,N_9622,N_9351);
and UO_976 (O_976,N_9373,N_9947);
nand UO_977 (O_977,N_9186,N_7532);
or UO_978 (O_978,N_8031,N_7515);
or UO_979 (O_979,N_9235,N_8001);
nand UO_980 (O_980,N_9162,N_7624);
and UO_981 (O_981,N_7787,N_8612);
nor UO_982 (O_982,N_7785,N_8189);
and UO_983 (O_983,N_9538,N_9427);
or UO_984 (O_984,N_9022,N_8523);
nor UO_985 (O_985,N_8044,N_9192);
or UO_986 (O_986,N_9330,N_9699);
nor UO_987 (O_987,N_8375,N_8796);
nand UO_988 (O_988,N_7782,N_7803);
nand UO_989 (O_989,N_9257,N_9205);
nand UO_990 (O_990,N_8849,N_9828);
or UO_991 (O_991,N_7526,N_8911);
or UO_992 (O_992,N_7824,N_9480);
and UO_993 (O_993,N_8128,N_7635);
nand UO_994 (O_994,N_9187,N_9875);
xnor UO_995 (O_995,N_9896,N_9045);
and UO_996 (O_996,N_8086,N_8203);
xor UO_997 (O_997,N_7940,N_9670);
nand UO_998 (O_998,N_9048,N_9211);
nand UO_999 (O_999,N_9611,N_7500);
nor UO_1000 (O_1000,N_7579,N_7583);
nor UO_1001 (O_1001,N_8624,N_9016);
nand UO_1002 (O_1002,N_9322,N_8833);
or UO_1003 (O_1003,N_9255,N_9428);
nand UO_1004 (O_1004,N_8331,N_9791);
nand UO_1005 (O_1005,N_8560,N_9589);
nor UO_1006 (O_1006,N_8786,N_9240);
xor UO_1007 (O_1007,N_8130,N_7908);
or UO_1008 (O_1008,N_8879,N_7679);
nand UO_1009 (O_1009,N_8226,N_7794);
and UO_1010 (O_1010,N_8469,N_9579);
nor UO_1011 (O_1011,N_9180,N_8335);
nand UO_1012 (O_1012,N_7545,N_8183);
and UO_1013 (O_1013,N_8556,N_9485);
nand UO_1014 (O_1014,N_9219,N_8599);
nor UO_1015 (O_1015,N_8988,N_9806);
or UO_1016 (O_1016,N_8831,N_8419);
and UO_1017 (O_1017,N_8333,N_9668);
and UO_1018 (O_1018,N_8657,N_8450);
or UO_1019 (O_1019,N_8163,N_8715);
and UO_1020 (O_1020,N_8383,N_7510);
nand UO_1021 (O_1021,N_8168,N_7901);
nor UO_1022 (O_1022,N_9334,N_9417);
or UO_1023 (O_1023,N_9404,N_7987);
nor UO_1024 (O_1024,N_8260,N_9994);
nor UO_1025 (O_1025,N_7633,N_8454);
or UO_1026 (O_1026,N_9072,N_8792);
and UO_1027 (O_1027,N_8304,N_9870);
nand UO_1028 (O_1028,N_8157,N_9008);
or UO_1029 (O_1029,N_7989,N_8277);
nor UO_1030 (O_1030,N_8596,N_9118);
nor UO_1031 (O_1031,N_9872,N_9759);
and UO_1032 (O_1032,N_8219,N_9302);
or UO_1033 (O_1033,N_8522,N_7544);
and UO_1034 (O_1034,N_8748,N_9934);
or UO_1035 (O_1035,N_8200,N_8518);
nand UO_1036 (O_1036,N_8685,N_9753);
nor UO_1037 (O_1037,N_9742,N_9196);
or UO_1038 (O_1038,N_8816,N_8554);
or UO_1039 (O_1039,N_9141,N_8162);
nand UO_1040 (O_1040,N_8623,N_8457);
nor UO_1041 (O_1041,N_8004,N_7756);
or UO_1042 (O_1042,N_9676,N_7902);
or UO_1043 (O_1043,N_9866,N_8899);
nand UO_1044 (O_1044,N_7680,N_8002);
and UO_1045 (O_1045,N_7809,N_7923);
nand UO_1046 (O_1046,N_9110,N_8063);
nor UO_1047 (O_1047,N_8524,N_8452);
and UO_1048 (O_1048,N_8527,N_9990);
nor UO_1049 (O_1049,N_8937,N_9725);
nand UO_1050 (O_1050,N_7865,N_7955);
nor UO_1051 (O_1051,N_9862,N_8973);
nand UO_1052 (O_1052,N_8686,N_9511);
or UO_1053 (O_1053,N_9439,N_9070);
and UO_1054 (O_1054,N_8838,N_9378);
or UO_1055 (O_1055,N_9051,N_7607);
nand UO_1056 (O_1056,N_8253,N_9857);
nor UO_1057 (O_1057,N_9158,N_8700);
nand UO_1058 (O_1058,N_7695,N_9476);
or UO_1059 (O_1059,N_8341,N_9628);
and UO_1060 (O_1060,N_9405,N_8538);
nor UO_1061 (O_1061,N_9001,N_7795);
xor UO_1062 (O_1062,N_7859,N_8395);
or UO_1063 (O_1063,N_7929,N_8016);
nand UO_1064 (O_1064,N_7619,N_9527);
or UO_1065 (O_1065,N_9613,N_7744);
or UO_1066 (O_1066,N_7885,N_9679);
and UO_1067 (O_1067,N_8090,N_8371);
nor UO_1068 (O_1068,N_8501,N_8439);
nor UO_1069 (O_1069,N_8694,N_7577);
or UO_1070 (O_1070,N_8468,N_9208);
nor UO_1071 (O_1071,N_8839,N_7660);
and UO_1072 (O_1072,N_8447,N_8006);
or UO_1073 (O_1073,N_9217,N_8818);
nor UO_1074 (O_1074,N_7738,N_8262);
and UO_1075 (O_1075,N_9594,N_9671);
or UO_1076 (O_1076,N_8482,N_7745);
and UO_1077 (O_1077,N_8192,N_9206);
nand UO_1078 (O_1078,N_7578,N_8907);
nor UO_1079 (O_1079,N_8111,N_9510);
nor UO_1080 (O_1080,N_8511,N_8667);
and UO_1081 (O_1081,N_7823,N_9371);
nand UO_1082 (O_1082,N_8041,N_8836);
nand UO_1083 (O_1083,N_9823,N_9193);
xor UO_1084 (O_1084,N_8822,N_9030);
and UO_1085 (O_1085,N_8995,N_9633);
and UO_1086 (O_1086,N_9272,N_8904);
or UO_1087 (O_1087,N_9421,N_8844);
nand UO_1088 (O_1088,N_8571,N_9238);
and UO_1089 (O_1089,N_8863,N_8014);
nand UO_1090 (O_1090,N_9261,N_9936);
nand UO_1091 (O_1091,N_7781,N_9836);
nand UO_1092 (O_1092,N_9999,N_9904);
nor UO_1093 (O_1093,N_9292,N_8711);
and UO_1094 (O_1094,N_8313,N_8837);
and UO_1095 (O_1095,N_7845,N_9328);
and UO_1096 (O_1096,N_9891,N_7972);
or UO_1097 (O_1097,N_8704,N_8976);
nand UO_1098 (O_1098,N_9625,N_9066);
or UO_1099 (O_1099,N_9276,N_7892);
nand UO_1100 (O_1100,N_8735,N_9076);
or UO_1101 (O_1101,N_9656,N_9603);
nand UO_1102 (O_1102,N_7626,N_8880);
or UO_1103 (O_1103,N_9609,N_9835);
and UO_1104 (O_1104,N_9027,N_9978);
nand UO_1105 (O_1105,N_8750,N_8229);
or UO_1106 (O_1106,N_8933,N_8201);
nand UO_1107 (O_1107,N_7927,N_7640);
nor UO_1108 (O_1108,N_9536,N_9121);
and UO_1109 (O_1109,N_8504,N_8108);
and UO_1110 (O_1110,N_9663,N_8350);
or UO_1111 (O_1111,N_7986,N_7864);
and UO_1112 (O_1112,N_8581,N_8803);
or UO_1113 (O_1113,N_7869,N_9629);
and UO_1114 (O_1114,N_9279,N_9650);
and UO_1115 (O_1115,N_8573,N_8578);
and UO_1116 (O_1116,N_8492,N_9865);
nor UO_1117 (O_1117,N_9403,N_9924);
nor UO_1118 (O_1118,N_7605,N_9512);
nor UO_1119 (O_1119,N_8059,N_7841);
nand UO_1120 (O_1120,N_9111,N_8602);
nand UO_1121 (O_1121,N_8507,N_7968);
and UO_1122 (O_1122,N_7698,N_9367);
or UO_1123 (O_1123,N_9805,N_9700);
nor UO_1124 (O_1124,N_9086,N_9487);
nor UO_1125 (O_1125,N_9359,N_8169);
or UO_1126 (O_1126,N_7630,N_9057);
and UO_1127 (O_1127,N_9054,N_9365);
and UO_1128 (O_1128,N_9094,N_9017);
nand UO_1129 (O_1129,N_9765,N_9737);
or UO_1130 (O_1130,N_8580,N_9881);
and UO_1131 (O_1131,N_9311,N_9068);
nor UO_1132 (O_1132,N_8345,N_9478);
nand UO_1133 (O_1133,N_8370,N_9447);
and UO_1134 (O_1134,N_8225,N_7947);
or UO_1135 (O_1135,N_9840,N_8372);
nor UO_1136 (O_1136,N_8390,N_9906);
nor UO_1137 (O_1137,N_8517,N_8550);
nor UO_1138 (O_1138,N_9940,N_7773);
nor UO_1139 (O_1139,N_9104,N_7887);
nor UO_1140 (O_1140,N_9645,N_9930);
nand UO_1141 (O_1141,N_8221,N_8605);
nor UO_1142 (O_1142,N_8164,N_8207);
and UO_1143 (O_1143,N_8114,N_8467);
nor UO_1144 (O_1144,N_9705,N_7696);
and UO_1145 (O_1145,N_8464,N_8052);
and UO_1146 (O_1146,N_9271,N_9533);
nor UO_1147 (O_1147,N_9911,N_7761);
or UO_1148 (O_1148,N_9163,N_9972);
nand UO_1149 (O_1149,N_8312,N_9660);
or UO_1150 (O_1150,N_8690,N_7866);
xor UO_1151 (O_1151,N_9020,N_7993);
nand UO_1152 (O_1152,N_9793,N_9383);
nor UO_1153 (O_1153,N_7799,N_9075);
or UO_1154 (O_1154,N_9687,N_9289);
xnor UO_1155 (O_1155,N_8915,N_9221);
nor UO_1156 (O_1156,N_9824,N_9722);
or UO_1157 (O_1157,N_7639,N_7628);
nand UO_1158 (O_1158,N_8676,N_9667);
nor UO_1159 (O_1159,N_7595,N_8042);
and UO_1160 (O_1160,N_7563,N_8806);
nor UO_1161 (O_1161,N_9976,N_9488);
nand UO_1162 (O_1162,N_9226,N_8150);
or UO_1163 (O_1163,N_9578,N_8713);
nand UO_1164 (O_1164,N_9385,N_9655);
nor UO_1165 (O_1165,N_9708,N_9399);
xor UO_1166 (O_1166,N_7915,N_8366);
and UO_1167 (O_1167,N_8416,N_8840);
or UO_1168 (O_1168,N_8388,N_8251);
or UO_1169 (O_1169,N_8881,N_9849);
and UO_1170 (O_1170,N_8347,N_9449);
nand UO_1171 (O_1171,N_8089,N_9293);
nor UO_1172 (O_1172,N_7777,N_7574);
and UO_1173 (O_1173,N_9281,N_8639);
and UO_1174 (O_1174,N_9601,N_8320);
and UO_1175 (O_1175,N_7922,N_8616);
and UO_1176 (O_1176,N_7959,N_8779);
and UO_1177 (O_1177,N_9032,N_8427);
or UO_1178 (O_1178,N_9247,N_9077);
or UO_1179 (O_1179,N_9816,N_8660);
nand UO_1180 (O_1180,N_8986,N_8291);
nor UO_1181 (O_1181,N_9437,N_8654);
nand UO_1182 (O_1182,N_7801,N_7858);
and UO_1183 (O_1183,N_7611,N_8541);
or UO_1184 (O_1184,N_9265,N_8188);
nor UO_1185 (O_1185,N_7702,N_7867);
and UO_1186 (O_1186,N_8555,N_7610);
nand UO_1187 (O_1187,N_9117,N_9169);
nor UO_1188 (O_1188,N_8215,N_8971);
and UO_1189 (O_1189,N_7796,N_8828);
nand UO_1190 (O_1190,N_8387,N_8733);
nor UO_1191 (O_1191,N_7827,N_9530);
or UO_1192 (O_1192,N_7527,N_9864);
nor UO_1193 (O_1193,N_9752,N_7772);
nand UO_1194 (O_1194,N_7953,N_7592);
nor UO_1195 (O_1195,N_8549,N_8272);
nand UO_1196 (O_1196,N_9814,N_7669);
nor UO_1197 (O_1197,N_9785,N_7503);
nand UO_1198 (O_1198,N_8081,N_9827);
nor UO_1199 (O_1199,N_8361,N_7651);
and UO_1200 (O_1200,N_9119,N_9847);
nand UO_1201 (O_1201,N_7877,N_8187);
and UO_1202 (O_1202,N_8895,N_8759);
nor UO_1203 (O_1203,N_9769,N_8845);
nor UO_1204 (O_1204,N_9860,N_9892);
and UO_1205 (O_1205,N_8497,N_8776);
and UO_1206 (O_1206,N_8645,N_8813);
and UO_1207 (O_1207,N_8944,N_7551);
nand UO_1208 (O_1208,N_9606,N_7878);
nor UO_1209 (O_1209,N_8088,N_9353);
nor UO_1210 (O_1210,N_9402,N_9254);
nor UO_1211 (O_1211,N_9653,N_9802);
and UO_1212 (O_1212,N_9125,N_7822);
nor UO_1213 (O_1213,N_8810,N_8058);
nand UO_1214 (O_1214,N_9003,N_8728);
nor UO_1215 (O_1215,N_9136,N_8949);
and UO_1216 (O_1216,N_9160,N_8180);
nor UO_1217 (O_1217,N_8683,N_9507);
nor UO_1218 (O_1218,N_7748,N_9283);
nor UO_1219 (O_1219,N_8934,N_7905);
nor UO_1220 (O_1220,N_8209,N_9457);
nor UO_1221 (O_1221,N_9544,N_7784);
xor UO_1222 (O_1222,N_7701,N_7839);
or UO_1223 (O_1223,N_9790,N_7967);
nand UO_1224 (O_1224,N_9915,N_9720);
nand UO_1225 (O_1225,N_7536,N_8883);
or UO_1226 (O_1226,N_8270,N_8514);
nor UO_1227 (O_1227,N_9745,N_9634);
nor UO_1228 (O_1228,N_9610,N_9620);
and UO_1229 (O_1229,N_7717,N_9776);
or UO_1230 (O_1230,N_7798,N_7889);
nand UO_1231 (O_1231,N_8636,N_8076);
nor UO_1232 (O_1232,N_7810,N_8265);
or UO_1233 (O_1233,N_8173,N_9326);
or UO_1234 (O_1234,N_9448,N_9630);
nor UO_1235 (O_1235,N_8471,N_7874);
nor UO_1236 (O_1236,N_9588,N_9552);
and UO_1237 (O_1237,N_8848,N_8379);
nand UO_1238 (O_1238,N_8515,N_7751);
and UO_1239 (O_1239,N_9624,N_8681);
nor UO_1240 (O_1240,N_9486,N_8021);
nand UO_1241 (O_1241,N_9188,N_9091);
and UO_1242 (O_1242,N_7759,N_7828);
nand UO_1243 (O_1243,N_7637,N_8196);
and UO_1244 (O_1244,N_9013,N_8797);
or UO_1245 (O_1245,N_8932,N_8358);
and UO_1246 (O_1246,N_9135,N_9581);
and UO_1247 (O_1247,N_7530,N_9945);
nand UO_1248 (O_1248,N_7996,N_8048);
and UO_1249 (O_1249,N_8132,N_7933);
or UO_1250 (O_1250,N_7528,N_9409);
nor UO_1251 (O_1251,N_8955,N_7820);
nand UO_1252 (O_1252,N_8539,N_7723);
nand UO_1253 (O_1253,N_8205,N_7550);
nand UO_1254 (O_1254,N_7892,N_9830);
nand UO_1255 (O_1255,N_9800,N_9049);
nand UO_1256 (O_1256,N_9715,N_8054);
and UO_1257 (O_1257,N_9519,N_7933);
nor UO_1258 (O_1258,N_9757,N_9251);
xnor UO_1259 (O_1259,N_9227,N_9353);
nand UO_1260 (O_1260,N_7535,N_8185);
nand UO_1261 (O_1261,N_9589,N_9598);
and UO_1262 (O_1262,N_8965,N_8352);
nor UO_1263 (O_1263,N_8016,N_9193);
nor UO_1264 (O_1264,N_8229,N_9478);
or UO_1265 (O_1265,N_8371,N_7955);
nand UO_1266 (O_1266,N_8246,N_8018);
nand UO_1267 (O_1267,N_9969,N_8155);
and UO_1268 (O_1268,N_7869,N_8324);
nand UO_1269 (O_1269,N_8523,N_7522);
or UO_1270 (O_1270,N_8927,N_8591);
or UO_1271 (O_1271,N_9748,N_7704);
nand UO_1272 (O_1272,N_9717,N_8788);
or UO_1273 (O_1273,N_8388,N_8988);
nand UO_1274 (O_1274,N_9185,N_9286);
or UO_1275 (O_1275,N_8082,N_9380);
and UO_1276 (O_1276,N_8543,N_9782);
or UO_1277 (O_1277,N_9820,N_9329);
nand UO_1278 (O_1278,N_9105,N_9048);
nor UO_1279 (O_1279,N_9468,N_9622);
nor UO_1280 (O_1280,N_8669,N_9494);
nand UO_1281 (O_1281,N_9489,N_7743);
nor UO_1282 (O_1282,N_8783,N_7823);
or UO_1283 (O_1283,N_9829,N_8104);
and UO_1284 (O_1284,N_8520,N_9812);
nand UO_1285 (O_1285,N_9446,N_8852);
nand UO_1286 (O_1286,N_8283,N_9694);
nor UO_1287 (O_1287,N_8431,N_8343);
nand UO_1288 (O_1288,N_9367,N_9052);
nor UO_1289 (O_1289,N_9051,N_8461);
nor UO_1290 (O_1290,N_8056,N_8200);
nand UO_1291 (O_1291,N_8499,N_9679);
nor UO_1292 (O_1292,N_9297,N_9581);
xnor UO_1293 (O_1293,N_8047,N_9904);
or UO_1294 (O_1294,N_8995,N_9035);
nor UO_1295 (O_1295,N_9820,N_9906);
nor UO_1296 (O_1296,N_7747,N_9368);
and UO_1297 (O_1297,N_8608,N_7600);
nand UO_1298 (O_1298,N_9378,N_8041);
nor UO_1299 (O_1299,N_8698,N_9098);
or UO_1300 (O_1300,N_8019,N_9288);
nor UO_1301 (O_1301,N_9836,N_8238);
nand UO_1302 (O_1302,N_8941,N_7885);
nand UO_1303 (O_1303,N_7868,N_8504);
nor UO_1304 (O_1304,N_7508,N_8859);
and UO_1305 (O_1305,N_8122,N_8081);
or UO_1306 (O_1306,N_8486,N_8667);
or UO_1307 (O_1307,N_9880,N_8177);
nor UO_1308 (O_1308,N_9193,N_7791);
nand UO_1309 (O_1309,N_9585,N_8192);
nor UO_1310 (O_1310,N_8696,N_9436);
and UO_1311 (O_1311,N_7510,N_7601);
or UO_1312 (O_1312,N_7740,N_9235);
nand UO_1313 (O_1313,N_9365,N_7677);
nor UO_1314 (O_1314,N_9126,N_8386);
or UO_1315 (O_1315,N_8129,N_9739);
or UO_1316 (O_1316,N_8470,N_9576);
nor UO_1317 (O_1317,N_9043,N_8214);
nor UO_1318 (O_1318,N_8323,N_8574);
nand UO_1319 (O_1319,N_7623,N_8140);
and UO_1320 (O_1320,N_7591,N_9285);
nand UO_1321 (O_1321,N_9244,N_8169);
nor UO_1322 (O_1322,N_7537,N_8806);
and UO_1323 (O_1323,N_8064,N_8656);
and UO_1324 (O_1324,N_7869,N_8490);
or UO_1325 (O_1325,N_8202,N_8847);
nand UO_1326 (O_1326,N_7619,N_9846);
nor UO_1327 (O_1327,N_7992,N_8738);
or UO_1328 (O_1328,N_8024,N_7926);
and UO_1329 (O_1329,N_8432,N_8677);
nor UO_1330 (O_1330,N_9541,N_8046);
or UO_1331 (O_1331,N_8353,N_8688);
nand UO_1332 (O_1332,N_8760,N_7998);
or UO_1333 (O_1333,N_8454,N_8500);
nor UO_1334 (O_1334,N_9197,N_9698);
or UO_1335 (O_1335,N_9068,N_9940);
nand UO_1336 (O_1336,N_9234,N_8392);
nand UO_1337 (O_1337,N_8506,N_9061);
and UO_1338 (O_1338,N_8982,N_7590);
or UO_1339 (O_1339,N_9175,N_8557);
nor UO_1340 (O_1340,N_8232,N_7995);
and UO_1341 (O_1341,N_8339,N_9451);
nand UO_1342 (O_1342,N_8589,N_8708);
nor UO_1343 (O_1343,N_9738,N_7595);
and UO_1344 (O_1344,N_8671,N_7660);
nand UO_1345 (O_1345,N_9780,N_8445);
nor UO_1346 (O_1346,N_9877,N_9381);
and UO_1347 (O_1347,N_8006,N_9955);
nand UO_1348 (O_1348,N_7977,N_7567);
or UO_1349 (O_1349,N_8187,N_8600);
nor UO_1350 (O_1350,N_9744,N_9508);
nand UO_1351 (O_1351,N_8673,N_7955);
or UO_1352 (O_1352,N_8068,N_8815);
nor UO_1353 (O_1353,N_8325,N_7873);
or UO_1354 (O_1354,N_8274,N_9235);
nor UO_1355 (O_1355,N_8991,N_8975);
or UO_1356 (O_1356,N_9196,N_8125);
nand UO_1357 (O_1357,N_9579,N_8882);
and UO_1358 (O_1358,N_9994,N_9133);
and UO_1359 (O_1359,N_8493,N_8977);
nand UO_1360 (O_1360,N_9676,N_8588);
and UO_1361 (O_1361,N_9460,N_8318);
nand UO_1362 (O_1362,N_8475,N_9465);
nor UO_1363 (O_1363,N_8478,N_7859);
and UO_1364 (O_1364,N_9545,N_9869);
and UO_1365 (O_1365,N_9810,N_7555);
nor UO_1366 (O_1366,N_8665,N_9724);
nand UO_1367 (O_1367,N_8432,N_9733);
nor UO_1368 (O_1368,N_9095,N_9033);
and UO_1369 (O_1369,N_9696,N_9193);
nor UO_1370 (O_1370,N_7609,N_8835);
and UO_1371 (O_1371,N_9016,N_8244);
nand UO_1372 (O_1372,N_8278,N_9012);
nor UO_1373 (O_1373,N_8368,N_7535);
nor UO_1374 (O_1374,N_8603,N_8277);
nand UO_1375 (O_1375,N_8089,N_9028);
nor UO_1376 (O_1376,N_9163,N_9937);
and UO_1377 (O_1377,N_7883,N_8045);
nor UO_1378 (O_1378,N_8066,N_9300);
and UO_1379 (O_1379,N_9305,N_9896);
or UO_1380 (O_1380,N_9626,N_9258);
nand UO_1381 (O_1381,N_8683,N_7677);
and UO_1382 (O_1382,N_9715,N_7779);
or UO_1383 (O_1383,N_7772,N_8855);
nand UO_1384 (O_1384,N_9548,N_9269);
nor UO_1385 (O_1385,N_9328,N_8057);
nand UO_1386 (O_1386,N_8641,N_9537);
and UO_1387 (O_1387,N_9036,N_8356);
nor UO_1388 (O_1388,N_8040,N_8799);
and UO_1389 (O_1389,N_7959,N_8738);
nor UO_1390 (O_1390,N_9507,N_9085);
nor UO_1391 (O_1391,N_8589,N_7626);
or UO_1392 (O_1392,N_7989,N_9016);
nand UO_1393 (O_1393,N_8000,N_7731);
or UO_1394 (O_1394,N_9308,N_9382);
and UO_1395 (O_1395,N_8335,N_8035);
nand UO_1396 (O_1396,N_9872,N_9463);
nand UO_1397 (O_1397,N_8053,N_7649);
and UO_1398 (O_1398,N_8042,N_7885);
nor UO_1399 (O_1399,N_9334,N_8641);
and UO_1400 (O_1400,N_9761,N_8806);
or UO_1401 (O_1401,N_9682,N_8757);
or UO_1402 (O_1402,N_7723,N_7503);
or UO_1403 (O_1403,N_8126,N_9063);
nor UO_1404 (O_1404,N_9675,N_8573);
nor UO_1405 (O_1405,N_8389,N_9174);
or UO_1406 (O_1406,N_9676,N_9463);
or UO_1407 (O_1407,N_8232,N_9836);
nand UO_1408 (O_1408,N_9182,N_9630);
nor UO_1409 (O_1409,N_8909,N_7686);
nor UO_1410 (O_1410,N_8780,N_7748);
nor UO_1411 (O_1411,N_8894,N_7889);
and UO_1412 (O_1412,N_7699,N_8336);
nor UO_1413 (O_1413,N_9437,N_9862);
nor UO_1414 (O_1414,N_8922,N_8748);
and UO_1415 (O_1415,N_7882,N_9021);
or UO_1416 (O_1416,N_8812,N_8464);
or UO_1417 (O_1417,N_9073,N_7508);
nand UO_1418 (O_1418,N_8375,N_7638);
nand UO_1419 (O_1419,N_9749,N_8254);
or UO_1420 (O_1420,N_8322,N_8540);
and UO_1421 (O_1421,N_8296,N_8534);
nand UO_1422 (O_1422,N_9610,N_7974);
nor UO_1423 (O_1423,N_7606,N_9102);
nor UO_1424 (O_1424,N_9212,N_9894);
nor UO_1425 (O_1425,N_9875,N_8773);
nor UO_1426 (O_1426,N_8662,N_9844);
nor UO_1427 (O_1427,N_8305,N_9307);
and UO_1428 (O_1428,N_9865,N_8195);
and UO_1429 (O_1429,N_9259,N_8529);
and UO_1430 (O_1430,N_7672,N_8307);
and UO_1431 (O_1431,N_9376,N_9460);
or UO_1432 (O_1432,N_7773,N_9341);
and UO_1433 (O_1433,N_9466,N_9994);
or UO_1434 (O_1434,N_9568,N_8278);
and UO_1435 (O_1435,N_9288,N_8805);
nand UO_1436 (O_1436,N_9615,N_9192);
or UO_1437 (O_1437,N_7654,N_8578);
or UO_1438 (O_1438,N_9485,N_8471);
or UO_1439 (O_1439,N_7510,N_8463);
and UO_1440 (O_1440,N_9600,N_9192);
and UO_1441 (O_1441,N_7888,N_9410);
nor UO_1442 (O_1442,N_7795,N_8262);
or UO_1443 (O_1443,N_8215,N_9081);
or UO_1444 (O_1444,N_8378,N_8172);
nand UO_1445 (O_1445,N_9388,N_9728);
and UO_1446 (O_1446,N_8799,N_8804);
nand UO_1447 (O_1447,N_7768,N_9717);
nor UO_1448 (O_1448,N_9892,N_8176);
or UO_1449 (O_1449,N_9240,N_9621);
nand UO_1450 (O_1450,N_8832,N_8922);
nand UO_1451 (O_1451,N_8373,N_7664);
or UO_1452 (O_1452,N_9454,N_8619);
nand UO_1453 (O_1453,N_9313,N_9608);
nor UO_1454 (O_1454,N_7732,N_9045);
or UO_1455 (O_1455,N_8674,N_8346);
nand UO_1456 (O_1456,N_8429,N_8616);
and UO_1457 (O_1457,N_8873,N_8199);
and UO_1458 (O_1458,N_7719,N_9203);
and UO_1459 (O_1459,N_7676,N_9135);
and UO_1460 (O_1460,N_8445,N_9927);
or UO_1461 (O_1461,N_7663,N_7642);
nand UO_1462 (O_1462,N_9017,N_7804);
nor UO_1463 (O_1463,N_7829,N_9257);
nand UO_1464 (O_1464,N_9801,N_8305);
nor UO_1465 (O_1465,N_9877,N_7651);
nand UO_1466 (O_1466,N_7532,N_7556);
and UO_1467 (O_1467,N_9937,N_8588);
nand UO_1468 (O_1468,N_9158,N_8694);
nand UO_1469 (O_1469,N_8652,N_9760);
nand UO_1470 (O_1470,N_8500,N_8981);
and UO_1471 (O_1471,N_9050,N_8035);
nand UO_1472 (O_1472,N_9940,N_7863);
or UO_1473 (O_1473,N_7716,N_7929);
or UO_1474 (O_1474,N_9349,N_9687);
or UO_1475 (O_1475,N_9378,N_8868);
nand UO_1476 (O_1476,N_8441,N_7916);
nor UO_1477 (O_1477,N_9152,N_7610);
nor UO_1478 (O_1478,N_8660,N_7896);
xnor UO_1479 (O_1479,N_9986,N_8722);
nand UO_1480 (O_1480,N_7629,N_7749);
nor UO_1481 (O_1481,N_9096,N_9020);
nor UO_1482 (O_1482,N_9390,N_9578);
xnor UO_1483 (O_1483,N_7562,N_8872);
or UO_1484 (O_1484,N_7850,N_9729);
or UO_1485 (O_1485,N_8839,N_9590);
nand UO_1486 (O_1486,N_9021,N_9294);
nor UO_1487 (O_1487,N_7617,N_8978);
or UO_1488 (O_1488,N_9530,N_7646);
or UO_1489 (O_1489,N_9189,N_7634);
and UO_1490 (O_1490,N_7730,N_9013);
and UO_1491 (O_1491,N_9067,N_8838);
nand UO_1492 (O_1492,N_8531,N_8855);
and UO_1493 (O_1493,N_8274,N_9736);
or UO_1494 (O_1494,N_8505,N_8542);
nand UO_1495 (O_1495,N_8867,N_8019);
nand UO_1496 (O_1496,N_9927,N_9950);
or UO_1497 (O_1497,N_7562,N_8933);
nor UO_1498 (O_1498,N_7979,N_7539);
nor UO_1499 (O_1499,N_8697,N_8945);
endmodule