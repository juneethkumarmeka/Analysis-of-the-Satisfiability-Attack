module basic_500_3000_500_30_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_378,In_340);
nand U1 (N_1,In_383,In_55);
xor U2 (N_2,In_140,In_363);
xor U3 (N_3,In_145,In_352);
and U4 (N_4,In_394,In_281);
xor U5 (N_5,In_477,In_336);
xor U6 (N_6,In_97,In_123);
nor U7 (N_7,In_331,In_486);
and U8 (N_8,In_358,In_445);
or U9 (N_9,In_479,In_343);
nand U10 (N_10,In_471,In_34);
xnor U11 (N_11,In_236,In_231);
or U12 (N_12,In_195,In_206);
nor U13 (N_13,In_210,In_414);
nor U14 (N_14,In_440,In_308);
nand U15 (N_15,In_277,In_256);
xnor U16 (N_16,In_95,In_133);
nor U17 (N_17,In_487,In_332);
or U18 (N_18,In_230,In_125);
xnor U19 (N_19,In_238,In_135);
nor U20 (N_20,In_404,In_385);
and U21 (N_21,In_166,In_320);
nor U22 (N_22,In_398,In_49);
and U23 (N_23,In_262,In_401);
xor U24 (N_24,In_172,In_190);
nand U25 (N_25,In_196,In_251);
xor U26 (N_26,In_76,In_204);
or U27 (N_27,In_453,In_311);
and U28 (N_28,In_214,In_60);
and U29 (N_29,In_327,In_420);
nor U30 (N_30,In_284,In_261);
and U31 (N_31,In_211,In_490);
nand U32 (N_32,In_424,In_244);
xnor U33 (N_33,In_104,In_397);
nor U34 (N_34,In_351,In_83);
nand U35 (N_35,In_456,In_136);
and U36 (N_36,In_80,In_285);
and U37 (N_37,In_380,In_313);
or U38 (N_38,In_485,In_30);
or U39 (N_39,In_442,In_81);
or U40 (N_40,In_291,In_37);
nand U41 (N_41,In_310,In_213);
nor U42 (N_42,In_433,In_434);
or U43 (N_43,In_186,In_240);
nor U44 (N_44,In_402,In_268);
nor U45 (N_45,In_447,In_316);
and U46 (N_46,In_149,In_259);
and U47 (N_47,In_342,In_146);
nor U48 (N_48,In_232,In_499);
and U49 (N_49,In_130,In_163);
nand U50 (N_50,In_274,In_33);
and U51 (N_51,In_105,In_208);
or U52 (N_52,In_198,In_319);
and U53 (N_53,In_188,In_241);
xor U54 (N_54,In_314,In_35);
and U55 (N_55,In_164,In_432);
and U56 (N_56,In_39,In_267);
and U57 (N_57,In_318,In_295);
or U58 (N_58,In_21,In_229);
xnor U59 (N_59,In_496,In_252);
or U60 (N_60,In_405,In_67);
nor U61 (N_61,In_148,In_386);
nand U62 (N_62,In_367,In_138);
or U63 (N_63,In_132,In_32);
nor U64 (N_64,In_181,In_297);
nand U65 (N_65,In_11,In_45);
and U66 (N_66,In_107,In_278);
nor U67 (N_67,In_171,In_79);
nand U68 (N_68,In_73,In_40);
xnor U69 (N_69,In_403,In_92);
and U70 (N_70,In_333,In_36);
and U71 (N_71,In_41,In_482);
or U72 (N_72,In_392,In_247);
or U73 (N_73,In_1,In_430);
and U74 (N_74,In_271,In_20);
nand U75 (N_75,In_476,In_377);
nor U76 (N_76,In_239,In_473);
nand U77 (N_77,In_234,In_279);
nor U78 (N_78,In_459,In_300);
and U79 (N_79,In_14,In_417);
nand U80 (N_80,In_187,In_156);
nand U81 (N_81,In_480,In_109);
nor U82 (N_82,In_154,In_461);
nand U83 (N_83,In_167,In_418);
nor U84 (N_84,In_365,In_68);
nand U85 (N_85,In_99,In_263);
and U86 (N_86,In_458,In_349);
xnor U87 (N_87,In_235,In_326);
or U88 (N_88,In_63,In_307);
nor U89 (N_89,In_406,In_15);
nand U90 (N_90,In_91,In_56);
and U91 (N_91,In_29,In_137);
and U92 (N_92,In_191,In_131);
xor U93 (N_93,In_346,In_493);
nor U94 (N_94,In_86,In_160);
and U95 (N_95,In_157,In_302);
and U96 (N_96,In_175,In_360);
and U97 (N_97,In_162,In_246);
nand U98 (N_98,In_457,In_151);
xor U99 (N_99,In_180,In_118);
or U100 (N_100,In_87,N_81);
nand U101 (N_101,In_23,In_395);
nand U102 (N_102,In_89,In_257);
nand U103 (N_103,N_78,In_357);
nand U104 (N_104,In_350,In_142);
xor U105 (N_105,N_77,In_225);
nand U106 (N_106,In_321,In_498);
nor U107 (N_107,In_84,In_483);
nand U108 (N_108,N_5,N_41);
nand U109 (N_109,In_373,In_269);
xnor U110 (N_110,In_304,In_48);
nor U111 (N_111,N_23,In_19);
or U112 (N_112,In_389,N_17);
or U113 (N_113,N_68,N_8);
or U114 (N_114,N_10,In_169);
and U115 (N_115,In_75,In_42);
nand U116 (N_116,In_280,In_301);
nand U117 (N_117,In_335,N_55);
xnor U118 (N_118,In_429,In_384);
nand U119 (N_119,In_64,In_98);
nor U120 (N_120,In_464,In_115);
nand U121 (N_121,In_345,In_382);
or U122 (N_122,In_286,In_255);
nor U123 (N_123,In_158,In_428);
or U124 (N_124,In_359,In_62);
or U125 (N_125,N_46,In_147);
or U126 (N_126,In_2,In_354);
and U127 (N_127,In_283,N_50);
nand U128 (N_128,In_159,In_66);
and U129 (N_129,In_243,In_24);
nand U130 (N_130,In_116,In_412);
or U131 (N_131,In_47,In_128);
nand U132 (N_132,In_381,In_144);
and U133 (N_133,N_99,N_57);
nor U134 (N_134,In_455,N_59);
or U135 (N_135,N_65,In_51);
or U136 (N_136,In_177,N_88);
or U137 (N_137,In_150,In_423);
xor U138 (N_138,N_28,In_452);
nor U139 (N_139,N_42,N_79);
or U140 (N_140,In_454,In_481);
and U141 (N_141,In_43,N_84);
or U142 (N_142,In_113,In_100);
nor U143 (N_143,In_366,In_117);
nor U144 (N_144,N_83,In_218);
or U145 (N_145,N_61,In_216);
nand U146 (N_146,N_82,In_96);
xor U147 (N_147,In_391,In_303);
or U148 (N_148,In_10,In_450);
nor U149 (N_149,In_400,In_441);
nand U150 (N_150,In_155,N_94);
nand U151 (N_151,In_178,N_51);
or U152 (N_152,N_1,N_16);
nand U153 (N_153,In_339,In_226);
xnor U154 (N_154,In_361,In_112);
and U155 (N_155,N_2,In_469);
and U156 (N_156,N_9,In_416);
nand U157 (N_157,In_82,In_396);
nor U158 (N_158,In_497,In_435);
nand U159 (N_159,N_31,In_78);
and U160 (N_160,In_431,In_266);
or U161 (N_161,In_224,In_170);
xor U162 (N_162,N_36,In_347);
xor U163 (N_163,N_6,In_119);
or U164 (N_164,In_356,In_201);
and U165 (N_165,N_14,In_426);
nand U166 (N_166,N_97,In_227);
nand U167 (N_167,In_368,In_94);
xnor U168 (N_168,In_338,In_182);
nor U169 (N_169,In_489,In_444);
and U170 (N_170,In_468,N_66);
xnor U171 (N_171,In_463,In_449);
nand U172 (N_172,In_179,In_353);
nand U173 (N_173,In_419,In_219);
xor U174 (N_174,In_451,In_122);
xnor U175 (N_175,In_324,In_44);
and U176 (N_176,In_273,In_120);
nor U177 (N_177,N_18,In_31);
or U178 (N_178,In_4,N_40);
nor U179 (N_179,In_103,In_0);
nor U180 (N_180,In_296,In_495);
nor U181 (N_181,In_312,In_293);
xor U182 (N_182,In_38,N_67);
nor U183 (N_183,In_334,In_292);
nand U184 (N_184,In_376,In_189);
nor U185 (N_185,In_298,In_448);
xor U186 (N_186,N_74,N_12);
or U187 (N_187,In_58,In_446);
or U188 (N_188,In_165,N_19);
nor U189 (N_189,In_379,In_460);
and U190 (N_190,In_106,N_69);
xor U191 (N_191,In_484,In_248);
and U192 (N_192,In_372,In_197);
or U193 (N_193,In_212,N_38);
or U194 (N_194,N_75,In_16);
and U195 (N_195,In_8,In_194);
xor U196 (N_196,N_48,In_121);
xor U197 (N_197,In_299,N_54);
nand U198 (N_198,In_330,In_69);
xnor U199 (N_199,N_35,N_49);
and U200 (N_200,N_104,In_413);
nand U201 (N_201,N_106,In_26);
xor U202 (N_202,In_85,N_171);
and U203 (N_203,N_155,N_195);
or U204 (N_204,In_233,In_111);
nand U205 (N_205,N_85,N_90);
or U206 (N_206,N_52,In_70);
and U207 (N_207,In_5,N_26);
nand U208 (N_208,In_393,In_478);
and U209 (N_209,In_375,N_113);
and U210 (N_210,N_130,N_157);
and U211 (N_211,N_165,In_223);
nor U212 (N_212,In_306,N_107);
or U213 (N_213,N_63,In_364);
nand U214 (N_214,In_409,N_76);
nor U215 (N_215,N_71,N_91);
xnor U216 (N_216,In_288,In_242);
or U217 (N_217,In_466,N_72);
nand U218 (N_218,In_46,N_179);
xnor U219 (N_219,In_126,In_17);
and U220 (N_220,In_264,In_249);
and U221 (N_221,N_124,N_169);
nand U222 (N_222,N_73,In_57);
nand U223 (N_223,N_156,In_390);
nand U224 (N_224,In_470,In_102);
xnor U225 (N_225,N_7,In_174);
and U226 (N_226,In_52,In_438);
and U227 (N_227,In_411,In_25);
nand U228 (N_228,N_153,N_119);
nand U229 (N_229,N_13,N_0);
xor U230 (N_230,In_93,In_315);
and U231 (N_231,In_415,In_475);
and U232 (N_232,In_183,N_143);
and U233 (N_233,N_123,In_427);
and U234 (N_234,In_407,N_140);
nor U235 (N_235,In_205,N_181);
and U236 (N_236,N_178,N_149);
xor U237 (N_237,In_65,In_253);
and U238 (N_238,N_129,In_207);
and U239 (N_239,N_45,N_92);
and U240 (N_240,In_348,N_160);
nand U241 (N_241,N_60,In_309);
or U242 (N_242,In_3,N_150);
nor U243 (N_243,N_33,In_370);
or U244 (N_244,In_408,In_488);
and U245 (N_245,N_131,N_20);
nor U246 (N_246,N_112,In_168);
nor U247 (N_247,N_64,N_70);
nand U248 (N_248,In_422,In_77);
or U249 (N_249,In_491,N_199);
and U250 (N_250,In_101,N_167);
nand U251 (N_251,In_108,N_183);
nor U252 (N_252,N_174,N_164);
xor U253 (N_253,N_11,In_317);
xor U254 (N_254,N_122,In_323);
and U255 (N_255,N_159,In_492);
nor U256 (N_256,N_194,In_369);
nand U257 (N_257,In_437,In_250);
and U258 (N_258,N_110,N_141);
nand U259 (N_259,In_71,N_62);
and U260 (N_260,N_21,In_467);
and U261 (N_261,N_145,In_289);
xor U262 (N_262,In_388,N_189);
nor U263 (N_263,In_193,N_170);
nor U264 (N_264,In_209,In_27);
and U265 (N_265,In_287,N_32);
xor U266 (N_266,N_148,N_136);
nand U267 (N_267,In_152,N_29);
nor U268 (N_268,N_126,In_341);
or U269 (N_269,In_220,In_329);
or U270 (N_270,N_146,In_276);
and U271 (N_271,N_44,In_28);
or U272 (N_272,N_89,N_133);
nand U273 (N_273,In_200,In_237);
xnor U274 (N_274,N_177,N_161);
nor U275 (N_275,N_27,N_132);
or U276 (N_276,In_114,N_24);
xnor U277 (N_277,In_124,N_93);
or U278 (N_278,N_105,N_144);
and U279 (N_279,N_34,In_18);
nor U280 (N_280,N_182,In_258);
or U281 (N_281,N_43,In_290);
xnor U282 (N_282,In_110,N_188);
xor U283 (N_283,N_186,N_98);
nor U284 (N_284,In_355,N_173);
or U285 (N_285,N_139,N_58);
xnor U286 (N_286,In_387,In_221);
nand U287 (N_287,In_228,In_74);
xnor U288 (N_288,N_142,In_143);
nand U289 (N_289,In_72,N_101);
xnor U290 (N_290,N_197,In_139);
nor U291 (N_291,N_100,In_90);
nand U292 (N_292,In_344,In_53);
nand U293 (N_293,N_96,In_6);
or U294 (N_294,N_86,N_151);
nor U295 (N_295,N_154,In_275);
xor U296 (N_296,N_125,N_102);
and U297 (N_297,In_127,In_59);
or U298 (N_298,In_472,In_399);
and U299 (N_299,N_172,N_37);
and U300 (N_300,N_241,In_362);
nor U301 (N_301,In_161,In_22);
and U302 (N_302,N_279,N_296);
or U303 (N_303,N_135,N_214);
xnor U304 (N_304,N_207,N_251);
or U305 (N_305,N_289,In_465);
and U306 (N_306,N_243,In_260);
and U307 (N_307,N_286,In_9);
and U308 (N_308,N_206,N_212);
nand U309 (N_309,N_208,In_337);
nor U310 (N_310,N_288,In_173);
nor U311 (N_311,N_266,In_325);
nand U312 (N_312,N_265,N_147);
xor U313 (N_313,In_272,In_141);
or U314 (N_314,N_163,N_111);
or U315 (N_315,In_134,In_474);
and U316 (N_316,N_267,N_15);
and U317 (N_317,In_436,N_261);
or U318 (N_318,N_264,N_87);
nand U319 (N_319,In_13,N_56);
nand U320 (N_320,In_425,N_120);
or U321 (N_321,In_305,N_176);
nand U322 (N_322,In_88,N_269);
xnor U323 (N_323,N_268,In_322);
nand U324 (N_324,N_294,In_203);
and U325 (N_325,N_128,N_168);
and U326 (N_326,N_256,N_257);
nor U327 (N_327,N_273,N_205);
xor U328 (N_328,N_250,N_225);
and U329 (N_329,N_229,N_185);
xnor U330 (N_330,N_222,N_245);
and U331 (N_331,N_263,N_246);
xnor U332 (N_332,N_191,N_184);
nor U333 (N_333,N_237,N_200);
nor U334 (N_334,N_30,N_4);
nor U335 (N_335,N_213,N_293);
nand U336 (N_336,In_294,N_127);
and U337 (N_337,N_275,N_210);
xor U338 (N_338,N_244,N_219);
nor U339 (N_339,N_236,N_240);
and U340 (N_340,N_249,N_121);
nand U341 (N_341,N_80,In_222);
nand U342 (N_342,N_137,N_270);
or U343 (N_343,N_228,N_162);
nand U344 (N_344,N_231,N_248);
nor U345 (N_345,N_223,N_259);
nor U346 (N_346,N_282,N_152);
nand U347 (N_347,In_282,N_277);
nand U348 (N_348,N_138,N_108);
nand U349 (N_349,N_258,In_328);
nor U350 (N_350,N_217,N_290);
or U351 (N_351,N_252,N_297);
and U352 (N_352,N_287,N_22);
xor U353 (N_353,In_54,N_280);
nand U354 (N_354,N_272,N_230);
and U355 (N_355,In_494,In_202);
nor U356 (N_356,N_253,N_234);
nor U357 (N_357,N_103,N_285);
xor U358 (N_358,In_371,N_242);
nand U359 (N_359,In_129,In_410);
and U360 (N_360,N_255,N_109);
xor U361 (N_361,In_462,N_220);
xor U362 (N_362,N_215,N_218);
nor U363 (N_363,In_50,N_134);
and U364 (N_364,N_202,N_274);
and U365 (N_365,N_204,In_176);
xnor U366 (N_366,N_187,N_116);
xor U367 (N_367,N_115,N_281);
or U368 (N_368,In_443,N_95);
nor U369 (N_369,N_192,N_247);
xor U370 (N_370,N_211,In_245);
xnor U371 (N_371,N_232,In_192);
nand U372 (N_372,N_118,In_184);
and U373 (N_373,In_12,N_190);
or U374 (N_374,In_254,N_193);
or U375 (N_375,N_226,N_295);
nand U376 (N_376,N_203,N_235);
xnor U377 (N_377,N_271,N_216);
and U378 (N_378,N_117,In_265);
nand U379 (N_379,N_221,N_39);
nand U380 (N_380,N_238,In_421);
nand U381 (N_381,N_227,N_53);
and U382 (N_382,N_158,In_439);
or U383 (N_383,N_233,N_276);
and U384 (N_384,In_199,In_7);
or U385 (N_385,N_3,In_217);
nand U386 (N_386,N_298,N_224);
nor U387 (N_387,N_209,N_166);
nand U388 (N_388,In_374,N_196);
xnor U389 (N_389,N_260,In_185);
xor U390 (N_390,N_201,N_114);
xnor U391 (N_391,In_215,N_278);
and U392 (N_392,N_292,N_47);
nor U393 (N_393,N_198,In_153);
nor U394 (N_394,N_239,N_175);
and U395 (N_395,N_291,N_284);
and U396 (N_396,N_25,N_180);
xnor U397 (N_397,In_270,N_299);
nand U398 (N_398,In_61,N_254);
and U399 (N_399,N_262,N_283);
and U400 (N_400,N_353,N_327);
nand U401 (N_401,N_337,N_385);
nand U402 (N_402,N_397,N_305);
xnor U403 (N_403,N_300,N_311);
or U404 (N_404,N_306,N_315);
or U405 (N_405,N_363,N_392);
nand U406 (N_406,N_398,N_302);
or U407 (N_407,N_345,N_395);
nor U408 (N_408,N_304,N_333);
nand U409 (N_409,N_346,N_377);
xnor U410 (N_410,N_382,N_341);
or U411 (N_411,N_351,N_321);
or U412 (N_412,N_354,N_347);
xor U413 (N_413,N_376,N_322);
nor U414 (N_414,N_331,N_393);
xnor U415 (N_415,N_334,N_355);
and U416 (N_416,N_375,N_352);
xnor U417 (N_417,N_301,N_390);
nor U418 (N_418,N_344,N_316);
nand U419 (N_419,N_325,N_380);
xnor U420 (N_420,N_383,N_371);
nand U421 (N_421,N_336,N_313);
or U422 (N_422,N_328,N_317);
and U423 (N_423,N_358,N_326);
nor U424 (N_424,N_307,N_378);
nand U425 (N_425,N_396,N_384);
nor U426 (N_426,N_339,N_362);
xor U427 (N_427,N_324,N_356);
xnor U428 (N_428,N_370,N_359);
or U429 (N_429,N_309,N_364);
nand U430 (N_430,N_386,N_310);
and U431 (N_431,N_388,N_373);
or U432 (N_432,N_319,N_394);
nor U433 (N_433,N_348,N_357);
nand U434 (N_434,N_308,N_312);
nand U435 (N_435,N_389,N_340);
and U436 (N_436,N_361,N_374);
and U437 (N_437,N_332,N_366);
and U438 (N_438,N_318,N_372);
nor U439 (N_439,N_369,N_335);
nand U440 (N_440,N_320,N_303);
nand U441 (N_441,N_379,N_367);
nor U442 (N_442,N_360,N_349);
nor U443 (N_443,N_350,N_399);
nor U444 (N_444,N_342,N_314);
nand U445 (N_445,N_381,N_368);
xnor U446 (N_446,N_330,N_387);
xor U447 (N_447,N_365,N_338);
and U448 (N_448,N_323,N_329);
xor U449 (N_449,N_391,N_343);
nand U450 (N_450,N_356,N_361);
or U451 (N_451,N_381,N_305);
nor U452 (N_452,N_379,N_312);
xnor U453 (N_453,N_386,N_359);
xor U454 (N_454,N_382,N_334);
and U455 (N_455,N_332,N_396);
and U456 (N_456,N_332,N_328);
and U457 (N_457,N_322,N_355);
nand U458 (N_458,N_327,N_368);
xor U459 (N_459,N_393,N_347);
xor U460 (N_460,N_387,N_345);
and U461 (N_461,N_332,N_347);
or U462 (N_462,N_389,N_397);
or U463 (N_463,N_311,N_331);
nor U464 (N_464,N_329,N_377);
and U465 (N_465,N_330,N_388);
and U466 (N_466,N_324,N_381);
or U467 (N_467,N_357,N_318);
nand U468 (N_468,N_306,N_369);
nand U469 (N_469,N_363,N_329);
xor U470 (N_470,N_348,N_340);
nor U471 (N_471,N_326,N_309);
nand U472 (N_472,N_345,N_342);
nor U473 (N_473,N_337,N_302);
and U474 (N_474,N_387,N_392);
nand U475 (N_475,N_388,N_319);
and U476 (N_476,N_380,N_383);
nand U477 (N_477,N_352,N_363);
xnor U478 (N_478,N_343,N_396);
or U479 (N_479,N_365,N_348);
nand U480 (N_480,N_374,N_377);
nand U481 (N_481,N_321,N_361);
nor U482 (N_482,N_390,N_338);
nand U483 (N_483,N_336,N_348);
nor U484 (N_484,N_386,N_314);
xor U485 (N_485,N_337,N_365);
nor U486 (N_486,N_384,N_367);
nor U487 (N_487,N_365,N_352);
and U488 (N_488,N_397,N_304);
nor U489 (N_489,N_358,N_392);
or U490 (N_490,N_379,N_358);
xnor U491 (N_491,N_348,N_352);
or U492 (N_492,N_362,N_359);
nand U493 (N_493,N_317,N_329);
nor U494 (N_494,N_338,N_360);
nor U495 (N_495,N_346,N_357);
xnor U496 (N_496,N_318,N_313);
or U497 (N_497,N_392,N_338);
and U498 (N_498,N_348,N_339);
nand U499 (N_499,N_384,N_373);
nor U500 (N_500,N_428,N_410);
nand U501 (N_501,N_485,N_483);
xnor U502 (N_502,N_480,N_430);
nand U503 (N_503,N_461,N_425);
nor U504 (N_504,N_446,N_487);
nor U505 (N_505,N_454,N_409);
and U506 (N_506,N_453,N_497);
or U507 (N_507,N_494,N_421);
nand U508 (N_508,N_404,N_438);
xor U509 (N_509,N_420,N_441);
nor U510 (N_510,N_402,N_481);
and U511 (N_511,N_408,N_426);
nand U512 (N_512,N_484,N_417);
or U513 (N_513,N_433,N_434);
xnor U514 (N_514,N_492,N_444);
nor U515 (N_515,N_455,N_401);
nor U516 (N_516,N_488,N_464);
and U517 (N_517,N_469,N_472);
and U518 (N_518,N_448,N_449);
nand U519 (N_519,N_457,N_479);
nand U520 (N_520,N_412,N_423);
or U521 (N_521,N_499,N_456);
and U522 (N_522,N_443,N_470);
xnor U523 (N_523,N_427,N_450);
or U524 (N_524,N_491,N_498);
or U525 (N_525,N_493,N_451);
xor U526 (N_526,N_432,N_471);
or U527 (N_527,N_406,N_478);
xnor U528 (N_528,N_400,N_473);
and U529 (N_529,N_403,N_436);
and U530 (N_530,N_486,N_465);
nand U531 (N_531,N_424,N_407);
and U532 (N_532,N_496,N_431);
or U533 (N_533,N_415,N_489);
xor U534 (N_534,N_459,N_467);
xor U535 (N_535,N_411,N_445);
nand U536 (N_536,N_468,N_490);
or U537 (N_537,N_429,N_419);
nand U538 (N_538,N_439,N_437);
and U539 (N_539,N_422,N_418);
xor U540 (N_540,N_463,N_475);
and U541 (N_541,N_477,N_413);
and U542 (N_542,N_440,N_442);
or U543 (N_543,N_416,N_474);
and U544 (N_544,N_447,N_460);
xor U545 (N_545,N_452,N_405);
xnor U546 (N_546,N_462,N_458);
and U547 (N_547,N_495,N_435);
xnor U548 (N_548,N_466,N_476);
or U549 (N_549,N_414,N_482);
nand U550 (N_550,N_452,N_408);
xor U551 (N_551,N_413,N_419);
and U552 (N_552,N_445,N_457);
and U553 (N_553,N_440,N_463);
nand U554 (N_554,N_400,N_463);
nand U555 (N_555,N_441,N_480);
xnor U556 (N_556,N_404,N_427);
xnor U557 (N_557,N_429,N_482);
nand U558 (N_558,N_407,N_414);
or U559 (N_559,N_435,N_476);
and U560 (N_560,N_457,N_418);
xnor U561 (N_561,N_431,N_429);
nand U562 (N_562,N_486,N_424);
and U563 (N_563,N_465,N_480);
xnor U564 (N_564,N_440,N_453);
or U565 (N_565,N_479,N_448);
and U566 (N_566,N_430,N_444);
nand U567 (N_567,N_453,N_457);
xor U568 (N_568,N_402,N_451);
nor U569 (N_569,N_453,N_495);
xor U570 (N_570,N_401,N_418);
or U571 (N_571,N_495,N_488);
xnor U572 (N_572,N_438,N_455);
nor U573 (N_573,N_426,N_444);
nand U574 (N_574,N_473,N_489);
nand U575 (N_575,N_458,N_423);
nor U576 (N_576,N_478,N_463);
nand U577 (N_577,N_429,N_488);
nand U578 (N_578,N_417,N_475);
nor U579 (N_579,N_480,N_482);
xor U580 (N_580,N_419,N_448);
nor U581 (N_581,N_467,N_430);
or U582 (N_582,N_458,N_420);
nand U583 (N_583,N_479,N_451);
or U584 (N_584,N_483,N_476);
or U585 (N_585,N_449,N_402);
nand U586 (N_586,N_433,N_493);
or U587 (N_587,N_487,N_481);
and U588 (N_588,N_467,N_441);
xnor U589 (N_589,N_498,N_476);
xor U590 (N_590,N_426,N_462);
and U591 (N_591,N_406,N_425);
nand U592 (N_592,N_476,N_426);
nand U593 (N_593,N_439,N_493);
nand U594 (N_594,N_454,N_411);
nor U595 (N_595,N_488,N_467);
and U596 (N_596,N_491,N_473);
or U597 (N_597,N_403,N_416);
or U598 (N_598,N_401,N_470);
or U599 (N_599,N_404,N_489);
nand U600 (N_600,N_501,N_542);
nor U601 (N_601,N_543,N_584);
nor U602 (N_602,N_582,N_589);
and U603 (N_603,N_522,N_503);
nand U604 (N_604,N_512,N_573);
and U605 (N_605,N_572,N_570);
xor U606 (N_606,N_586,N_556);
or U607 (N_607,N_544,N_557);
or U608 (N_608,N_587,N_525);
xnor U609 (N_609,N_599,N_576);
xor U610 (N_610,N_554,N_541);
nand U611 (N_611,N_555,N_546);
or U612 (N_612,N_514,N_538);
or U613 (N_613,N_545,N_517);
nor U614 (N_614,N_547,N_500);
xor U615 (N_615,N_561,N_595);
or U616 (N_616,N_575,N_533);
nor U617 (N_617,N_578,N_524);
nor U618 (N_618,N_559,N_574);
nor U619 (N_619,N_564,N_529);
nand U620 (N_620,N_571,N_532);
xnor U621 (N_621,N_560,N_539);
and U622 (N_622,N_506,N_523);
nor U623 (N_623,N_536,N_558);
xor U624 (N_624,N_567,N_511);
xor U625 (N_625,N_566,N_530);
or U626 (N_626,N_513,N_552);
nor U627 (N_627,N_568,N_548);
xor U628 (N_628,N_594,N_509);
nor U629 (N_629,N_592,N_553);
or U630 (N_630,N_504,N_585);
nand U631 (N_631,N_597,N_593);
nand U632 (N_632,N_596,N_515);
nand U633 (N_633,N_535,N_526);
nor U634 (N_634,N_588,N_521);
nor U635 (N_635,N_540,N_510);
xnor U636 (N_636,N_563,N_565);
and U637 (N_637,N_508,N_598);
xor U638 (N_638,N_516,N_583);
and U639 (N_639,N_519,N_591);
nand U640 (N_640,N_562,N_505);
or U641 (N_641,N_537,N_527);
or U642 (N_642,N_577,N_581);
and U643 (N_643,N_569,N_518);
and U644 (N_644,N_528,N_551);
and U645 (N_645,N_534,N_502);
and U646 (N_646,N_579,N_550);
xor U647 (N_647,N_520,N_531);
and U648 (N_648,N_590,N_549);
nand U649 (N_649,N_507,N_580);
nor U650 (N_650,N_544,N_518);
and U651 (N_651,N_516,N_592);
xnor U652 (N_652,N_529,N_538);
xor U653 (N_653,N_531,N_549);
and U654 (N_654,N_519,N_513);
and U655 (N_655,N_515,N_501);
and U656 (N_656,N_562,N_573);
xnor U657 (N_657,N_508,N_567);
nand U658 (N_658,N_550,N_594);
nor U659 (N_659,N_583,N_566);
nor U660 (N_660,N_529,N_579);
xnor U661 (N_661,N_511,N_579);
nor U662 (N_662,N_526,N_552);
or U663 (N_663,N_599,N_555);
nor U664 (N_664,N_502,N_514);
and U665 (N_665,N_505,N_513);
or U666 (N_666,N_553,N_535);
xor U667 (N_667,N_514,N_565);
and U668 (N_668,N_512,N_582);
xor U669 (N_669,N_522,N_537);
nor U670 (N_670,N_575,N_540);
nand U671 (N_671,N_550,N_575);
and U672 (N_672,N_589,N_519);
nor U673 (N_673,N_580,N_518);
or U674 (N_674,N_561,N_518);
xnor U675 (N_675,N_571,N_522);
or U676 (N_676,N_540,N_544);
nor U677 (N_677,N_593,N_537);
or U678 (N_678,N_553,N_556);
nor U679 (N_679,N_500,N_540);
or U680 (N_680,N_578,N_564);
and U681 (N_681,N_521,N_563);
or U682 (N_682,N_518,N_571);
and U683 (N_683,N_589,N_588);
or U684 (N_684,N_582,N_525);
nand U685 (N_685,N_594,N_581);
xnor U686 (N_686,N_500,N_544);
nor U687 (N_687,N_519,N_599);
nand U688 (N_688,N_594,N_582);
and U689 (N_689,N_549,N_573);
nor U690 (N_690,N_582,N_584);
xnor U691 (N_691,N_573,N_502);
nor U692 (N_692,N_525,N_559);
or U693 (N_693,N_524,N_522);
or U694 (N_694,N_586,N_532);
nand U695 (N_695,N_528,N_545);
or U696 (N_696,N_575,N_544);
or U697 (N_697,N_523,N_588);
nand U698 (N_698,N_564,N_519);
or U699 (N_699,N_578,N_577);
or U700 (N_700,N_616,N_699);
xnor U701 (N_701,N_676,N_696);
or U702 (N_702,N_662,N_625);
xor U703 (N_703,N_621,N_689);
or U704 (N_704,N_612,N_698);
nor U705 (N_705,N_617,N_648);
nor U706 (N_706,N_661,N_618);
or U707 (N_707,N_629,N_695);
xnor U708 (N_708,N_620,N_645);
or U709 (N_709,N_670,N_659);
nand U710 (N_710,N_655,N_614);
nand U711 (N_711,N_631,N_680);
and U712 (N_712,N_624,N_690);
nor U713 (N_713,N_669,N_691);
and U714 (N_714,N_678,N_627);
or U715 (N_715,N_644,N_665);
or U716 (N_716,N_675,N_677);
nand U717 (N_717,N_652,N_600);
nand U718 (N_718,N_609,N_672);
nor U719 (N_719,N_651,N_615);
xor U720 (N_720,N_607,N_632);
or U721 (N_721,N_673,N_637);
and U722 (N_722,N_692,N_602);
or U723 (N_723,N_608,N_643);
and U724 (N_724,N_639,N_606);
or U725 (N_725,N_635,N_623);
or U726 (N_726,N_656,N_664);
xnor U727 (N_727,N_647,N_681);
or U728 (N_728,N_610,N_697);
nor U729 (N_729,N_693,N_634);
nor U730 (N_730,N_622,N_694);
and U731 (N_731,N_613,N_605);
nand U732 (N_732,N_653,N_650);
or U733 (N_733,N_619,N_658);
or U734 (N_734,N_649,N_671);
or U735 (N_735,N_601,N_630);
xor U736 (N_736,N_667,N_638);
or U737 (N_737,N_603,N_626);
and U738 (N_738,N_683,N_666);
or U739 (N_739,N_657,N_687);
nor U740 (N_740,N_685,N_636);
nor U741 (N_741,N_668,N_663);
or U742 (N_742,N_604,N_641);
nand U743 (N_743,N_688,N_611);
and U744 (N_744,N_640,N_654);
xor U745 (N_745,N_679,N_684);
nand U746 (N_746,N_633,N_642);
xor U747 (N_747,N_646,N_674);
or U748 (N_748,N_628,N_686);
nand U749 (N_749,N_682,N_660);
nand U750 (N_750,N_605,N_654);
or U751 (N_751,N_604,N_633);
nand U752 (N_752,N_696,N_681);
nor U753 (N_753,N_642,N_639);
and U754 (N_754,N_695,N_622);
nand U755 (N_755,N_675,N_648);
nand U756 (N_756,N_652,N_651);
or U757 (N_757,N_635,N_645);
nand U758 (N_758,N_661,N_615);
xor U759 (N_759,N_641,N_600);
or U760 (N_760,N_641,N_633);
xnor U761 (N_761,N_642,N_652);
nand U762 (N_762,N_693,N_610);
and U763 (N_763,N_641,N_681);
nand U764 (N_764,N_656,N_619);
and U765 (N_765,N_605,N_694);
or U766 (N_766,N_627,N_606);
xnor U767 (N_767,N_621,N_639);
and U768 (N_768,N_699,N_618);
or U769 (N_769,N_687,N_695);
and U770 (N_770,N_619,N_691);
xor U771 (N_771,N_641,N_601);
or U772 (N_772,N_663,N_682);
nand U773 (N_773,N_619,N_685);
xor U774 (N_774,N_620,N_626);
nand U775 (N_775,N_643,N_684);
nor U776 (N_776,N_622,N_634);
nor U777 (N_777,N_625,N_687);
nor U778 (N_778,N_655,N_652);
nor U779 (N_779,N_665,N_657);
nor U780 (N_780,N_670,N_680);
nand U781 (N_781,N_683,N_682);
and U782 (N_782,N_636,N_607);
and U783 (N_783,N_664,N_642);
nor U784 (N_784,N_695,N_605);
and U785 (N_785,N_647,N_636);
xor U786 (N_786,N_613,N_604);
or U787 (N_787,N_664,N_662);
or U788 (N_788,N_686,N_601);
nor U789 (N_789,N_606,N_616);
and U790 (N_790,N_626,N_624);
nand U791 (N_791,N_647,N_642);
xnor U792 (N_792,N_641,N_685);
nor U793 (N_793,N_609,N_677);
or U794 (N_794,N_663,N_603);
nand U795 (N_795,N_655,N_647);
and U796 (N_796,N_623,N_687);
nor U797 (N_797,N_619,N_625);
and U798 (N_798,N_655,N_613);
or U799 (N_799,N_663,N_690);
nor U800 (N_800,N_734,N_767);
nor U801 (N_801,N_788,N_709);
xnor U802 (N_802,N_745,N_781);
or U803 (N_803,N_713,N_750);
or U804 (N_804,N_756,N_730);
nand U805 (N_805,N_772,N_744);
and U806 (N_806,N_711,N_741);
or U807 (N_807,N_752,N_755);
nor U808 (N_808,N_776,N_719);
and U809 (N_809,N_733,N_712);
or U810 (N_810,N_770,N_739);
xnor U811 (N_811,N_717,N_722);
and U812 (N_812,N_738,N_701);
nor U813 (N_813,N_779,N_715);
xnor U814 (N_814,N_725,N_736);
nand U815 (N_815,N_758,N_797);
xor U816 (N_816,N_787,N_792);
nor U817 (N_817,N_791,N_740);
or U818 (N_818,N_794,N_746);
xnor U819 (N_819,N_714,N_751);
nand U820 (N_820,N_793,N_798);
xor U821 (N_821,N_773,N_768);
and U822 (N_822,N_769,N_726);
or U823 (N_823,N_729,N_749);
nor U824 (N_824,N_783,N_735);
nor U825 (N_825,N_766,N_778);
and U826 (N_826,N_782,N_796);
or U827 (N_827,N_720,N_742);
nand U828 (N_828,N_759,N_732);
nor U829 (N_829,N_723,N_774);
and U830 (N_830,N_789,N_762);
or U831 (N_831,N_703,N_771);
xor U832 (N_832,N_761,N_799);
xor U833 (N_833,N_702,N_737);
xor U834 (N_834,N_748,N_775);
xnor U835 (N_835,N_753,N_710);
or U836 (N_836,N_777,N_707);
nand U837 (N_837,N_747,N_786);
nor U838 (N_838,N_706,N_760);
and U839 (N_839,N_757,N_727);
or U840 (N_840,N_764,N_705);
and U841 (N_841,N_718,N_716);
xor U842 (N_842,N_724,N_795);
nor U843 (N_843,N_790,N_763);
and U844 (N_844,N_708,N_784);
xor U845 (N_845,N_728,N_765);
xor U846 (N_846,N_731,N_754);
nor U847 (N_847,N_704,N_785);
or U848 (N_848,N_743,N_780);
nor U849 (N_849,N_700,N_721);
xnor U850 (N_850,N_788,N_780);
xor U851 (N_851,N_717,N_748);
xnor U852 (N_852,N_712,N_768);
or U853 (N_853,N_793,N_770);
or U854 (N_854,N_711,N_769);
nor U855 (N_855,N_725,N_721);
xnor U856 (N_856,N_735,N_740);
and U857 (N_857,N_742,N_709);
and U858 (N_858,N_775,N_709);
nor U859 (N_859,N_763,N_731);
nand U860 (N_860,N_792,N_741);
or U861 (N_861,N_757,N_728);
xnor U862 (N_862,N_787,N_786);
nand U863 (N_863,N_730,N_721);
or U864 (N_864,N_788,N_784);
and U865 (N_865,N_749,N_722);
or U866 (N_866,N_754,N_737);
xnor U867 (N_867,N_754,N_778);
or U868 (N_868,N_786,N_705);
nand U869 (N_869,N_715,N_751);
nor U870 (N_870,N_742,N_743);
nor U871 (N_871,N_782,N_771);
xnor U872 (N_872,N_758,N_735);
xor U873 (N_873,N_749,N_741);
or U874 (N_874,N_793,N_721);
nand U875 (N_875,N_740,N_743);
or U876 (N_876,N_729,N_734);
xnor U877 (N_877,N_725,N_795);
nor U878 (N_878,N_777,N_714);
and U879 (N_879,N_792,N_711);
or U880 (N_880,N_728,N_791);
nand U881 (N_881,N_725,N_744);
nand U882 (N_882,N_716,N_711);
xnor U883 (N_883,N_707,N_763);
nor U884 (N_884,N_769,N_744);
or U885 (N_885,N_772,N_737);
and U886 (N_886,N_760,N_769);
or U887 (N_887,N_718,N_711);
and U888 (N_888,N_760,N_795);
and U889 (N_889,N_707,N_792);
and U890 (N_890,N_714,N_700);
and U891 (N_891,N_736,N_740);
or U892 (N_892,N_744,N_700);
nor U893 (N_893,N_770,N_776);
or U894 (N_894,N_795,N_706);
or U895 (N_895,N_719,N_796);
nand U896 (N_896,N_781,N_705);
and U897 (N_897,N_732,N_772);
and U898 (N_898,N_722,N_718);
or U899 (N_899,N_740,N_705);
nor U900 (N_900,N_800,N_841);
or U901 (N_901,N_856,N_837);
nand U902 (N_902,N_876,N_882);
xnor U903 (N_903,N_858,N_803);
and U904 (N_904,N_849,N_813);
or U905 (N_905,N_854,N_801);
or U906 (N_906,N_896,N_884);
and U907 (N_907,N_843,N_853);
nand U908 (N_908,N_822,N_833);
or U909 (N_909,N_814,N_870);
and U910 (N_910,N_834,N_869);
or U911 (N_911,N_802,N_805);
nand U912 (N_912,N_825,N_865);
xor U913 (N_913,N_809,N_880);
nand U914 (N_914,N_894,N_844);
nand U915 (N_915,N_828,N_892);
or U916 (N_916,N_845,N_835);
xor U917 (N_917,N_857,N_860);
nor U918 (N_918,N_872,N_831);
or U919 (N_919,N_887,N_846);
and U920 (N_920,N_879,N_851);
or U921 (N_921,N_836,N_818);
nor U922 (N_922,N_895,N_890);
and U923 (N_923,N_859,N_889);
and U924 (N_924,N_830,N_866);
or U925 (N_925,N_863,N_823);
and U926 (N_926,N_810,N_815);
nand U927 (N_927,N_886,N_839);
nand U928 (N_928,N_867,N_838);
nand U929 (N_929,N_899,N_832);
nor U930 (N_930,N_883,N_807);
nand U931 (N_931,N_855,N_874);
nor U932 (N_932,N_881,N_861);
or U933 (N_933,N_868,N_864);
xor U934 (N_934,N_873,N_824);
nor U935 (N_935,N_885,N_804);
or U936 (N_936,N_875,N_847);
and U937 (N_937,N_898,N_820);
xor U938 (N_938,N_897,N_842);
or U939 (N_939,N_871,N_852);
or U940 (N_940,N_808,N_806);
xor U941 (N_941,N_817,N_878);
xor U942 (N_942,N_850,N_826);
or U943 (N_943,N_893,N_840);
nand U944 (N_944,N_812,N_891);
or U945 (N_945,N_829,N_862);
xor U946 (N_946,N_827,N_811);
nor U947 (N_947,N_888,N_816);
and U948 (N_948,N_819,N_821);
xor U949 (N_949,N_877,N_848);
and U950 (N_950,N_872,N_886);
nand U951 (N_951,N_862,N_818);
nor U952 (N_952,N_870,N_873);
xnor U953 (N_953,N_896,N_857);
nand U954 (N_954,N_883,N_816);
xnor U955 (N_955,N_814,N_880);
and U956 (N_956,N_884,N_889);
nand U957 (N_957,N_883,N_840);
xnor U958 (N_958,N_815,N_852);
or U959 (N_959,N_812,N_845);
xnor U960 (N_960,N_809,N_810);
and U961 (N_961,N_899,N_884);
nand U962 (N_962,N_843,N_866);
nor U963 (N_963,N_865,N_848);
or U964 (N_964,N_865,N_891);
xor U965 (N_965,N_818,N_841);
nor U966 (N_966,N_843,N_841);
xnor U967 (N_967,N_831,N_815);
nor U968 (N_968,N_894,N_860);
and U969 (N_969,N_840,N_839);
and U970 (N_970,N_896,N_809);
nand U971 (N_971,N_846,N_879);
nand U972 (N_972,N_861,N_848);
xor U973 (N_973,N_821,N_834);
or U974 (N_974,N_845,N_898);
nor U975 (N_975,N_890,N_891);
or U976 (N_976,N_859,N_808);
or U977 (N_977,N_895,N_827);
or U978 (N_978,N_871,N_846);
nor U979 (N_979,N_834,N_820);
xnor U980 (N_980,N_800,N_879);
nor U981 (N_981,N_884,N_853);
nor U982 (N_982,N_899,N_882);
and U983 (N_983,N_863,N_890);
nor U984 (N_984,N_863,N_831);
or U985 (N_985,N_835,N_828);
nor U986 (N_986,N_814,N_833);
nor U987 (N_987,N_852,N_837);
xor U988 (N_988,N_844,N_813);
or U989 (N_989,N_892,N_885);
and U990 (N_990,N_828,N_846);
xor U991 (N_991,N_830,N_826);
or U992 (N_992,N_886,N_815);
xnor U993 (N_993,N_881,N_830);
xor U994 (N_994,N_864,N_847);
or U995 (N_995,N_888,N_889);
or U996 (N_996,N_838,N_811);
or U997 (N_997,N_838,N_816);
nand U998 (N_998,N_894,N_815);
or U999 (N_999,N_866,N_818);
and U1000 (N_1000,N_993,N_956);
nand U1001 (N_1001,N_997,N_982);
or U1002 (N_1002,N_947,N_935);
nor U1003 (N_1003,N_964,N_925);
nor U1004 (N_1004,N_910,N_962);
nor U1005 (N_1005,N_995,N_950);
xor U1006 (N_1006,N_971,N_907);
nor U1007 (N_1007,N_954,N_920);
xor U1008 (N_1008,N_932,N_970);
nor U1009 (N_1009,N_980,N_938);
or U1010 (N_1010,N_974,N_972);
xor U1011 (N_1011,N_923,N_922);
or U1012 (N_1012,N_904,N_916);
and U1013 (N_1013,N_912,N_988);
and U1014 (N_1014,N_983,N_967);
and U1015 (N_1015,N_986,N_944);
xnor U1016 (N_1016,N_943,N_991);
xor U1017 (N_1017,N_978,N_900);
and U1018 (N_1018,N_939,N_945);
nor U1019 (N_1019,N_946,N_994);
xnor U1020 (N_1020,N_917,N_968);
nand U1021 (N_1021,N_975,N_998);
and U1022 (N_1022,N_941,N_958);
or U1023 (N_1023,N_934,N_985);
xor U1024 (N_1024,N_911,N_973);
or U1025 (N_1025,N_955,N_931);
nor U1026 (N_1026,N_908,N_927);
or U1027 (N_1027,N_928,N_996);
and U1028 (N_1028,N_942,N_914);
nand U1029 (N_1029,N_913,N_953);
and U1030 (N_1030,N_905,N_919);
xor U1031 (N_1031,N_940,N_948);
nor U1032 (N_1032,N_992,N_930);
xor U1033 (N_1033,N_933,N_989);
or U1034 (N_1034,N_987,N_960);
nand U1035 (N_1035,N_952,N_961);
nand U1036 (N_1036,N_924,N_909);
or U1037 (N_1037,N_921,N_918);
xor U1038 (N_1038,N_929,N_984);
xor U1039 (N_1039,N_959,N_915);
and U1040 (N_1040,N_963,N_965);
or U1041 (N_1041,N_999,N_949);
nand U1042 (N_1042,N_957,N_926);
nand U1043 (N_1043,N_976,N_990);
and U1044 (N_1044,N_937,N_966);
and U1045 (N_1045,N_981,N_936);
or U1046 (N_1046,N_969,N_906);
or U1047 (N_1047,N_977,N_979);
nor U1048 (N_1048,N_901,N_903);
and U1049 (N_1049,N_902,N_951);
xor U1050 (N_1050,N_907,N_982);
and U1051 (N_1051,N_937,N_916);
nor U1052 (N_1052,N_992,N_957);
xor U1053 (N_1053,N_985,N_994);
xnor U1054 (N_1054,N_983,N_923);
and U1055 (N_1055,N_921,N_957);
and U1056 (N_1056,N_905,N_950);
or U1057 (N_1057,N_970,N_949);
xor U1058 (N_1058,N_939,N_973);
and U1059 (N_1059,N_987,N_929);
nor U1060 (N_1060,N_970,N_990);
nor U1061 (N_1061,N_950,N_971);
nand U1062 (N_1062,N_914,N_924);
and U1063 (N_1063,N_904,N_939);
nor U1064 (N_1064,N_983,N_950);
nand U1065 (N_1065,N_941,N_966);
or U1066 (N_1066,N_968,N_907);
or U1067 (N_1067,N_931,N_919);
xnor U1068 (N_1068,N_995,N_912);
or U1069 (N_1069,N_958,N_927);
and U1070 (N_1070,N_957,N_960);
or U1071 (N_1071,N_930,N_974);
xor U1072 (N_1072,N_999,N_950);
or U1073 (N_1073,N_952,N_984);
xor U1074 (N_1074,N_982,N_996);
and U1075 (N_1075,N_921,N_919);
nor U1076 (N_1076,N_975,N_928);
nor U1077 (N_1077,N_960,N_918);
nor U1078 (N_1078,N_950,N_917);
and U1079 (N_1079,N_917,N_980);
or U1080 (N_1080,N_937,N_985);
nand U1081 (N_1081,N_952,N_960);
and U1082 (N_1082,N_938,N_978);
nor U1083 (N_1083,N_964,N_953);
nand U1084 (N_1084,N_924,N_935);
or U1085 (N_1085,N_931,N_959);
and U1086 (N_1086,N_971,N_973);
and U1087 (N_1087,N_983,N_982);
and U1088 (N_1088,N_982,N_954);
nor U1089 (N_1089,N_940,N_966);
or U1090 (N_1090,N_961,N_920);
or U1091 (N_1091,N_944,N_912);
nor U1092 (N_1092,N_904,N_994);
or U1093 (N_1093,N_930,N_958);
or U1094 (N_1094,N_921,N_996);
and U1095 (N_1095,N_957,N_915);
xor U1096 (N_1096,N_967,N_969);
nor U1097 (N_1097,N_922,N_987);
or U1098 (N_1098,N_988,N_914);
or U1099 (N_1099,N_998,N_990);
xnor U1100 (N_1100,N_1092,N_1020);
or U1101 (N_1101,N_1038,N_1067);
or U1102 (N_1102,N_1028,N_1061);
xor U1103 (N_1103,N_1065,N_1095);
xor U1104 (N_1104,N_1001,N_1085);
or U1105 (N_1105,N_1052,N_1046);
nor U1106 (N_1106,N_1081,N_1023);
nand U1107 (N_1107,N_1073,N_1053);
xnor U1108 (N_1108,N_1074,N_1014);
or U1109 (N_1109,N_1041,N_1033);
xnor U1110 (N_1110,N_1083,N_1003);
nor U1111 (N_1111,N_1031,N_1090);
nand U1112 (N_1112,N_1040,N_1034);
xnor U1113 (N_1113,N_1025,N_1070);
xnor U1114 (N_1114,N_1068,N_1088);
xnor U1115 (N_1115,N_1050,N_1045);
or U1116 (N_1116,N_1086,N_1036);
or U1117 (N_1117,N_1013,N_1079);
nand U1118 (N_1118,N_1099,N_1048);
nor U1119 (N_1119,N_1010,N_1017);
nor U1120 (N_1120,N_1032,N_1080);
xor U1121 (N_1121,N_1026,N_1043);
nor U1122 (N_1122,N_1063,N_1098);
and U1123 (N_1123,N_1071,N_1066);
xor U1124 (N_1124,N_1054,N_1089);
nand U1125 (N_1125,N_1024,N_1042);
nor U1126 (N_1126,N_1057,N_1072);
nand U1127 (N_1127,N_1064,N_1058);
and U1128 (N_1128,N_1047,N_1044);
xor U1129 (N_1129,N_1075,N_1007);
xor U1130 (N_1130,N_1097,N_1027);
xnor U1131 (N_1131,N_1078,N_1082);
xnor U1132 (N_1132,N_1018,N_1002);
nand U1133 (N_1133,N_1091,N_1029);
nand U1134 (N_1134,N_1076,N_1004);
xnor U1135 (N_1135,N_1016,N_1060);
nor U1136 (N_1136,N_1062,N_1000);
or U1137 (N_1137,N_1077,N_1015);
and U1138 (N_1138,N_1051,N_1039);
nand U1139 (N_1139,N_1009,N_1035);
or U1140 (N_1140,N_1059,N_1093);
xor U1141 (N_1141,N_1008,N_1096);
xor U1142 (N_1142,N_1055,N_1019);
or U1143 (N_1143,N_1030,N_1056);
or U1144 (N_1144,N_1022,N_1087);
or U1145 (N_1145,N_1021,N_1011);
and U1146 (N_1146,N_1037,N_1084);
or U1147 (N_1147,N_1094,N_1049);
xor U1148 (N_1148,N_1005,N_1012);
nor U1149 (N_1149,N_1006,N_1069);
or U1150 (N_1150,N_1011,N_1043);
or U1151 (N_1151,N_1048,N_1057);
and U1152 (N_1152,N_1044,N_1030);
nor U1153 (N_1153,N_1003,N_1052);
nor U1154 (N_1154,N_1051,N_1002);
nor U1155 (N_1155,N_1015,N_1085);
and U1156 (N_1156,N_1013,N_1072);
xor U1157 (N_1157,N_1042,N_1099);
or U1158 (N_1158,N_1011,N_1098);
and U1159 (N_1159,N_1045,N_1071);
or U1160 (N_1160,N_1043,N_1073);
nand U1161 (N_1161,N_1068,N_1052);
xor U1162 (N_1162,N_1000,N_1049);
xnor U1163 (N_1163,N_1083,N_1044);
nor U1164 (N_1164,N_1027,N_1005);
nand U1165 (N_1165,N_1004,N_1010);
and U1166 (N_1166,N_1024,N_1098);
nor U1167 (N_1167,N_1042,N_1041);
and U1168 (N_1168,N_1060,N_1028);
nand U1169 (N_1169,N_1083,N_1059);
nand U1170 (N_1170,N_1061,N_1011);
xnor U1171 (N_1171,N_1056,N_1058);
nor U1172 (N_1172,N_1018,N_1011);
and U1173 (N_1173,N_1000,N_1045);
nand U1174 (N_1174,N_1010,N_1058);
and U1175 (N_1175,N_1004,N_1021);
and U1176 (N_1176,N_1057,N_1010);
nor U1177 (N_1177,N_1081,N_1075);
nor U1178 (N_1178,N_1011,N_1053);
nand U1179 (N_1179,N_1073,N_1067);
nor U1180 (N_1180,N_1056,N_1051);
nor U1181 (N_1181,N_1002,N_1026);
xor U1182 (N_1182,N_1091,N_1013);
or U1183 (N_1183,N_1067,N_1072);
xor U1184 (N_1184,N_1026,N_1036);
and U1185 (N_1185,N_1098,N_1043);
and U1186 (N_1186,N_1008,N_1054);
and U1187 (N_1187,N_1025,N_1017);
and U1188 (N_1188,N_1016,N_1014);
nand U1189 (N_1189,N_1092,N_1063);
nand U1190 (N_1190,N_1020,N_1046);
or U1191 (N_1191,N_1016,N_1088);
nor U1192 (N_1192,N_1034,N_1061);
xnor U1193 (N_1193,N_1092,N_1031);
nor U1194 (N_1194,N_1047,N_1000);
xnor U1195 (N_1195,N_1033,N_1035);
nor U1196 (N_1196,N_1081,N_1009);
nor U1197 (N_1197,N_1050,N_1025);
or U1198 (N_1198,N_1059,N_1096);
nor U1199 (N_1199,N_1073,N_1027);
and U1200 (N_1200,N_1153,N_1149);
and U1201 (N_1201,N_1113,N_1126);
and U1202 (N_1202,N_1105,N_1160);
nor U1203 (N_1203,N_1145,N_1142);
or U1204 (N_1204,N_1106,N_1127);
xor U1205 (N_1205,N_1118,N_1128);
nor U1206 (N_1206,N_1159,N_1176);
or U1207 (N_1207,N_1165,N_1107);
or U1208 (N_1208,N_1136,N_1100);
or U1209 (N_1209,N_1111,N_1148);
nand U1210 (N_1210,N_1190,N_1140);
xnor U1211 (N_1211,N_1110,N_1166);
xnor U1212 (N_1212,N_1169,N_1121);
nand U1213 (N_1213,N_1180,N_1115);
nand U1214 (N_1214,N_1151,N_1167);
nand U1215 (N_1215,N_1132,N_1137);
nor U1216 (N_1216,N_1173,N_1189);
or U1217 (N_1217,N_1187,N_1161);
xnor U1218 (N_1218,N_1184,N_1181);
nor U1219 (N_1219,N_1168,N_1102);
and U1220 (N_1220,N_1114,N_1122);
or U1221 (N_1221,N_1163,N_1125);
xnor U1222 (N_1222,N_1141,N_1119);
or U1223 (N_1223,N_1124,N_1199);
xor U1224 (N_1224,N_1195,N_1157);
nand U1225 (N_1225,N_1175,N_1108);
nand U1226 (N_1226,N_1154,N_1133);
and U1227 (N_1227,N_1117,N_1155);
xor U1228 (N_1228,N_1150,N_1183);
or U1229 (N_1229,N_1129,N_1179);
and U1230 (N_1230,N_1198,N_1112);
nand U1231 (N_1231,N_1177,N_1156);
xnor U1232 (N_1232,N_1186,N_1101);
and U1233 (N_1233,N_1146,N_1162);
xor U1234 (N_1234,N_1109,N_1196);
nor U1235 (N_1235,N_1130,N_1123);
and U1236 (N_1236,N_1116,N_1143);
nand U1237 (N_1237,N_1194,N_1171);
nor U1238 (N_1238,N_1164,N_1131);
nand U1239 (N_1239,N_1158,N_1104);
xnor U1240 (N_1240,N_1193,N_1135);
nor U1241 (N_1241,N_1192,N_1188);
and U1242 (N_1242,N_1185,N_1152);
nand U1243 (N_1243,N_1134,N_1174);
xnor U1244 (N_1244,N_1178,N_1170);
nand U1245 (N_1245,N_1147,N_1138);
nor U1246 (N_1246,N_1144,N_1172);
nand U1247 (N_1247,N_1182,N_1139);
and U1248 (N_1248,N_1197,N_1103);
nand U1249 (N_1249,N_1191,N_1120);
nand U1250 (N_1250,N_1127,N_1144);
xnor U1251 (N_1251,N_1164,N_1105);
nor U1252 (N_1252,N_1119,N_1163);
and U1253 (N_1253,N_1122,N_1127);
or U1254 (N_1254,N_1138,N_1167);
nor U1255 (N_1255,N_1151,N_1103);
xnor U1256 (N_1256,N_1197,N_1143);
nand U1257 (N_1257,N_1183,N_1130);
and U1258 (N_1258,N_1169,N_1109);
or U1259 (N_1259,N_1179,N_1170);
xnor U1260 (N_1260,N_1157,N_1142);
or U1261 (N_1261,N_1103,N_1167);
and U1262 (N_1262,N_1104,N_1175);
nand U1263 (N_1263,N_1191,N_1100);
and U1264 (N_1264,N_1178,N_1189);
or U1265 (N_1265,N_1177,N_1158);
nand U1266 (N_1266,N_1139,N_1148);
xnor U1267 (N_1267,N_1176,N_1178);
nor U1268 (N_1268,N_1176,N_1135);
xnor U1269 (N_1269,N_1164,N_1151);
and U1270 (N_1270,N_1192,N_1118);
xor U1271 (N_1271,N_1116,N_1162);
xor U1272 (N_1272,N_1159,N_1130);
nor U1273 (N_1273,N_1162,N_1137);
xnor U1274 (N_1274,N_1177,N_1175);
nand U1275 (N_1275,N_1122,N_1181);
or U1276 (N_1276,N_1160,N_1122);
nor U1277 (N_1277,N_1181,N_1183);
and U1278 (N_1278,N_1103,N_1190);
or U1279 (N_1279,N_1144,N_1197);
nand U1280 (N_1280,N_1160,N_1140);
and U1281 (N_1281,N_1136,N_1183);
xor U1282 (N_1282,N_1171,N_1163);
and U1283 (N_1283,N_1166,N_1142);
nor U1284 (N_1284,N_1130,N_1179);
or U1285 (N_1285,N_1169,N_1135);
or U1286 (N_1286,N_1141,N_1132);
xor U1287 (N_1287,N_1104,N_1174);
and U1288 (N_1288,N_1172,N_1195);
xnor U1289 (N_1289,N_1159,N_1106);
nor U1290 (N_1290,N_1180,N_1133);
nand U1291 (N_1291,N_1197,N_1113);
or U1292 (N_1292,N_1193,N_1103);
nor U1293 (N_1293,N_1160,N_1121);
and U1294 (N_1294,N_1102,N_1158);
nand U1295 (N_1295,N_1193,N_1154);
nand U1296 (N_1296,N_1137,N_1143);
xnor U1297 (N_1297,N_1153,N_1138);
and U1298 (N_1298,N_1156,N_1112);
nand U1299 (N_1299,N_1183,N_1169);
and U1300 (N_1300,N_1270,N_1236);
and U1301 (N_1301,N_1211,N_1255);
and U1302 (N_1302,N_1220,N_1275);
and U1303 (N_1303,N_1210,N_1205);
xnor U1304 (N_1304,N_1250,N_1268);
nand U1305 (N_1305,N_1269,N_1285);
or U1306 (N_1306,N_1291,N_1249);
or U1307 (N_1307,N_1243,N_1217);
and U1308 (N_1308,N_1200,N_1231);
or U1309 (N_1309,N_1296,N_1224);
xnor U1310 (N_1310,N_1203,N_1218);
or U1311 (N_1311,N_1276,N_1264);
and U1312 (N_1312,N_1265,N_1233);
and U1313 (N_1313,N_1204,N_1207);
nand U1314 (N_1314,N_1241,N_1214);
nor U1315 (N_1315,N_1242,N_1295);
or U1316 (N_1316,N_1212,N_1286);
and U1317 (N_1317,N_1202,N_1253);
xnor U1318 (N_1318,N_1280,N_1279);
nor U1319 (N_1319,N_1260,N_1299);
nor U1320 (N_1320,N_1201,N_1257);
xor U1321 (N_1321,N_1283,N_1219);
xnor U1322 (N_1322,N_1235,N_1262);
nand U1323 (N_1323,N_1272,N_1254);
and U1324 (N_1324,N_1267,N_1290);
xnor U1325 (N_1325,N_1232,N_1245);
nor U1326 (N_1326,N_1208,N_1282);
nand U1327 (N_1327,N_1263,N_1225);
and U1328 (N_1328,N_1281,N_1251);
nand U1329 (N_1329,N_1237,N_1256);
or U1330 (N_1330,N_1221,N_1216);
xnor U1331 (N_1331,N_1238,N_1229);
nor U1332 (N_1332,N_1252,N_1215);
or U1333 (N_1333,N_1234,N_1209);
and U1334 (N_1334,N_1248,N_1230);
or U1335 (N_1335,N_1259,N_1293);
and U1336 (N_1336,N_1261,N_1222);
xor U1337 (N_1337,N_1289,N_1223);
xnor U1338 (N_1338,N_1298,N_1297);
and U1339 (N_1339,N_1240,N_1206);
xnor U1340 (N_1340,N_1294,N_1239);
or U1341 (N_1341,N_1244,N_1247);
or U1342 (N_1342,N_1274,N_1226);
and U1343 (N_1343,N_1277,N_1266);
nor U1344 (N_1344,N_1213,N_1288);
nand U1345 (N_1345,N_1284,N_1271);
xor U1346 (N_1346,N_1227,N_1287);
xnor U1347 (N_1347,N_1228,N_1292);
and U1348 (N_1348,N_1258,N_1278);
xnor U1349 (N_1349,N_1273,N_1246);
nor U1350 (N_1350,N_1226,N_1230);
nor U1351 (N_1351,N_1267,N_1231);
xnor U1352 (N_1352,N_1278,N_1274);
and U1353 (N_1353,N_1274,N_1299);
or U1354 (N_1354,N_1261,N_1283);
nand U1355 (N_1355,N_1281,N_1270);
or U1356 (N_1356,N_1236,N_1264);
xnor U1357 (N_1357,N_1223,N_1214);
or U1358 (N_1358,N_1214,N_1244);
xnor U1359 (N_1359,N_1275,N_1274);
nand U1360 (N_1360,N_1233,N_1253);
and U1361 (N_1361,N_1203,N_1240);
nand U1362 (N_1362,N_1247,N_1233);
nor U1363 (N_1363,N_1250,N_1274);
nor U1364 (N_1364,N_1278,N_1247);
or U1365 (N_1365,N_1215,N_1238);
or U1366 (N_1366,N_1249,N_1258);
or U1367 (N_1367,N_1214,N_1269);
and U1368 (N_1368,N_1266,N_1202);
nor U1369 (N_1369,N_1243,N_1233);
nand U1370 (N_1370,N_1244,N_1237);
xor U1371 (N_1371,N_1297,N_1256);
nor U1372 (N_1372,N_1276,N_1214);
nor U1373 (N_1373,N_1290,N_1220);
xnor U1374 (N_1374,N_1203,N_1260);
and U1375 (N_1375,N_1265,N_1242);
nand U1376 (N_1376,N_1279,N_1276);
xnor U1377 (N_1377,N_1251,N_1298);
nand U1378 (N_1378,N_1248,N_1259);
and U1379 (N_1379,N_1234,N_1211);
nand U1380 (N_1380,N_1214,N_1275);
and U1381 (N_1381,N_1219,N_1236);
and U1382 (N_1382,N_1207,N_1279);
nand U1383 (N_1383,N_1210,N_1266);
nor U1384 (N_1384,N_1293,N_1278);
or U1385 (N_1385,N_1268,N_1296);
nor U1386 (N_1386,N_1246,N_1295);
or U1387 (N_1387,N_1297,N_1224);
nor U1388 (N_1388,N_1299,N_1289);
and U1389 (N_1389,N_1236,N_1282);
xor U1390 (N_1390,N_1219,N_1235);
nor U1391 (N_1391,N_1241,N_1294);
and U1392 (N_1392,N_1238,N_1288);
or U1393 (N_1393,N_1295,N_1293);
xor U1394 (N_1394,N_1285,N_1290);
and U1395 (N_1395,N_1266,N_1271);
xor U1396 (N_1396,N_1287,N_1232);
and U1397 (N_1397,N_1235,N_1296);
xnor U1398 (N_1398,N_1273,N_1255);
xor U1399 (N_1399,N_1200,N_1224);
xnor U1400 (N_1400,N_1364,N_1353);
and U1401 (N_1401,N_1342,N_1370);
nor U1402 (N_1402,N_1328,N_1367);
and U1403 (N_1403,N_1340,N_1394);
xnor U1404 (N_1404,N_1351,N_1376);
and U1405 (N_1405,N_1321,N_1339);
or U1406 (N_1406,N_1338,N_1361);
or U1407 (N_1407,N_1385,N_1331);
nand U1408 (N_1408,N_1382,N_1397);
nor U1409 (N_1409,N_1379,N_1345);
or U1410 (N_1410,N_1332,N_1365);
xor U1411 (N_1411,N_1343,N_1347);
nor U1412 (N_1412,N_1325,N_1395);
nand U1413 (N_1413,N_1399,N_1320);
and U1414 (N_1414,N_1388,N_1381);
xnor U1415 (N_1415,N_1363,N_1375);
nand U1416 (N_1416,N_1369,N_1373);
xnor U1417 (N_1417,N_1359,N_1358);
nor U1418 (N_1418,N_1344,N_1306);
or U1419 (N_1419,N_1315,N_1313);
nor U1420 (N_1420,N_1322,N_1312);
or U1421 (N_1421,N_1329,N_1391);
and U1422 (N_1422,N_1310,N_1304);
or U1423 (N_1423,N_1303,N_1371);
xor U1424 (N_1424,N_1333,N_1305);
and U1425 (N_1425,N_1360,N_1316);
xnor U1426 (N_1426,N_1348,N_1318);
xnor U1427 (N_1427,N_1387,N_1380);
nand U1428 (N_1428,N_1311,N_1384);
nor U1429 (N_1429,N_1393,N_1354);
nor U1430 (N_1430,N_1386,N_1337);
nand U1431 (N_1431,N_1330,N_1366);
xor U1432 (N_1432,N_1341,N_1368);
or U1433 (N_1433,N_1349,N_1355);
nand U1434 (N_1434,N_1357,N_1389);
nand U1435 (N_1435,N_1356,N_1335);
nand U1436 (N_1436,N_1362,N_1323);
nor U1437 (N_1437,N_1300,N_1326);
xor U1438 (N_1438,N_1383,N_1392);
nor U1439 (N_1439,N_1377,N_1398);
or U1440 (N_1440,N_1374,N_1317);
and U1441 (N_1441,N_1324,N_1302);
xor U1442 (N_1442,N_1308,N_1390);
xnor U1443 (N_1443,N_1334,N_1327);
nor U1444 (N_1444,N_1396,N_1319);
nand U1445 (N_1445,N_1309,N_1346);
nor U1446 (N_1446,N_1307,N_1372);
nand U1447 (N_1447,N_1350,N_1301);
nor U1448 (N_1448,N_1378,N_1352);
nand U1449 (N_1449,N_1314,N_1336);
nor U1450 (N_1450,N_1364,N_1308);
and U1451 (N_1451,N_1332,N_1358);
xnor U1452 (N_1452,N_1395,N_1340);
xor U1453 (N_1453,N_1324,N_1343);
xor U1454 (N_1454,N_1337,N_1370);
nor U1455 (N_1455,N_1346,N_1396);
and U1456 (N_1456,N_1335,N_1366);
xor U1457 (N_1457,N_1344,N_1349);
xor U1458 (N_1458,N_1393,N_1346);
and U1459 (N_1459,N_1314,N_1371);
xor U1460 (N_1460,N_1303,N_1360);
or U1461 (N_1461,N_1353,N_1320);
xnor U1462 (N_1462,N_1354,N_1332);
nand U1463 (N_1463,N_1315,N_1382);
nor U1464 (N_1464,N_1350,N_1362);
nand U1465 (N_1465,N_1301,N_1341);
or U1466 (N_1466,N_1308,N_1328);
or U1467 (N_1467,N_1398,N_1302);
nand U1468 (N_1468,N_1357,N_1305);
nand U1469 (N_1469,N_1382,N_1342);
and U1470 (N_1470,N_1359,N_1355);
and U1471 (N_1471,N_1358,N_1322);
and U1472 (N_1472,N_1329,N_1387);
or U1473 (N_1473,N_1383,N_1342);
xor U1474 (N_1474,N_1393,N_1333);
nor U1475 (N_1475,N_1336,N_1391);
or U1476 (N_1476,N_1319,N_1348);
nor U1477 (N_1477,N_1335,N_1397);
or U1478 (N_1478,N_1333,N_1331);
or U1479 (N_1479,N_1353,N_1360);
nor U1480 (N_1480,N_1377,N_1383);
and U1481 (N_1481,N_1398,N_1330);
and U1482 (N_1482,N_1341,N_1326);
nor U1483 (N_1483,N_1316,N_1350);
or U1484 (N_1484,N_1395,N_1345);
nor U1485 (N_1485,N_1333,N_1346);
xnor U1486 (N_1486,N_1332,N_1341);
nor U1487 (N_1487,N_1388,N_1310);
nor U1488 (N_1488,N_1385,N_1398);
xor U1489 (N_1489,N_1314,N_1332);
xnor U1490 (N_1490,N_1345,N_1388);
nand U1491 (N_1491,N_1368,N_1375);
nand U1492 (N_1492,N_1352,N_1364);
and U1493 (N_1493,N_1352,N_1340);
or U1494 (N_1494,N_1350,N_1305);
xnor U1495 (N_1495,N_1301,N_1316);
nand U1496 (N_1496,N_1397,N_1318);
and U1497 (N_1497,N_1308,N_1355);
nor U1498 (N_1498,N_1307,N_1316);
and U1499 (N_1499,N_1350,N_1369);
nor U1500 (N_1500,N_1412,N_1408);
xnor U1501 (N_1501,N_1419,N_1458);
nand U1502 (N_1502,N_1478,N_1403);
nor U1503 (N_1503,N_1496,N_1415);
nor U1504 (N_1504,N_1426,N_1452);
xnor U1505 (N_1505,N_1407,N_1421);
nand U1506 (N_1506,N_1498,N_1460);
or U1507 (N_1507,N_1405,N_1409);
or U1508 (N_1508,N_1427,N_1440);
or U1509 (N_1509,N_1453,N_1446);
or U1510 (N_1510,N_1471,N_1406);
nand U1511 (N_1511,N_1492,N_1431);
nand U1512 (N_1512,N_1455,N_1475);
and U1513 (N_1513,N_1410,N_1459);
xnor U1514 (N_1514,N_1423,N_1424);
and U1515 (N_1515,N_1472,N_1464);
xnor U1516 (N_1516,N_1429,N_1479);
nand U1517 (N_1517,N_1400,N_1468);
xnor U1518 (N_1518,N_1473,N_1488);
nand U1519 (N_1519,N_1476,N_1461);
or U1520 (N_1520,N_1442,N_1436);
nor U1521 (N_1521,N_1493,N_1495);
or U1522 (N_1522,N_1404,N_1469);
xnor U1523 (N_1523,N_1413,N_1448);
or U1524 (N_1524,N_1430,N_1402);
and U1525 (N_1525,N_1420,N_1482);
or U1526 (N_1526,N_1474,N_1457);
or U1527 (N_1527,N_1450,N_1490);
nor U1528 (N_1528,N_1483,N_1484);
or U1529 (N_1529,N_1491,N_1422);
xnor U1530 (N_1530,N_1494,N_1447);
xor U1531 (N_1531,N_1451,N_1480);
xnor U1532 (N_1532,N_1449,N_1443);
nor U1533 (N_1533,N_1425,N_1437);
nand U1534 (N_1534,N_1489,N_1465);
nor U1535 (N_1535,N_1418,N_1456);
nor U1536 (N_1536,N_1435,N_1485);
or U1537 (N_1537,N_1477,N_1433);
nor U1538 (N_1538,N_1487,N_1463);
nor U1539 (N_1539,N_1411,N_1401);
or U1540 (N_1540,N_1434,N_1445);
nand U1541 (N_1541,N_1444,N_1439);
and U1542 (N_1542,N_1470,N_1432);
nor U1543 (N_1543,N_1499,N_1481);
or U1544 (N_1544,N_1466,N_1438);
nor U1545 (N_1545,N_1441,N_1454);
xnor U1546 (N_1546,N_1467,N_1416);
nor U1547 (N_1547,N_1462,N_1486);
nor U1548 (N_1548,N_1497,N_1414);
nor U1549 (N_1549,N_1417,N_1428);
xor U1550 (N_1550,N_1400,N_1486);
or U1551 (N_1551,N_1495,N_1444);
xnor U1552 (N_1552,N_1452,N_1489);
or U1553 (N_1553,N_1427,N_1497);
xnor U1554 (N_1554,N_1427,N_1418);
and U1555 (N_1555,N_1450,N_1421);
or U1556 (N_1556,N_1433,N_1473);
nand U1557 (N_1557,N_1449,N_1462);
nand U1558 (N_1558,N_1465,N_1406);
nand U1559 (N_1559,N_1497,N_1404);
nand U1560 (N_1560,N_1426,N_1403);
and U1561 (N_1561,N_1472,N_1480);
nor U1562 (N_1562,N_1486,N_1413);
nor U1563 (N_1563,N_1451,N_1432);
nor U1564 (N_1564,N_1440,N_1412);
nand U1565 (N_1565,N_1485,N_1413);
and U1566 (N_1566,N_1452,N_1427);
nor U1567 (N_1567,N_1415,N_1436);
nand U1568 (N_1568,N_1475,N_1458);
xor U1569 (N_1569,N_1401,N_1450);
or U1570 (N_1570,N_1484,N_1454);
nor U1571 (N_1571,N_1443,N_1421);
nand U1572 (N_1572,N_1419,N_1428);
xor U1573 (N_1573,N_1495,N_1476);
xor U1574 (N_1574,N_1428,N_1407);
xor U1575 (N_1575,N_1471,N_1470);
nor U1576 (N_1576,N_1417,N_1483);
and U1577 (N_1577,N_1480,N_1407);
nand U1578 (N_1578,N_1430,N_1476);
nor U1579 (N_1579,N_1437,N_1401);
and U1580 (N_1580,N_1488,N_1410);
or U1581 (N_1581,N_1485,N_1453);
nand U1582 (N_1582,N_1454,N_1409);
or U1583 (N_1583,N_1493,N_1430);
nand U1584 (N_1584,N_1428,N_1471);
nor U1585 (N_1585,N_1432,N_1456);
nand U1586 (N_1586,N_1495,N_1406);
or U1587 (N_1587,N_1420,N_1435);
and U1588 (N_1588,N_1416,N_1466);
or U1589 (N_1589,N_1444,N_1414);
xnor U1590 (N_1590,N_1465,N_1474);
and U1591 (N_1591,N_1428,N_1421);
nand U1592 (N_1592,N_1497,N_1421);
and U1593 (N_1593,N_1468,N_1441);
nand U1594 (N_1594,N_1406,N_1497);
or U1595 (N_1595,N_1492,N_1472);
and U1596 (N_1596,N_1480,N_1421);
or U1597 (N_1597,N_1427,N_1400);
xnor U1598 (N_1598,N_1426,N_1449);
and U1599 (N_1599,N_1477,N_1495);
or U1600 (N_1600,N_1537,N_1577);
nand U1601 (N_1601,N_1544,N_1557);
nor U1602 (N_1602,N_1506,N_1563);
and U1603 (N_1603,N_1581,N_1573);
xnor U1604 (N_1604,N_1535,N_1553);
xor U1605 (N_1605,N_1599,N_1527);
xor U1606 (N_1606,N_1546,N_1592);
nand U1607 (N_1607,N_1572,N_1585);
xor U1608 (N_1608,N_1554,N_1565);
nor U1609 (N_1609,N_1528,N_1548);
xnor U1610 (N_1610,N_1501,N_1559);
xnor U1611 (N_1611,N_1543,N_1584);
or U1612 (N_1612,N_1530,N_1590);
and U1613 (N_1613,N_1510,N_1545);
nand U1614 (N_1614,N_1583,N_1570);
xor U1615 (N_1615,N_1560,N_1551);
or U1616 (N_1616,N_1550,N_1507);
nor U1617 (N_1617,N_1520,N_1533);
xor U1618 (N_1618,N_1591,N_1549);
xor U1619 (N_1619,N_1566,N_1569);
xnor U1620 (N_1620,N_1532,N_1503);
and U1621 (N_1621,N_1568,N_1594);
nand U1622 (N_1622,N_1523,N_1516);
nand U1623 (N_1623,N_1522,N_1539);
or U1624 (N_1624,N_1515,N_1517);
xor U1625 (N_1625,N_1531,N_1540);
and U1626 (N_1626,N_1575,N_1508);
xnor U1627 (N_1627,N_1580,N_1597);
nor U1628 (N_1628,N_1525,N_1509);
or U1629 (N_1629,N_1555,N_1547);
and U1630 (N_1630,N_1558,N_1562);
xor U1631 (N_1631,N_1598,N_1518);
or U1632 (N_1632,N_1578,N_1534);
nor U1633 (N_1633,N_1513,N_1561);
and U1634 (N_1634,N_1587,N_1582);
nand U1635 (N_1635,N_1526,N_1538);
or U1636 (N_1636,N_1511,N_1567);
and U1637 (N_1637,N_1505,N_1574);
nand U1638 (N_1638,N_1556,N_1536);
xor U1639 (N_1639,N_1595,N_1576);
and U1640 (N_1640,N_1529,N_1541);
nor U1641 (N_1641,N_1588,N_1596);
and U1642 (N_1642,N_1524,N_1593);
xor U1643 (N_1643,N_1542,N_1514);
xnor U1644 (N_1644,N_1579,N_1504);
xnor U1645 (N_1645,N_1500,N_1502);
or U1646 (N_1646,N_1519,N_1589);
xor U1647 (N_1647,N_1564,N_1512);
nand U1648 (N_1648,N_1586,N_1521);
or U1649 (N_1649,N_1571,N_1552);
xnor U1650 (N_1650,N_1520,N_1574);
nor U1651 (N_1651,N_1519,N_1568);
xnor U1652 (N_1652,N_1596,N_1574);
or U1653 (N_1653,N_1524,N_1519);
nand U1654 (N_1654,N_1537,N_1585);
xor U1655 (N_1655,N_1529,N_1572);
nor U1656 (N_1656,N_1531,N_1563);
xnor U1657 (N_1657,N_1537,N_1530);
nand U1658 (N_1658,N_1581,N_1576);
nor U1659 (N_1659,N_1571,N_1510);
nor U1660 (N_1660,N_1529,N_1551);
xnor U1661 (N_1661,N_1544,N_1583);
or U1662 (N_1662,N_1584,N_1576);
or U1663 (N_1663,N_1515,N_1528);
and U1664 (N_1664,N_1511,N_1525);
or U1665 (N_1665,N_1571,N_1520);
or U1666 (N_1666,N_1569,N_1546);
nand U1667 (N_1667,N_1511,N_1522);
nand U1668 (N_1668,N_1505,N_1522);
nor U1669 (N_1669,N_1570,N_1594);
nor U1670 (N_1670,N_1547,N_1568);
and U1671 (N_1671,N_1527,N_1552);
xor U1672 (N_1672,N_1599,N_1506);
or U1673 (N_1673,N_1503,N_1527);
xnor U1674 (N_1674,N_1588,N_1565);
nor U1675 (N_1675,N_1507,N_1501);
or U1676 (N_1676,N_1548,N_1571);
and U1677 (N_1677,N_1516,N_1598);
nor U1678 (N_1678,N_1597,N_1540);
or U1679 (N_1679,N_1533,N_1537);
nand U1680 (N_1680,N_1515,N_1545);
and U1681 (N_1681,N_1553,N_1594);
xor U1682 (N_1682,N_1530,N_1545);
nor U1683 (N_1683,N_1562,N_1575);
and U1684 (N_1684,N_1536,N_1572);
and U1685 (N_1685,N_1596,N_1598);
nand U1686 (N_1686,N_1593,N_1560);
nor U1687 (N_1687,N_1579,N_1569);
nor U1688 (N_1688,N_1534,N_1514);
nor U1689 (N_1689,N_1595,N_1522);
and U1690 (N_1690,N_1501,N_1537);
and U1691 (N_1691,N_1574,N_1556);
nand U1692 (N_1692,N_1517,N_1537);
xor U1693 (N_1693,N_1547,N_1503);
and U1694 (N_1694,N_1548,N_1565);
nand U1695 (N_1695,N_1599,N_1519);
xnor U1696 (N_1696,N_1566,N_1504);
nand U1697 (N_1697,N_1565,N_1552);
and U1698 (N_1698,N_1579,N_1589);
xnor U1699 (N_1699,N_1596,N_1568);
or U1700 (N_1700,N_1678,N_1668);
nand U1701 (N_1701,N_1618,N_1660);
nand U1702 (N_1702,N_1639,N_1694);
xnor U1703 (N_1703,N_1649,N_1609);
nor U1704 (N_1704,N_1653,N_1656);
or U1705 (N_1705,N_1600,N_1697);
nand U1706 (N_1706,N_1691,N_1698);
or U1707 (N_1707,N_1657,N_1635);
xnor U1708 (N_1708,N_1651,N_1652);
xor U1709 (N_1709,N_1684,N_1699);
and U1710 (N_1710,N_1648,N_1619);
xnor U1711 (N_1711,N_1661,N_1630);
or U1712 (N_1712,N_1682,N_1692);
nand U1713 (N_1713,N_1620,N_1695);
or U1714 (N_1714,N_1642,N_1672);
and U1715 (N_1715,N_1647,N_1632);
or U1716 (N_1716,N_1627,N_1637);
nor U1717 (N_1717,N_1607,N_1640);
and U1718 (N_1718,N_1686,N_1665);
and U1719 (N_1719,N_1666,N_1689);
or U1720 (N_1720,N_1621,N_1623);
or U1721 (N_1721,N_1693,N_1674);
nand U1722 (N_1722,N_1671,N_1625);
xor U1723 (N_1723,N_1679,N_1662);
xnor U1724 (N_1724,N_1663,N_1631);
or U1725 (N_1725,N_1683,N_1617);
nor U1726 (N_1726,N_1624,N_1622);
nor U1727 (N_1727,N_1615,N_1658);
or U1728 (N_1728,N_1626,N_1638);
nand U1729 (N_1729,N_1603,N_1633);
nand U1730 (N_1730,N_1685,N_1629);
and U1731 (N_1731,N_1645,N_1664);
and U1732 (N_1732,N_1634,N_1628);
nor U1733 (N_1733,N_1650,N_1601);
or U1734 (N_1734,N_1687,N_1676);
or U1735 (N_1735,N_1667,N_1680);
nand U1736 (N_1736,N_1696,N_1681);
xor U1737 (N_1737,N_1641,N_1673);
nand U1738 (N_1738,N_1654,N_1604);
nor U1739 (N_1739,N_1616,N_1606);
xor U1740 (N_1740,N_1655,N_1636);
and U1741 (N_1741,N_1610,N_1646);
nor U1742 (N_1742,N_1669,N_1611);
xnor U1743 (N_1743,N_1677,N_1675);
xor U1744 (N_1744,N_1659,N_1643);
or U1745 (N_1745,N_1644,N_1670);
xnor U1746 (N_1746,N_1614,N_1612);
nor U1747 (N_1747,N_1602,N_1613);
and U1748 (N_1748,N_1688,N_1605);
xor U1749 (N_1749,N_1608,N_1690);
or U1750 (N_1750,N_1678,N_1624);
and U1751 (N_1751,N_1695,N_1676);
nand U1752 (N_1752,N_1603,N_1629);
nand U1753 (N_1753,N_1612,N_1673);
nand U1754 (N_1754,N_1679,N_1625);
and U1755 (N_1755,N_1652,N_1621);
or U1756 (N_1756,N_1679,N_1674);
and U1757 (N_1757,N_1690,N_1692);
and U1758 (N_1758,N_1600,N_1602);
or U1759 (N_1759,N_1627,N_1601);
and U1760 (N_1760,N_1662,N_1650);
xor U1761 (N_1761,N_1619,N_1629);
or U1762 (N_1762,N_1625,N_1627);
or U1763 (N_1763,N_1695,N_1640);
and U1764 (N_1764,N_1649,N_1647);
xor U1765 (N_1765,N_1663,N_1636);
nand U1766 (N_1766,N_1619,N_1682);
nor U1767 (N_1767,N_1687,N_1624);
and U1768 (N_1768,N_1645,N_1648);
xnor U1769 (N_1769,N_1607,N_1645);
xor U1770 (N_1770,N_1636,N_1603);
or U1771 (N_1771,N_1652,N_1688);
or U1772 (N_1772,N_1624,N_1662);
xor U1773 (N_1773,N_1693,N_1683);
and U1774 (N_1774,N_1630,N_1650);
xnor U1775 (N_1775,N_1609,N_1691);
or U1776 (N_1776,N_1611,N_1664);
and U1777 (N_1777,N_1689,N_1672);
nand U1778 (N_1778,N_1672,N_1607);
nor U1779 (N_1779,N_1692,N_1679);
xnor U1780 (N_1780,N_1655,N_1684);
or U1781 (N_1781,N_1649,N_1619);
and U1782 (N_1782,N_1616,N_1656);
xor U1783 (N_1783,N_1697,N_1696);
and U1784 (N_1784,N_1694,N_1699);
and U1785 (N_1785,N_1604,N_1648);
nor U1786 (N_1786,N_1636,N_1617);
nor U1787 (N_1787,N_1653,N_1688);
xnor U1788 (N_1788,N_1640,N_1604);
or U1789 (N_1789,N_1652,N_1681);
nor U1790 (N_1790,N_1647,N_1618);
nor U1791 (N_1791,N_1647,N_1631);
nand U1792 (N_1792,N_1630,N_1675);
nor U1793 (N_1793,N_1662,N_1689);
nand U1794 (N_1794,N_1602,N_1667);
or U1795 (N_1795,N_1674,N_1620);
and U1796 (N_1796,N_1672,N_1653);
and U1797 (N_1797,N_1630,N_1606);
nand U1798 (N_1798,N_1635,N_1642);
nor U1799 (N_1799,N_1618,N_1696);
nor U1800 (N_1800,N_1781,N_1739);
xnor U1801 (N_1801,N_1719,N_1753);
xnor U1802 (N_1802,N_1791,N_1758);
nor U1803 (N_1803,N_1782,N_1707);
nor U1804 (N_1804,N_1773,N_1701);
or U1805 (N_1805,N_1738,N_1769);
and U1806 (N_1806,N_1780,N_1730);
nand U1807 (N_1807,N_1712,N_1720);
and U1808 (N_1808,N_1795,N_1793);
and U1809 (N_1809,N_1749,N_1733);
xor U1810 (N_1810,N_1755,N_1754);
and U1811 (N_1811,N_1737,N_1783);
xor U1812 (N_1812,N_1774,N_1747);
and U1813 (N_1813,N_1703,N_1771);
nand U1814 (N_1814,N_1721,N_1728);
nand U1815 (N_1815,N_1777,N_1722);
or U1816 (N_1816,N_1752,N_1792);
nand U1817 (N_1817,N_1756,N_1702);
nor U1818 (N_1818,N_1772,N_1776);
xor U1819 (N_1819,N_1710,N_1763);
or U1820 (N_1820,N_1742,N_1779);
xor U1821 (N_1821,N_1785,N_1757);
nor U1822 (N_1822,N_1770,N_1735);
nand U1823 (N_1823,N_1706,N_1726);
or U1824 (N_1824,N_1711,N_1798);
nand U1825 (N_1825,N_1723,N_1744);
and U1826 (N_1826,N_1748,N_1797);
xor U1827 (N_1827,N_1768,N_1740);
nand U1828 (N_1828,N_1751,N_1760);
or U1829 (N_1829,N_1732,N_1746);
nor U1830 (N_1830,N_1741,N_1765);
and U1831 (N_1831,N_1775,N_1705);
or U1832 (N_1832,N_1717,N_1750);
nand U1833 (N_1833,N_1734,N_1764);
nor U1834 (N_1834,N_1708,N_1784);
xor U1835 (N_1835,N_1704,N_1759);
nor U1836 (N_1836,N_1790,N_1799);
and U1837 (N_1837,N_1786,N_1745);
nand U1838 (N_1838,N_1729,N_1766);
xnor U1839 (N_1839,N_1731,N_1715);
xnor U1840 (N_1840,N_1787,N_1762);
xor U1841 (N_1841,N_1718,N_1709);
or U1842 (N_1842,N_1767,N_1743);
nor U1843 (N_1843,N_1778,N_1796);
or U1844 (N_1844,N_1789,N_1788);
xnor U1845 (N_1845,N_1736,N_1724);
xnor U1846 (N_1846,N_1725,N_1714);
and U1847 (N_1847,N_1700,N_1761);
and U1848 (N_1848,N_1794,N_1713);
nand U1849 (N_1849,N_1716,N_1727);
and U1850 (N_1850,N_1787,N_1734);
nor U1851 (N_1851,N_1794,N_1765);
nor U1852 (N_1852,N_1734,N_1775);
or U1853 (N_1853,N_1718,N_1771);
nand U1854 (N_1854,N_1736,N_1748);
nand U1855 (N_1855,N_1768,N_1736);
nor U1856 (N_1856,N_1770,N_1711);
nor U1857 (N_1857,N_1749,N_1747);
and U1858 (N_1858,N_1783,N_1787);
xor U1859 (N_1859,N_1782,N_1710);
nor U1860 (N_1860,N_1795,N_1737);
or U1861 (N_1861,N_1766,N_1719);
nor U1862 (N_1862,N_1780,N_1737);
nand U1863 (N_1863,N_1786,N_1720);
nor U1864 (N_1864,N_1796,N_1723);
xor U1865 (N_1865,N_1764,N_1787);
or U1866 (N_1866,N_1752,N_1775);
or U1867 (N_1867,N_1729,N_1733);
and U1868 (N_1868,N_1703,N_1795);
or U1869 (N_1869,N_1725,N_1746);
nor U1870 (N_1870,N_1745,N_1719);
nor U1871 (N_1871,N_1753,N_1725);
nor U1872 (N_1872,N_1795,N_1781);
or U1873 (N_1873,N_1798,N_1747);
nor U1874 (N_1874,N_1786,N_1742);
or U1875 (N_1875,N_1728,N_1790);
xnor U1876 (N_1876,N_1777,N_1783);
xor U1877 (N_1877,N_1788,N_1761);
xor U1878 (N_1878,N_1709,N_1748);
nand U1879 (N_1879,N_1725,N_1795);
and U1880 (N_1880,N_1778,N_1736);
nor U1881 (N_1881,N_1707,N_1777);
and U1882 (N_1882,N_1773,N_1776);
xor U1883 (N_1883,N_1773,N_1766);
or U1884 (N_1884,N_1726,N_1732);
and U1885 (N_1885,N_1750,N_1757);
and U1886 (N_1886,N_1720,N_1776);
and U1887 (N_1887,N_1734,N_1737);
xnor U1888 (N_1888,N_1745,N_1726);
or U1889 (N_1889,N_1721,N_1704);
nor U1890 (N_1890,N_1732,N_1795);
and U1891 (N_1891,N_1752,N_1773);
or U1892 (N_1892,N_1788,N_1742);
and U1893 (N_1893,N_1769,N_1736);
or U1894 (N_1894,N_1782,N_1754);
nor U1895 (N_1895,N_1712,N_1725);
nand U1896 (N_1896,N_1763,N_1762);
and U1897 (N_1897,N_1753,N_1717);
nand U1898 (N_1898,N_1786,N_1703);
nor U1899 (N_1899,N_1768,N_1702);
xnor U1900 (N_1900,N_1844,N_1892);
xnor U1901 (N_1901,N_1883,N_1886);
xor U1902 (N_1902,N_1874,N_1849);
nand U1903 (N_1903,N_1878,N_1855);
and U1904 (N_1904,N_1802,N_1839);
or U1905 (N_1905,N_1847,N_1853);
nor U1906 (N_1906,N_1829,N_1828);
or U1907 (N_1907,N_1825,N_1811);
nand U1908 (N_1908,N_1864,N_1818);
and U1909 (N_1909,N_1804,N_1834);
nor U1910 (N_1910,N_1887,N_1876);
and U1911 (N_1911,N_1841,N_1879);
and U1912 (N_1912,N_1801,N_1872);
or U1913 (N_1913,N_1836,N_1896);
nand U1914 (N_1914,N_1899,N_1816);
nand U1915 (N_1915,N_1880,N_1803);
or U1916 (N_1916,N_1813,N_1865);
or U1917 (N_1917,N_1831,N_1840);
and U1918 (N_1918,N_1805,N_1861);
or U1919 (N_1919,N_1822,N_1815);
and U1920 (N_1920,N_1893,N_1835);
xnor U1921 (N_1921,N_1823,N_1848);
or U1922 (N_1922,N_1888,N_1807);
and U1923 (N_1923,N_1809,N_1808);
or U1924 (N_1924,N_1856,N_1830);
nor U1925 (N_1925,N_1860,N_1898);
xnor U1926 (N_1926,N_1859,N_1867);
and U1927 (N_1927,N_1843,N_1881);
nand U1928 (N_1928,N_1870,N_1824);
and U1929 (N_1929,N_1842,N_1891);
xnor U1930 (N_1930,N_1871,N_1838);
nor U1931 (N_1931,N_1889,N_1897);
nor U1932 (N_1932,N_1826,N_1854);
nor U1933 (N_1933,N_1858,N_1885);
and U1934 (N_1934,N_1837,N_1857);
nor U1935 (N_1935,N_1832,N_1894);
xnor U1936 (N_1936,N_1884,N_1820);
nor U1937 (N_1937,N_1800,N_1806);
nor U1938 (N_1938,N_1862,N_1882);
nand U1939 (N_1939,N_1846,N_1817);
nor U1940 (N_1940,N_1875,N_1890);
xnor U1941 (N_1941,N_1833,N_1869);
xor U1942 (N_1942,N_1851,N_1895);
and U1943 (N_1943,N_1850,N_1873);
or U1944 (N_1944,N_1812,N_1866);
nor U1945 (N_1945,N_1819,N_1868);
and U1946 (N_1946,N_1852,N_1810);
xor U1947 (N_1947,N_1877,N_1814);
nand U1948 (N_1948,N_1827,N_1845);
and U1949 (N_1949,N_1863,N_1821);
and U1950 (N_1950,N_1817,N_1850);
and U1951 (N_1951,N_1859,N_1878);
nand U1952 (N_1952,N_1860,N_1817);
nand U1953 (N_1953,N_1831,N_1864);
nand U1954 (N_1954,N_1810,N_1803);
xor U1955 (N_1955,N_1847,N_1848);
nor U1956 (N_1956,N_1819,N_1818);
or U1957 (N_1957,N_1872,N_1851);
xnor U1958 (N_1958,N_1858,N_1891);
nand U1959 (N_1959,N_1884,N_1893);
xor U1960 (N_1960,N_1815,N_1810);
nor U1961 (N_1961,N_1861,N_1830);
and U1962 (N_1962,N_1808,N_1873);
and U1963 (N_1963,N_1832,N_1819);
xor U1964 (N_1964,N_1880,N_1810);
or U1965 (N_1965,N_1810,N_1840);
xor U1966 (N_1966,N_1837,N_1831);
and U1967 (N_1967,N_1885,N_1823);
nand U1968 (N_1968,N_1885,N_1843);
nand U1969 (N_1969,N_1878,N_1829);
or U1970 (N_1970,N_1826,N_1808);
nand U1971 (N_1971,N_1893,N_1851);
or U1972 (N_1972,N_1805,N_1833);
nor U1973 (N_1973,N_1815,N_1823);
xnor U1974 (N_1974,N_1845,N_1886);
or U1975 (N_1975,N_1840,N_1811);
or U1976 (N_1976,N_1863,N_1857);
xor U1977 (N_1977,N_1810,N_1877);
nor U1978 (N_1978,N_1845,N_1855);
or U1979 (N_1979,N_1842,N_1874);
nor U1980 (N_1980,N_1867,N_1886);
or U1981 (N_1981,N_1862,N_1856);
and U1982 (N_1982,N_1836,N_1887);
or U1983 (N_1983,N_1862,N_1891);
and U1984 (N_1984,N_1841,N_1807);
and U1985 (N_1985,N_1881,N_1846);
nor U1986 (N_1986,N_1866,N_1818);
or U1987 (N_1987,N_1898,N_1873);
nor U1988 (N_1988,N_1832,N_1856);
xnor U1989 (N_1989,N_1838,N_1821);
nand U1990 (N_1990,N_1817,N_1820);
and U1991 (N_1991,N_1800,N_1809);
nor U1992 (N_1992,N_1855,N_1841);
and U1993 (N_1993,N_1845,N_1812);
nor U1994 (N_1994,N_1874,N_1885);
nand U1995 (N_1995,N_1858,N_1871);
xor U1996 (N_1996,N_1832,N_1855);
and U1997 (N_1997,N_1878,N_1808);
or U1998 (N_1998,N_1850,N_1858);
nor U1999 (N_1999,N_1832,N_1896);
nand U2000 (N_2000,N_1933,N_1993);
nand U2001 (N_2001,N_1900,N_1984);
nor U2002 (N_2002,N_1927,N_1968);
or U2003 (N_2003,N_1985,N_1967);
nor U2004 (N_2004,N_1988,N_1981);
nor U2005 (N_2005,N_1969,N_1955);
xor U2006 (N_2006,N_1920,N_1937);
nor U2007 (N_2007,N_1919,N_1952);
xnor U2008 (N_2008,N_1997,N_1973);
nor U2009 (N_2009,N_1922,N_1979);
or U2010 (N_2010,N_1926,N_1915);
nor U2011 (N_2011,N_1990,N_1991);
or U2012 (N_2012,N_1939,N_1998);
xor U2013 (N_2013,N_1902,N_1944);
or U2014 (N_2014,N_1951,N_1965);
nand U2015 (N_2015,N_1962,N_1982);
nor U2016 (N_2016,N_1942,N_1932);
nand U2017 (N_2017,N_1972,N_1921);
or U2018 (N_2018,N_1961,N_1960);
and U2019 (N_2019,N_1918,N_1916);
xnor U2020 (N_2020,N_1948,N_1911);
xnor U2021 (N_2021,N_1912,N_1974);
and U2022 (N_2022,N_1947,N_1923);
nand U2023 (N_2023,N_1971,N_1977);
or U2024 (N_2024,N_1975,N_1956);
xnor U2025 (N_2025,N_1940,N_1949);
nand U2026 (N_2026,N_1992,N_1954);
or U2027 (N_2027,N_1953,N_1966);
nand U2028 (N_2028,N_1917,N_1930);
or U2029 (N_2029,N_1928,N_1929);
or U2030 (N_2030,N_1901,N_1959);
nor U2031 (N_2031,N_1957,N_1935);
nor U2032 (N_2032,N_1913,N_1907);
nand U2033 (N_2033,N_1936,N_1941);
and U2034 (N_2034,N_1986,N_1999);
nand U2035 (N_2035,N_1945,N_1996);
nand U2036 (N_2036,N_1931,N_1925);
nand U2037 (N_2037,N_1938,N_1904);
and U2038 (N_2038,N_1934,N_1983);
nand U2039 (N_2039,N_1976,N_1924);
and U2040 (N_2040,N_1978,N_1909);
xor U2041 (N_2041,N_1970,N_1995);
xor U2042 (N_2042,N_1943,N_1963);
and U2043 (N_2043,N_1910,N_1980);
xor U2044 (N_2044,N_1964,N_1906);
nor U2045 (N_2045,N_1987,N_1905);
or U2046 (N_2046,N_1994,N_1950);
nand U2047 (N_2047,N_1989,N_1908);
nor U2048 (N_2048,N_1946,N_1914);
and U2049 (N_2049,N_1903,N_1958);
nand U2050 (N_2050,N_1945,N_1901);
or U2051 (N_2051,N_1982,N_1953);
or U2052 (N_2052,N_1921,N_1992);
and U2053 (N_2053,N_1935,N_1973);
xnor U2054 (N_2054,N_1913,N_1995);
and U2055 (N_2055,N_1927,N_1904);
and U2056 (N_2056,N_1902,N_1973);
xnor U2057 (N_2057,N_1939,N_1951);
nand U2058 (N_2058,N_1921,N_1952);
xnor U2059 (N_2059,N_1953,N_1903);
and U2060 (N_2060,N_1964,N_1924);
nand U2061 (N_2061,N_1917,N_1983);
nor U2062 (N_2062,N_1990,N_1945);
and U2063 (N_2063,N_1929,N_1948);
xor U2064 (N_2064,N_1922,N_1901);
or U2065 (N_2065,N_1939,N_1917);
nand U2066 (N_2066,N_1958,N_1975);
xnor U2067 (N_2067,N_1900,N_1986);
nand U2068 (N_2068,N_1949,N_1900);
and U2069 (N_2069,N_1997,N_1986);
and U2070 (N_2070,N_1930,N_1955);
nor U2071 (N_2071,N_1933,N_1974);
nand U2072 (N_2072,N_1957,N_1984);
or U2073 (N_2073,N_1929,N_1923);
xnor U2074 (N_2074,N_1995,N_1916);
nand U2075 (N_2075,N_1941,N_1911);
xor U2076 (N_2076,N_1901,N_1987);
and U2077 (N_2077,N_1912,N_1924);
nand U2078 (N_2078,N_1974,N_1989);
nand U2079 (N_2079,N_1978,N_1924);
nor U2080 (N_2080,N_1963,N_1928);
nand U2081 (N_2081,N_1952,N_1982);
and U2082 (N_2082,N_1977,N_1919);
or U2083 (N_2083,N_1957,N_1902);
nand U2084 (N_2084,N_1990,N_1984);
nor U2085 (N_2085,N_1939,N_1931);
nor U2086 (N_2086,N_1950,N_1984);
nand U2087 (N_2087,N_1988,N_1922);
or U2088 (N_2088,N_1999,N_1917);
nand U2089 (N_2089,N_1973,N_1929);
nand U2090 (N_2090,N_1908,N_1966);
and U2091 (N_2091,N_1934,N_1976);
and U2092 (N_2092,N_1900,N_1988);
xor U2093 (N_2093,N_1917,N_1907);
nor U2094 (N_2094,N_1978,N_1917);
xor U2095 (N_2095,N_1920,N_1990);
xor U2096 (N_2096,N_1990,N_1908);
xor U2097 (N_2097,N_1968,N_1909);
xor U2098 (N_2098,N_1918,N_1993);
or U2099 (N_2099,N_1909,N_1928);
nor U2100 (N_2100,N_2005,N_2030);
nor U2101 (N_2101,N_2089,N_2022);
nor U2102 (N_2102,N_2085,N_2019);
nand U2103 (N_2103,N_2098,N_2084);
and U2104 (N_2104,N_2015,N_2055);
nand U2105 (N_2105,N_2042,N_2028);
or U2106 (N_2106,N_2049,N_2059);
and U2107 (N_2107,N_2020,N_2046);
or U2108 (N_2108,N_2025,N_2070);
nor U2109 (N_2109,N_2039,N_2043);
and U2110 (N_2110,N_2040,N_2051);
nand U2111 (N_2111,N_2003,N_2000);
nand U2112 (N_2112,N_2047,N_2038);
nor U2113 (N_2113,N_2094,N_2027);
xnor U2114 (N_2114,N_2054,N_2052);
xor U2115 (N_2115,N_2012,N_2083);
nor U2116 (N_2116,N_2087,N_2018);
xnor U2117 (N_2117,N_2065,N_2023);
and U2118 (N_2118,N_2037,N_2082);
xor U2119 (N_2119,N_2058,N_2066);
or U2120 (N_2120,N_2061,N_2076);
and U2121 (N_2121,N_2035,N_2088);
and U2122 (N_2122,N_2095,N_2048);
and U2123 (N_2123,N_2093,N_2034);
xnor U2124 (N_2124,N_2002,N_2014);
nor U2125 (N_2125,N_2045,N_2060);
and U2126 (N_2126,N_2078,N_2079);
and U2127 (N_2127,N_2024,N_2032);
nand U2128 (N_2128,N_2016,N_2062);
nand U2129 (N_2129,N_2067,N_2004);
nand U2130 (N_2130,N_2071,N_2007);
and U2131 (N_2131,N_2081,N_2026);
and U2132 (N_2132,N_2068,N_2090);
xor U2133 (N_2133,N_2033,N_2092);
nor U2134 (N_2134,N_2096,N_2001);
nor U2135 (N_2135,N_2077,N_2074);
nand U2136 (N_2136,N_2009,N_2064);
nand U2137 (N_2137,N_2097,N_2006);
or U2138 (N_2138,N_2063,N_2053);
and U2139 (N_2139,N_2057,N_2041);
or U2140 (N_2140,N_2010,N_2044);
and U2141 (N_2141,N_2036,N_2099);
nor U2142 (N_2142,N_2080,N_2073);
and U2143 (N_2143,N_2069,N_2091);
nand U2144 (N_2144,N_2031,N_2013);
nor U2145 (N_2145,N_2086,N_2056);
nor U2146 (N_2146,N_2021,N_2072);
nor U2147 (N_2147,N_2008,N_2017);
or U2148 (N_2148,N_2050,N_2029);
or U2149 (N_2149,N_2011,N_2075);
nor U2150 (N_2150,N_2003,N_2039);
and U2151 (N_2151,N_2097,N_2018);
and U2152 (N_2152,N_2066,N_2064);
xor U2153 (N_2153,N_2060,N_2096);
xor U2154 (N_2154,N_2006,N_2040);
nor U2155 (N_2155,N_2091,N_2039);
or U2156 (N_2156,N_2079,N_2090);
or U2157 (N_2157,N_2011,N_2089);
xor U2158 (N_2158,N_2056,N_2099);
and U2159 (N_2159,N_2042,N_2009);
and U2160 (N_2160,N_2057,N_2023);
or U2161 (N_2161,N_2096,N_2029);
nand U2162 (N_2162,N_2053,N_2078);
xnor U2163 (N_2163,N_2026,N_2065);
nor U2164 (N_2164,N_2077,N_2096);
and U2165 (N_2165,N_2030,N_2057);
and U2166 (N_2166,N_2069,N_2095);
or U2167 (N_2167,N_2038,N_2077);
nor U2168 (N_2168,N_2029,N_2018);
xor U2169 (N_2169,N_2093,N_2035);
nor U2170 (N_2170,N_2049,N_2061);
or U2171 (N_2171,N_2095,N_2018);
nand U2172 (N_2172,N_2044,N_2067);
or U2173 (N_2173,N_2059,N_2019);
or U2174 (N_2174,N_2025,N_2029);
xor U2175 (N_2175,N_2018,N_2049);
or U2176 (N_2176,N_2063,N_2030);
nand U2177 (N_2177,N_2004,N_2042);
and U2178 (N_2178,N_2019,N_2054);
and U2179 (N_2179,N_2023,N_2093);
and U2180 (N_2180,N_2032,N_2042);
nor U2181 (N_2181,N_2067,N_2055);
or U2182 (N_2182,N_2068,N_2078);
nand U2183 (N_2183,N_2029,N_2005);
nor U2184 (N_2184,N_2023,N_2070);
xor U2185 (N_2185,N_2047,N_2041);
xor U2186 (N_2186,N_2086,N_2018);
nand U2187 (N_2187,N_2022,N_2056);
xnor U2188 (N_2188,N_2034,N_2031);
xnor U2189 (N_2189,N_2046,N_2096);
and U2190 (N_2190,N_2069,N_2020);
or U2191 (N_2191,N_2081,N_2096);
nand U2192 (N_2192,N_2013,N_2014);
xnor U2193 (N_2193,N_2054,N_2051);
xor U2194 (N_2194,N_2089,N_2070);
nand U2195 (N_2195,N_2092,N_2029);
and U2196 (N_2196,N_2019,N_2062);
xor U2197 (N_2197,N_2073,N_2021);
xnor U2198 (N_2198,N_2005,N_2080);
and U2199 (N_2199,N_2028,N_2011);
nor U2200 (N_2200,N_2107,N_2147);
or U2201 (N_2201,N_2189,N_2174);
or U2202 (N_2202,N_2162,N_2136);
nor U2203 (N_2203,N_2130,N_2151);
and U2204 (N_2204,N_2171,N_2138);
and U2205 (N_2205,N_2182,N_2183);
xor U2206 (N_2206,N_2194,N_2170);
nand U2207 (N_2207,N_2191,N_2111);
or U2208 (N_2208,N_2115,N_2181);
and U2209 (N_2209,N_2167,N_2118);
and U2210 (N_2210,N_2166,N_2192);
nand U2211 (N_2211,N_2148,N_2173);
nand U2212 (N_2212,N_2129,N_2196);
and U2213 (N_2213,N_2133,N_2108);
nand U2214 (N_2214,N_2197,N_2158);
or U2215 (N_2215,N_2176,N_2131);
nor U2216 (N_2216,N_2113,N_2145);
nand U2217 (N_2217,N_2112,N_2154);
nor U2218 (N_2218,N_2184,N_2114);
xor U2219 (N_2219,N_2100,N_2140);
or U2220 (N_2220,N_2124,N_2103);
nand U2221 (N_2221,N_2142,N_2199);
xor U2222 (N_2222,N_2119,N_2101);
or U2223 (N_2223,N_2120,N_2116);
nand U2224 (N_2224,N_2149,N_2195);
and U2225 (N_2225,N_2164,N_2186);
nand U2226 (N_2226,N_2190,N_2127);
nand U2227 (N_2227,N_2185,N_2163);
and U2228 (N_2228,N_2104,N_2122);
nand U2229 (N_2229,N_2161,N_2177);
nand U2230 (N_2230,N_2152,N_2141);
xnor U2231 (N_2231,N_2172,N_2169);
xor U2232 (N_2232,N_2146,N_2160);
nor U2233 (N_2233,N_2155,N_2143);
xor U2234 (N_2234,N_2165,N_2144);
and U2235 (N_2235,N_2102,N_2150);
xnor U2236 (N_2236,N_2134,N_2137);
nand U2237 (N_2237,N_2175,N_2105);
xnor U2238 (N_2238,N_2106,N_2117);
xnor U2239 (N_2239,N_2135,N_2180);
nor U2240 (N_2240,N_2159,N_2123);
nand U2241 (N_2241,N_2109,N_2188);
nor U2242 (N_2242,N_2157,N_2125);
and U2243 (N_2243,N_2128,N_2110);
xnor U2244 (N_2244,N_2121,N_2198);
nand U2245 (N_2245,N_2178,N_2179);
and U2246 (N_2246,N_2132,N_2193);
nor U2247 (N_2247,N_2156,N_2168);
and U2248 (N_2248,N_2153,N_2187);
or U2249 (N_2249,N_2139,N_2126);
nor U2250 (N_2250,N_2171,N_2144);
nand U2251 (N_2251,N_2155,N_2160);
and U2252 (N_2252,N_2189,N_2181);
or U2253 (N_2253,N_2106,N_2129);
nor U2254 (N_2254,N_2180,N_2194);
nand U2255 (N_2255,N_2154,N_2125);
xor U2256 (N_2256,N_2100,N_2137);
nor U2257 (N_2257,N_2163,N_2113);
nand U2258 (N_2258,N_2145,N_2148);
and U2259 (N_2259,N_2101,N_2158);
xor U2260 (N_2260,N_2196,N_2113);
or U2261 (N_2261,N_2193,N_2182);
nor U2262 (N_2262,N_2165,N_2130);
and U2263 (N_2263,N_2116,N_2113);
xnor U2264 (N_2264,N_2108,N_2115);
nand U2265 (N_2265,N_2192,N_2176);
xnor U2266 (N_2266,N_2167,N_2172);
or U2267 (N_2267,N_2140,N_2156);
and U2268 (N_2268,N_2199,N_2138);
nand U2269 (N_2269,N_2122,N_2155);
and U2270 (N_2270,N_2113,N_2194);
or U2271 (N_2271,N_2121,N_2154);
or U2272 (N_2272,N_2137,N_2166);
or U2273 (N_2273,N_2114,N_2172);
nand U2274 (N_2274,N_2146,N_2183);
nand U2275 (N_2275,N_2135,N_2137);
xnor U2276 (N_2276,N_2127,N_2108);
or U2277 (N_2277,N_2169,N_2149);
nor U2278 (N_2278,N_2137,N_2192);
or U2279 (N_2279,N_2148,N_2192);
or U2280 (N_2280,N_2157,N_2152);
xnor U2281 (N_2281,N_2146,N_2123);
nor U2282 (N_2282,N_2136,N_2125);
or U2283 (N_2283,N_2145,N_2182);
nand U2284 (N_2284,N_2164,N_2123);
or U2285 (N_2285,N_2176,N_2115);
xor U2286 (N_2286,N_2132,N_2168);
xor U2287 (N_2287,N_2131,N_2133);
xor U2288 (N_2288,N_2130,N_2182);
nor U2289 (N_2289,N_2191,N_2132);
or U2290 (N_2290,N_2134,N_2164);
xor U2291 (N_2291,N_2108,N_2130);
xor U2292 (N_2292,N_2187,N_2145);
xnor U2293 (N_2293,N_2157,N_2186);
nand U2294 (N_2294,N_2128,N_2118);
xnor U2295 (N_2295,N_2159,N_2112);
xor U2296 (N_2296,N_2168,N_2176);
xor U2297 (N_2297,N_2111,N_2110);
and U2298 (N_2298,N_2142,N_2145);
or U2299 (N_2299,N_2145,N_2114);
xor U2300 (N_2300,N_2270,N_2275);
nor U2301 (N_2301,N_2236,N_2296);
or U2302 (N_2302,N_2283,N_2293);
or U2303 (N_2303,N_2226,N_2209);
nor U2304 (N_2304,N_2281,N_2203);
xnor U2305 (N_2305,N_2250,N_2218);
xnor U2306 (N_2306,N_2277,N_2205);
nor U2307 (N_2307,N_2278,N_2238);
nand U2308 (N_2308,N_2260,N_2267);
and U2309 (N_2309,N_2279,N_2257);
and U2310 (N_2310,N_2262,N_2255);
or U2311 (N_2311,N_2265,N_2216);
nand U2312 (N_2312,N_2219,N_2256);
and U2313 (N_2313,N_2230,N_2286);
or U2314 (N_2314,N_2239,N_2240);
nor U2315 (N_2315,N_2291,N_2284);
and U2316 (N_2316,N_2220,N_2259);
nand U2317 (N_2317,N_2212,N_2208);
and U2318 (N_2318,N_2251,N_2298);
nand U2319 (N_2319,N_2292,N_2294);
or U2320 (N_2320,N_2225,N_2272);
and U2321 (N_2321,N_2252,N_2223);
nor U2322 (N_2322,N_2213,N_2276);
xor U2323 (N_2323,N_2200,N_2235);
xnor U2324 (N_2324,N_2210,N_2228);
xnor U2325 (N_2325,N_2268,N_2269);
and U2326 (N_2326,N_2207,N_2201);
nand U2327 (N_2327,N_2206,N_2282);
nor U2328 (N_2328,N_2271,N_2280);
nand U2329 (N_2329,N_2244,N_2263);
nor U2330 (N_2330,N_2287,N_2288);
nand U2331 (N_2331,N_2247,N_2224);
xor U2332 (N_2332,N_2295,N_2204);
and U2333 (N_2333,N_2249,N_2297);
and U2334 (N_2334,N_2229,N_2266);
xnor U2335 (N_2335,N_2274,N_2258);
and U2336 (N_2336,N_2242,N_2233);
nand U2337 (N_2337,N_2202,N_2234);
and U2338 (N_2338,N_2232,N_2241);
or U2339 (N_2339,N_2246,N_2243);
and U2340 (N_2340,N_2248,N_2231);
or U2341 (N_2341,N_2211,N_2290);
xor U2342 (N_2342,N_2285,N_2245);
or U2343 (N_2343,N_2253,N_2261);
and U2344 (N_2344,N_2299,N_2214);
and U2345 (N_2345,N_2227,N_2222);
and U2346 (N_2346,N_2221,N_2289);
xnor U2347 (N_2347,N_2215,N_2273);
xor U2348 (N_2348,N_2254,N_2264);
nand U2349 (N_2349,N_2217,N_2237);
and U2350 (N_2350,N_2248,N_2224);
or U2351 (N_2351,N_2248,N_2227);
nand U2352 (N_2352,N_2234,N_2291);
and U2353 (N_2353,N_2280,N_2235);
xnor U2354 (N_2354,N_2229,N_2264);
or U2355 (N_2355,N_2251,N_2292);
nor U2356 (N_2356,N_2254,N_2238);
nand U2357 (N_2357,N_2216,N_2271);
xor U2358 (N_2358,N_2264,N_2223);
or U2359 (N_2359,N_2293,N_2297);
and U2360 (N_2360,N_2247,N_2263);
xor U2361 (N_2361,N_2295,N_2293);
or U2362 (N_2362,N_2231,N_2278);
xnor U2363 (N_2363,N_2259,N_2216);
xnor U2364 (N_2364,N_2213,N_2284);
nand U2365 (N_2365,N_2270,N_2219);
xor U2366 (N_2366,N_2261,N_2225);
and U2367 (N_2367,N_2289,N_2242);
and U2368 (N_2368,N_2250,N_2213);
nand U2369 (N_2369,N_2247,N_2231);
and U2370 (N_2370,N_2290,N_2272);
xnor U2371 (N_2371,N_2248,N_2275);
nor U2372 (N_2372,N_2204,N_2221);
or U2373 (N_2373,N_2296,N_2298);
xor U2374 (N_2374,N_2264,N_2268);
and U2375 (N_2375,N_2254,N_2248);
nor U2376 (N_2376,N_2201,N_2285);
or U2377 (N_2377,N_2282,N_2224);
or U2378 (N_2378,N_2286,N_2223);
nand U2379 (N_2379,N_2259,N_2245);
xor U2380 (N_2380,N_2228,N_2254);
or U2381 (N_2381,N_2232,N_2207);
and U2382 (N_2382,N_2298,N_2263);
and U2383 (N_2383,N_2218,N_2236);
xor U2384 (N_2384,N_2236,N_2214);
and U2385 (N_2385,N_2203,N_2247);
xnor U2386 (N_2386,N_2299,N_2222);
nand U2387 (N_2387,N_2259,N_2278);
nand U2388 (N_2388,N_2296,N_2277);
nor U2389 (N_2389,N_2236,N_2255);
nor U2390 (N_2390,N_2255,N_2268);
nand U2391 (N_2391,N_2274,N_2253);
xor U2392 (N_2392,N_2249,N_2207);
nand U2393 (N_2393,N_2215,N_2282);
nand U2394 (N_2394,N_2290,N_2289);
nand U2395 (N_2395,N_2236,N_2274);
xnor U2396 (N_2396,N_2268,N_2213);
xnor U2397 (N_2397,N_2208,N_2275);
xnor U2398 (N_2398,N_2265,N_2297);
nand U2399 (N_2399,N_2268,N_2286);
or U2400 (N_2400,N_2330,N_2310);
and U2401 (N_2401,N_2390,N_2367);
nand U2402 (N_2402,N_2350,N_2384);
nand U2403 (N_2403,N_2395,N_2338);
nor U2404 (N_2404,N_2357,N_2381);
xor U2405 (N_2405,N_2364,N_2361);
nor U2406 (N_2406,N_2368,N_2349);
nand U2407 (N_2407,N_2318,N_2340);
or U2408 (N_2408,N_2378,N_2375);
nand U2409 (N_2409,N_2328,N_2380);
nor U2410 (N_2410,N_2351,N_2302);
nor U2411 (N_2411,N_2333,N_2391);
and U2412 (N_2412,N_2358,N_2341);
or U2413 (N_2413,N_2305,N_2336);
and U2414 (N_2414,N_2342,N_2388);
or U2415 (N_2415,N_2314,N_2376);
or U2416 (N_2416,N_2300,N_2306);
xnor U2417 (N_2417,N_2379,N_2335);
and U2418 (N_2418,N_2392,N_2370);
xnor U2419 (N_2419,N_2382,N_2354);
xnor U2420 (N_2420,N_2309,N_2319);
xor U2421 (N_2421,N_2346,N_2313);
or U2422 (N_2422,N_2396,N_2345);
xnor U2423 (N_2423,N_2389,N_2334);
nand U2424 (N_2424,N_2308,N_2348);
nand U2425 (N_2425,N_2356,N_2366);
xnor U2426 (N_2426,N_2371,N_2365);
and U2427 (N_2427,N_2377,N_2355);
and U2428 (N_2428,N_2304,N_2337);
nor U2429 (N_2429,N_2327,N_2373);
and U2430 (N_2430,N_2397,N_2363);
or U2431 (N_2431,N_2369,N_2344);
and U2432 (N_2432,N_2325,N_2312);
or U2433 (N_2433,N_2347,N_2387);
xnor U2434 (N_2434,N_2326,N_2317);
xor U2435 (N_2435,N_2301,N_2372);
or U2436 (N_2436,N_2360,N_2321);
nand U2437 (N_2437,N_2339,N_2324);
nor U2438 (N_2438,N_2374,N_2353);
and U2439 (N_2439,N_2362,N_2303);
nand U2440 (N_2440,N_2311,N_2320);
xnor U2441 (N_2441,N_2385,N_2331);
and U2442 (N_2442,N_2315,N_2307);
xor U2443 (N_2443,N_2393,N_2399);
nand U2444 (N_2444,N_2383,N_2343);
nor U2445 (N_2445,N_2332,N_2398);
xnor U2446 (N_2446,N_2359,N_2329);
and U2447 (N_2447,N_2352,N_2316);
nor U2448 (N_2448,N_2323,N_2322);
nor U2449 (N_2449,N_2386,N_2394);
and U2450 (N_2450,N_2351,N_2343);
nor U2451 (N_2451,N_2335,N_2380);
nor U2452 (N_2452,N_2365,N_2370);
xor U2453 (N_2453,N_2323,N_2334);
xor U2454 (N_2454,N_2345,N_2304);
nor U2455 (N_2455,N_2374,N_2321);
nand U2456 (N_2456,N_2348,N_2373);
xnor U2457 (N_2457,N_2379,N_2309);
and U2458 (N_2458,N_2394,N_2351);
xor U2459 (N_2459,N_2361,N_2323);
xor U2460 (N_2460,N_2300,N_2356);
nor U2461 (N_2461,N_2356,N_2318);
xor U2462 (N_2462,N_2395,N_2391);
nor U2463 (N_2463,N_2334,N_2387);
xnor U2464 (N_2464,N_2335,N_2327);
nand U2465 (N_2465,N_2312,N_2396);
nand U2466 (N_2466,N_2393,N_2337);
nor U2467 (N_2467,N_2391,N_2376);
xnor U2468 (N_2468,N_2390,N_2384);
nor U2469 (N_2469,N_2315,N_2309);
nor U2470 (N_2470,N_2326,N_2306);
or U2471 (N_2471,N_2308,N_2362);
nor U2472 (N_2472,N_2307,N_2334);
and U2473 (N_2473,N_2335,N_2354);
or U2474 (N_2474,N_2369,N_2350);
and U2475 (N_2475,N_2338,N_2357);
or U2476 (N_2476,N_2395,N_2309);
and U2477 (N_2477,N_2327,N_2345);
xor U2478 (N_2478,N_2315,N_2308);
xnor U2479 (N_2479,N_2387,N_2354);
nor U2480 (N_2480,N_2306,N_2358);
nor U2481 (N_2481,N_2335,N_2358);
or U2482 (N_2482,N_2364,N_2333);
xor U2483 (N_2483,N_2356,N_2345);
nor U2484 (N_2484,N_2384,N_2305);
or U2485 (N_2485,N_2371,N_2315);
nand U2486 (N_2486,N_2384,N_2322);
xnor U2487 (N_2487,N_2306,N_2397);
xnor U2488 (N_2488,N_2347,N_2339);
nor U2489 (N_2489,N_2303,N_2378);
nor U2490 (N_2490,N_2312,N_2380);
or U2491 (N_2491,N_2332,N_2386);
nand U2492 (N_2492,N_2331,N_2399);
and U2493 (N_2493,N_2388,N_2353);
or U2494 (N_2494,N_2330,N_2314);
nand U2495 (N_2495,N_2351,N_2306);
nand U2496 (N_2496,N_2329,N_2384);
and U2497 (N_2497,N_2324,N_2333);
and U2498 (N_2498,N_2334,N_2393);
xnor U2499 (N_2499,N_2363,N_2390);
nand U2500 (N_2500,N_2462,N_2475);
and U2501 (N_2501,N_2482,N_2401);
and U2502 (N_2502,N_2485,N_2466);
and U2503 (N_2503,N_2440,N_2409);
nor U2504 (N_2504,N_2406,N_2473);
nand U2505 (N_2505,N_2452,N_2492);
xor U2506 (N_2506,N_2484,N_2402);
or U2507 (N_2507,N_2428,N_2453);
and U2508 (N_2508,N_2488,N_2418);
nor U2509 (N_2509,N_2408,N_2480);
and U2510 (N_2510,N_2432,N_2496);
nand U2511 (N_2511,N_2443,N_2400);
nor U2512 (N_2512,N_2416,N_2490);
xnor U2513 (N_2513,N_2470,N_2438);
nor U2514 (N_2514,N_2436,N_2413);
xnor U2515 (N_2515,N_2429,N_2446);
nand U2516 (N_2516,N_2468,N_2476);
and U2517 (N_2517,N_2449,N_2494);
nor U2518 (N_2518,N_2405,N_2447);
nand U2519 (N_2519,N_2469,N_2442);
nor U2520 (N_2520,N_2487,N_2495);
nand U2521 (N_2521,N_2419,N_2444);
nand U2522 (N_2522,N_2435,N_2499);
and U2523 (N_2523,N_2407,N_2422);
or U2524 (N_2524,N_2493,N_2421);
or U2525 (N_2525,N_2486,N_2403);
or U2526 (N_2526,N_2424,N_2481);
xor U2527 (N_2527,N_2431,N_2474);
or U2528 (N_2528,N_2415,N_2441);
or U2529 (N_2529,N_2450,N_2437);
nor U2530 (N_2530,N_2478,N_2434);
xnor U2531 (N_2531,N_2464,N_2433);
nor U2532 (N_2532,N_2498,N_2456);
and U2533 (N_2533,N_2427,N_2439);
xnor U2534 (N_2534,N_2425,N_2420);
and U2535 (N_2535,N_2491,N_2471);
xor U2536 (N_2536,N_2412,N_2458);
xnor U2537 (N_2537,N_2451,N_2489);
nor U2538 (N_2538,N_2479,N_2463);
nor U2539 (N_2539,N_2472,N_2461);
nor U2540 (N_2540,N_2423,N_2455);
nand U2541 (N_2541,N_2404,N_2426);
and U2542 (N_2542,N_2465,N_2454);
xnor U2543 (N_2543,N_2414,N_2477);
nand U2544 (N_2544,N_2411,N_2445);
and U2545 (N_2545,N_2467,N_2457);
xnor U2546 (N_2546,N_2410,N_2430);
and U2547 (N_2547,N_2448,N_2483);
or U2548 (N_2548,N_2460,N_2497);
xnor U2549 (N_2549,N_2459,N_2417);
and U2550 (N_2550,N_2447,N_2461);
and U2551 (N_2551,N_2473,N_2447);
nor U2552 (N_2552,N_2448,N_2434);
nand U2553 (N_2553,N_2484,N_2423);
and U2554 (N_2554,N_2405,N_2400);
nand U2555 (N_2555,N_2478,N_2406);
or U2556 (N_2556,N_2467,N_2459);
xor U2557 (N_2557,N_2464,N_2484);
nor U2558 (N_2558,N_2475,N_2414);
and U2559 (N_2559,N_2498,N_2430);
or U2560 (N_2560,N_2417,N_2478);
nand U2561 (N_2561,N_2491,N_2444);
or U2562 (N_2562,N_2409,N_2430);
nor U2563 (N_2563,N_2474,N_2452);
or U2564 (N_2564,N_2448,N_2409);
or U2565 (N_2565,N_2445,N_2444);
nor U2566 (N_2566,N_2484,N_2483);
or U2567 (N_2567,N_2470,N_2449);
nor U2568 (N_2568,N_2401,N_2423);
and U2569 (N_2569,N_2485,N_2445);
and U2570 (N_2570,N_2458,N_2423);
nor U2571 (N_2571,N_2447,N_2469);
xnor U2572 (N_2572,N_2489,N_2462);
nor U2573 (N_2573,N_2474,N_2418);
nand U2574 (N_2574,N_2427,N_2419);
xnor U2575 (N_2575,N_2482,N_2484);
nor U2576 (N_2576,N_2403,N_2423);
or U2577 (N_2577,N_2436,N_2485);
nor U2578 (N_2578,N_2426,N_2424);
or U2579 (N_2579,N_2427,N_2452);
nand U2580 (N_2580,N_2477,N_2444);
or U2581 (N_2581,N_2499,N_2419);
xnor U2582 (N_2582,N_2429,N_2458);
nand U2583 (N_2583,N_2450,N_2489);
and U2584 (N_2584,N_2406,N_2499);
nand U2585 (N_2585,N_2458,N_2452);
nand U2586 (N_2586,N_2438,N_2440);
and U2587 (N_2587,N_2430,N_2431);
or U2588 (N_2588,N_2485,N_2448);
xor U2589 (N_2589,N_2459,N_2414);
xor U2590 (N_2590,N_2436,N_2456);
nand U2591 (N_2591,N_2429,N_2413);
or U2592 (N_2592,N_2495,N_2499);
xnor U2593 (N_2593,N_2454,N_2410);
xnor U2594 (N_2594,N_2455,N_2483);
nor U2595 (N_2595,N_2422,N_2490);
nor U2596 (N_2596,N_2449,N_2499);
xnor U2597 (N_2597,N_2421,N_2404);
xnor U2598 (N_2598,N_2422,N_2418);
xor U2599 (N_2599,N_2456,N_2405);
and U2600 (N_2600,N_2595,N_2507);
or U2601 (N_2601,N_2597,N_2505);
or U2602 (N_2602,N_2536,N_2551);
nand U2603 (N_2603,N_2532,N_2514);
nand U2604 (N_2604,N_2559,N_2552);
or U2605 (N_2605,N_2577,N_2580);
nand U2606 (N_2606,N_2569,N_2541);
xnor U2607 (N_2607,N_2581,N_2556);
nand U2608 (N_2608,N_2570,N_2501);
nand U2609 (N_2609,N_2535,N_2589);
nand U2610 (N_2610,N_2546,N_2578);
xor U2611 (N_2611,N_2526,N_2565);
and U2612 (N_2612,N_2567,N_2531);
and U2613 (N_2613,N_2518,N_2524);
nand U2614 (N_2614,N_2575,N_2545);
nand U2615 (N_2615,N_2530,N_2538);
nor U2616 (N_2616,N_2516,N_2522);
nor U2617 (N_2617,N_2592,N_2515);
and U2618 (N_2618,N_2568,N_2594);
nor U2619 (N_2619,N_2503,N_2563);
nor U2620 (N_2620,N_2555,N_2521);
xor U2621 (N_2621,N_2502,N_2561);
and U2622 (N_2622,N_2579,N_2558);
or U2623 (N_2623,N_2533,N_2504);
or U2624 (N_2624,N_2510,N_2571);
or U2625 (N_2625,N_2525,N_2509);
or U2626 (N_2626,N_2523,N_2599);
xnor U2627 (N_2627,N_2591,N_2553);
xor U2628 (N_2628,N_2564,N_2585);
and U2629 (N_2629,N_2583,N_2574);
nor U2630 (N_2630,N_2598,N_2572);
xor U2631 (N_2631,N_2517,N_2547);
xnor U2632 (N_2632,N_2543,N_2550);
nand U2633 (N_2633,N_2539,N_2588);
nor U2634 (N_2634,N_2529,N_2542);
or U2635 (N_2635,N_2500,N_2520);
xnor U2636 (N_2636,N_2593,N_2548);
xnor U2637 (N_2637,N_2590,N_2527);
or U2638 (N_2638,N_2544,N_2554);
and U2639 (N_2639,N_2596,N_2537);
or U2640 (N_2640,N_2557,N_2549);
and U2641 (N_2641,N_2519,N_2513);
xnor U2642 (N_2642,N_2512,N_2576);
xor U2643 (N_2643,N_2511,N_2540);
xor U2644 (N_2644,N_2528,N_2584);
and U2645 (N_2645,N_2587,N_2582);
nor U2646 (N_2646,N_2534,N_2560);
nor U2647 (N_2647,N_2586,N_2506);
and U2648 (N_2648,N_2562,N_2566);
nand U2649 (N_2649,N_2573,N_2508);
or U2650 (N_2650,N_2531,N_2509);
nor U2651 (N_2651,N_2516,N_2547);
or U2652 (N_2652,N_2533,N_2532);
and U2653 (N_2653,N_2523,N_2568);
nor U2654 (N_2654,N_2538,N_2578);
and U2655 (N_2655,N_2540,N_2535);
xor U2656 (N_2656,N_2586,N_2575);
and U2657 (N_2657,N_2535,N_2549);
xor U2658 (N_2658,N_2585,N_2583);
nand U2659 (N_2659,N_2525,N_2543);
xor U2660 (N_2660,N_2532,N_2528);
nand U2661 (N_2661,N_2593,N_2573);
xor U2662 (N_2662,N_2562,N_2594);
nor U2663 (N_2663,N_2519,N_2594);
xnor U2664 (N_2664,N_2552,N_2568);
or U2665 (N_2665,N_2572,N_2538);
nand U2666 (N_2666,N_2535,N_2570);
nand U2667 (N_2667,N_2544,N_2514);
xnor U2668 (N_2668,N_2569,N_2572);
nor U2669 (N_2669,N_2585,N_2586);
xor U2670 (N_2670,N_2527,N_2559);
nand U2671 (N_2671,N_2541,N_2582);
or U2672 (N_2672,N_2507,N_2582);
xnor U2673 (N_2673,N_2561,N_2587);
nor U2674 (N_2674,N_2536,N_2522);
nand U2675 (N_2675,N_2573,N_2556);
and U2676 (N_2676,N_2562,N_2592);
nand U2677 (N_2677,N_2585,N_2567);
or U2678 (N_2678,N_2505,N_2501);
nand U2679 (N_2679,N_2529,N_2587);
or U2680 (N_2680,N_2544,N_2536);
xor U2681 (N_2681,N_2570,N_2565);
xnor U2682 (N_2682,N_2539,N_2500);
or U2683 (N_2683,N_2523,N_2518);
or U2684 (N_2684,N_2510,N_2560);
xor U2685 (N_2685,N_2573,N_2558);
xor U2686 (N_2686,N_2537,N_2577);
nand U2687 (N_2687,N_2596,N_2598);
xor U2688 (N_2688,N_2551,N_2510);
xor U2689 (N_2689,N_2506,N_2589);
xnor U2690 (N_2690,N_2596,N_2568);
nand U2691 (N_2691,N_2565,N_2571);
or U2692 (N_2692,N_2552,N_2502);
or U2693 (N_2693,N_2520,N_2503);
and U2694 (N_2694,N_2572,N_2563);
xor U2695 (N_2695,N_2576,N_2519);
xor U2696 (N_2696,N_2520,N_2516);
nand U2697 (N_2697,N_2579,N_2527);
or U2698 (N_2698,N_2574,N_2534);
nand U2699 (N_2699,N_2537,N_2543);
and U2700 (N_2700,N_2631,N_2688);
xor U2701 (N_2701,N_2601,N_2694);
xnor U2702 (N_2702,N_2639,N_2604);
or U2703 (N_2703,N_2676,N_2690);
and U2704 (N_2704,N_2669,N_2625);
nand U2705 (N_2705,N_2695,N_2657);
or U2706 (N_2706,N_2611,N_2693);
xnor U2707 (N_2707,N_2612,N_2624);
or U2708 (N_2708,N_2615,N_2618);
and U2709 (N_2709,N_2671,N_2643);
nand U2710 (N_2710,N_2633,N_2614);
or U2711 (N_2711,N_2609,N_2683);
or U2712 (N_2712,N_2617,N_2621);
xor U2713 (N_2713,N_2650,N_2642);
nor U2714 (N_2714,N_2634,N_2678);
or U2715 (N_2715,N_2663,N_2619);
and U2716 (N_2716,N_2685,N_2666);
nand U2717 (N_2717,N_2682,N_2659);
and U2718 (N_2718,N_2641,N_2689);
and U2719 (N_2719,N_2616,N_2674);
nand U2720 (N_2720,N_2662,N_2654);
nand U2721 (N_2721,N_2600,N_2629);
xnor U2722 (N_2722,N_2635,N_2658);
nor U2723 (N_2723,N_2675,N_2627);
and U2724 (N_2724,N_2607,N_2605);
or U2725 (N_2725,N_2656,N_2687);
or U2726 (N_2726,N_2680,N_2679);
xnor U2727 (N_2727,N_2626,N_2636);
nand U2728 (N_2728,N_2699,N_2630);
or U2729 (N_2729,N_2681,N_2670);
and U2730 (N_2730,N_2603,N_2613);
or U2731 (N_2731,N_2655,N_2660);
nor U2732 (N_2732,N_2645,N_2623);
nor U2733 (N_2733,N_2691,N_2696);
and U2734 (N_2734,N_2672,N_2637);
nand U2735 (N_2735,N_2644,N_2664);
xnor U2736 (N_2736,N_2665,N_2661);
or U2737 (N_2737,N_2602,N_2648);
and U2738 (N_2738,N_2697,N_2686);
or U2739 (N_2739,N_2620,N_2652);
nor U2740 (N_2740,N_2698,N_2640);
xnor U2741 (N_2741,N_2628,N_2673);
nand U2742 (N_2742,N_2651,N_2684);
or U2743 (N_2743,N_2638,N_2646);
xor U2744 (N_2744,N_2668,N_2632);
and U2745 (N_2745,N_2622,N_2667);
and U2746 (N_2746,N_2608,N_2677);
nor U2747 (N_2747,N_2606,N_2692);
and U2748 (N_2748,N_2647,N_2649);
nand U2749 (N_2749,N_2610,N_2653);
xor U2750 (N_2750,N_2625,N_2651);
and U2751 (N_2751,N_2688,N_2679);
xor U2752 (N_2752,N_2665,N_2635);
xnor U2753 (N_2753,N_2623,N_2653);
or U2754 (N_2754,N_2641,N_2630);
nor U2755 (N_2755,N_2688,N_2677);
nand U2756 (N_2756,N_2655,N_2686);
and U2757 (N_2757,N_2622,N_2694);
or U2758 (N_2758,N_2689,N_2651);
or U2759 (N_2759,N_2636,N_2625);
nand U2760 (N_2760,N_2660,N_2662);
and U2761 (N_2761,N_2641,N_2636);
or U2762 (N_2762,N_2652,N_2693);
and U2763 (N_2763,N_2690,N_2685);
nand U2764 (N_2764,N_2679,N_2608);
or U2765 (N_2765,N_2622,N_2615);
nor U2766 (N_2766,N_2617,N_2649);
xor U2767 (N_2767,N_2677,N_2601);
nand U2768 (N_2768,N_2670,N_2677);
or U2769 (N_2769,N_2610,N_2671);
or U2770 (N_2770,N_2639,N_2664);
and U2771 (N_2771,N_2654,N_2649);
and U2772 (N_2772,N_2685,N_2640);
and U2773 (N_2773,N_2617,N_2608);
nor U2774 (N_2774,N_2646,N_2620);
nor U2775 (N_2775,N_2642,N_2654);
or U2776 (N_2776,N_2660,N_2639);
nor U2777 (N_2777,N_2683,N_2634);
nand U2778 (N_2778,N_2634,N_2609);
or U2779 (N_2779,N_2624,N_2617);
nand U2780 (N_2780,N_2627,N_2631);
xnor U2781 (N_2781,N_2627,N_2601);
nand U2782 (N_2782,N_2606,N_2630);
xor U2783 (N_2783,N_2674,N_2680);
or U2784 (N_2784,N_2631,N_2653);
and U2785 (N_2785,N_2612,N_2639);
nand U2786 (N_2786,N_2636,N_2631);
or U2787 (N_2787,N_2609,N_2635);
nand U2788 (N_2788,N_2683,N_2680);
nand U2789 (N_2789,N_2612,N_2673);
nor U2790 (N_2790,N_2641,N_2686);
nand U2791 (N_2791,N_2637,N_2680);
xnor U2792 (N_2792,N_2605,N_2614);
xor U2793 (N_2793,N_2689,N_2688);
and U2794 (N_2794,N_2602,N_2622);
or U2795 (N_2795,N_2683,N_2636);
xnor U2796 (N_2796,N_2685,N_2691);
nand U2797 (N_2797,N_2677,N_2653);
nand U2798 (N_2798,N_2655,N_2693);
or U2799 (N_2799,N_2696,N_2659);
or U2800 (N_2800,N_2745,N_2716);
or U2801 (N_2801,N_2706,N_2786);
nand U2802 (N_2802,N_2740,N_2784);
xor U2803 (N_2803,N_2730,N_2764);
or U2804 (N_2804,N_2700,N_2792);
nand U2805 (N_2805,N_2747,N_2749);
xnor U2806 (N_2806,N_2783,N_2780);
or U2807 (N_2807,N_2717,N_2720);
or U2808 (N_2808,N_2714,N_2728);
nor U2809 (N_2809,N_2776,N_2766);
xor U2810 (N_2810,N_2769,N_2713);
xor U2811 (N_2811,N_2782,N_2775);
xnor U2812 (N_2812,N_2771,N_2762);
and U2813 (N_2813,N_2778,N_2772);
nor U2814 (N_2814,N_2754,N_2753);
or U2815 (N_2815,N_2742,N_2722);
and U2816 (N_2816,N_2768,N_2732);
nand U2817 (N_2817,N_2734,N_2736);
nand U2818 (N_2818,N_2723,N_2733);
or U2819 (N_2819,N_2712,N_2773);
and U2820 (N_2820,N_2703,N_2727);
or U2821 (N_2821,N_2788,N_2798);
nand U2822 (N_2822,N_2708,N_2755);
or U2823 (N_2823,N_2789,N_2793);
or U2824 (N_2824,N_2731,N_2715);
or U2825 (N_2825,N_2719,N_2781);
xor U2826 (N_2826,N_2758,N_2756);
nand U2827 (N_2827,N_2761,N_2701);
xnor U2828 (N_2828,N_2718,N_2744);
nor U2829 (N_2829,N_2726,N_2737);
xor U2830 (N_2830,N_2738,N_2709);
and U2831 (N_2831,N_2704,N_2741);
xor U2832 (N_2832,N_2710,N_2777);
nor U2833 (N_2833,N_2785,N_2795);
nor U2834 (N_2834,N_2735,N_2770);
nor U2835 (N_2835,N_2721,N_2746);
nor U2836 (N_2836,N_2724,N_2743);
and U2837 (N_2837,N_2759,N_2748);
or U2838 (N_2838,N_2729,N_2791);
or U2839 (N_2839,N_2797,N_2796);
nor U2840 (N_2840,N_2705,N_2707);
xor U2841 (N_2841,N_2760,N_2767);
xnor U2842 (N_2842,N_2799,N_2702);
nor U2843 (N_2843,N_2774,N_2765);
or U2844 (N_2844,N_2750,N_2725);
and U2845 (N_2845,N_2779,N_2787);
and U2846 (N_2846,N_2752,N_2763);
and U2847 (N_2847,N_2711,N_2794);
nor U2848 (N_2848,N_2757,N_2751);
xor U2849 (N_2849,N_2739,N_2790);
nand U2850 (N_2850,N_2706,N_2720);
nor U2851 (N_2851,N_2768,N_2747);
xor U2852 (N_2852,N_2739,N_2769);
and U2853 (N_2853,N_2770,N_2701);
and U2854 (N_2854,N_2784,N_2738);
and U2855 (N_2855,N_2737,N_2752);
nand U2856 (N_2856,N_2760,N_2750);
nand U2857 (N_2857,N_2716,N_2720);
and U2858 (N_2858,N_2763,N_2749);
or U2859 (N_2859,N_2704,N_2772);
xor U2860 (N_2860,N_2718,N_2767);
nor U2861 (N_2861,N_2785,N_2764);
xor U2862 (N_2862,N_2753,N_2723);
or U2863 (N_2863,N_2792,N_2723);
and U2864 (N_2864,N_2718,N_2733);
nand U2865 (N_2865,N_2783,N_2793);
nand U2866 (N_2866,N_2719,N_2756);
xnor U2867 (N_2867,N_2715,N_2789);
xnor U2868 (N_2868,N_2758,N_2796);
nor U2869 (N_2869,N_2709,N_2784);
nor U2870 (N_2870,N_2797,N_2733);
nor U2871 (N_2871,N_2763,N_2751);
xor U2872 (N_2872,N_2754,N_2777);
and U2873 (N_2873,N_2737,N_2711);
nand U2874 (N_2874,N_2763,N_2788);
nor U2875 (N_2875,N_2799,N_2767);
nor U2876 (N_2876,N_2716,N_2711);
or U2877 (N_2877,N_2748,N_2711);
nor U2878 (N_2878,N_2707,N_2724);
and U2879 (N_2879,N_2789,N_2772);
nand U2880 (N_2880,N_2720,N_2765);
and U2881 (N_2881,N_2702,N_2772);
and U2882 (N_2882,N_2762,N_2743);
nor U2883 (N_2883,N_2736,N_2778);
or U2884 (N_2884,N_2705,N_2718);
nand U2885 (N_2885,N_2740,N_2778);
and U2886 (N_2886,N_2782,N_2771);
nor U2887 (N_2887,N_2784,N_2771);
and U2888 (N_2888,N_2761,N_2749);
nor U2889 (N_2889,N_2719,N_2714);
nor U2890 (N_2890,N_2724,N_2711);
nor U2891 (N_2891,N_2742,N_2765);
and U2892 (N_2892,N_2757,N_2719);
nor U2893 (N_2893,N_2784,N_2714);
and U2894 (N_2894,N_2761,N_2711);
nor U2895 (N_2895,N_2763,N_2767);
nand U2896 (N_2896,N_2776,N_2798);
nand U2897 (N_2897,N_2753,N_2710);
nor U2898 (N_2898,N_2789,N_2756);
xnor U2899 (N_2899,N_2703,N_2715);
and U2900 (N_2900,N_2815,N_2889);
xnor U2901 (N_2901,N_2806,N_2820);
nand U2902 (N_2902,N_2816,N_2845);
xor U2903 (N_2903,N_2800,N_2812);
or U2904 (N_2904,N_2857,N_2896);
or U2905 (N_2905,N_2855,N_2814);
or U2906 (N_2906,N_2831,N_2848);
and U2907 (N_2907,N_2866,N_2849);
xnor U2908 (N_2908,N_2832,N_2830);
or U2909 (N_2909,N_2876,N_2861);
nand U2910 (N_2910,N_2827,N_2894);
and U2911 (N_2911,N_2893,N_2883);
or U2912 (N_2912,N_2881,N_2825);
and U2913 (N_2913,N_2898,N_2890);
or U2914 (N_2914,N_2859,N_2874);
xnor U2915 (N_2915,N_2873,N_2877);
xnor U2916 (N_2916,N_2836,N_2875);
nor U2917 (N_2917,N_2810,N_2835);
nand U2918 (N_2918,N_2805,N_2853);
and U2919 (N_2919,N_2838,N_2884);
nor U2920 (N_2920,N_2870,N_2887);
nor U2921 (N_2921,N_2868,N_2844);
nor U2922 (N_2922,N_2897,N_2839);
nor U2923 (N_2923,N_2801,N_2811);
nand U2924 (N_2924,N_2864,N_2886);
or U2925 (N_2925,N_2809,N_2860);
and U2926 (N_2926,N_2823,N_2888);
and U2927 (N_2927,N_2854,N_2841);
nor U2928 (N_2928,N_2872,N_2802);
nand U2929 (N_2929,N_2899,N_2895);
or U2930 (N_2930,N_2818,N_2813);
nor U2931 (N_2931,N_2847,N_2850);
nand U2932 (N_2932,N_2843,N_2882);
nand U2933 (N_2933,N_2807,N_2826);
nor U2934 (N_2934,N_2858,N_2892);
or U2935 (N_2935,N_2829,N_2846);
nand U2936 (N_2936,N_2834,N_2803);
nor U2937 (N_2937,N_2819,N_2822);
xnor U2938 (N_2938,N_2862,N_2851);
or U2939 (N_2939,N_2865,N_2828);
and U2940 (N_2940,N_2891,N_2842);
and U2941 (N_2941,N_2837,N_2852);
or U2942 (N_2942,N_2833,N_2863);
and U2943 (N_2943,N_2804,N_2879);
and U2944 (N_2944,N_2817,N_2840);
or U2945 (N_2945,N_2808,N_2871);
or U2946 (N_2946,N_2885,N_2824);
nor U2947 (N_2947,N_2869,N_2821);
and U2948 (N_2948,N_2878,N_2856);
xnor U2949 (N_2949,N_2867,N_2880);
or U2950 (N_2950,N_2892,N_2888);
xnor U2951 (N_2951,N_2844,N_2831);
nor U2952 (N_2952,N_2810,N_2858);
xnor U2953 (N_2953,N_2897,N_2835);
and U2954 (N_2954,N_2822,N_2895);
nor U2955 (N_2955,N_2880,N_2816);
or U2956 (N_2956,N_2805,N_2827);
nand U2957 (N_2957,N_2815,N_2856);
or U2958 (N_2958,N_2824,N_2842);
and U2959 (N_2959,N_2849,N_2816);
xor U2960 (N_2960,N_2880,N_2832);
nor U2961 (N_2961,N_2873,N_2897);
nand U2962 (N_2962,N_2820,N_2836);
nor U2963 (N_2963,N_2864,N_2806);
or U2964 (N_2964,N_2814,N_2819);
or U2965 (N_2965,N_2861,N_2879);
or U2966 (N_2966,N_2873,N_2867);
or U2967 (N_2967,N_2889,N_2882);
and U2968 (N_2968,N_2840,N_2877);
and U2969 (N_2969,N_2833,N_2818);
or U2970 (N_2970,N_2864,N_2869);
or U2971 (N_2971,N_2812,N_2877);
xor U2972 (N_2972,N_2857,N_2878);
nand U2973 (N_2973,N_2825,N_2819);
nand U2974 (N_2974,N_2811,N_2867);
and U2975 (N_2975,N_2805,N_2871);
or U2976 (N_2976,N_2853,N_2883);
nor U2977 (N_2977,N_2805,N_2845);
and U2978 (N_2978,N_2856,N_2889);
or U2979 (N_2979,N_2869,N_2823);
and U2980 (N_2980,N_2814,N_2894);
nor U2981 (N_2981,N_2810,N_2861);
nor U2982 (N_2982,N_2889,N_2820);
xnor U2983 (N_2983,N_2839,N_2867);
nand U2984 (N_2984,N_2897,N_2860);
or U2985 (N_2985,N_2899,N_2841);
xor U2986 (N_2986,N_2895,N_2804);
nor U2987 (N_2987,N_2826,N_2810);
nand U2988 (N_2988,N_2830,N_2898);
or U2989 (N_2989,N_2873,N_2864);
nand U2990 (N_2990,N_2816,N_2839);
or U2991 (N_2991,N_2855,N_2852);
nand U2992 (N_2992,N_2864,N_2877);
nor U2993 (N_2993,N_2874,N_2835);
nor U2994 (N_2994,N_2829,N_2838);
nand U2995 (N_2995,N_2810,N_2893);
and U2996 (N_2996,N_2870,N_2843);
and U2997 (N_2997,N_2835,N_2863);
nor U2998 (N_2998,N_2888,N_2840);
and U2999 (N_2999,N_2805,N_2821);
xnor UO_0 (O_0,N_2937,N_2939);
nor UO_1 (O_1,N_2959,N_2915);
or UO_2 (O_2,N_2921,N_2918);
and UO_3 (O_3,N_2982,N_2947);
and UO_4 (O_4,N_2944,N_2957);
nand UO_5 (O_5,N_2953,N_2994);
or UO_6 (O_6,N_2930,N_2988);
nor UO_7 (O_7,N_2903,N_2902);
xnor UO_8 (O_8,N_2901,N_2911);
and UO_9 (O_9,N_2990,N_2907);
xnor UO_10 (O_10,N_2931,N_2934);
nand UO_11 (O_11,N_2908,N_2912);
xnor UO_12 (O_12,N_2932,N_2987);
and UO_13 (O_13,N_2964,N_2967);
nor UO_14 (O_14,N_2913,N_2972);
xor UO_15 (O_15,N_2979,N_2941);
nor UO_16 (O_16,N_2976,N_2996);
nor UO_17 (O_17,N_2991,N_2949);
or UO_18 (O_18,N_2951,N_2927);
xnor UO_19 (O_19,N_2943,N_2998);
nand UO_20 (O_20,N_2954,N_2929);
or UO_21 (O_21,N_2922,N_2905);
and UO_22 (O_22,N_2935,N_2983);
and UO_23 (O_23,N_2970,N_2936);
nor UO_24 (O_24,N_2933,N_2963);
xor UO_25 (O_25,N_2993,N_2909);
xor UO_26 (O_26,N_2985,N_2975);
or UO_27 (O_27,N_2956,N_2984);
nor UO_28 (O_28,N_2960,N_2950);
xnor UO_29 (O_29,N_2992,N_2952);
nor UO_30 (O_30,N_2978,N_2955);
xnor UO_31 (O_31,N_2904,N_2923);
nor UO_32 (O_32,N_2958,N_2977);
nor UO_33 (O_33,N_2919,N_2914);
nand UO_34 (O_34,N_2948,N_2968);
xnor UO_35 (O_35,N_2946,N_2969);
or UO_36 (O_36,N_2974,N_2962);
nor UO_37 (O_37,N_2980,N_2999);
and UO_38 (O_38,N_2906,N_2986);
xor UO_39 (O_39,N_2910,N_2925);
nand UO_40 (O_40,N_2973,N_2989);
nor UO_41 (O_41,N_2965,N_2916);
or UO_42 (O_42,N_2940,N_2995);
nor UO_43 (O_43,N_2926,N_2961);
xnor UO_44 (O_44,N_2966,N_2997);
xor UO_45 (O_45,N_2938,N_2981);
and UO_46 (O_46,N_2971,N_2942);
xor UO_47 (O_47,N_2920,N_2917);
and UO_48 (O_48,N_2945,N_2928);
and UO_49 (O_49,N_2924,N_2900);
and UO_50 (O_50,N_2998,N_2997);
nand UO_51 (O_51,N_2911,N_2994);
nand UO_52 (O_52,N_2946,N_2941);
or UO_53 (O_53,N_2957,N_2963);
or UO_54 (O_54,N_2928,N_2969);
and UO_55 (O_55,N_2920,N_2945);
nor UO_56 (O_56,N_2905,N_2924);
and UO_57 (O_57,N_2902,N_2909);
and UO_58 (O_58,N_2968,N_2956);
xnor UO_59 (O_59,N_2963,N_2922);
or UO_60 (O_60,N_2907,N_2951);
nor UO_61 (O_61,N_2912,N_2913);
nor UO_62 (O_62,N_2970,N_2915);
or UO_63 (O_63,N_2945,N_2994);
and UO_64 (O_64,N_2957,N_2955);
nor UO_65 (O_65,N_2959,N_2938);
and UO_66 (O_66,N_2941,N_2915);
nor UO_67 (O_67,N_2954,N_2946);
and UO_68 (O_68,N_2939,N_2948);
nand UO_69 (O_69,N_2911,N_2950);
or UO_70 (O_70,N_2992,N_2923);
or UO_71 (O_71,N_2995,N_2955);
or UO_72 (O_72,N_2983,N_2907);
and UO_73 (O_73,N_2950,N_2930);
or UO_74 (O_74,N_2926,N_2942);
nor UO_75 (O_75,N_2977,N_2973);
nand UO_76 (O_76,N_2905,N_2981);
xnor UO_77 (O_77,N_2973,N_2903);
xnor UO_78 (O_78,N_2946,N_2998);
nor UO_79 (O_79,N_2974,N_2970);
nand UO_80 (O_80,N_2905,N_2961);
nor UO_81 (O_81,N_2906,N_2937);
xor UO_82 (O_82,N_2912,N_2970);
nand UO_83 (O_83,N_2968,N_2946);
or UO_84 (O_84,N_2934,N_2982);
nand UO_85 (O_85,N_2901,N_2939);
or UO_86 (O_86,N_2944,N_2914);
or UO_87 (O_87,N_2926,N_2918);
nor UO_88 (O_88,N_2958,N_2926);
xor UO_89 (O_89,N_2956,N_2980);
nor UO_90 (O_90,N_2946,N_2945);
nand UO_91 (O_91,N_2929,N_2938);
nand UO_92 (O_92,N_2921,N_2957);
nor UO_93 (O_93,N_2915,N_2967);
or UO_94 (O_94,N_2919,N_2999);
nor UO_95 (O_95,N_2978,N_2986);
or UO_96 (O_96,N_2970,N_2983);
nand UO_97 (O_97,N_2943,N_2932);
or UO_98 (O_98,N_2922,N_2989);
nand UO_99 (O_99,N_2922,N_2995);
or UO_100 (O_100,N_2947,N_2952);
and UO_101 (O_101,N_2997,N_2967);
and UO_102 (O_102,N_2917,N_2963);
nor UO_103 (O_103,N_2917,N_2950);
or UO_104 (O_104,N_2922,N_2964);
or UO_105 (O_105,N_2946,N_2901);
xor UO_106 (O_106,N_2912,N_2999);
xnor UO_107 (O_107,N_2951,N_2972);
xnor UO_108 (O_108,N_2972,N_2911);
or UO_109 (O_109,N_2954,N_2969);
nand UO_110 (O_110,N_2907,N_2955);
nand UO_111 (O_111,N_2976,N_2973);
xnor UO_112 (O_112,N_2954,N_2930);
and UO_113 (O_113,N_2992,N_2901);
xnor UO_114 (O_114,N_2909,N_2986);
nor UO_115 (O_115,N_2942,N_2918);
and UO_116 (O_116,N_2994,N_2904);
and UO_117 (O_117,N_2961,N_2984);
nor UO_118 (O_118,N_2954,N_2918);
or UO_119 (O_119,N_2946,N_2966);
or UO_120 (O_120,N_2936,N_2988);
and UO_121 (O_121,N_2951,N_2934);
and UO_122 (O_122,N_2937,N_2940);
nand UO_123 (O_123,N_2940,N_2931);
nand UO_124 (O_124,N_2983,N_2932);
nor UO_125 (O_125,N_2909,N_2918);
and UO_126 (O_126,N_2913,N_2998);
or UO_127 (O_127,N_2903,N_2943);
nor UO_128 (O_128,N_2964,N_2921);
or UO_129 (O_129,N_2905,N_2901);
nand UO_130 (O_130,N_2949,N_2901);
and UO_131 (O_131,N_2914,N_2907);
or UO_132 (O_132,N_2930,N_2953);
or UO_133 (O_133,N_2978,N_2946);
or UO_134 (O_134,N_2941,N_2916);
or UO_135 (O_135,N_2920,N_2978);
nand UO_136 (O_136,N_2943,N_2907);
and UO_137 (O_137,N_2932,N_2914);
xor UO_138 (O_138,N_2991,N_2956);
and UO_139 (O_139,N_2926,N_2931);
nand UO_140 (O_140,N_2956,N_2954);
and UO_141 (O_141,N_2989,N_2929);
or UO_142 (O_142,N_2938,N_2917);
or UO_143 (O_143,N_2995,N_2983);
and UO_144 (O_144,N_2986,N_2905);
and UO_145 (O_145,N_2945,N_2921);
xor UO_146 (O_146,N_2918,N_2929);
nand UO_147 (O_147,N_2947,N_2937);
xor UO_148 (O_148,N_2963,N_2939);
or UO_149 (O_149,N_2971,N_2978);
and UO_150 (O_150,N_2918,N_2986);
and UO_151 (O_151,N_2955,N_2929);
xnor UO_152 (O_152,N_2905,N_2900);
xor UO_153 (O_153,N_2954,N_2989);
nand UO_154 (O_154,N_2920,N_2977);
xnor UO_155 (O_155,N_2958,N_2951);
xnor UO_156 (O_156,N_2913,N_2999);
nand UO_157 (O_157,N_2921,N_2936);
and UO_158 (O_158,N_2965,N_2926);
xnor UO_159 (O_159,N_2965,N_2978);
and UO_160 (O_160,N_2965,N_2920);
xnor UO_161 (O_161,N_2996,N_2997);
nor UO_162 (O_162,N_2955,N_2994);
nand UO_163 (O_163,N_2982,N_2930);
nor UO_164 (O_164,N_2930,N_2906);
nor UO_165 (O_165,N_2909,N_2938);
xnor UO_166 (O_166,N_2994,N_2995);
and UO_167 (O_167,N_2931,N_2918);
xnor UO_168 (O_168,N_2911,N_2977);
xor UO_169 (O_169,N_2984,N_2910);
and UO_170 (O_170,N_2939,N_2981);
or UO_171 (O_171,N_2907,N_2973);
xor UO_172 (O_172,N_2965,N_2957);
nor UO_173 (O_173,N_2922,N_2973);
or UO_174 (O_174,N_2976,N_2931);
nand UO_175 (O_175,N_2918,N_2966);
xnor UO_176 (O_176,N_2999,N_2966);
nand UO_177 (O_177,N_2958,N_2942);
or UO_178 (O_178,N_2995,N_2977);
and UO_179 (O_179,N_2963,N_2931);
nand UO_180 (O_180,N_2981,N_2920);
or UO_181 (O_181,N_2978,N_2932);
and UO_182 (O_182,N_2982,N_2975);
nor UO_183 (O_183,N_2955,N_2963);
or UO_184 (O_184,N_2916,N_2901);
or UO_185 (O_185,N_2936,N_2956);
or UO_186 (O_186,N_2976,N_2987);
xor UO_187 (O_187,N_2976,N_2948);
nor UO_188 (O_188,N_2993,N_2945);
xor UO_189 (O_189,N_2905,N_2934);
xnor UO_190 (O_190,N_2923,N_2902);
xor UO_191 (O_191,N_2931,N_2990);
or UO_192 (O_192,N_2948,N_2965);
xor UO_193 (O_193,N_2958,N_2914);
and UO_194 (O_194,N_2963,N_2999);
nor UO_195 (O_195,N_2952,N_2900);
nand UO_196 (O_196,N_2945,N_2960);
nand UO_197 (O_197,N_2989,N_2953);
nor UO_198 (O_198,N_2981,N_2906);
or UO_199 (O_199,N_2925,N_2931);
nand UO_200 (O_200,N_2949,N_2926);
nor UO_201 (O_201,N_2904,N_2953);
and UO_202 (O_202,N_2954,N_2953);
or UO_203 (O_203,N_2933,N_2907);
xor UO_204 (O_204,N_2927,N_2982);
and UO_205 (O_205,N_2948,N_2904);
nand UO_206 (O_206,N_2929,N_2921);
or UO_207 (O_207,N_2965,N_2947);
xnor UO_208 (O_208,N_2910,N_2922);
or UO_209 (O_209,N_2973,N_2947);
and UO_210 (O_210,N_2983,N_2939);
xor UO_211 (O_211,N_2955,N_2973);
and UO_212 (O_212,N_2972,N_2971);
or UO_213 (O_213,N_2985,N_2938);
nand UO_214 (O_214,N_2935,N_2990);
nor UO_215 (O_215,N_2913,N_2947);
or UO_216 (O_216,N_2965,N_2968);
and UO_217 (O_217,N_2952,N_2924);
or UO_218 (O_218,N_2918,N_2913);
nand UO_219 (O_219,N_2990,N_2975);
nor UO_220 (O_220,N_2949,N_2932);
or UO_221 (O_221,N_2946,N_2902);
nand UO_222 (O_222,N_2994,N_2903);
nor UO_223 (O_223,N_2960,N_2947);
or UO_224 (O_224,N_2916,N_2913);
nand UO_225 (O_225,N_2966,N_2962);
or UO_226 (O_226,N_2974,N_2997);
xor UO_227 (O_227,N_2971,N_2975);
nor UO_228 (O_228,N_2935,N_2952);
and UO_229 (O_229,N_2979,N_2910);
nand UO_230 (O_230,N_2967,N_2944);
and UO_231 (O_231,N_2983,N_2962);
or UO_232 (O_232,N_2960,N_2928);
nand UO_233 (O_233,N_2906,N_2913);
nor UO_234 (O_234,N_2932,N_2918);
or UO_235 (O_235,N_2967,N_2994);
or UO_236 (O_236,N_2969,N_2964);
nor UO_237 (O_237,N_2905,N_2948);
nor UO_238 (O_238,N_2975,N_2963);
nand UO_239 (O_239,N_2940,N_2958);
xor UO_240 (O_240,N_2963,N_2992);
xnor UO_241 (O_241,N_2994,N_2926);
nand UO_242 (O_242,N_2901,N_2935);
nand UO_243 (O_243,N_2951,N_2906);
and UO_244 (O_244,N_2994,N_2988);
nor UO_245 (O_245,N_2984,N_2948);
or UO_246 (O_246,N_2907,N_2977);
nand UO_247 (O_247,N_2902,N_2940);
xnor UO_248 (O_248,N_2911,N_2979);
xor UO_249 (O_249,N_2993,N_2995);
and UO_250 (O_250,N_2970,N_2940);
nor UO_251 (O_251,N_2931,N_2979);
or UO_252 (O_252,N_2928,N_2918);
xor UO_253 (O_253,N_2960,N_2988);
xor UO_254 (O_254,N_2924,N_2922);
nor UO_255 (O_255,N_2912,N_2906);
nand UO_256 (O_256,N_2975,N_2980);
or UO_257 (O_257,N_2952,N_2986);
and UO_258 (O_258,N_2903,N_2984);
nor UO_259 (O_259,N_2927,N_2977);
and UO_260 (O_260,N_2984,N_2955);
or UO_261 (O_261,N_2922,N_2987);
or UO_262 (O_262,N_2900,N_2989);
nor UO_263 (O_263,N_2951,N_2910);
xnor UO_264 (O_264,N_2921,N_2914);
or UO_265 (O_265,N_2939,N_2993);
xor UO_266 (O_266,N_2900,N_2933);
nand UO_267 (O_267,N_2953,N_2957);
or UO_268 (O_268,N_2954,N_2912);
nor UO_269 (O_269,N_2954,N_2992);
xnor UO_270 (O_270,N_2926,N_2973);
and UO_271 (O_271,N_2903,N_2926);
nand UO_272 (O_272,N_2902,N_2959);
nor UO_273 (O_273,N_2998,N_2992);
or UO_274 (O_274,N_2927,N_2985);
nor UO_275 (O_275,N_2982,N_2937);
or UO_276 (O_276,N_2985,N_2965);
and UO_277 (O_277,N_2916,N_2966);
xnor UO_278 (O_278,N_2909,N_2968);
nor UO_279 (O_279,N_2900,N_2987);
xnor UO_280 (O_280,N_2907,N_2949);
nand UO_281 (O_281,N_2922,N_2985);
xnor UO_282 (O_282,N_2915,N_2906);
nand UO_283 (O_283,N_2900,N_2930);
xor UO_284 (O_284,N_2916,N_2972);
nand UO_285 (O_285,N_2928,N_2942);
or UO_286 (O_286,N_2945,N_2988);
and UO_287 (O_287,N_2914,N_2900);
and UO_288 (O_288,N_2979,N_2933);
nor UO_289 (O_289,N_2911,N_2939);
or UO_290 (O_290,N_2977,N_2952);
xor UO_291 (O_291,N_2946,N_2952);
nor UO_292 (O_292,N_2996,N_2958);
nand UO_293 (O_293,N_2934,N_2987);
xor UO_294 (O_294,N_2901,N_2970);
and UO_295 (O_295,N_2991,N_2911);
nor UO_296 (O_296,N_2941,N_2957);
nor UO_297 (O_297,N_2931,N_2947);
nor UO_298 (O_298,N_2954,N_2983);
nor UO_299 (O_299,N_2996,N_2989);
xnor UO_300 (O_300,N_2945,N_2944);
nor UO_301 (O_301,N_2971,N_2969);
nand UO_302 (O_302,N_2947,N_2904);
nand UO_303 (O_303,N_2982,N_2998);
nor UO_304 (O_304,N_2900,N_2967);
nand UO_305 (O_305,N_2927,N_2934);
or UO_306 (O_306,N_2935,N_2961);
nor UO_307 (O_307,N_2906,N_2969);
or UO_308 (O_308,N_2994,N_2966);
or UO_309 (O_309,N_2949,N_2980);
or UO_310 (O_310,N_2935,N_2930);
nor UO_311 (O_311,N_2909,N_2941);
or UO_312 (O_312,N_2921,N_2941);
xor UO_313 (O_313,N_2974,N_2950);
or UO_314 (O_314,N_2914,N_2983);
and UO_315 (O_315,N_2920,N_2975);
xnor UO_316 (O_316,N_2967,N_2943);
xnor UO_317 (O_317,N_2960,N_2983);
nand UO_318 (O_318,N_2998,N_2957);
or UO_319 (O_319,N_2961,N_2999);
nor UO_320 (O_320,N_2934,N_2992);
xor UO_321 (O_321,N_2999,N_2921);
and UO_322 (O_322,N_2912,N_2997);
xnor UO_323 (O_323,N_2902,N_2977);
nand UO_324 (O_324,N_2905,N_2959);
nand UO_325 (O_325,N_2908,N_2905);
xor UO_326 (O_326,N_2934,N_2917);
nor UO_327 (O_327,N_2946,N_2920);
or UO_328 (O_328,N_2951,N_2990);
nor UO_329 (O_329,N_2932,N_2937);
or UO_330 (O_330,N_2944,N_2973);
nand UO_331 (O_331,N_2923,N_2956);
nand UO_332 (O_332,N_2936,N_2945);
nor UO_333 (O_333,N_2962,N_2905);
nand UO_334 (O_334,N_2905,N_2943);
or UO_335 (O_335,N_2985,N_2915);
nor UO_336 (O_336,N_2961,N_2909);
nor UO_337 (O_337,N_2992,N_2981);
and UO_338 (O_338,N_2925,N_2971);
or UO_339 (O_339,N_2957,N_2929);
xnor UO_340 (O_340,N_2930,N_2911);
and UO_341 (O_341,N_2909,N_2991);
nor UO_342 (O_342,N_2995,N_2907);
or UO_343 (O_343,N_2932,N_2948);
xor UO_344 (O_344,N_2912,N_2903);
xor UO_345 (O_345,N_2902,N_2991);
nor UO_346 (O_346,N_2908,N_2982);
or UO_347 (O_347,N_2994,N_2987);
nor UO_348 (O_348,N_2960,N_2965);
or UO_349 (O_349,N_2943,N_2939);
and UO_350 (O_350,N_2907,N_2945);
nand UO_351 (O_351,N_2931,N_2915);
nand UO_352 (O_352,N_2948,N_2933);
and UO_353 (O_353,N_2919,N_2943);
nor UO_354 (O_354,N_2916,N_2930);
nand UO_355 (O_355,N_2941,N_2905);
and UO_356 (O_356,N_2911,N_2995);
or UO_357 (O_357,N_2957,N_2974);
nor UO_358 (O_358,N_2906,N_2997);
nand UO_359 (O_359,N_2951,N_2903);
xor UO_360 (O_360,N_2960,N_2944);
and UO_361 (O_361,N_2957,N_2988);
and UO_362 (O_362,N_2983,N_2924);
or UO_363 (O_363,N_2992,N_2920);
or UO_364 (O_364,N_2935,N_2944);
nor UO_365 (O_365,N_2958,N_2964);
and UO_366 (O_366,N_2915,N_2990);
xor UO_367 (O_367,N_2950,N_2970);
nand UO_368 (O_368,N_2993,N_2959);
xnor UO_369 (O_369,N_2991,N_2993);
and UO_370 (O_370,N_2974,N_2978);
and UO_371 (O_371,N_2907,N_2994);
xor UO_372 (O_372,N_2993,N_2964);
nand UO_373 (O_373,N_2995,N_2981);
nor UO_374 (O_374,N_2943,N_2971);
and UO_375 (O_375,N_2938,N_2933);
nand UO_376 (O_376,N_2971,N_2986);
xnor UO_377 (O_377,N_2988,N_2980);
xor UO_378 (O_378,N_2976,N_2979);
or UO_379 (O_379,N_2902,N_2918);
or UO_380 (O_380,N_2902,N_2978);
nand UO_381 (O_381,N_2963,N_2934);
or UO_382 (O_382,N_2985,N_2947);
xnor UO_383 (O_383,N_2979,N_2996);
xor UO_384 (O_384,N_2900,N_2973);
nand UO_385 (O_385,N_2912,N_2992);
nor UO_386 (O_386,N_2954,N_2924);
or UO_387 (O_387,N_2969,N_2949);
xor UO_388 (O_388,N_2957,N_2985);
and UO_389 (O_389,N_2930,N_2914);
and UO_390 (O_390,N_2940,N_2987);
nand UO_391 (O_391,N_2923,N_2962);
and UO_392 (O_392,N_2974,N_2938);
or UO_393 (O_393,N_2901,N_2969);
and UO_394 (O_394,N_2953,N_2915);
nor UO_395 (O_395,N_2998,N_2954);
nand UO_396 (O_396,N_2933,N_2951);
xor UO_397 (O_397,N_2900,N_2942);
nor UO_398 (O_398,N_2991,N_2908);
nor UO_399 (O_399,N_2962,N_2995);
nor UO_400 (O_400,N_2974,N_2910);
nand UO_401 (O_401,N_2943,N_2969);
and UO_402 (O_402,N_2982,N_2996);
nor UO_403 (O_403,N_2930,N_2904);
nand UO_404 (O_404,N_2950,N_2942);
and UO_405 (O_405,N_2953,N_2944);
xor UO_406 (O_406,N_2956,N_2900);
xor UO_407 (O_407,N_2981,N_2911);
xnor UO_408 (O_408,N_2976,N_2949);
or UO_409 (O_409,N_2996,N_2941);
nand UO_410 (O_410,N_2967,N_2966);
xor UO_411 (O_411,N_2965,N_2941);
and UO_412 (O_412,N_2915,N_2945);
and UO_413 (O_413,N_2931,N_2920);
xor UO_414 (O_414,N_2936,N_2937);
xnor UO_415 (O_415,N_2923,N_2950);
and UO_416 (O_416,N_2930,N_2961);
xor UO_417 (O_417,N_2928,N_2922);
nor UO_418 (O_418,N_2967,N_2914);
xnor UO_419 (O_419,N_2983,N_2994);
or UO_420 (O_420,N_2909,N_2945);
xnor UO_421 (O_421,N_2912,N_2994);
nor UO_422 (O_422,N_2952,N_2917);
or UO_423 (O_423,N_2909,N_2965);
or UO_424 (O_424,N_2956,N_2994);
or UO_425 (O_425,N_2994,N_2915);
nand UO_426 (O_426,N_2933,N_2944);
nand UO_427 (O_427,N_2927,N_2912);
nand UO_428 (O_428,N_2982,N_2949);
nand UO_429 (O_429,N_2978,N_2985);
xnor UO_430 (O_430,N_2949,N_2910);
nor UO_431 (O_431,N_2937,N_2983);
xor UO_432 (O_432,N_2954,N_2933);
nor UO_433 (O_433,N_2910,N_2973);
and UO_434 (O_434,N_2948,N_2987);
xnor UO_435 (O_435,N_2948,N_2954);
xnor UO_436 (O_436,N_2973,N_2939);
or UO_437 (O_437,N_2944,N_2936);
and UO_438 (O_438,N_2954,N_2985);
nand UO_439 (O_439,N_2920,N_2995);
xnor UO_440 (O_440,N_2947,N_2964);
or UO_441 (O_441,N_2909,N_2911);
and UO_442 (O_442,N_2998,N_2903);
and UO_443 (O_443,N_2994,N_2976);
or UO_444 (O_444,N_2904,N_2990);
and UO_445 (O_445,N_2948,N_2972);
nor UO_446 (O_446,N_2937,N_2975);
nor UO_447 (O_447,N_2979,N_2921);
or UO_448 (O_448,N_2910,N_2985);
or UO_449 (O_449,N_2970,N_2945);
and UO_450 (O_450,N_2973,N_2942);
nor UO_451 (O_451,N_2903,N_2955);
nand UO_452 (O_452,N_2910,N_2950);
nor UO_453 (O_453,N_2962,N_2997);
nand UO_454 (O_454,N_2992,N_2910);
and UO_455 (O_455,N_2970,N_2955);
and UO_456 (O_456,N_2919,N_2985);
nor UO_457 (O_457,N_2920,N_2967);
nand UO_458 (O_458,N_2992,N_2911);
or UO_459 (O_459,N_2912,N_2931);
xor UO_460 (O_460,N_2999,N_2975);
nand UO_461 (O_461,N_2997,N_2960);
or UO_462 (O_462,N_2977,N_2901);
or UO_463 (O_463,N_2991,N_2969);
xor UO_464 (O_464,N_2984,N_2967);
nand UO_465 (O_465,N_2931,N_2987);
xor UO_466 (O_466,N_2916,N_2943);
and UO_467 (O_467,N_2944,N_2925);
xor UO_468 (O_468,N_2982,N_2944);
xor UO_469 (O_469,N_2942,N_2909);
nand UO_470 (O_470,N_2977,N_2968);
or UO_471 (O_471,N_2909,N_2960);
nor UO_472 (O_472,N_2951,N_2941);
or UO_473 (O_473,N_2921,N_2975);
xor UO_474 (O_474,N_2914,N_2954);
and UO_475 (O_475,N_2941,N_2986);
or UO_476 (O_476,N_2939,N_2975);
nand UO_477 (O_477,N_2904,N_2961);
nor UO_478 (O_478,N_2936,N_2913);
or UO_479 (O_479,N_2913,N_2965);
or UO_480 (O_480,N_2970,N_2985);
and UO_481 (O_481,N_2949,N_2986);
nand UO_482 (O_482,N_2929,N_2967);
nor UO_483 (O_483,N_2980,N_2906);
or UO_484 (O_484,N_2954,N_2972);
nand UO_485 (O_485,N_2912,N_2969);
nand UO_486 (O_486,N_2918,N_2969);
and UO_487 (O_487,N_2990,N_2949);
xnor UO_488 (O_488,N_2925,N_2964);
and UO_489 (O_489,N_2921,N_2950);
and UO_490 (O_490,N_2911,N_2998);
nand UO_491 (O_491,N_2900,N_2978);
or UO_492 (O_492,N_2967,N_2985);
nand UO_493 (O_493,N_2965,N_2914);
xor UO_494 (O_494,N_2935,N_2946);
nand UO_495 (O_495,N_2950,N_2906);
nand UO_496 (O_496,N_2901,N_2966);
nor UO_497 (O_497,N_2922,N_2933);
xnor UO_498 (O_498,N_2946,N_2971);
nand UO_499 (O_499,N_2993,N_2982);
endmodule