module basic_500_3000_500_3_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_293,In_217);
or U1 (N_1,In_104,In_341);
or U2 (N_2,In_330,In_162);
nor U3 (N_3,In_347,In_172);
or U4 (N_4,In_411,In_321);
nand U5 (N_5,In_19,In_451);
or U6 (N_6,In_18,In_353);
and U7 (N_7,In_359,In_138);
and U8 (N_8,In_32,In_443);
or U9 (N_9,In_350,In_251);
nor U10 (N_10,In_54,In_439);
or U11 (N_11,In_271,In_144);
and U12 (N_12,In_399,In_346);
nor U13 (N_13,In_7,In_100);
nand U14 (N_14,In_35,In_428);
nand U15 (N_15,In_235,In_364);
or U16 (N_16,In_420,In_63);
nand U17 (N_17,In_183,In_328);
and U18 (N_18,In_177,In_272);
and U19 (N_19,In_440,In_64);
and U20 (N_20,In_351,In_381);
nand U21 (N_21,In_91,In_3);
and U22 (N_22,In_355,In_415);
nand U23 (N_23,In_65,In_260);
nand U24 (N_24,In_462,In_15);
and U25 (N_25,In_202,In_273);
nand U26 (N_26,In_14,In_228);
nor U27 (N_27,In_250,In_120);
and U28 (N_28,In_157,In_30);
and U29 (N_29,In_173,In_188);
nand U30 (N_30,In_189,In_2);
or U31 (N_31,In_145,In_392);
and U32 (N_32,In_71,In_77);
nand U33 (N_33,In_236,In_418);
or U34 (N_34,In_487,In_195);
and U35 (N_35,In_69,In_301);
and U36 (N_36,In_221,In_36);
nand U37 (N_37,In_17,In_51);
and U38 (N_38,In_52,In_86);
or U39 (N_39,In_410,In_229);
and U40 (N_40,In_267,In_115);
nor U41 (N_41,In_467,In_327);
nand U42 (N_42,In_149,In_358);
nand U43 (N_43,In_231,In_498);
nor U44 (N_44,In_155,In_174);
nand U45 (N_45,In_372,In_222);
nor U46 (N_46,In_335,In_279);
or U47 (N_47,In_13,In_471);
xnor U48 (N_48,In_6,In_331);
nor U49 (N_49,In_401,In_170);
nand U50 (N_50,In_379,In_31);
or U51 (N_51,In_227,In_389);
xor U52 (N_52,In_181,In_48);
or U53 (N_53,In_299,In_218);
or U54 (N_54,In_322,In_388);
or U55 (N_55,In_429,In_316);
and U56 (N_56,In_340,In_306);
xnor U57 (N_57,In_323,In_94);
and U58 (N_58,In_239,In_484);
nand U59 (N_59,In_412,In_101);
and U60 (N_60,In_194,In_404);
nand U61 (N_61,In_375,In_332);
nand U62 (N_62,In_191,In_414);
nand U63 (N_63,In_461,In_313);
nand U64 (N_64,In_24,In_136);
nand U65 (N_65,In_481,In_395);
and U66 (N_66,In_445,In_489);
or U67 (N_67,In_234,In_40);
nor U68 (N_68,In_394,In_454);
or U69 (N_69,In_465,In_84);
and U70 (N_70,In_113,In_344);
or U71 (N_71,In_237,In_102);
or U72 (N_72,In_9,In_249);
or U73 (N_73,In_44,In_472);
nor U74 (N_74,In_232,In_396);
nor U75 (N_75,In_413,In_374);
or U76 (N_76,In_49,In_398);
nor U77 (N_77,In_20,In_238);
nor U78 (N_78,In_407,In_466);
nand U79 (N_79,In_391,In_284);
nor U80 (N_80,In_342,In_380);
nor U81 (N_81,In_349,In_473);
or U82 (N_82,In_304,In_432);
nand U83 (N_83,In_156,In_494);
nand U84 (N_84,In_108,In_208);
nor U85 (N_85,In_85,In_285);
and U86 (N_86,In_290,In_164);
nor U87 (N_87,In_452,In_400);
and U88 (N_88,In_421,In_79);
nor U89 (N_89,In_135,In_456);
nor U90 (N_90,In_103,In_282);
and U91 (N_91,In_226,In_146);
and U92 (N_92,In_53,In_55);
and U93 (N_93,In_444,In_387);
and U94 (N_94,In_329,In_60);
nand U95 (N_95,In_58,In_72);
or U96 (N_96,In_75,In_118);
and U97 (N_97,In_447,In_204);
or U98 (N_98,In_325,In_38);
and U99 (N_99,In_46,In_165);
and U100 (N_100,In_116,In_326);
and U101 (N_101,In_270,In_169);
and U102 (N_102,In_119,In_151);
nand U103 (N_103,In_266,In_491);
nor U104 (N_104,In_434,In_121);
nor U105 (N_105,In_76,In_5);
and U106 (N_106,In_367,In_393);
or U107 (N_107,In_47,In_132);
nor U108 (N_108,In_314,In_89);
and U109 (N_109,In_348,In_8);
and U110 (N_110,In_137,In_496);
nor U111 (N_111,In_261,In_470);
and U112 (N_112,In_493,In_245);
nor U113 (N_113,In_406,In_219);
nand U114 (N_114,In_281,In_297);
and U115 (N_115,In_286,In_483);
or U116 (N_116,In_463,In_209);
and U117 (N_117,In_29,In_338);
and U118 (N_118,In_275,In_74);
or U119 (N_119,In_106,In_167);
nand U120 (N_120,In_424,In_438);
or U121 (N_121,In_128,In_111);
xor U122 (N_122,In_190,In_324);
and U123 (N_123,In_433,In_4);
nor U124 (N_124,In_10,In_259);
nor U125 (N_125,In_130,In_230);
nand U126 (N_126,In_223,In_352);
nor U127 (N_127,In_214,In_198);
nor U128 (N_128,In_246,In_311);
nor U129 (N_129,In_366,In_478);
or U130 (N_130,In_277,In_403);
and U131 (N_131,In_252,In_129);
nor U132 (N_132,In_464,In_337);
nand U133 (N_133,In_154,In_288);
nand U134 (N_134,In_436,In_303);
or U135 (N_135,In_240,In_242);
and U136 (N_136,In_1,In_215);
nand U137 (N_137,In_354,In_186);
nor U138 (N_138,In_482,In_131);
nor U139 (N_139,In_446,In_110);
and U140 (N_140,In_107,In_320);
or U141 (N_141,In_253,In_25);
nor U142 (N_142,In_203,In_365);
nor U143 (N_143,In_370,In_345);
nand U144 (N_144,In_161,In_216);
or U145 (N_145,In_264,In_268);
or U146 (N_146,In_476,In_402);
nand U147 (N_147,In_37,In_112);
nor U148 (N_148,In_114,In_90);
nor U149 (N_149,In_417,In_81);
and U150 (N_150,In_133,In_180);
nor U151 (N_151,In_12,In_93);
xor U152 (N_152,In_41,In_178);
or U153 (N_153,In_298,In_276);
or U154 (N_154,In_166,In_39);
nand U155 (N_155,In_66,In_373);
nor U156 (N_156,In_459,In_96);
nand U157 (N_157,In_117,In_175);
nor U158 (N_158,In_453,In_88);
nand U159 (N_159,In_292,In_333);
nand U160 (N_160,In_125,In_159);
and U161 (N_161,In_274,In_300);
and U162 (N_162,In_254,In_458);
and U163 (N_163,In_312,In_23);
nor U164 (N_164,In_139,In_184);
nand U165 (N_165,In_62,In_278);
nor U166 (N_166,In_416,In_83);
nor U167 (N_167,In_295,In_196);
nand U168 (N_168,In_449,In_78);
or U169 (N_169,In_307,In_361);
nand U170 (N_170,In_182,In_95);
nor U171 (N_171,In_435,In_386);
or U172 (N_172,In_80,In_422);
nor U173 (N_173,In_124,In_442);
nor U174 (N_174,In_244,In_360);
and U175 (N_175,In_34,In_98);
nand U176 (N_176,In_16,In_213);
and U177 (N_177,In_153,In_134);
nor U178 (N_178,In_187,In_423);
nand U179 (N_179,In_225,In_158);
and U180 (N_180,In_357,In_233);
or U181 (N_181,In_105,In_280);
and U182 (N_182,In_455,In_475);
and U183 (N_183,In_371,In_384);
nand U184 (N_184,In_368,In_287);
nor U185 (N_185,In_152,In_148);
and U186 (N_186,In_61,In_450);
nand U187 (N_187,In_383,In_241);
nand U188 (N_188,In_163,In_362);
and U189 (N_189,In_22,In_431);
and U190 (N_190,In_283,In_97);
and U191 (N_191,In_59,In_390);
nor U192 (N_192,In_457,In_206);
nand U193 (N_193,In_0,In_302);
nand U194 (N_194,In_140,In_210);
and U195 (N_195,In_319,In_176);
nor U196 (N_196,In_334,In_42);
nor U197 (N_197,In_123,In_356);
nand U198 (N_198,In_317,In_27);
nand U199 (N_199,In_171,In_291);
nor U200 (N_200,In_199,In_382);
and U201 (N_201,In_397,In_33);
and U202 (N_202,In_419,In_486);
nor U203 (N_203,In_220,In_305);
nand U204 (N_204,In_207,In_247);
xor U205 (N_205,In_426,In_50);
nand U206 (N_206,In_310,In_70);
nor U207 (N_207,In_243,In_99);
or U208 (N_208,In_309,In_460);
nand U209 (N_209,In_289,In_127);
nor U210 (N_210,In_212,In_211);
and U211 (N_211,In_109,In_67);
nor U212 (N_212,In_269,In_87);
and U213 (N_213,In_262,In_409);
or U214 (N_214,In_57,In_474);
nor U215 (N_215,In_160,In_255);
or U216 (N_216,In_92,In_318);
or U217 (N_217,In_425,In_485);
and U218 (N_218,In_448,In_480);
nor U219 (N_219,In_315,In_378);
or U220 (N_220,In_224,In_477);
and U221 (N_221,In_256,In_492);
nor U222 (N_222,In_197,In_263);
nand U223 (N_223,In_248,In_192);
and U224 (N_224,In_82,In_408);
or U225 (N_225,In_430,In_339);
nor U226 (N_226,In_490,In_308);
or U227 (N_227,In_495,In_68);
and U228 (N_228,In_343,In_168);
nor U229 (N_229,In_265,In_126);
nand U230 (N_230,In_258,In_437);
or U231 (N_231,In_179,In_143);
or U232 (N_232,In_193,In_376);
nor U233 (N_233,In_369,In_56);
or U234 (N_234,In_405,In_499);
nand U235 (N_235,In_296,In_43);
nor U236 (N_236,In_205,In_363);
nand U237 (N_237,In_497,In_257);
nand U238 (N_238,In_441,In_201);
nand U239 (N_239,In_150,In_385);
or U240 (N_240,In_73,In_469);
nand U241 (N_241,In_21,In_26);
or U242 (N_242,In_28,In_336);
and U243 (N_243,In_479,In_488);
and U244 (N_244,In_294,In_142);
nand U245 (N_245,In_141,In_122);
nand U246 (N_246,In_468,In_377);
nor U247 (N_247,In_147,In_427);
nand U248 (N_248,In_45,In_200);
nor U249 (N_249,In_185,In_11);
nor U250 (N_250,In_406,In_37);
nand U251 (N_251,In_406,In_239);
or U252 (N_252,In_418,In_35);
or U253 (N_253,In_486,In_62);
or U254 (N_254,In_86,In_189);
nor U255 (N_255,In_63,In_452);
and U256 (N_256,In_29,In_437);
nand U257 (N_257,In_72,In_438);
and U258 (N_258,In_161,In_482);
nand U259 (N_259,In_117,In_13);
and U260 (N_260,In_247,In_70);
nor U261 (N_261,In_475,In_221);
nor U262 (N_262,In_321,In_253);
and U263 (N_263,In_113,In_473);
nand U264 (N_264,In_161,In_360);
and U265 (N_265,In_21,In_369);
or U266 (N_266,In_432,In_429);
xor U267 (N_267,In_468,In_126);
nand U268 (N_268,In_481,In_68);
and U269 (N_269,In_491,In_254);
and U270 (N_270,In_363,In_459);
or U271 (N_271,In_360,In_455);
nand U272 (N_272,In_286,In_452);
and U273 (N_273,In_403,In_390);
and U274 (N_274,In_181,In_120);
or U275 (N_275,In_46,In_182);
nor U276 (N_276,In_172,In_59);
nor U277 (N_277,In_134,In_104);
and U278 (N_278,In_174,In_151);
nand U279 (N_279,In_238,In_4);
and U280 (N_280,In_148,In_468);
nor U281 (N_281,In_184,In_322);
or U282 (N_282,In_453,In_169);
nor U283 (N_283,In_148,In_341);
nand U284 (N_284,In_124,In_486);
nand U285 (N_285,In_74,In_25);
xnor U286 (N_286,In_111,In_236);
nand U287 (N_287,In_348,In_95);
and U288 (N_288,In_78,In_62);
nand U289 (N_289,In_309,In_228);
or U290 (N_290,In_120,In_45);
or U291 (N_291,In_120,In_153);
and U292 (N_292,In_158,In_470);
nor U293 (N_293,In_75,In_417);
nor U294 (N_294,In_186,In_65);
and U295 (N_295,In_297,In_164);
nor U296 (N_296,In_348,In_244);
nand U297 (N_297,In_31,In_496);
and U298 (N_298,In_227,In_64);
and U299 (N_299,In_339,In_273);
nor U300 (N_300,In_100,In_239);
or U301 (N_301,In_47,In_308);
and U302 (N_302,In_392,In_495);
and U303 (N_303,In_296,In_411);
nand U304 (N_304,In_345,In_273);
or U305 (N_305,In_133,In_424);
nand U306 (N_306,In_477,In_482);
and U307 (N_307,In_310,In_65);
nand U308 (N_308,In_104,In_292);
and U309 (N_309,In_255,In_295);
nand U310 (N_310,In_390,In_107);
nor U311 (N_311,In_269,In_93);
nor U312 (N_312,In_248,In_314);
nand U313 (N_313,In_384,In_499);
or U314 (N_314,In_194,In_99);
nor U315 (N_315,In_24,In_458);
nor U316 (N_316,In_351,In_408);
nand U317 (N_317,In_420,In_174);
or U318 (N_318,In_331,In_439);
or U319 (N_319,In_334,In_212);
nand U320 (N_320,In_468,In_74);
or U321 (N_321,In_497,In_465);
nor U322 (N_322,In_228,In_357);
nor U323 (N_323,In_228,In_54);
or U324 (N_324,In_271,In_326);
nand U325 (N_325,In_208,In_98);
and U326 (N_326,In_67,In_180);
and U327 (N_327,In_138,In_71);
nor U328 (N_328,In_400,In_31);
or U329 (N_329,In_242,In_90);
nor U330 (N_330,In_322,In_193);
or U331 (N_331,In_319,In_137);
and U332 (N_332,In_60,In_227);
and U333 (N_333,In_76,In_171);
and U334 (N_334,In_399,In_417);
or U335 (N_335,In_182,In_16);
and U336 (N_336,In_378,In_167);
or U337 (N_337,In_441,In_444);
nand U338 (N_338,In_354,In_258);
or U339 (N_339,In_143,In_180);
nor U340 (N_340,In_62,In_100);
and U341 (N_341,In_480,In_110);
xnor U342 (N_342,In_384,In_226);
and U343 (N_343,In_353,In_55);
and U344 (N_344,In_450,In_275);
and U345 (N_345,In_164,In_243);
nand U346 (N_346,In_276,In_299);
or U347 (N_347,In_453,In_474);
and U348 (N_348,In_30,In_294);
nor U349 (N_349,In_180,In_127);
nor U350 (N_350,In_30,In_20);
nor U351 (N_351,In_24,In_326);
nand U352 (N_352,In_489,In_380);
or U353 (N_353,In_189,In_139);
and U354 (N_354,In_315,In_30);
nor U355 (N_355,In_322,In_248);
nor U356 (N_356,In_52,In_449);
nand U357 (N_357,In_460,In_0);
nor U358 (N_358,In_468,In_212);
nor U359 (N_359,In_101,In_462);
nor U360 (N_360,In_472,In_405);
nor U361 (N_361,In_383,In_498);
nor U362 (N_362,In_340,In_446);
and U363 (N_363,In_284,In_222);
nand U364 (N_364,In_284,In_10);
nand U365 (N_365,In_344,In_458);
and U366 (N_366,In_260,In_111);
nand U367 (N_367,In_50,In_22);
nand U368 (N_368,In_468,In_201);
nand U369 (N_369,In_145,In_316);
or U370 (N_370,In_121,In_368);
and U371 (N_371,In_90,In_380);
and U372 (N_372,In_407,In_79);
xor U373 (N_373,In_65,In_229);
and U374 (N_374,In_202,In_380);
or U375 (N_375,In_302,In_400);
and U376 (N_376,In_126,In_469);
nand U377 (N_377,In_274,In_398);
nor U378 (N_378,In_319,In_455);
or U379 (N_379,In_23,In_153);
and U380 (N_380,In_307,In_29);
or U381 (N_381,In_441,In_221);
and U382 (N_382,In_161,In_63);
nand U383 (N_383,In_207,In_97);
or U384 (N_384,In_72,In_390);
or U385 (N_385,In_341,In_161);
and U386 (N_386,In_377,In_46);
or U387 (N_387,In_75,In_217);
and U388 (N_388,In_344,In_0);
nor U389 (N_389,In_457,In_489);
nand U390 (N_390,In_338,In_435);
nand U391 (N_391,In_298,In_145);
and U392 (N_392,In_183,In_139);
nor U393 (N_393,In_392,In_277);
or U394 (N_394,In_80,In_206);
nand U395 (N_395,In_92,In_46);
and U396 (N_396,In_181,In_1);
and U397 (N_397,In_175,In_447);
nor U398 (N_398,In_326,In_390);
nand U399 (N_399,In_460,In_338);
nor U400 (N_400,In_351,In_199);
or U401 (N_401,In_80,In_425);
and U402 (N_402,In_5,In_177);
or U403 (N_403,In_428,In_400);
nand U404 (N_404,In_100,In_184);
or U405 (N_405,In_322,In_453);
and U406 (N_406,In_435,In_243);
xor U407 (N_407,In_383,In_328);
nand U408 (N_408,In_162,In_394);
and U409 (N_409,In_493,In_210);
nor U410 (N_410,In_238,In_170);
and U411 (N_411,In_206,In_276);
or U412 (N_412,In_209,In_121);
nand U413 (N_413,In_158,In_355);
nand U414 (N_414,In_341,In_394);
nand U415 (N_415,In_358,In_287);
or U416 (N_416,In_257,In_265);
nor U417 (N_417,In_150,In_369);
or U418 (N_418,In_451,In_336);
or U419 (N_419,In_472,In_5);
or U420 (N_420,In_156,In_469);
nor U421 (N_421,In_258,In_169);
or U422 (N_422,In_162,In_495);
nor U423 (N_423,In_473,In_329);
xnor U424 (N_424,In_474,In_40);
nand U425 (N_425,In_393,In_394);
and U426 (N_426,In_399,In_345);
and U427 (N_427,In_146,In_178);
or U428 (N_428,In_299,In_294);
and U429 (N_429,In_395,In_262);
or U430 (N_430,In_82,In_170);
nand U431 (N_431,In_168,In_405);
or U432 (N_432,In_329,In_52);
nand U433 (N_433,In_233,In_179);
and U434 (N_434,In_1,In_15);
nand U435 (N_435,In_492,In_438);
or U436 (N_436,In_62,In_194);
nand U437 (N_437,In_472,In_436);
and U438 (N_438,In_424,In_37);
and U439 (N_439,In_109,In_476);
or U440 (N_440,In_170,In_249);
xor U441 (N_441,In_294,In_88);
nor U442 (N_442,In_303,In_496);
nand U443 (N_443,In_367,In_312);
or U444 (N_444,In_379,In_218);
and U445 (N_445,In_350,In_102);
xor U446 (N_446,In_392,In_149);
nand U447 (N_447,In_390,In_445);
nor U448 (N_448,In_120,In_279);
and U449 (N_449,In_24,In_396);
nor U450 (N_450,In_352,In_40);
and U451 (N_451,In_321,In_456);
and U452 (N_452,In_478,In_298);
nand U453 (N_453,In_189,In_277);
and U454 (N_454,In_47,In_150);
nand U455 (N_455,In_124,In_301);
or U456 (N_456,In_239,In_154);
or U457 (N_457,In_22,In_62);
or U458 (N_458,In_8,In_376);
or U459 (N_459,In_225,In_469);
and U460 (N_460,In_101,In_323);
nor U461 (N_461,In_446,In_434);
nand U462 (N_462,In_16,In_68);
or U463 (N_463,In_490,In_128);
or U464 (N_464,In_364,In_71);
nand U465 (N_465,In_412,In_417);
nand U466 (N_466,In_263,In_462);
and U467 (N_467,In_304,In_248);
and U468 (N_468,In_418,In_188);
or U469 (N_469,In_207,In_128);
nor U470 (N_470,In_159,In_407);
nor U471 (N_471,In_10,In_463);
or U472 (N_472,In_306,In_178);
or U473 (N_473,In_189,In_357);
or U474 (N_474,In_278,In_67);
nand U475 (N_475,In_48,In_212);
or U476 (N_476,In_140,In_474);
or U477 (N_477,In_487,In_54);
or U478 (N_478,In_190,In_111);
and U479 (N_479,In_229,In_0);
nor U480 (N_480,In_129,In_411);
nand U481 (N_481,In_387,In_168);
nor U482 (N_482,In_279,In_322);
nand U483 (N_483,In_303,In_297);
or U484 (N_484,In_351,In_204);
and U485 (N_485,In_362,In_368);
or U486 (N_486,In_167,In_350);
or U487 (N_487,In_217,In_498);
or U488 (N_488,In_127,In_25);
xnor U489 (N_489,In_71,In_447);
and U490 (N_490,In_126,In_49);
nand U491 (N_491,In_13,In_414);
and U492 (N_492,In_345,In_66);
and U493 (N_493,In_14,In_46);
or U494 (N_494,In_440,In_292);
nor U495 (N_495,In_468,In_242);
and U496 (N_496,In_11,In_338);
or U497 (N_497,In_7,In_48);
and U498 (N_498,In_328,In_219);
and U499 (N_499,In_39,In_211);
and U500 (N_500,In_200,In_21);
and U501 (N_501,In_235,In_44);
nand U502 (N_502,In_243,In_416);
nand U503 (N_503,In_271,In_372);
or U504 (N_504,In_410,In_102);
nor U505 (N_505,In_177,In_319);
xor U506 (N_506,In_110,In_476);
nand U507 (N_507,In_313,In_372);
nand U508 (N_508,In_315,In_17);
nand U509 (N_509,In_143,In_470);
or U510 (N_510,In_443,In_42);
nor U511 (N_511,In_345,In_258);
nand U512 (N_512,In_12,In_269);
or U513 (N_513,In_423,In_369);
nand U514 (N_514,In_210,In_388);
nand U515 (N_515,In_0,In_221);
nand U516 (N_516,In_294,In_249);
nor U517 (N_517,In_195,In_208);
or U518 (N_518,In_127,In_440);
and U519 (N_519,In_169,In_385);
nor U520 (N_520,In_87,In_303);
or U521 (N_521,In_336,In_52);
nor U522 (N_522,In_232,In_235);
nand U523 (N_523,In_53,In_90);
nor U524 (N_524,In_343,In_231);
or U525 (N_525,In_375,In_135);
or U526 (N_526,In_248,In_494);
and U527 (N_527,In_18,In_0);
nor U528 (N_528,In_153,In_371);
nand U529 (N_529,In_437,In_471);
xor U530 (N_530,In_182,In_384);
nor U531 (N_531,In_478,In_428);
nand U532 (N_532,In_92,In_34);
nand U533 (N_533,In_231,In_97);
nand U534 (N_534,In_6,In_439);
nand U535 (N_535,In_205,In_253);
nor U536 (N_536,In_26,In_119);
and U537 (N_537,In_143,In_397);
or U538 (N_538,In_308,In_321);
nand U539 (N_539,In_335,In_467);
and U540 (N_540,In_248,In_232);
nor U541 (N_541,In_497,In_106);
or U542 (N_542,In_99,In_179);
and U543 (N_543,In_110,In_190);
and U544 (N_544,In_373,In_309);
or U545 (N_545,In_413,In_340);
and U546 (N_546,In_386,In_233);
xnor U547 (N_547,In_439,In_307);
or U548 (N_548,In_9,In_119);
nor U549 (N_549,In_331,In_15);
and U550 (N_550,In_478,In_121);
nand U551 (N_551,In_341,In_9);
nor U552 (N_552,In_345,In_189);
or U553 (N_553,In_204,In_239);
or U554 (N_554,In_282,In_493);
and U555 (N_555,In_482,In_421);
nor U556 (N_556,In_213,In_94);
nand U557 (N_557,In_104,In_41);
nand U558 (N_558,In_11,In_266);
nand U559 (N_559,In_12,In_106);
nand U560 (N_560,In_209,In_479);
nand U561 (N_561,In_15,In_386);
and U562 (N_562,In_315,In_207);
or U563 (N_563,In_77,In_369);
and U564 (N_564,In_361,In_388);
or U565 (N_565,In_243,In_246);
nand U566 (N_566,In_263,In_332);
and U567 (N_567,In_44,In_303);
or U568 (N_568,In_103,In_267);
nor U569 (N_569,In_342,In_278);
nand U570 (N_570,In_142,In_53);
nand U571 (N_571,In_391,In_54);
nor U572 (N_572,In_116,In_240);
or U573 (N_573,In_438,In_434);
and U574 (N_574,In_66,In_79);
xnor U575 (N_575,In_204,In_426);
or U576 (N_576,In_225,In_125);
nor U577 (N_577,In_216,In_109);
nor U578 (N_578,In_201,In_492);
or U579 (N_579,In_450,In_4);
and U580 (N_580,In_319,In_439);
nor U581 (N_581,In_109,In_346);
nor U582 (N_582,In_150,In_33);
and U583 (N_583,In_51,In_309);
and U584 (N_584,In_247,In_66);
nor U585 (N_585,In_179,In_261);
nor U586 (N_586,In_278,In_417);
or U587 (N_587,In_274,In_96);
or U588 (N_588,In_454,In_279);
or U589 (N_589,In_79,In_142);
or U590 (N_590,In_3,In_300);
nor U591 (N_591,In_471,In_195);
or U592 (N_592,In_249,In_413);
nor U593 (N_593,In_131,In_98);
nor U594 (N_594,In_110,In_131);
and U595 (N_595,In_498,In_443);
nor U596 (N_596,In_166,In_388);
nand U597 (N_597,In_282,In_445);
or U598 (N_598,In_162,In_396);
xor U599 (N_599,In_319,In_401);
or U600 (N_600,In_334,In_398);
nand U601 (N_601,In_205,In_383);
nor U602 (N_602,In_163,In_481);
or U603 (N_603,In_234,In_142);
or U604 (N_604,In_55,In_40);
and U605 (N_605,In_171,In_237);
or U606 (N_606,In_459,In_499);
or U607 (N_607,In_367,In_327);
or U608 (N_608,In_33,In_496);
or U609 (N_609,In_225,In_27);
nand U610 (N_610,In_24,In_455);
and U611 (N_611,In_393,In_338);
nor U612 (N_612,In_22,In_234);
nand U613 (N_613,In_179,In_81);
nand U614 (N_614,In_275,In_199);
and U615 (N_615,In_270,In_275);
and U616 (N_616,In_312,In_88);
nor U617 (N_617,In_344,In_269);
nand U618 (N_618,In_365,In_209);
or U619 (N_619,In_239,In_368);
and U620 (N_620,In_362,In_431);
nand U621 (N_621,In_227,In_180);
nand U622 (N_622,In_288,In_80);
nand U623 (N_623,In_118,In_200);
nand U624 (N_624,In_106,In_137);
nor U625 (N_625,In_298,In_3);
and U626 (N_626,In_493,In_235);
or U627 (N_627,In_122,In_91);
and U628 (N_628,In_478,In_24);
or U629 (N_629,In_356,In_252);
and U630 (N_630,In_192,In_478);
and U631 (N_631,In_183,In_184);
nor U632 (N_632,In_416,In_201);
or U633 (N_633,In_472,In_322);
or U634 (N_634,In_198,In_209);
nor U635 (N_635,In_188,In_26);
or U636 (N_636,In_368,In_241);
or U637 (N_637,In_282,In_218);
and U638 (N_638,In_61,In_475);
nor U639 (N_639,In_435,In_127);
nand U640 (N_640,In_463,In_303);
or U641 (N_641,In_425,In_491);
nor U642 (N_642,In_171,In_495);
and U643 (N_643,In_313,In_222);
and U644 (N_644,In_180,In_445);
nand U645 (N_645,In_125,In_460);
or U646 (N_646,In_274,In_452);
and U647 (N_647,In_469,In_214);
and U648 (N_648,In_420,In_5);
nand U649 (N_649,In_91,In_472);
or U650 (N_650,In_174,In_394);
nand U651 (N_651,In_110,In_209);
and U652 (N_652,In_140,In_403);
nand U653 (N_653,In_55,In_219);
and U654 (N_654,In_439,In_427);
nor U655 (N_655,In_325,In_201);
or U656 (N_656,In_113,In_132);
nand U657 (N_657,In_179,In_368);
nor U658 (N_658,In_149,In_402);
nand U659 (N_659,In_33,In_395);
nor U660 (N_660,In_59,In_208);
and U661 (N_661,In_95,In_443);
nand U662 (N_662,In_316,In_351);
or U663 (N_663,In_1,In_275);
nor U664 (N_664,In_25,In_472);
nand U665 (N_665,In_20,In_388);
or U666 (N_666,In_328,In_411);
and U667 (N_667,In_119,In_397);
nor U668 (N_668,In_101,In_183);
nand U669 (N_669,In_149,In_147);
nor U670 (N_670,In_356,In_376);
or U671 (N_671,In_478,In_350);
nor U672 (N_672,In_316,In_123);
and U673 (N_673,In_166,In_120);
nor U674 (N_674,In_9,In_173);
nor U675 (N_675,In_223,In_47);
nand U676 (N_676,In_347,In_320);
nor U677 (N_677,In_91,In_65);
nand U678 (N_678,In_249,In_27);
or U679 (N_679,In_454,In_287);
nand U680 (N_680,In_296,In_119);
nand U681 (N_681,In_242,In_50);
and U682 (N_682,In_165,In_63);
or U683 (N_683,In_425,In_471);
and U684 (N_684,In_477,In_114);
nand U685 (N_685,In_123,In_208);
nor U686 (N_686,In_221,In_25);
and U687 (N_687,In_116,In_291);
and U688 (N_688,In_128,In_109);
nor U689 (N_689,In_493,In_37);
and U690 (N_690,In_260,In_151);
and U691 (N_691,In_199,In_363);
and U692 (N_692,In_20,In_342);
or U693 (N_693,In_156,In_414);
nand U694 (N_694,In_337,In_173);
nor U695 (N_695,In_99,In_402);
nor U696 (N_696,In_388,In_493);
and U697 (N_697,In_428,In_87);
nor U698 (N_698,In_177,In_61);
nand U699 (N_699,In_169,In_243);
and U700 (N_700,In_244,In_367);
or U701 (N_701,In_478,In_169);
and U702 (N_702,In_205,In_73);
or U703 (N_703,In_250,In_381);
nand U704 (N_704,In_427,In_113);
nand U705 (N_705,In_445,In_399);
and U706 (N_706,In_86,In_139);
nand U707 (N_707,In_414,In_75);
or U708 (N_708,In_57,In_214);
nor U709 (N_709,In_225,In_11);
nand U710 (N_710,In_53,In_215);
or U711 (N_711,In_48,In_443);
nand U712 (N_712,In_50,In_74);
or U713 (N_713,In_282,In_456);
nor U714 (N_714,In_208,In_20);
nand U715 (N_715,In_91,In_66);
and U716 (N_716,In_349,In_460);
nand U717 (N_717,In_351,In_237);
nor U718 (N_718,In_200,In_179);
or U719 (N_719,In_232,In_200);
nand U720 (N_720,In_328,In_47);
or U721 (N_721,In_374,In_184);
and U722 (N_722,In_402,In_50);
and U723 (N_723,In_382,In_16);
and U724 (N_724,In_246,In_156);
or U725 (N_725,In_242,In_207);
and U726 (N_726,In_395,In_482);
xnor U727 (N_727,In_75,In_403);
nand U728 (N_728,In_451,In_265);
or U729 (N_729,In_170,In_340);
or U730 (N_730,In_52,In_231);
or U731 (N_731,In_100,In_148);
or U732 (N_732,In_150,In_149);
and U733 (N_733,In_370,In_492);
and U734 (N_734,In_443,In_316);
and U735 (N_735,In_323,In_236);
nand U736 (N_736,In_257,In_393);
or U737 (N_737,In_248,In_108);
nand U738 (N_738,In_426,In_272);
nand U739 (N_739,In_331,In_12);
nor U740 (N_740,In_283,In_57);
nor U741 (N_741,In_196,In_486);
and U742 (N_742,In_428,In_256);
nor U743 (N_743,In_213,In_135);
and U744 (N_744,In_116,In_90);
or U745 (N_745,In_19,In_270);
and U746 (N_746,In_128,In_2);
nor U747 (N_747,In_277,In_95);
nor U748 (N_748,In_497,In_335);
and U749 (N_749,In_263,In_215);
and U750 (N_750,In_284,In_193);
nand U751 (N_751,In_452,In_407);
nand U752 (N_752,In_169,In_259);
nor U753 (N_753,In_371,In_60);
or U754 (N_754,In_105,In_256);
nand U755 (N_755,In_396,In_156);
xor U756 (N_756,In_159,In_417);
or U757 (N_757,In_307,In_167);
nor U758 (N_758,In_91,In_6);
nor U759 (N_759,In_249,In_162);
and U760 (N_760,In_490,In_307);
nor U761 (N_761,In_418,In_164);
nor U762 (N_762,In_284,In_221);
or U763 (N_763,In_61,In_272);
and U764 (N_764,In_88,In_216);
nand U765 (N_765,In_492,In_331);
or U766 (N_766,In_466,In_344);
nor U767 (N_767,In_423,In_169);
or U768 (N_768,In_423,In_315);
and U769 (N_769,In_404,In_407);
nor U770 (N_770,In_63,In_483);
nor U771 (N_771,In_141,In_261);
nand U772 (N_772,In_214,In_479);
and U773 (N_773,In_22,In_425);
nor U774 (N_774,In_372,In_311);
nand U775 (N_775,In_267,In_131);
nor U776 (N_776,In_351,In_56);
and U777 (N_777,In_222,In_377);
or U778 (N_778,In_250,In_201);
nor U779 (N_779,In_368,In_198);
and U780 (N_780,In_366,In_464);
nor U781 (N_781,In_239,In_186);
and U782 (N_782,In_185,In_382);
xor U783 (N_783,In_229,In_47);
or U784 (N_784,In_282,In_307);
nor U785 (N_785,In_239,In_196);
and U786 (N_786,In_427,In_127);
nand U787 (N_787,In_115,In_292);
nand U788 (N_788,In_324,In_442);
and U789 (N_789,In_201,In_388);
nor U790 (N_790,In_485,In_52);
or U791 (N_791,In_75,In_232);
or U792 (N_792,In_404,In_116);
and U793 (N_793,In_131,In_203);
and U794 (N_794,In_436,In_20);
or U795 (N_795,In_141,In_221);
nor U796 (N_796,In_9,In_298);
nand U797 (N_797,In_355,In_188);
nor U798 (N_798,In_333,In_486);
and U799 (N_799,In_189,In_71);
or U800 (N_800,In_392,In_400);
nor U801 (N_801,In_429,In_10);
or U802 (N_802,In_26,In_156);
nand U803 (N_803,In_481,In_492);
nor U804 (N_804,In_217,In_129);
nor U805 (N_805,In_207,In_311);
nand U806 (N_806,In_56,In_477);
and U807 (N_807,In_256,In_197);
nand U808 (N_808,In_469,In_370);
or U809 (N_809,In_450,In_86);
or U810 (N_810,In_311,In_453);
or U811 (N_811,In_392,In_254);
or U812 (N_812,In_50,In_380);
nor U813 (N_813,In_153,In_341);
and U814 (N_814,In_199,In_198);
nor U815 (N_815,In_463,In_230);
and U816 (N_816,In_133,In_83);
nor U817 (N_817,In_125,In_39);
nand U818 (N_818,In_332,In_102);
and U819 (N_819,In_310,In_157);
nand U820 (N_820,In_257,In_97);
nor U821 (N_821,In_81,In_498);
and U822 (N_822,In_104,In_270);
nand U823 (N_823,In_263,In_367);
nor U824 (N_824,In_288,In_436);
xor U825 (N_825,In_32,In_307);
nand U826 (N_826,In_233,In_171);
nor U827 (N_827,In_459,In_216);
and U828 (N_828,In_390,In_275);
nand U829 (N_829,In_383,In_294);
or U830 (N_830,In_6,In_40);
or U831 (N_831,In_178,In_276);
nand U832 (N_832,In_84,In_225);
and U833 (N_833,In_415,In_116);
nand U834 (N_834,In_446,In_271);
and U835 (N_835,In_284,In_273);
and U836 (N_836,In_316,In_147);
nor U837 (N_837,In_223,In_99);
or U838 (N_838,In_298,In_390);
or U839 (N_839,In_157,In_371);
nand U840 (N_840,In_190,In_131);
nor U841 (N_841,In_185,In_120);
or U842 (N_842,In_203,In_118);
nand U843 (N_843,In_287,In_109);
nand U844 (N_844,In_440,In_272);
or U845 (N_845,In_290,In_395);
and U846 (N_846,In_116,In_247);
nand U847 (N_847,In_56,In_154);
or U848 (N_848,In_213,In_332);
nor U849 (N_849,In_160,In_403);
nand U850 (N_850,In_336,In_159);
and U851 (N_851,In_77,In_151);
nor U852 (N_852,In_164,In_44);
nor U853 (N_853,In_150,In_276);
or U854 (N_854,In_201,In_341);
and U855 (N_855,In_385,In_262);
nor U856 (N_856,In_248,In_185);
or U857 (N_857,In_290,In_77);
or U858 (N_858,In_269,In_373);
and U859 (N_859,In_210,In_399);
and U860 (N_860,In_494,In_451);
nor U861 (N_861,In_404,In_95);
and U862 (N_862,In_6,In_94);
xnor U863 (N_863,In_380,In_140);
nand U864 (N_864,In_269,In_496);
or U865 (N_865,In_347,In_465);
and U866 (N_866,In_174,In_378);
nor U867 (N_867,In_224,In_350);
nand U868 (N_868,In_62,In_364);
nand U869 (N_869,In_279,In_476);
nand U870 (N_870,In_138,In_70);
or U871 (N_871,In_244,In_51);
or U872 (N_872,In_257,In_480);
nor U873 (N_873,In_87,In_172);
nor U874 (N_874,In_215,In_448);
nand U875 (N_875,In_72,In_176);
xnor U876 (N_876,In_368,In_277);
and U877 (N_877,In_458,In_55);
nand U878 (N_878,In_274,In_286);
or U879 (N_879,In_263,In_239);
nand U880 (N_880,In_329,In_494);
or U881 (N_881,In_311,In_274);
and U882 (N_882,In_279,In_137);
and U883 (N_883,In_110,In_177);
nor U884 (N_884,In_107,In_203);
and U885 (N_885,In_442,In_92);
nor U886 (N_886,In_417,In_195);
nand U887 (N_887,In_334,In_417);
nor U888 (N_888,In_405,In_448);
xnor U889 (N_889,In_49,In_421);
nand U890 (N_890,In_379,In_289);
or U891 (N_891,In_433,In_381);
nand U892 (N_892,In_172,In_71);
nand U893 (N_893,In_46,In_227);
nor U894 (N_894,In_154,In_355);
or U895 (N_895,In_407,In_310);
nor U896 (N_896,In_94,In_375);
nor U897 (N_897,In_395,In_492);
nor U898 (N_898,In_333,In_367);
nand U899 (N_899,In_140,In_325);
nand U900 (N_900,In_72,In_393);
nand U901 (N_901,In_256,In_458);
and U902 (N_902,In_334,In_102);
nor U903 (N_903,In_376,In_422);
nor U904 (N_904,In_98,In_422);
or U905 (N_905,In_118,In_77);
and U906 (N_906,In_456,In_85);
and U907 (N_907,In_96,In_395);
nor U908 (N_908,In_190,In_380);
or U909 (N_909,In_269,In_194);
nor U910 (N_910,In_437,In_207);
and U911 (N_911,In_414,In_242);
nor U912 (N_912,In_208,In_143);
nor U913 (N_913,In_439,In_116);
nand U914 (N_914,In_370,In_437);
or U915 (N_915,In_282,In_361);
or U916 (N_916,In_81,In_359);
and U917 (N_917,In_273,In_245);
xnor U918 (N_918,In_84,In_277);
xor U919 (N_919,In_398,In_484);
and U920 (N_920,In_118,In_479);
or U921 (N_921,In_223,In_30);
or U922 (N_922,In_171,In_281);
and U923 (N_923,In_115,In_259);
nor U924 (N_924,In_250,In_133);
or U925 (N_925,In_210,In_127);
nor U926 (N_926,In_20,In_183);
and U927 (N_927,In_98,In_319);
and U928 (N_928,In_330,In_154);
and U929 (N_929,In_128,In_208);
nor U930 (N_930,In_323,In_283);
or U931 (N_931,In_258,In_18);
nand U932 (N_932,In_456,In_382);
nand U933 (N_933,In_425,In_132);
or U934 (N_934,In_260,In_75);
nand U935 (N_935,In_394,In_469);
and U936 (N_936,In_234,In_112);
nor U937 (N_937,In_171,In_63);
nand U938 (N_938,In_151,In_329);
or U939 (N_939,In_20,In_493);
or U940 (N_940,In_308,In_287);
nor U941 (N_941,In_474,In_360);
nand U942 (N_942,In_456,In_262);
and U943 (N_943,In_483,In_219);
or U944 (N_944,In_149,In_450);
nor U945 (N_945,In_207,In_276);
nand U946 (N_946,In_70,In_345);
or U947 (N_947,In_146,In_250);
nand U948 (N_948,In_426,In_318);
nor U949 (N_949,In_19,In_466);
and U950 (N_950,In_412,In_419);
nand U951 (N_951,In_74,In_288);
nand U952 (N_952,In_185,In_17);
nand U953 (N_953,In_461,In_466);
nor U954 (N_954,In_363,In_175);
or U955 (N_955,In_132,In_458);
nand U956 (N_956,In_174,In_206);
nand U957 (N_957,In_55,In_110);
or U958 (N_958,In_261,In_64);
nor U959 (N_959,In_343,In_405);
and U960 (N_960,In_168,In_302);
nand U961 (N_961,In_171,In_496);
nand U962 (N_962,In_232,In_24);
and U963 (N_963,In_233,In_1);
nand U964 (N_964,In_377,In_66);
xor U965 (N_965,In_432,In_359);
nand U966 (N_966,In_337,In_395);
nor U967 (N_967,In_309,In_54);
and U968 (N_968,In_101,In_400);
nand U969 (N_969,In_304,In_449);
and U970 (N_970,In_337,In_416);
nand U971 (N_971,In_154,In_404);
nand U972 (N_972,In_124,In_416);
or U973 (N_973,In_320,In_408);
nand U974 (N_974,In_373,In_442);
nand U975 (N_975,In_87,In_402);
and U976 (N_976,In_305,In_178);
or U977 (N_977,In_104,In_9);
nor U978 (N_978,In_363,In_125);
nand U979 (N_979,In_244,In_125);
xnor U980 (N_980,In_397,In_268);
nand U981 (N_981,In_413,In_198);
xor U982 (N_982,In_150,In_200);
nand U983 (N_983,In_187,In_160);
nand U984 (N_984,In_1,In_103);
nand U985 (N_985,In_223,In_373);
nor U986 (N_986,In_310,In_371);
nor U987 (N_987,In_191,In_60);
and U988 (N_988,In_168,In_20);
or U989 (N_989,In_416,In_24);
or U990 (N_990,In_492,In_214);
and U991 (N_991,In_186,In_12);
and U992 (N_992,In_252,In_257);
nor U993 (N_993,In_482,In_282);
nand U994 (N_994,In_360,In_421);
or U995 (N_995,In_483,In_273);
or U996 (N_996,In_433,In_271);
and U997 (N_997,In_234,In_154);
or U998 (N_998,In_356,In_408);
and U999 (N_999,In_190,In_117);
nand U1000 (N_1000,N_834,N_742);
or U1001 (N_1001,N_387,N_660);
and U1002 (N_1002,N_167,N_195);
nand U1003 (N_1003,N_526,N_373);
nand U1004 (N_1004,N_412,N_897);
and U1005 (N_1005,N_44,N_908);
or U1006 (N_1006,N_108,N_497);
nor U1007 (N_1007,N_164,N_629);
and U1008 (N_1008,N_615,N_792);
and U1009 (N_1009,N_348,N_93);
and U1010 (N_1010,N_817,N_544);
and U1011 (N_1011,N_643,N_559);
and U1012 (N_1012,N_881,N_621);
nand U1013 (N_1013,N_449,N_860);
nand U1014 (N_1014,N_966,N_504);
or U1015 (N_1015,N_435,N_539);
nand U1016 (N_1016,N_40,N_852);
or U1017 (N_1017,N_177,N_809);
nor U1018 (N_1018,N_142,N_13);
nor U1019 (N_1019,N_196,N_406);
nand U1020 (N_1020,N_439,N_148);
or U1021 (N_1021,N_851,N_156);
nor U1022 (N_1022,N_998,N_807);
nor U1023 (N_1023,N_285,N_224);
nand U1024 (N_1024,N_231,N_457);
nand U1025 (N_1025,N_268,N_941);
and U1026 (N_1026,N_447,N_181);
or U1027 (N_1027,N_855,N_613);
or U1028 (N_1028,N_124,N_172);
or U1029 (N_1029,N_70,N_741);
or U1030 (N_1030,N_498,N_996);
nand U1031 (N_1031,N_596,N_991);
and U1032 (N_1032,N_135,N_915);
nor U1033 (N_1033,N_843,N_485);
nor U1034 (N_1034,N_714,N_434);
nor U1035 (N_1035,N_948,N_607);
nand U1036 (N_1036,N_975,N_969);
nand U1037 (N_1037,N_598,N_747);
nor U1038 (N_1038,N_116,N_475);
and U1039 (N_1039,N_166,N_17);
and U1040 (N_1040,N_756,N_345);
nor U1041 (N_1041,N_674,N_324);
nor U1042 (N_1042,N_865,N_540);
or U1043 (N_1043,N_317,N_654);
xor U1044 (N_1044,N_191,N_401);
and U1045 (N_1045,N_242,N_913);
or U1046 (N_1046,N_678,N_636);
xor U1047 (N_1047,N_986,N_637);
nor U1048 (N_1048,N_105,N_237);
and U1049 (N_1049,N_858,N_154);
and U1050 (N_1050,N_123,N_14);
and U1051 (N_1051,N_261,N_735);
and U1052 (N_1052,N_152,N_985);
nor U1053 (N_1053,N_66,N_980);
or U1054 (N_1054,N_733,N_689);
nor U1055 (N_1055,N_266,N_850);
nand U1056 (N_1056,N_194,N_667);
nand U1057 (N_1057,N_787,N_63);
or U1058 (N_1058,N_483,N_983);
or U1059 (N_1059,N_472,N_369);
nor U1060 (N_1060,N_833,N_803);
nor U1061 (N_1061,N_724,N_647);
nor U1062 (N_1062,N_357,N_698);
nand U1063 (N_1063,N_665,N_290);
nand U1064 (N_1064,N_664,N_928);
or U1065 (N_1065,N_604,N_397);
nor U1066 (N_1066,N_750,N_147);
and U1067 (N_1067,N_22,N_137);
and U1068 (N_1068,N_879,N_611);
and U1069 (N_1069,N_829,N_994);
or U1070 (N_1070,N_512,N_549);
nor U1071 (N_1071,N_715,N_326);
nand U1072 (N_1072,N_86,N_593);
nor U1073 (N_1073,N_443,N_788);
xnor U1074 (N_1074,N_107,N_849);
and U1075 (N_1075,N_28,N_46);
and U1076 (N_1076,N_377,N_354);
nand U1077 (N_1077,N_269,N_918);
nor U1078 (N_1078,N_365,N_20);
and U1079 (N_1079,N_130,N_478);
nor U1080 (N_1080,N_917,N_565);
and U1081 (N_1081,N_911,N_694);
or U1082 (N_1082,N_458,N_537);
nand U1083 (N_1083,N_572,N_614);
nor U1084 (N_1084,N_276,N_819);
nor U1085 (N_1085,N_892,N_555);
or U1086 (N_1086,N_704,N_119);
nor U1087 (N_1087,N_836,N_902);
or U1088 (N_1088,N_837,N_853);
nor U1089 (N_1089,N_518,N_620);
or U1090 (N_1090,N_971,N_525);
and U1091 (N_1091,N_366,N_600);
and U1092 (N_1092,N_721,N_372);
nand U1093 (N_1093,N_554,N_486);
nand U1094 (N_1094,N_198,N_552);
nor U1095 (N_1095,N_474,N_146);
or U1096 (N_1096,N_36,N_205);
xor U1097 (N_1097,N_482,N_591);
or U1098 (N_1098,N_15,N_779);
nor U1099 (N_1099,N_305,N_333);
nor U1100 (N_1100,N_690,N_592);
and U1101 (N_1101,N_81,N_111);
and U1102 (N_1102,N_679,N_249);
and U1103 (N_1103,N_113,N_220);
nand U1104 (N_1104,N_736,N_876);
nor U1105 (N_1105,N_255,N_293);
nand U1106 (N_1106,N_404,N_649);
or U1107 (N_1107,N_529,N_362);
nor U1108 (N_1108,N_956,N_110);
nand U1109 (N_1109,N_306,N_327);
and U1110 (N_1110,N_386,N_687);
or U1111 (N_1111,N_453,N_634);
or U1112 (N_1112,N_120,N_257);
nor U1113 (N_1113,N_244,N_981);
nand U1114 (N_1114,N_589,N_831);
nand U1115 (N_1115,N_378,N_646);
and U1116 (N_1116,N_188,N_605);
nand U1117 (N_1117,N_309,N_153);
nand U1118 (N_1118,N_891,N_511);
nor U1119 (N_1119,N_251,N_612);
nand U1120 (N_1120,N_417,N_184);
and U1121 (N_1121,N_294,N_127);
nor U1122 (N_1122,N_574,N_77);
and U1123 (N_1123,N_631,N_914);
and U1124 (N_1124,N_466,N_661);
nand U1125 (N_1125,N_568,N_382);
nand U1126 (N_1126,N_932,N_3);
and U1127 (N_1127,N_701,N_173);
nor U1128 (N_1128,N_757,N_601);
nor U1129 (N_1129,N_909,N_199);
nand U1130 (N_1130,N_313,N_633);
or U1131 (N_1131,N_463,N_754);
and U1132 (N_1132,N_54,N_502);
nor U1133 (N_1133,N_250,N_946);
nand U1134 (N_1134,N_118,N_424);
and U1135 (N_1135,N_558,N_197);
nand U1136 (N_1136,N_877,N_630);
xnor U1137 (N_1137,N_542,N_955);
nand U1138 (N_1138,N_332,N_616);
nor U1139 (N_1139,N_626,N_639);
or U1140 (N_1140,N_984,N_562);
and U1141 (N_1141,N_346,N_273);
and U1142 (N_1142,N_494,N_95);
nor U1143 (N_1143,N_150,N_812);
nand U1144 (N_1144,N_936,N_274);
nor U1145 (N_1145,N_24,N_784);
or U1146 (N_1146,N_929,N_218);
nor U1147 (N_1147,N_978,N_945);
or U1148 (N_1148,N_61,N_490);
nor U1149 (N_1149,N_210,N_450);
nor U1150 (N_1150,N_997,N_115);
or U1151 (N_1151,N_712,N_872);
or U1152 (N_1152,N_58,N_312);
nor U1153 (N_1153,N_92,N_182);
and U1154 (N_1154,N_193,N_436);
and U1155 (N_1155,N_441,N_260);
and U1156 (N_1156,N_638,N_253);
nor U1157 (N_1157,N_64,N_43);
and U1158 (N_1158,N_433,N_532);
nor U1159 (N_1159,N_726,N_960);
and U1160 (N_1160,N_10,N_295);
nor U1161 (N_1161,N_265,N_376);
and U1162 (N_1162,N_318,N_45);
and U1163 (N_1163,N_597,N_245);
nor U1164 (N_1164,N_533,N_924);
or U1165 (N_1165,N_155,N_781);
and U1166 (N_1166,N_415,N_145);
or U1167 (N_1167,N_780,N_506);
nor U1168 (N_1168,N_297,N_964);
or U1169 (N_1169,N_190,N_6);
nand U1170 (N_1170,N_144,N_768);
nand U1171 (N_1171,N_53,N_323);
and U1172 (N_1172,N_527,N_758);
and U1173 (N_1173,N_947,N_395);
or U1174 (N_1174,N_888,N_514);
and U1175 (N_1175,N_625,N_684);
and U1176 (N_1176,N_753,N_728);
nor U1177 (N_1177,N_185,N_503);
xor U1178 (N_1178,N_931,N_96);
or U1179 (N_1179,N_222,N_692);
nand U1180 (N_1180,N_41,N_666);
or U1181 (N_1181,N_4,N_774);
nor U1182 (N_1182,N_825,N_577);
nor U1183 (N_1183,N_423,N_740);
or U1184 (N_1184,N_229,N_765);
or U1185 (N_1185,N_460,N_1);
or U1186 (N_1186,N_428,N_990);
or U1187 (N_1187,N_448,N_248);
nor U1188 (N_1188,N_99,N_283);
nor U1189 (N_1189,N_921,N_828);
and U1190 (N_1190,N_949,N_430);
or U1191 (N_1191,N_968,N_481);
nand U1192 (N_1192,N_487,N_233);
and U1193 (N_1193,N_800,N_48);
and U1194 (N_1194,N_916,N_886);
nor U1195 (N_1195,N_520,N_353);
and U1196 (N_1196,N_937,N_957);
nand U1197 (N_1197,N_341,N_685);
nor U1198 (N_1198,N_737,N_141);
nand U1199 (N_1199,N_82,N_743);
or U1200 (N_1200,N_303,N_240);
and U1201 (N_1201,N_848,N_839);
and U1202 (N_1202,N_489,N_374);
nand U1203 (N_1203,N_923,N_73);
and U1204 (N_1204,N_717,N_109);
nand U1205 (N_1205,N_920,N_296);
nor U1206 (N_1206,N_659,N_700);
and U1207 (N_1207,N_962,N_223);
or U1208 (N_1208,N_885,N_575);
nor U1209 (N_1209,N_650,N_408);
nor U1210 (N_1210,N_557,N_820);
nor U1211 (N_1211,N_379,N_68);
nor U1212 (N_1212,N_361,N_479);
and U1213 (N_1213,N_356,N_720);
or U1214 (N_1214,N_319,N_965);
and U1215 (N_1215,N_484,N_236);
or U1216 (N_1216,N_579,N_139);
or U1217 (N_1217,N_846,N_31);
and U1218 (N_1218,N_950,N_573);
and U1219 (N_1219,N_183,N_880);
nor U1220 (N_1220,N_103,N_791);
or U1221 (N_1221,N_603,N_873);
nor U1222 (N_1222,N_169,N_322);
nand U1223 (N_1223,N_898,N_777);
xnor U1224 (N_1224,N_651,N_288);
nand U1225 (N_1225,N_627,N_778);
or U1226 (N_1226,N_905,N_904);
or U1227 (N_1227,N_396,N_522);
or U1228 (N_1228,N_360,N_707);
and U1229 (N_1229,N_708,N_286);
and U1230 (N_1230,N_827,N_763);
or U1231 (N_1231,N_783,N_595);
and U1232 (N_1232,N_355,N_927);
nand U1233 (N_1233,N_88,N_462);
nand U1234 (N_1234,N_215,N_519);
xnor U1235 (N_1235,N_775,N_350);
nor U1236 (N_1236,N_782,N_870);
nor U1237 (N_1237,N_940,N_938);
and U1238 (N_1238,N_582,N_821);
or U1239 (N_1239,N_238,N_217);
nand U1240 (N_1240,N_531,N_746);
or U1241 (N_1241,N_822,N_57);
nand U1242 (N_1242,N_953,N_926);
or U1243 (N_1243,N_934,N_392);
or U1244 (N_1244,N_551,N_344);
nor U1245 (N_1245,N_263,N_7);
nand U1246 (N_1246,N_944,N_307);
nor U1247 (N_1247,N_583,N_468);
and U1248 (N_1248,N_213,N_545);
or U1249 (N_1249,N_19,N_202);
or U1250 (N_1250,N_727,N_566);
or U1251 (N_1251,N_586,N_246);
nor U1252 (N_1252,N_959,N_221);
or U1253 (N_1253,N_208,N_799);
nor U1254 (N_1254,N_570,N_102);
or U1255 (N_1255,N_770,N_422);
or U1256 (N_1256,N_806,N_52);
nand U1257 (N_1257,N_939,N_899);
and U1258 (N_1258,N_187,N_561);
and U1259 (N_1259,N_546,N_168);
and U1260 (N_1260,N_25,N_55);
or U1261 (N_1261,N_79,N_162);
and U1262 (N_1262,N_399,N_624);
nand U1263 (N_1263,N_608,N_206);
or U1264 (N_1264,N_919,N_772);
nand U1265 (N_1265,N_342,N_21);
and U1266 (N_1266,N_445,N_710);
nand U1267 (N_1267,N_718,N_830);
nor U1268 (N_1268,N_644,N_764);
nor U1269 (N_1269,N_451,N_730);
nor U1270 (N_1270,N_845,N_992);
or U1271 (N_1271,N_30,N_270);
nor U1272 (N_1272,N_693,N_691);
nor U1273 (N_1273,N_722,N_477);
nor U1274 (N_1274,N_90,N_321);
nor U1275 (N_1275,N_804,N_391);
or U1276 (N_1276,N_869,N_761);
and U1277 (N_1277,N_363,N_907);
nand U1278 (N_1278,N_653,N_427);
nand U1279 (N_1279,N_910,N_211);
and U1280 (N_1280,N_461,N_16);
nor U1281 (N_1281,N_576,N_696);
xor U1282 (N_1282,N_35,N_844);
nor U1283 (N_1283,N_553,N_56);
or U1284 (N_1284,N_227,N_219);
nor U1285 (N_1285,N_330,N_446);
nor U1286 (N_1286,N_706,N_767);
nand U1287 (N_1287,N_200,N_398);
nand U1288 (N_1288,N_226,N_534);
and U1289 (N_1289,N_337,N_509);
or U1290 (N_1290,N_178,N_359);
nand U1291 (N_1291,N_381,N_935);
nand U1292 (N_1292,N_622,N_287);
or U1293 (N_1293,N_982,N_241);
or U1294 (N_1294,N_254,N_411);
or U1295 (N_1295,N_496,N_871);
or U1296 (N_1296,N_138,N_94);
nor U1297 (N_1297,N_671,N_413);
nor U1298 (N_1298,N_74,N_203);
nand U1299 (N_1299,N_835,N_635);
or U1300 (N_1300,N_403,N_49);
and U1301 (N_1301,N_655,N_495);
nand U1302 (N_1302,N_501,N_672);
nand U1303 (N_1303,N_958,N_32);
nor U1304 (N_1304,N_906,N_340);
nand U1305 (N_1305,N_745,N_122);
xor U1306 (N_1306,N_272,N_569);
nand U1307 (N_1307,N_98,N_394);
nor U1308 (N_1308,N_771,N_862);
nand U1309 (N_1309,N_400,N_977);
and U1310 (N_1310,N_65,N_785);
and U1311 (N_1311,N_289,N_517);
or U1312 (N_1312,N_414,N_857);
nor U1313 (N_1313,N_71,N_963);
and U1314 (N_1314,N_69,N_389);
nor U1315 (N_1315,N_328,N_599);
nand U1316 (N_1316,N_874,N_29);
nand U1317 (N_1317,N_838,N_252);
and U1318 (N_1318,N_987,N_314);
and U1319 (N_1319,N_171,N_75);
nand U1320 (N_1320,N_352,N_912);
and U1321 (N_1321,N_731,N_11);
nand U1322 (N_1322,N_160,N_465);
and U1323 (N_1323,N_429,N_39);
nor U1324 (N_1324,N_444,N_349);
nand U1325 (N_1325,N_967,N_158);
and U1326 (N_1326,N_204,N_170);
nand U1327 (N_1327,N_284,N_292);
nand U1328 (N_1328,N_578,N_331);
xnor U1329 (N_1329,N_890,N_640);
nor U1330 (N_1330,N_673,N_87);
nand U1331 (N_1331,N_675,N_723);
or U1332 (N_1332,N_680,N_681);
nand U1333 (N_1333,N_459,N_464);
nand U1334 (N_1334,N_507,N_895);
nor U1335 (N_1335,N_970,N_530);
or U1336 (N_1336,N_278,N_59);
nor U1337 (N_1337,N_480,N_523);
and U1338 (N_1338,N_824,N_2);
nor U1339 (N_1339,N_471,N_100);
and U1340 (N_1340,N_861,N_364);
and U1341 (N_1341,N_62,N_390);
or U1342 (N_1342,N_33,N_709);
or U1343 (N_1343,N_499,N_473);
and U1344 (N_1344,N_662,N_755);
or U1345 (N_1345,N_407,N_329);
or U1346 (N_1346,N_143,N_793);
nand U1347 (N_1347,N_973,N_452);
and U1348 (N_1348,N_856,N_8);
or U1349 (N_1349,N_894,N_409);
or U1350 (N_1350,N_808,N_277);
nor U1351 (N_1351,N_488,N_766);
and U1352 (N_1352,N_47,N_201);
nor U1353 (N_1353,N_797,N_590);
nor U1354 (N_1354,N_121,N_697);
and U1355 (N_1355,N_128,N_311);
nor U1356 (N_1356,N_440,N_711);
and U1357 (N_1357,N_567,N_734);
nand U1358 (N_1358,N_281,N_425);
nand U1359 (N_1359,N_802,N_789);
and U1360 (N_1360,N_393,N_585);
and U1361 (N_1361,N_256,N_581);
or U1362 (N_1362,N_628,N_536);
or U1363 (N_1363,N_882,N_426);
nand U1364 (N_1364,N_420,N_713);
or U1365 (N_1365,N_584,N_505);
and U1366 (N_1366,N_338,N_161);
nand U1367 (N_1367,N_794,N_132);
xor U1368 (N_1368,N_719,N_686);
and U1369 (N_1369,N_149,N_104);
nor U1370 (N_1370,N_903,N_832);
or U1371 (N_1371,N_816,N_887);
nand U1372 (N_1372,N_126,N_974);
nor U1373 (N_1373,N_619,N_541);
and U1374 (N_1374,N_267,N_656);
and U1375 (N_1375,N_275,N_648);
nor U1376 (N_1376,N_469,N_952);
nand U1377 (N_1377,N_900,N_216);
and U1378 (N_1378,N_493,N_840);
nor U1379 (N_1379,N_106,N_34);
nand U1380 (N_1380,N_112,N_370);
nand U1381 (N_1381,N_176,N_602);
nand U1382 (N_1382,N_37,N_842);
nand U1383 (N_1383,N_878,N_528);
and U1384 (N_1384,N_560,N_159);
nor U1385 (N_1385,N_438,N_27);
and U1386 (N_1386,N_491,N_658);
and U1387 (N_1387,N_385,N_470);
nor U1388 (N_1388,N_212,N_405);
nor U1389 (N_1389,N_23,N_232);
or U1390 (N_1390,N_933,N_214);
or U1391 (N_1391,N_308,N_773);
nor U1392 (N_1392,N_535,N_26);
xor U1393 (N_1393,N_186,N_442);
nand U1394 (N_1394,N_988,N_78);
nor U1395 (N_1395,N_699,N_371);
nand U1396 (N_1396,N_418,N_140);
nand U1397 (N_1397,N_677,N_500);
and U1398 (N_1398,N_642,N_606);
nand U1399 (N_1399,N_760,N_85);
or U1400 (N_1400,N_716,N_863);
and U1401 (N_1401,N_60,N_291);
or U1402 (N_1402,N_796,N_437);
nor U1403 (N_1403,N_50,N_347);
and U1404 (N_1404,N_38,N_367);
nor U1405 (N_1405,N_264,N_84);
nor U1406 (N_1406,N_930,N_375);
nor U1407 (N_1407,N_883,N_91);
nand U1408 (N_1408,N_189,N_83);
nand U1409 (N_1409,N_587,N_641);
or U1410 (N_1410,N_165,N_610);
nand U1411 (N_1411,N_618,N_133);
nand U1412 (N_1412,N_645,N_823);
and U1413 (N_1413,N_209,N_688);
or U1414 (N_1414,N_258,N_383);
nand U1415 (N_1415,N_335,N_456);
nor U1416 (N_1416,N_663,N_97);
or U1417 (N_1417,N_492,N_151);
nor U1418 (N_1418,N_368,N_225);
and U1419 (N_1419,N_623,N_0);
or U1420 (N_1420,N_738,N_682);
and U1421 (N_1421,N_790,N_739);
nor U1422 (N_1422,N_744,N_247);
nand U1423 (N_1423,N_669,N_798);
nand U1424 (N_1424,N_163,N_230);
or U1425 (N_1425,N_548,N_652);
and U1426 (N_1426,N_751,N_801);
nand U1427 (N_1427,N_795,N_925);
or U1428 (N_1428,N_814,N_228);
nor U1429 (N_1429,N_513,N_380);
and U1430 (N_1430,N_543,N_703);
nor U1431 (N_1431,N_358,N_732);
or U1432 (N_1432,N_676,N_351);
nand U1433 (N_1433,N_259,N_334);
or U1434 (N_1434,N_125,N_174);
or U1435 (N_1435,N_841,N_759);
nand U1436 (N_1436,N_76,N_826);
and U1437 (N_1437,N_410,N_901);
nor U1438 (N_1438,N_454,N_813);
nor U1439 (N_1439,N_563,N_310);
or U1440 (N_1440,N_609,N_134);
nand U1441 (N_1441,N_301,N_864);
nand U1442 (N_1442,N_657,N_951);
or U1443 (N_1443,N_131,N_776);
and U1444 (N_1444,N_136,N_476);
or U1445 (N_1445,N_416,N_868);
or U1446 (N_1446,N_954,N_67);
or U1447 (N_1447,N_180,N_695);
nand U1448 (N_1448,N_302,N_976);
and U1449 (N_1449,N_325,N_234);
or U1450 (N_1450,N_300,N_538);
nand U1451 (N_1451,N_972,N_875);
and U1452 (N_1452,N_282,N_670);
nor U1453 (N_1453,N_668,N_705);
and U1454 (N_1454,N_725,N_179);
nand U1455 (N_1455,N_979,N_42);
nand U1456 (N_1456,N_889,N_943);
nand U1457 (N_1457,N_298,N_854);
or U1458 (N_1458,N_114,N_243);
and U1459 (N_1459,N_508,N_805);
nand U1460 (N_1460,N_995,N_175);
xnor U1461 (N_1461,N_556,N_455);
nand U1462 (N_1462,N_12,N_942);
and U1463 (N_1463,N_280,N_431);
nand U1464 (N_1464,N_993,N_884);
nand U1465 (N_1465,N_632,N_810);
or U1466 (N_1466,N_524,N_580);
and U1467 (N_1467,N_402,N_683);
nand U1468 (N_1468,N_769,N_550);
nand U1469 (N_1469,N_388,N_101);
and U1470 (N_1470,N_235,N_320);
or U1471 (N_1471,N_547,N_343);
nand U1472 (N_1472,N_588,N_9);
nand U1473 (N_1473,N_157,N_702);
nor U1474 (N_1474,N_896,N_419);
and U1475 (N_1475,N_239,N_515);
xnor U1476 (N_1476,N_594,N_336);
xnor U1477 (N_1477,N_18,N_299);
and U1478 (N_1478,N_818,N_339);
nand U1479 (N_1479,N_207,N_729);
nor U1480 (N_1480,N_316,N_271);
nand U1481 (N_1481,N_859,N_617);
and U1482 (N_1482,N_304,N_421);
nand U1483 (N_1483,N_752,N_80);
and U1484 (N_1484,N_516,N_262);
nand U1485 (N_1485,N_72,N_89);
nand U1486 (N_1486,N_521,N_847);
or U1487 (N_1487,N_192,N_989);
or U1488 (N_1488,N_467,N_279);
and U1489 (N_1489,N_129,N_384);
or U1490 (N_1490,N_749,N_786);
nor U1491 (N_1491,N_748,N_51);
nand U1492 (N_1492,N_867,N_893);
nor U1493 (N_1493,N_999,N_564);
nor U1494 (N_1494,N_5,N_315);
nor U1495 (N_1495,N_815,N_117);
or U1496 (N_1496,N_811,N_571);
or U1497 (N_1497,N_922,N_432);
nand U1498 (N_1498,N_762,N_510);
nor U1499 (N_1499,N_961,N_866);
or U1500 (N_1500,N_329,N_932);
nand U1501 (N_1501,N_167,N_251);
nor U1502 (N_1502,N_63,N_596);
nor U1503 (N_1503,N_397,N_952);
or U1504 (N_1504,N_360,N_879);
nor U1505 (N_1505,N_325,N_913);
nor U1506 (N_1506,N_189,N_944);
xor U1507 (N_1507,N_106,N_524);
and U1508 (N_1508,N_251,N_659);
nor U1509 (N_1509,N_31,N_199);
nor U1510 (N_1510,N_769,N_319);
nand U1511 (N_1511,N_898,N_377);
nor U1512 (N_1512,N_909,N_177);
nand U1513 (N_1513,N_499,N_204);
nand U1514 (N_1514,N_525,N_422);
nand U1515 (N_1515,N_268,N_674);
nor U1516 (N_1516,N_54,N_747);
or U1517 (N_1517,N_650,N_977);
and U1518 (N_1518,N_943,N_249);
and U1519 (N_1519,N_192,N_906);
or U1520 (N_1520,N_478,N_452);
or U1521 (N_1521,N_484,N_359);
or U1522 (N_1522,N_999,N_75);
or U1523 (N_1523,N_126,N_807);
nor U1524 (N_1524,N_147,N_357);
and U1525 (N_1525,N_617,N_789);
nor U1526 (N_1526,N_565,N_798);
or U1527 (N_1527,N_0,N_853);
nand U1528 (N_1528,N_679,N_601);
nand U1529 (N_1529,N_329,N_386);
nor U1530 (N_1530,N_250,N_823);
nand U1531 (N_1531,N_489,N_207);
or U1532 (N_1532,N_521,N_206);
nand U1533 (N_1533,N_533,N_660);
nand U1534 (N_1534,N_372,N_977);
nor U1535 (N_1535,N_768,N_127);
or U1536 (N_1536,N_347,N_141);
nand U1537 (N_1537,N_896,N_238);
or U1538 (N_1538,N_863,N_770);
nand U1539 (N_1539,N_791,N_735);
and U1540 (N_1540,N_701,N_275);
or U1541 (N_1541,N_15,N_976);
nor U1542 (N_1542,N_688,N_744);
nor U1543 (N_1543,N_719,N_42);
nor U1544 (N_1544,N_859,N_240);
and U1545 (N_1545,N_625,N_275);
or U1546 (N_1546,N_281,N_816);
or U1547 (N_1547,N_678,N_837);
nor U1548 (N_1548,N_808,N_195);
nand U1549 (N_1549,N_275,N_744);
nor U1550 (N_1550,N_625,N_678);
nor U1551 (N_1551,N_480,N_300);
nor U1552 (N_1552,N_249,N_693);
nand U1553 (N_1553,N_285,N_696);
nor U1554 (N_1554,N_435,N_63);
and U1555 (N_1555,N_194,N_421);
nor U1556 (N_1556,N_704,N_527);
or U1557 (N_1557,N_5,N_166);
nor U1558 (N_1558,N_496,N_656);
and U1559 (N_1559,N_982,N_980);
xor U1560 (N_1560,N_671,N_660);
or U1561 (N_1561,N_985,N_46);
nand U1562 (N_1562,N_787,N_949);
nor U1563 (N_1563,N_484,N_3);
nor U1564 (N_1564,N_982,N_523);
nor U1565 (N_1565,N_820,N_670);
nand U1566 (N_1566,N_60,N_851);
or U1567 (N_1567,N_282,N_562);
nor U1568 (N_1568,N_644,N_735);
or U1569 (N_1569,N_795,N_542);
nand U1570 (N_1570,N_973,N_464);
nor U1571 (N_1571,N_321,N_492);
nand U1572 (N_1572,N_179,N_163);
and U1573 (N_1573,N_760,N_232);
and U1574 (N_1574,N_670,N_786);
or U1575 (N_1575,N_346,N_96);
and U1576 (N_1576,N_575,N_744);
nor U1577 (N_1577,N_764,N_276);
and U1578 (N_1578,N_517,N_452);
nor U1579 (N_1579,N_131,N_306);
nand U1580 (N_1580,N_574,N_237);
or U1581 (N_1581,N_410,N_594);
and U1582 (N_1582,N_786,N_746);
and U1583 (N_1583,N_826,N_416);
nand U1584 (N_1584,N_377,N_992);
and U1585 (N_1585,N_13,N_23);
xnor U1586 (N_1586,N_920,N_651);
nand U1587 (N_1587,N_468,N_301);
nor U1588 (N_1588,N_619,N_454);
nor U1589 (N_1589,N_316,N_703);
nor U1590 (N_1590,N_545,N_68);
and U1591 (N_1591,N_184,N_257);
and U1592 (N_1592,N_195,N_445);
or U1593 (N_1593,N_965,N_336);
nor U1594 (N_1594,N_25,N_96);
xor U1595 (N_1595,N_123,N_121);
nor U1596 (N_1596,N_814,N_358);
nand U1597 (N_1597,N_243,N_639);
xnor U1598 (N_1598,N_780,N_881);
nand U1599 (N_1599,N_702,N_792);
or U1600 (N_1600,N_915,N_285);
nor U1601 (N_1601,N_747,N_627);
nand U1602 (N_1602,N_399,N_588);
or U1603 (N_1603,N_277,N_853);
nor U1604 (N_1604,N_50,N_830);
nand U1605 (N_1605,N_558,N_883);
nor U1606 (N_1606,N_241,N_78);
nand U1607 (N_1607,N_124,N_251);
and U1608 (N_1608,N_735,N_753);
and U1609 (N_1609,N_871,N_592);
nand U1610 (N_1610,N_485,N_571);
and U1611 (N_1611,N_37,N_44);
or U1612 (N_1612,N_287,N_414);
or U1613 (N_1613,N_26,N_185);
or U1614 (N_1614,N_571,N_502);
nand U1615 (N_1615,N_824,N_799);
nand U1616 (N_1616,N_456,N_703);
and U1617 (N_1617,N_907,N_636);
nor U1618 (N_1618,N_140,N_243);
nand U1619 (N_1619,N_287,N_584);
and U1620 (N_1620,N_585,N_564);
or U1621 (N_1621,N_368,N_815);
or U1622 (N_1622,N_31,N_651);
or U1623 (N_1623,N_473,N_882);
nor U1624 (N_1624,N_694,N_51);
or U1625 (N_1625,N_477,N_139);
and U1626 (N_1626,N_565,N_145);
or U1627 (N_1627,N_923,N_713);
nand U1628 (N_1628,N_153,N_30);
and U1629 (N_1629,N_164,N_96);
and U1630 (N_1630,N_843,N_147);
or U1631 (N_1631,N_441,N_923);
nand U1632 (N_1632,N_74,N_702);
nor U1633 (N_1633,N_141,N_440);
or U1634 (N_1634,N_476,N_43);
and U1635 (N_1635,N_750,N_920);
and U1636 (N_1636,N_877,N_821);
nor U1637 (N_1637,N_821,N_559);
or U1638 (N_1638,N_46,N_121);
and U1639 (N_1639,N_271,N_297);
and U1640 (N_1640,N_537,N_261);
nor U1641 (N_1641,N_104,N_323);
or U1642 (N_1642,N_455,N_667);
and U1643 (N_1643,N_404,N_674);
nor U1644 (N_1644,N_982,N_852);
or U1645 (N_1645,N_884,N_705);
or U1646 (N_1646,N_433,N_353);
nand U1647 (N_1647,N_953,N_332);
nor U1648 (N_1648,N_933,N_382);
and U1649 (N_1649,N_11,N_850);
nor U1650 (N_1650,N_993,N_264);
or U1651 (N_1651,N_522,N_733);
nor U1652 (N_1652,N_846,N_738);
or U1653 (N_1653,N_446,N_401);
and U1654 (N_1654,N_741,N_505);
nor U1655 (N_1655,N_451,N_530);
nand U1656 (N_1656,N_504,N_623);
or U1657 (N_1657,N_228,N_308);
or U1658 (N_1658,N_216,N_297);
and U1659 (N_1659,N_931,N_405);
nor U1660 (N_1660,N_867,N_322);
and U1661 (N_1661,N_251,N_714);
nor U1662 (N_1662,N_352,N_838);
or U1663 (N_1663,N_435,N_336);
nor U1664 (N_1664,N_35,N_89);
or U1665 (N_1665,N_292,N_675);
and U1666 (N_1666,N_280,N_632);
nand U1667 (N_1667,N_153,N_270);
nor U1668 (N_1668,N_999,N_109);
nor U1669 (N_1669,N_84,N_224);
nand U1670 (N_1670,N_330,N_137);
and U1671 (N_1671,N_76,N_630);
nand U1672 (N_1672,N_555,N_900);
or U1673 (N_1673,N_861,N_293);
or U1674 (N_1674,N_621,N_328);
xnor U1675 (N_1675,N_240,N_843);
nand U1676 (N_1676,N_236,N_146);
nand U1677 (N_1677,N_698,N_97);
or U1678 (N_1678,N_137,N_704);
and U1679 (N_1679,N_355,N_334);
and U1680 (N_1680,N_433,N_876);
nand U1681 (N_1681,N_397,N_153);
nand U1682 (N_1682,N_978,N_188);
nand U1683 (N_1683,N_721,N_822);
or U1684 (N_1684,N_627,N_974);
or U1685 (N_1685,N_552,N_900);
nand U1686 (N_1686,N_721,N_498);
nand U1687 (N_1687,N_197,N_758);
nor U1688 (N_1688,N_671,N_451);
and U1689 (N_1689,N_422,N_995);
nor U1690 (N_1690,N_32,N_91);
and U1691 (N_1691,N_765,N_840);
nand U1692 (N_1692,N_909,N_855);
and U1693 (N_1693,N_236,N_715);
nand U1694 (N_1694,N_597,N_236);
or U1695 (N_1695,N_370,N_467);
nand U1696 (N_1696,N_124,N_875);
xnor U1697 (N_1697,N_323,N_568);
nand U1698 (N_1698,N_406,N_127);
and U1699 (N_1699,N_475,N_751);
or U1700 (N_1700,N_658,N_416);
and U1701 (N_1701,N_751,N_827);
and U1702 (N_1702,N_980,N_181);
or U1703 (N_1703,N_890,N_26);
or U1704 (N_1704,N_594,N_821);
nor U1705 (N_1705,N_667,N_419);
and U1706 (N_1706,N_626,N_718);
and U1707 (N_1707,N_230,N_291);
nor U1708 (N_1708,N_55,N_384);
nor U1709 (N_1709,N_451,N_874);
and U1710 (N_1710,N_901,N_374);
or U1711 (N_1711,N_129,N_70);
nand U1712 (N_1712,N_795,N_854);
nor U1713 (N_1713,N_193,N_281);
or U1714 (N_1714,N_152,N_325);
and U1715 (N_1715,N_789,N_350);
nor U1716 (N_1716,N_365,N_720);
or U1717 (N_1717,N_575,N_874);
and U1718 (N_1718,N_982,N_644);
or U1719 (N_1719,N_831,N_638);
and U1720 (N_1720,N_103,N_574);
nor U1721 (N_1721,N_94,N_230);
nand U1722 (N_1722,N_404,N_436);
nand U1723 (N_1723,N_665,N_624);
nor U1724 (N_1724,N_937,N_621);
or U1725 (N_1725,N_72,N_696);
and U1726 (N_1726,N_105,N_478);
and U1727 (N_1727,N_340,N_462);
and U1728 (N_1728,N_273,N_95);
or U1729 (N_1729,N_657,N_662);
or U1730 (N_1730,N_491,N_582);
or U1731 (N_1731,N_409,N_913);
and U1732 (N_1732,N_323,N_765);
nor U1733 (N_1733,N_10,N_535);
xnor U1734 (N_1734,N_564,N_905);
nand U1735 (N_1735,N_628,N_35);
and U1736 (N_1736,N_82,N_756);
and U1737 (N_1737,N_44,N_151);
and U1738 (N_1738,N_341,N_22);
nor U1739 (N_1739,N_165,N_600);
nand U1740 (N_1740,N_632,N_309);
nand U1741 (N_1741,N_635,N_876);
and U1742 (N_1742,N_948,N_940);
nor U1743 (N_1743,N_453,N_841);
or U1744 (N_1744,N_604,N_336);
nor U1745 (N_1745,N_283,N_780);
nand U1746 (N_1746,N_765,N_452);
xor U1747 (N_1747,N_944,N_757);
nand U1748 (N_1748,N_826,N_914);
nor U1749 (N_1749,N_888,N_387);
and U1750 (N_1750,N_290,N_168);
nand U1751 (N_1751,N_330,N_258);
or U1752 (N_1752,N_85,N_808);
xnor U1753 (N_1753,N_107,N_501);
nor U1754 (N_1754,N_677,N_816);
or U1755 (N_1755,N_53,N_507);
or U1756 (N_1756,N_872,N_476);
nand U1757 (N_1757,N_794,N_6);
and U1758 (N_1758,N_761,N_666);
nand U1759 (N_1759,N_78,N_719);
nor U1760 (N_1760,N_856,N_200);
nor U1761 (N_1761,N_88,N_845);
nand U1762 (N_1762,N_318,N_999);
nor U1763 (N_1763,N_398,N_565);
or U1764 (N_1764,N_580,N_555);
or U1765 (N_1765,N_112,N_154);
nand U1766 (N_1766,N_68,N_692);
and U1767 (N_1767,N_677,N_838);
nand U1768 (N_1768,N_150,N_764);
and U1769 (N_1769,N_655,N_720);
and U1770 (N_1770,N_324,N_98);
or U1771 (N_1771,N_546,N_592);
and U1772 (N_1772,N_949,N_578);
or U1773 (N_1773,N_615,N_425);
and U1774 (N_1774,N_934,N_395);
nand U1775 (N_1775,N_480,N_66);
nand U1776 (N_1776,N_290,N_758);
nor U1777 (N_1777,N_699,N_155);
nor U1778 (N_1778,N_401,N_878);
or U1779 (N_1779,N_165,N_0);
nor U1780 (N_1780,N_899,N_76);
or U1781 (N_1781,N_198,N_946);
and U1782 (N_1782,N_423,N_380);
or U1783 (N_1783,N_96,N_274);
and U1784 (N_1784,N_318,N_670);
nand U1785 (N_1785,N_62,N_835);
nor U1786 (N_1786,N_603,N_523);
nand U1787 (N_1787,N_807,N_800);
or U1788 (N_1788,N_30,N_637);
xnor U1789 (N_1789,N_401,N_107);
nand U1790 (N_1790,N_313,N_621);
or U1791 (N_1791,N_573,N_618);
xnor U1792 (N_1792,N_438,N_231);
and U1793 (N_1793,N_61,N_97);
and U1794 (N_1794,N_407,N_31);
nor U1795 (N_1795,N_236,N_40);
or U1796 (N_1796,N_947,N_542);
and U1797 (N_1797,N_491,N_208);
or U1798 (N_1798,N_574,N_540);
or U1799 (N_1799,N_802,N_251);
nand U1800 (N_1800,N_599,N_711);
or U1801 (N_1801,N_874,N_96);
nand U1802 (N_1802,N_821,N_940);
nor U1803 (N_1803,N_543,N_676);
or U1804 (N_1804,N_170,N_579);
nor U1805 (N_1805,N_875,N_485);
nor U1806 (N_1806,N_584,N_830);
or U1807 (N_1807,N_733,N_244);
and U1808 (N_1808,N_522,N_56);
nand U1809 (N_1809,N_219,N_923);
nand U1810 (N_1810,N_784,N_758);
nor U1811 (N_1811,N_423,N_299);
and U1812 (N_1812,N_848,N_203);
nor U1813 (N_1813,N_888,N_622);
or U1814 (N_1814,N_415,N_232);
nor U1815 (N_1815,N_607,N_153);
or U1816 (N_1816,N_392,N_764);
nand U1817 (N_1817,N_1,N_532);
nor U1818 (N_1818,N_373,N_731);
nand U1819 (N_1819,N_175,N_625);
nand U1820 (N_1820,N_44,N_427);
nor U1821 (N_1821,N_692,N_849);
or U1822 (N_1822,N_275,N_349);
nor U1823 (N_1823,N_466,N_294);
and U1824 (N_1824,N_419,N_495);
nor U1825 (N_1825,N_568,N_617);
and U1826 (N_1826,N_332,N_373);
nand U1827 (N_1827,N_675,N_529);
nor U1828 (N_1828,N_302,N_550);
nor U1829 (N_1829,N_573,N_965);
nand U1830 (N_1830,N_412,N_300);
nand U1831 (N_1831,N_498,N_914);
nand U1832 (N_1832,N_99,N_177);
nor U1833 (N_1833,N_907,N_735);
or U1834 (N_1834,N_655,N_588);
and U1835 (N_1835,N_321,N_984);
nand U1836 (N_1836,N_832,N_355);
and U1837 (N_1837,N_404,N_403);
or U1838 (N_1838,N_754,N_309);
and U1839 (N_1839,N_744,N_117);
nand U1840 (N_1840,N_330,N_235);
or U1841 (N_1841,N_576,N_217);
or U1842 (N_1842,N_590,N_392);
and U1843 (N_1843,N_365,N_942);
or U1844 (N_1844,N_44,N_675);
nor U1845 (N_1845,N_761,N_153);
or U1846 (N_1846,N_899,N_133);
nand U1847 (N_1847,N_820,N_666);
xnor U1848 (N_1848,N_502,N_559);
nor U1849 (N_1849,N_995,N_310);
and U1850 (N_1850,N_560,N_591);
xnor U1851 (N_1851,N_404,N_353);
nand U1852 (N_1852,N_946,N_477);
or U1853 (N_1853,N_370,N_67);
or U1854 (N_1854,N_181,N_434);
nand U1855 (N_1855,N_829,N_938);
nor U1856 (N_1856,N_114,N_593);
and U1857 (N_1857,N_44,N_107);
nor U1858 (N_1858,N_43,N_445);
nand U1859 (N_1859,N_436,N_673);
and U1860 (N_1860,N_328,N_805);
and U1861 (N_1861,N_148,N_681);
and U1862 (N_1862,N_331,N_111);
nor U1863 (N_1863,N_165,N_42);
nor U1864 (N_1864,N_591,N_732);
nor U1865 (N_1865,N_248,N_85);
or U1866 (N_1866,N_412,N_282);
nor U1867 (N_1867,N_566,N_449);
or U1868 (N_1868,N_853,N_363);
nand U1869 (N_1869,N_427,N_465);
nor U1870 (N_1870,N_77,N_142);
nand U1871 (N_1871,N_683,N_634);
and U1872 (N_1872,N_417,N_873);
and U1873 (N_1873,N_746,N_27);
nor U1874 (N_1874,N_838,N_980);
or U1875 (N_1875,N_698,N_479);
nor U1876 (N_1876,N_963,N_784);
nor U1877 (N_1877,N_886,N_120);
nand U1878 (N_1878,N_538,N_64);
nor U1879 (N_1879,N_518,N_926);
nor U1880 (N_1880,N_129,N_239);
nor U1881 (N_1881,N_818,N_115);
or U1882 (N_1882,N_137,N_906);
nor U1883 (N_1883,N_750,N_643);
nand U1884 (N_1884,N_201,N_989);
nand U1885 (N_1885,N_751,N_169);
nor U1886 (N_1886,N_637,N_50);
nor U1887 (N_1887,N_935,N_226);
and U1888 (N_1888,N_691,N_927);
or U1889 (N_1889,N_317,N_202);
nor U1890 (N_1890,N_467,N_670);
nand U1891 (N_1891,N_839,N_265);
or U1892 (N_1892,N_508,N_880);
or U1893 (N_1893,N_756,N_747);
nand U1894 (N_1894,N_781,N_837);
nor U1895 (N_1895,N_826,N_180);
nor U1896 (N_1896,N_683,N_799);
nor U1897 (N_1897,N_90,N_373);
nor U1898 (N_1898,N_319,N_730);
or U1899 (N_1899,N_979,N_78);
nand U1900 (N_1900,N_942,N_914);
nand U1901 (N_1901,N_70,N_969);
or U1902 (N_1902,N_411,N_46);
or U1903 (N_1903,N_115,N_397);
nand U1904 (N_1904,N_841,N_967);
nand U1905 (N_1905,N_893,N_413);
or U1906 (N_1906,N_269,N_929);
nor U1907 (N_1907,N_902,N_68);
and U1908 (N_1908,N_978,N_482);
nand U1909 (N_1909,N_854,N_365);
or U1910 (N_1910,N_70,N_650);
or U1911 (N_1911,N_774,N_19);
nand U1912 (N_1912,N_723,N_129);
nand U1913 (N_1913,N_267,N_192);
or U1914 (N_1914,N_746,N_111);
and U1915 (N_1915,N_128,N_143);
and U1916 (N_1916,N_125,N_724);
or U1917 (N_1917,N_594,N_492);
nand U1918 (N_1918,N_640,N_534);
nand U1919 (N_1919,N_314,N_737);
and U1920 (N_1920,N_839,N_287);
nand U1921 (N_1921,N_699,N_529);
nor U1922 (N_1922,N_279,N_448);
nand U1923 (N_1923,N_983,N_818);
nor U1924 (N_1924,N_450,N_49);
or U1925 (N_1925,N_960,N_856);
nand U1926 (N_1926,N_188,N_286);
nor U1927 (N_1927,N_207,N_393);
or U1928 (N_1928,N_247,N_467);
and U1929 (N_1929,N_3,N_302);
or U1930 (N_1930,N_496,N_911);
nand U1931 (N_1931,N_496,N_847);
nor U1932 (N_1932,N_561,N_543);
nand U1933 (N_1933,N_747,N_263);
or U1934 (N_1934,N_648,N_863);
nor U1935 (N_1935,N_530,N_292);
or U1936 (N_1936,N_95,N_475);
nand U1937 (N_1937,N_128,N_505);
xor U1938 (N_1938,N_78,N_819);
and U1939 (N_1939,N_633,N_818);
and U1940 (N_1940,N_433,N_986);
nand U1941 (N_1941,N_370,N_0);
and U1942 (N_1942,N_618,N_859);
or U1943 (N_1943,N_98,N_732);
and U1944 (N_1944,N_922,N_277);
and U1945 (N_1945,N_795,N_152);
and U1946 (N_1946,N_785,N_572);
nand U1947 (N_1947,N_185,N_307);
or U1948 (N_1948,N_890,N_911);
and U1949 (N_1949,N_551,N_918);
nand U1950 (N_1950,N_279,N_229);
nor U1951 (N_1951,N_645,N_678);
nor U1952 (N_1952,N_646,N_398);
nor U1953 (N_1953,N_382,N_288);
or U1954 (N_1954,N_484,N_625);
and U1955 (N_1955,N_675,N_534);
and U1956 (N_1956,N_949,N_600);
and U1957 (N_1957,N_851,N_253);
nand U1958 (N_1958,N_326,N_96);
or U1959 (N_1959,N_274,N_583);
nand U1960 (N_1960,N_264,N_271);
nor U1961 (N_1961,N_3,N_775);
nand U1962 (N_1962,N_164,N_806);
or U1963 (N_1963,N_291,N_670);
nand U1964 (N_1964,N_293,N_169);
or U1965 (N_1965,N_242,N_248);
or U1966 (N_1966,N_809,N_886);
nand U1967 (N_1967,N_373,N_493);
nor U1968 (N_1968,N_311,N_907);
nor U1969 (N_1969,N_705,N_979);
nor U1970 (N_1970,N_305,N_550);
nand U1971 (N_1971,N_755,N_859);
nand U1972 (N_1972,N_874,N_377);
and U1973 (N_1973,N_933,N_556);
or U1974 (N_1974,N_670,N_787);
nand U1975 (N_1975,N_576,N_203);
nand U1976 (N_1976,N_38,N_231);
or U1977 (N_1977,N_768,N_500);
and U1978 (N_1978,N_76,N_907);
nor U1979 (N_1979,N_754,N_921);
and U1980 (N_1980,N_849,N_347);
or U1981 (N_1981,N_309,N_83);
xor U1982 (N_1982,N_385,N_101);
or U1983 (N_1983,N_643,N_261);
and U1984 (N_1984,N_956,N_309);
nor U1985 (N_1985,N_357,N_303);
nand U1986 (N_1986,N_293,N_916);
nor U1987 (N_1987,N_733,N_253);
nor U1988 (N_1988,N_260,N_526);
or U1989 (N_1989,N_102,N_939);
nor U1990 (N_1990,N_559,N_475);
or U1991 (N_1991,N_969,N_588);
or U1992 (N_1992,N_913,N_666);
and U1993 (N_1993,N_812,N_892);
xnor U1994 (N_1994,N_168,N_38);
nor U1995 (N_1995,N_683,N_584);
nor U1996 (N_1996,N_768,N_677);
or U1997 (N_1997,N_929,N_719);
nand U1998 (N_1998,N_303,N_695);
nor U1999 (N_1999,N_876,N_918);
and U2000 (N_2000,N_1851,N_1633);
or U2001 (N_2001,N_1008,N_1291);
nand U2002 (N_2002,N_1528,N_1597);
nor U2003 (N_2003,N_1768,N_1019);
and U2004 (N_2004,N_1079,N_1563);
and U2005 (N_2005,N_1757,N_1083);
nor U2006 (N_2006,N_1846,N_1630);
and U2007 (N_2007,N_1461,N_1863);
and U2008 (N_2008,N_1705,N_1545);
or U2009 (N_2009,N_1660,N_1918);
or U2010 (N_2010,N_1895,N_1625);
or U2011 (N_2011,N_1653,N_1575);
nand U2012 (N_2012,N_1230,N_1915);
nor U2013 (N_2013,N_1685,N_1410);
nand U2014 (N_2014,N_1284,N_1960);
nand U2015 (N_2015,N_1654,N_1229);
nand U2016 (N_2016,N_1866,N_1560);
xnor U2017 (N_2017,N_1458,N_1295);
nor U2018 (N_2018,N_1692,N_1278);
nand U2019 (N_2019,N_1057,N_1704);
and U2020 (N_2020,N_1273,N_1418);
nand U2021 (N_2021,N_1210,N_1457);
xnor U2022 (N_2022,N_1700,N_1832);
nand U2023 (N_2023,N_1592,N_1228);
and U2024 (N_2024,N_1163,N_1894);
nand U2025 (N_2025,N_1996,N_1287);
or U2026 (N_2026,N_1344,N_1858);
and U2027 (N_2027,N_1060,N_1183);
or U2028 (N_2028,N_1932,N_1138);
nor U2029 (N_2029,N_1025,N_1076);
nor U2030 (N_2030,N_1486,N_1389);
and U2031 (N_2031,N_1154,N_1446);
or U2032 (N_2032,N_1999,N_1441);
nor U2033 (N_2033,N_1550,N_1316);
or U2034 (N_2034,N_1787,N_1107);
nand U2035 (N_2035,N_1725,N_1776);
or U2036 (N_2036,N_1641,N_1385);
nor U2037 (N_2037,N_1549,N_1392);
nand U2038 (N_2038,N_1507,N_1425);
and U2039 (N_2039,N_1595,N_1924);
or U2040 (N_2040,N_1506,N_1128);
or U2041 (N_2041,N_1017,N_1796);
nor U2042 (N_2042,N_1576,N_1394);
and U2043 (N_2043,N_1429,N_1515);
and U2044 (N_2044,N_1124,N_1369);
nand U2045 (N_2045,N_1845,N_1015);
or U2046 (N_2046,N_1783,N_1744);
or U2047 (N_2047,N_1161,N_1123);
or U2048 (N_2048,N_1728,N_1112);
or U2049 (N_2049,N_1979,N_1772);
nor U2050 (N_2050,N_1766,N_1255);
nand U2051 (N_2051,N_1187,N_1074);
nor U2052 (N_2052,N_1227,N_1340);
and U2053 (N_2053,N_1159,N_1212);
or U2054 (N_2054,N_1175,N_1946);
or U2055 (N_2055,N_1677,N_1105);
nand U2056 (N_2056,N_1906,N_1508);
nor U2057 (N_2057,N_1436,N_1140);
xnor U2058 (N_2058,N_1162,N_1405);
and U2059 (N_2059,N_1011,N_1988);
or U2060 (N_2060,N_1945,N_1075);
and U2061 (N_2061,N_1752,N_1192);
nor U2062 (N_2062,N_1839,N_1093);
and U2063 (N_2063,N_1543,N_1214);
nor U2064 (N_2064,N_1809,N_1463);
or U2065 (N_2065,N_1217,N_1880);
nand U2066 (N_2066,N_1044,N_1879);
xnor U2067 (N_2067,N_1817,N_1947);
and U2068 (N_2068,N_1579,N_1538);
and U2069 (N_2069,N_1141,N_1750);
nand U2070 (N_2070,N_1479,N_1155);
and U2071 (N_2071,N_1473,N_1202);
or U2072 (N_2072,N_1574,N_1178);
nand U2073 (N_2073,N_1424,N_1820);
nand U2074 (N_2074,N_1802,N_1968);
nand U2075 (N_2075,N_1353,N_1715);
and U2076 (N_2076,N_1456,N_1805);
nor U2077 (N_2077,N_1379,N_1514);
or U2078 (N_2078,N_1203,N_1050);
nor U2079 (N_2079,N_1673,N_1177);
nand U2080 (N_2080,N_1304,N_1421);
and U2081 (N_2081,N_1064,N_1337);
and U2082 (N_2082,N_1078,N_1559);
nor U2083 (N_2083,N_1836,N_1814);
nor U2084 (N_2084,N_1351,N_1070);
xnor U2085 (N_2085,N_1306,N_1554);
or U2086 (N_2086,N_1003,N_1002);
and U2087 (N_2087,N_1419,N_1738);
or U2088 (N_2088,N_1236,N_1955);
xor U2089 (N_2089,N_1697,N_1584);
or U2090 (N_2090,N_1330,N_1525);
nand U2091 (N_2091,N_1443,N_1849);
nand U2092 (N_2092,N_1620,N_1073);
and U2093 (N_2093,N_1072,N_1089);
nor U2094 (N_2094,N_1031,N_1838);
nand U2095 (N_2095,N_1701,N_1156);
or U2096 (N_2096,N_1961,N_1856);
nand U2097 (N_2097,N_1931,N_1029);
nand U2098 (N_2098,N_1577,N_1129);
and U2099 (N_2099,N_1908,N_1523);
nand U2100 (N_2100,N_1920,N_1611);
nand U2101 (N_2101,N_1748,N_1153);
or U2102 (N_2102,N_1695,N_1355);
nand U2103 (N_2103,N_1322,N_1157);
nor U2104 (N_2104,N_1771,N_1091);
and U2105 (N_2105,N_1669,N_1125);
xor U2106 (N_2106,N_1556,N_1169);
xor U2107 (N_2107,N_1827,N_1835);
nand U2108 (N_2108,N_1134,N_1135);
or U2109 (N_2109,N_1294,N_1813);
nor U2110 (N_2110,N_1784,N_1035);
or U2111 (N_2111,N_1415,N_1109);
and U2112 (N_2112,N_1609,N_1504);
nand U2113 (N_2113,N_1923,N_1742);
and U2114 (N_2114,N_1751,N_1586);
or U2115 (N_2115,N_1068,N_1100);
and U2116 (N_2116,N_1843,N_1948);
nor U2117 (N_2117,N_1220,N_1150);
or U2118 (N_2118,N_1873,N_1269);
nor U2119 (N_2119,N_1250,N_1483);
and U2120 (N_2120,N_1027,N_1264);
nand U2121 (N_2121,N_1088,N_1606);
nand U2122 (N_2122,N_1136,N_1148);
and U2123 (N_2123,N_1887,N_1071);
nand U2124 (N_2124,N_1607,N_1546);
nor U2125 (N_2125,N_1336,N_1434);
and U2126 (N_2126,N_1747,N_1343);
nor U2127 (N_2127,N_1581,N_1241);
or U2128 (N_2128,N_1855,N_1638);
nor U2129 (N_2129,N_1339,N_1235);
or U2130 (N_2130,N_1147,N_1262);
xor U2131 (N_2131,N_1475,N_1661);
nor U2132 (N_2132,N_1197,N_1536);
nand U2133 (N_2133,N_1464,N_1708);
and U2134 (N_2134,N_1867,N_1886);
nor U2135 (N_2135,N_1570,N_1341);
or U2136 (N_2136,N_1454,N_1520);
nand U2137 (N_2137,N_1232,N_1444);
nand U2138 (N_2138,N_1233,N_1553);
nand U2139 (N_2139,N_1094,N_1739);
nor U2140 (N_2140,N_1290,N_1335);
nand U2141 (N_2141,N_1213,N_1489);
xor U2142 (N_2142,N_1986,N_1216);
nand U2143 (N_2143,N_1307,N_1268);
and U2144 (N_2144,N_1300,N_1086);
nand U2145 (N_2145,N_1734,N_1830);
nand U2146 (N_2146,N_1604,N_1605);
nand U2147 (N_2147,N_1934,N_1621);
and U2148 (N_2148,N_1438,N_1758);
and U2149 (N_2149,N_1626,N_1859);
and U2150 (N_2150,N_1404,N_1181);
or U2151 (N_2151,N_1007,N_1608);
or U2152 (N_2152,N_1413,N_1723);
and U2153 (N_2153,N_1885,N_1769);
nand U2154 (N_2154,N_1126,N_1022);
nand U2155 (N_2155,N_1190,N_1451);
xor U2156 (N_2156,N_1234,N_1872);
and U2157 (N_2157,N_1713,N_1984);
nor U2158 (N_2158,N_1224,N_1939);
nand U2159 (N_2159,N_1555,N_1529);
nand U2160 (N_2160,N_1455,N_1569);
nand U2161 (N_2161,N_1816,N_1612);
nor U2162 (N_2162,N_1987,N_1670);
and U2163 (N_2163,N_1376,N_1430);
nand U2164 (N_2164,N_1797,N_1706);
nor U2165 (N_2165,N_1084,N_1703);
nor U2166 (N_2166,N_1943,N_1097);
and U2167 (N_2167,N_1737,N_1365);
nor U2168 (N_2168,N_1145,N_1219);
and U2169 (N_2169,N_1401,N_1082);
and U2170 (N_2170,N_1712,N_1285);
and U2171 (N_2171,N_1298,N_1358);
nand U2172 (N_2172,N_1590,N_1067);
or U2173 (N_2173,N_1326,N_1512);
nor U2174 (N_2174,N_1449,N_1477);
and U2175 (N_2175,N_1045,N_1840);
nand U2176 (N_2176,N_1402,N_1622);
nand U2177 (N_2177,N_1773,N_1266);
and U2178 (N_2178,N_1509,N_1791);
nor U2179 (N_2179,N_1874,N_1828);
nand U2180 (N_2180,N_1052,N_1786);
and U2181 (N_2181,N_1991,N_1499);
nand U2182 (N_2182,N_1599,N_1348);
nand U2183 (N_2183,N_1676,N_1938);
nor U2184 (N_2184,N_1994,N_1903);
nor U2185 (N_2185,N_1720,N_1727);
nor U2186 (N_2186,N_1465,N_1557);
nor U2187 (N_2187,N_1995,N_1912);
and U2188 (N_2188,N_1399,N_1790);
nand U2189 (N_2189,N_1117,N_1922);
and U2190 (N_2190,N_1686,N_1042);
and U2191 (N_2191,N_1884,N_1883);
xnor U2192 (N_2192,N_1977,N_1629);
and U2193 (N_2193,N_1598,N_1741);
nor U2194 (N_2194,N_1349,N_1239);
and U2195 (N_2195,N_1275,N_1591);
nand U2196 (N_2196,N_1716,N_1646);
and U2197 (N_2197,N_1146,N_1400);
nor U2198 (N_2198,N_1092,N_1619);
or U2199 (N_2199,N_1989,N_1667);
nand U2200 (N_2200,N_1637,N_1258);
and U2201 (N_2201,N_1039,N_1580);
and U2202 (N_2202,N_1852,N_1460);
or U2203 (N_2203,N_1485,N_1522);
nor U2204 (N_2204,N_1806,N_1829);
nor U2205 (N_2205,N_1675,N_1648);
nand U2206 (N_2206,N_1870,N_1286);
and U2207 (N_2207,N_1313,N_1253);
nor U2208 (N_2208,N_1770,N_1209);
nand U2209 (N_2209,N_1127,N_1936);
nor U2210 (N_2210,N_1910,N_1541);
and U2211 (N_2211,N_1502,N_1587);
or U2212 (N_2212,N_1009,N_1588);
nand U2213 (N_2213,N_1182,N_1831);
and U2214 (N_2214,N_1657,N_1311);
nor U2215 (N_2215,N_1414,N_1020);
nand U2216 (N_2216,N_1618,N_1833);
nand U2217 (N_2217,N_1482,N_1360);
nand U2218 (N_2218,N_1242,N_1412);
or U2219 (N_2219,N_1274,N_1186);
nor U2220 (N_2220,N_1005,N_1452);
and U2221 (N_2221,N_1564,N_1668);
and U2222 (N_2222,N_1199,N_1658);
or U2223 (N_2223,N_1717,N_1122);
and U2224 (N_2224,N_1530,N_1540);
nand U2225 (N_2225,N_1387,N_1571);
nand U2226 (N_2226,N_1892,N_1257);
and U2227 (N_2227,N_1171,N_1731);
nand U2228 (N_2228,N_1245,N_1659);
nor U2229 (N_2229,N_1665,N_1760);
nand U2230 (N_2230,N_1767,N_1282);
nor U2231 (N_2231,N_1299,N_1318);
nand U2232 (N_2232,N_1913,N_1811);
nand U2233 (N_2233,N_1280,N_1371);
or U2234 (N_2234,N_1423,N_1909);
or U2235 (N_2235,N_1108,N_1524);
or U2236 (N_2236,N_1860,N_1231);
nand U2237 (N_2237,N_1497,N_1959);
nor U2238 (N_2238,N_1868,N_1950);
and U2239 (N_2239,N_1098,N_1366);
or U2240 (N_2240,N_1062,N_1435);
nor U2241 (N_2241,N_1498,N_1222);
xnor U2242 (N_2242,N_1367,N_1370);
and U2243 (N_2243,N_1215,N_1680);
and U2244 (N_2244,N_1130,N_1188);
and U2245 (N_2245,N_1359,N_1848);
nand U2246 (N_2246,N_1777,N_1517);
or U2247 (N_2247,N_1121,N_1998);
or U2248 (N_2248,N_1303,N_1378);
nor U2249 (N_2249,N_1493,N_1753);
nor U2250 (N_2250,N_1864,N_1730);
or U2251 (N_2251,N_1940,N_1119);
nand U2252 (N_2252,N_1180,N_1539);
or U2253 (N_2253,N_1066,N_1671);
nor U2254 (N_2254,N_1890,N_1321);
nand U2255 (N_2255,N_1899,N_1201);
or U2256 (N_2256,N_1195,N_1925);
or U2257 (N_2257,N_1324,N_1778);
nor U2258 (N_2258,N_1645,N_1077);
or U2259 (N_2259,N_1519,N_1058);
and U2260 (N_2260,N_1647,N_1081);
nor U2261 (N_2261,N_1310,N_1755);
xor U2262 (N_2262,N_1568,N_1798);
nand U2263 (N_2263,N_1743,N_1032);
nand U2264 (N_2264,N_1143,N_1893);
and U2265 (N_2265,N_1678,N_1722);
or U2266 (N_2266,N_1476,N_1876);
and U2267 (N_2267,N_1963,N_1036);
and U2268 (N_2268,N_1942,N_1970);
and U2269 (N_2269,N_1320,N_1990);
nor U2270 (N_2270,N_1815,N_1226);
nor U2271 (N_2271,N_1779,N_1276);
nor U2272 (N_2272,N_1142,N_1118);
and U2273 (N_2273,N_1562,N_1432);
nand U2274 (N_2274,N_1634,N_1023);
nor U2275 (N_2275,N_1381,N_1347);
or U2276 (N_2276,N_1279,N_1302);
nor U2277 (N_2277,N_1930,N_1969);
and U2278 (N_2278,N_1496,N_1914);
nand U2279 (N_2279,N_1964,N_1333);
nor U2280 (N_2280,N_1377,N_1439);
or U2281 (N_2281,N_1249,N_1610);
or U2282 (N_2282,N_1566,N_1624);
nor U2283 (N_2283,N_1137,N_1762);
or U2284 (N_2284,N_1825,N_1131);
or U2285 (N_2285,N_1251,N_1211);
or U2286 (N_2286,N_1390,N_1733);
nand U2287 (N_2287,N_1782,N_1521);
or U2288 (N_2288,N_1847,N_1516);
nor U2289 (N_2289,N_1696,N_1308);
nand U2290 (N_2290,N_1325,N_1013);
nor U2291 (N_2291,N_1941,N_1189);
and U2292 (N_2292,N_1469,N_1967);
or U2293 (N_2293,N_1063,N_1099);
nand U2294 (N_2294,N_1411,N_1533);
and U2295 (N_2295,N_1921,N_1467);
or U2296 (N_2296,N_1972,N_1225);
nand U2297 (N_2297,N_1018,N_1904);
nor U2298 (N_2298,N_1875,N_1547);
nand U2299 (N_2299,N_1113,N_1652);
and U2300 (N_2300,N_1272,N_1398);
nor U2301 (N_2301,N_1822,N_1635);
nand U2302 (N_2302,N_1087,N_1926);
and U2303 (N_2303,N_1462,N_1780);
or U2304 (N_2304,N_1511,N_1288);
nor U2305 (N_2305,N_1103,N_1724);
or U2306 (N_2306,N_1132,N_1759);
and U2307 (N_2307,N_1763,N_1433);
or U2308 (N_2308,N_1596,N_1319);
nor U2309 (N_2309,N_1937,N_1297);
or U2310 (N_2310,N_1615,N_1080);
and U2311 (N_2311,N_1259,N_1247);
nor U2312 (N_2312,N_1927,N_1488);
or U2313 (N_2313,N_1204,N_1110);
nor U2314 (N_2314,N_1952,N_1649);
or U2315 (N_2315,N_1980,N_1283);
nand U2316 (N_2316,N_1567,N_1656);
or U2317 (N_2317,N_1983,N_1478);
or U2318 (N_2318,N_1957,N_1021);
nor U2319 (N_2319,N_1632,N_1740);
or U2320 (N_2320,N_1384,N_1601);
or U2321 (N_2321,N_1898,N_1480);
nor U2322 (N_2322,N_1417,N_1168);
and U2323 (N_2323,N_1391,N_1014);
nand U2324 (N_2324,N_1373,N_1674);
or U2325 (N_2325,N_1636,N_1881);
or U2326 (N_2326,N_1386,N_1537);
nand U2327 (N_2327,N_1526,N_1683);
or U2328 (N_2328,N_1012,N_1997);
and U2329 (N_2329,N_1244,N_1114);
and U2330 (N_2330,N_1749,N_1582);
nand U2331 (N_2331,N_1445,N_1949);
nand U2332 (N_2332,N_1403,N_1368);
or U2333 (N_2333,N_1055,N_1594);
and U2334 (N_2334,N_1223,N_1041);
and U2335 (N_2335,N_1407,N_1237);
nor U2336 (N_2336,N_1205,N_1650);
or U2337 (N_2337,N_1746,N_1795);
or U2338 (N_2338,N_1270,N_1312);
nor U2339 (N_2339,N_1929,N_1681);
or U2340 (N_2340,N_1069,N_1917);
and U2341 (N_2341,N_1714,N_1792);
or U2342 (N_2342,N_1573,N_1691);
nand U2343 (N_2343,N_1603,N_1719);
nand U2344 (N_2344,N_1732,N_1271);
xnor U2345 (N_2345,N_1356,N_1248);
or U2346 (N_2346,N_1267,N_1450);
and U2347 (N_2347,N_1643,N_1357);
xnor U2348 (N_2348,N_1170,N_1133);
and U2349 (N_2349,N_1172,N_1785);
nand U2350 (N_2350,N_1185,N_1552);
and U2351 (N_2351,N_1046,N_1718);
nor U2352 (N_2352,N_1470,N_1803);
and U2353 (N_2353,N_1971,N_1165);
and U2354 (N_2354,N_1933,N_1026);
nand U2355 (N_2355,N_1850,N_1854);
nand U2356 (N_2356,N_1487,N_1328);
and U2357 (N_2357,N_1702,N_1837);
nor U2358 (N_2358,N_1466,N_1289);
or U2359 (N_2359,N_1902,N_1754);
or U2360 (N_2360,N_1301,N_1561);
nor U2361 (N_2361,N_1048,N_1551);
nand U2362 (N_2362,N_1729,N_1196);
or U2363 (N_2363,N_1613,N_1982);
nand U2364 (N_2364,N_1651,N_1102);
xor U2365 (N_2365,N_1096,N_1388);
nand U2366 (N_2366,N_1954,N_1437);
nand U2367 (N_2367,N_1338,N_1167);
and U2368 (N_2368,N_1240,N_1260);
nor U2369 (N_2369,N_1207,N_1935);
and U2370 (N_2370,N_1544,N_1965);
nand U2371 (N_2371,N_1891,N_1472);
or U2372 (N_2372,N_1548,N_1642);
and U2373 (N_2373,N_1293,N_1687);
and U2374 (N_2374,N_1865,N_1054);
and U2375 (N_2375,N_1030,N_1166);
nor U2376 (N_2376,N_1558,N_1793);
nor U2377 (N_2377,N_1735,N_1916);
or U2378 (N_2378,N_1655,N_1422);
nand U2379 (N_2379,N_1495,N_1416);
nand U2380 (N_2380,N_1395,N_1628);
or U2381 (N_2381,N_1393,N_1664);
nand U2382 (N_2382,N_1028,N_1788);
or U2383 (N_2383,N_1382,N_1428);
nor U2384 (N_2384,N_1144,N_1765);
nor U2385 (N_2385,N_1174,N_1200);
nand U2386 (N_2386,N_1471,N_1871);
nand U2387 (N_2387,N_1907,N_1491);
and U2388 (N_2388,N_1900,N_1345);
or U2389 (N_2389,N_1263,N_1106);
nor U2390 (N_2390,N_1254,N_1789);
and U2391 (N_2391,N_1427,N_1024);
xnor U2392 (N_2392,N_1761,N_1616);
nor U2393 (N_2393,N_1206,N_1492);
nand U2394 (N_2394,N_1431,N_1101);
nand U2395 (N_2395,N_1694,N_1362);
nand U2396 (N_2396,N_1882,N_1572);
or U2397 (N_2397,N_1468,N_1823);
nand U2398 (N_2398,N_1420,N_1111);
or U2399 (N_2399,N_1578,N_1801);
or U2400 (N_2400,N_1061,N_1104);
nand U2401 (N_2401,N_1614,N_1490);
nand U2402 (N_2402,N_1006,N_1672);
or U2403 (N_2403,N_1966,N_1352);
xnor U2404 (N_2404,N_1243,N_1252);
and U2405 (N_2405,N_1447,N_1627);
nand U2406 (N_2406,N_1095,N_1409);
and U2407 (N_2407,N_1841,N_1756);
or U2408 (N_2408,N_1736,N_1040);
or U2409 (N_2409,N_1518,N_1292);
and U2410 (N_2410,N_1600,N_1975);
or U2411 (N_2411,N_1115,N_1459);
and U2412 (N_2412,N_1120,N_1296);
or U2413 (N_2413,N_1380,N_1152);
nor U2414 (N_2414,N_1047,N_1500);
and U2415 (N_2415,N_1256,N_1531);
or U2416 (N_2416,N_1710,N_1824);
nand U2417 (N_2417,N_1857,N_1602);
or U2418 (N_2418,N_1327,N_1265);
or U2419 (N_2419,N_1221,N_1346);
or U2420 (N_2420,N_1663,N_1993);
or U2421 (N_2421,N_1869,N_1781);
or U2422 (N_2422,N_1453,N_1375);
nand U2423 (N_2423,N_1363,N_1261);
nor U2424 (N_2424,N_1305,N_1342);
nand U2425 (N_2425,N_1775,N_1193);
nand U2426 (N_2426,N_1992,N_1208);
nand U2427 (N_2427,N_1944,N_1281);
or U2428 (N_2428,N_1238,N_1981);
or U2429 (N_2429,N_1583,N_1690);
or U2430 (N_2430,N_1426,N_1503);
xor U2431 (N_2431,N_1709,N_1494);
and U2432 (N_2432,N_1065,N_1361);
or U2433 (N_2433,N_1085,N_1818);
nor U2434 (N_2434,N_1976,N_1699);
and U2435 (N_2435,N_1139,N_1919);
nor U2436 (N_2436,N_1973,N_1593);
nand U2437 (N_2437,N_1034,N_1812);
xnor U2438 (N_2438,N_1090,N_1151);
nor U2439 (N_2439,N_1038,N_1484);
nor U2440 (N_2440,N_1149,N_1640);
nor U2441 (N_2441,N_1745,N_1277);
or U2442 (N_2442,N_1049,N_1534);
and U2443 (N_2443,N_1956,N_1354);
nand U2444 (N_2444,N_1684,N_1510);
nand U2445 (N_2445,N_1897,N_1037);
nand U2446 (N_2446,N_1158,N_1331);
nor U2447 (N_2447,N_1440,N_1707);
or U2448 (N_2448,N_1623,N_1666);
or U2449 (N_2449,N_1928,N_1905);
nand U2450 (N_2450,N_1501,N_1689);
nor U2451 (N_2451,N_1323,N_1059);
nand U2452 (N_2452,N_1315,N_1826);
or U2453 (N_2453,N_1978,N_1764);
and U2454 (N_2454,N_1191,N_1682);
or U2455 (N_2455,N_1198,N_1819);
and U2456 (N_2456,N_1053,N_1962);
nor U2457 (N_2457,N_1821,N_1406);
and U2458 (N_2458,N_1179,N_1116);
and U2459 (N_2459,N_1721,N_1314);
and U2460 (N_2460,N_1834,N_1794);
xnor U2461 (N_2461,N_1810,N_1888);
or U2462 (N_2462,N_1246,N_1218);
nand U2463 (N_2463,N_1505,N_1862);
nor U2464 (N_2464,N_1016,N_1442);
nand U2465 (N_2465,N_1033,N_1662);
nand U2466 (N_2466,N_1951,N_1688);
or U2467 (N_2467,N_1176,N_1585);
or U2468 (N_2468,N_1808,N_1953);
nor U2469 (N_2469,N_1527,N_1974);
nor U2470 (N_2470,N_1901,N_1408);
nor U2471 (N_2471,N_1958,N_1004);
or U2472 (N_2472,N_1164,N_1396);
and U2473 (N_2473,N_1774,N_1542);
nor U2474 (N_2474,N_1056,N_1374);
and U2475 (N_2475,N_1807,N_1448);
or U2476 (N_2476,N_1535,N_1364);
nand U2477 (N_2477,N_1481,N_1160);
nor U2478 (N_2478,N_1513,N_1001);
and U2479 (N_2479,N_1184,N_1726);
nand U2480 (N_2480,N_1861,N_1589);
nor U2481 (N_2481,N_1332,N_1985);
nor U2482 (N_2482,N_1173,N_1693);
or U2483 (N_2483,N_1698,N_1397);
and U2484 (N_2484,N_1631,N_1800);
nor U2485 (N_2485,N_1334,N_1043);
and U2486 (N_2486,N_1889,N_1383);
and U2487 (N_2487,N_1372,N_1804);
and U2488 (N_2488,N_1194,N_1842);
nor U2489 (N_2489,N_1679,N_1844);
nor U2490 (N_2490,N_1896,N_1532);
or U2491 (N_2491,N_1617,N_1911);
nor U2492 (N_2492,N_1711,N_1000);
nor U2493 (N_2493,N_1309,N_1317);
nand U2494 (N_2494,N_1853,N_1639);
nor U2495 (N_2495,N_1329,N_1051);
or U2496 (N_2496,N_1878,N_1010);
and U2497 (N_2497,N_1644,N_1877);
nor U2498 (N_2498,N_1350,N_1474);
or U2499 (N_2499,N_1565,N_1799);
or U2500 (N_2500,N_1091,N_1742);
and U2501 (N_2501,N_1383,N_1118);
or U2502 (N_2502,N_1235,N_1543);
or U2503 (N_2503,N_1539,N_1107);
and U2504 (N_2504,N_1539,N_1844);
or U2505 (N_2505,N_1258,N_1483);
xor U2506 (N_2506,N_1773,N_1906);
or U2507 (N_2507,N_1344,N_1301);
and U2508 (N_2508,N_1305,N_1527);
nor U2509 (N_2509,N_1422,N_1531);
nor U2510 (N_2510,N_1769,N_1350);
nor U2511 (N_2511,N_1953,N_1678);
and U2512 (N_2512,N_1062,N_1056);
nor U2513 (N_2513,N_1345,N_1670);
and U2514 (N_2514,N_1181,N_1528);
and U2515 (N_2515,N_1381,N_1965);
nor U2516 (N_2516,N_1456,N_1636);
and U2517 (N_2517,N_1923,N_1031);
and U2518 (N_2518,N_1248,N_1467);
or U2519 (N_2519,N_1196,N_1596);
or U2520 (N_2520,N_1870,N_1507);
nor U2521 (N_2521,N_1857,N_1649);
and U2522 (N_2522,N_1462,N_1125);
nand U2523 (N_2523,N_1381,N_1830);
and U2524 (N_2524,N_1957,N_1438);
or U2525 (N_2525,N_1521,N_1629);
or U2526 (N_2526,N_1827,N_1884);
nand U2527 (N_2527,N_1208,N_1953);
nor U2528 (N_2528,N_1978,N_1087);
nand U2529 (N_2529,N_1078,N_1045);
or U2530 (N_2530,N_1613,N_1807);
nand U2531 (N_2531,N_1536,N_1787);
nand U2532 (N_2532,N_1040,N_1707);
or U2533 (N_2533,N_1458,N_1552);
and U2534 (N_2534,N_1849,N_1716);
nor U2535 (N_2535,N_1626,N_1337);
nor U2536 (N_2536,N_1836,N_1040);
or U2537 (N_2537,N_1989,N_1473);
nand U2538 (N_2538,N_1582,N_1580);
nor U2539 (N_2539,N_1901,N_1547);
nor U2540 (N_2540,N_1590,N_1830);
or U2541 (N_2541,N_1370,N_1467);
nand U2542 (N_2542,N_1060,N_1854);
or U2543 (N_2543,N_1588,N_1931);
or U2544 (N_2544,N_1282,N_1332);
and U2545 (N_2545,N_1681,N_1190);
nand U2546 (N_2546,N_1022,N_1894);
or U2547 (N_2547,N_1238,N_1384);
or U2548 (N_2548,N_1433,N_1776);
or U2549 (N_2549,N_1685,N_1440);
nor U2550 (N_2550,N_1132,N_1584);
or U2551 (N_2551,N_1463,N_1525);
or U2552 (N_2552,N_1486,N_1393);
and U2553 (N_2553,N_1654,N_1181);
nand U2554 (N_2554,N_1385,N_1195);
nor U2555 (N_2555,N_1622,N_1098);
or U2556 (N_2556,N_1978,N_1469);
or U2557 (N_2557,N_1218,N_1736);
nor U2558 (N_2558,N_1558,N_1864);
and U2559 (N_2559,N_1167,N_1403);
and U2560 (N_2560,N_1756,N_1989);
or U2561 (N_2561,N_1190,N_1826);
nand U2562 (N_2562,N_1484,N_1873);
and U2563 (N_2563,N_1994,N_1104);
and U2564 (N_2564,N_1804,N_1832);
nand U2565 (N_2565,N_1264,N_1786);
xor U2566 (N_2566,N_1326,N_1158);
and U2567 (N_2567,N_1811,N_1378);
and U2568 (N_2568,N_1463,N_1863);
nand U2569 (N_2569,N_1221,N_1982);
nand U2570 (N_2570,N_1383,N_1918);
nor U2571 (N_2571,N_1609,N_1223);
nand U2572 (N_2572,N_1235,N_1728);
and U2573 (N_2573,N_1528,N_1836);
or U2574 (N_2574,N_1405,N_1906);
nand U2575 (N_2575,N_1357,N_1470);
xnor U2576 (N_2576,N_1292,N_1411);
xor U2577 (N_2577,N_1336,N_1457);
and U2578 (N_2578,N_1169,N_1785);
nor U2579 (N_2579,N_1200,N_1869);
and U2580 (N_2580,N_1543,N_1503);
nor U2581 (N_2581,N_1899,N_1276);
and U2582 (N_2582,N_1238,N_1313);
nand U2583 (N_2583,N_1324,N_1951);
or U2584 (N_2584,N_1793,N_1589);
nor U2585 (N_2585,N_1350,N_1977);
nand U2586 (N_2586,N_1880,N_1479);
and U2587 (N_2587,N_1128,N_1919);
and U2588 (N_2588,N_1284,N_1916);
xor U2589 (N_2589,N_1861,N_1206);
nand U2590 (N_2590,N_1420,N_1266);
nor U2591 (N_2591,N_1077,N_1464);
or U2592 (N_2592,N_1034,N_1999);
nand U2593 (N_2593,N_1991,N_1732);
nand U2594 (N_2594,N_1338,N_1986);
and U2595 (N_2595,N_1806,N_1071);
or U2596 (N_2596,N_1594,N_1548);
and U2597 (N_2597,N_1198,N_1343);
nand U2598 (N_2598,N_1748,N_1292);
or U2599 (N_2599,N_1455,N_1000);
nand U2600 (N_2600,N_1765,N_1461);
nand U2601 (N_2601,N_1282,N_1488);
nand U2602 (N_2602,N_1748,N_1585);
nor U2603 (N_2603,N_1679,N_1974);
nand U2604 (N_2604,N_1766,N_1819);
nor U2605 (N_2605,N_1747,N_1024);
or U2606 (N_2606,N_1839,N_1948);
nor U2607 (N_2607,N_1847,N_1284);
nand U2608 (N_2608,N_1509,N_1278);
nor U2609 (N_2609,N_1667,N_1147);
or U2610 (N_2610,N_1273,N_1569);
nor U2611 (N_2611,N_1857,N_1604);
nor U2612 (N_2612,N_1241,N_1077);
and U2613 (N_2613,N_1046,N_1586);
nor U2614 (N_2614,N_1142,N_1445);
and U2615 (N_2615,N_1411,N_1714);
or U2616 (N_2616,N_1614,N_1568);
nor U2617 (N_2617,N_1979,N_1732);
nand U2618 (N_2618,N_1409,N_1377);
nor U2619 (N_2619,N_1751,N_1889);
and U2620 (N_2620,N_1382,N_1704);
nor U2621 (N_2621,N_1510,N_1986);
and U2622 (N_2622,N_1981,N_1604);
or U2623 (N_2623,N_1746,N_1185);
nor U2624 (N_2624,N_1426,N_1788);
nor U2625 (N_2625,N_1111,N_1492);
and U2626 (N_2626,N_1487,N_1450);
nor U2627 (N_2627,N_1093,N_1354);
nor U2628 (N_2628,N_1129,N_1468);
or U2629 (N_2629,N_1396,N_1762);
nor U2630 (N_2630,N_1783,N_1629);
or U2631 (N_2631,N_1030,N_1321);
nand U2632 (N_2632,N_1716,N_1833);
and U2633 (N_2633,N_1894,N_1018);
nand U2634 (N_2634,N_1122,N_1422);
and U2635 (N_2635,N_1578,N_1258);
nor U2636 (N_2636,N_1299,N_1145);
nand U2637 (N_2637,N_1086,N_1053);
nand U2638 (N_2638,N_1039,N_1974);
and U2639 (N_2639,N_1241,N_1032);
nor U2640 (N_2640,N_1107,N_1470);
nor U2641 (N_2641,N_1569,N_1939);
and U2642 (N_2642,N_1146,N_1578);
nand U2643 (N_2643,N_1252,N_1598);
nand U2644 (N_2644,N_1637,N_1536);
nand U2645 (N_2645,N_1524,N_1122);
nand U2646 (N_2646,N_1921,N_1450);
nand U2647 (N_2647,N_1139,N_1210);
and U2648 (N_2648,N_1237,N_1109);
nand U2649 (N_2649,N_1638,N_1557);
nor U2650 (N_2650,N_1735,N_1092);
nor U2651 (N_2651,N_1517,N_1427);
or U2652 (N_2652,N_1726,N_1725);
or U2653 (N_2653,N_1783,N_1984);
and U2654 (N_2654,N_1743,N_1440);
and U2655 (N_2655,N_1374,N_1994);
and U2656 (N_2656,N_1380,N_1270);
or U2657 (N_2657,N_1304,N_1371);
nor U2658 (N_2658,N_1963,N_1988);
and U2659 (N_2659,N_1025,N_1179);
and U2660 (N_2660,N_1247,N_1483);
nor U2661 (N_2661,N_1612,N_1874);
and U2662 (N_2662,N_1777,N_1675);
nand U2663 (N_2663,N_1160,N_1714);
and U2664 (N_2664,N_1430,N_1906);
nor U2665 (N_2665,N_1689,N_1495);
nor U2666 (N_2666,N_1317,N_1890);
nand U2667 (N_2667,N_1552,N_1376);
or U2668 (N_2668,N_1048,N_1654);
nand U2669 (N_2669,N_1467,N_1439);
nand U2670 (N_2670,N_1644,N_1277);
or U2671 (N_2671,N_1478,N_1090);
or U2672 (N_2672,N_1329,N_1043);
or U2673 (N_2673,N_1774,N_1334);
nand U2674 (N_2674,N_1537,N_1296);
or U2675 (N_2675,N_1179,N_1153);
or U2676 (N_2676,N_1560,N_1928);
xnor U2677 (N_2677,N_1872,N_1515);
nor U2678 (N_2678,N_1989,N_1067);
or U2679 (N_2679,N_1961,N_1212);
and U2680 (N_2680,N_1482,N_1143);
nand U2681 (N_2681,N_1472,N_1599);
nand U2682 (N_2682,N_1053,N_1626);
and U2683 (N_2683,N_1815,N_1750);
nor U2684 (N_2684,N_1074,N_1209);
and U2685 (N_2685,N_1253,N_1941);
nand U2686 (N_2686,N_1180,N_1844);
or U2687 (N_2687,N_1341,N_1556);
or U2688 (N_2688,N_1438,N_1730);
and U2689 (N_2689,N_1564,N_1919);
nor U2690 (N_2690,N_1026,N_1847);
nor U2691 (N_2691,N_1166,N_1624);
nor U2692 (N_2692,N_1527,N_1794);
and U2693 (N_2693,N_1543,N_1428);
and U2694 (N_2694,N_1457,N_1189);
nor U2695 (N_2695,N_1589,N_1864);
nor U2696 (N_2696,N_1112,N_1850);
and U2697 (N_2697,N_1274,N_1376);
nand U2698 (N_2698,N_1590,N_1315);
and U2699 (N_2699,N_1360,N_1495);
or U2700 (N_2700,N_1517,N_1042);
nand U2701 (N_2701,N_1514,N_1935);
nor U2702 (N_2702,N_1492,N_1781);
nand U2703 (N_2703,N_1363,N_1101);
nor U2704 (N_2704,N_1402,N_1888);
and U2705 (N_2705,N_1265,N_1954);
nand U2706 (N_2706,N_1690,N_1469);
and U2707 (N_2707,N_1188,N_1059);
nand U2708 (N_2708,N_1859,N_1903);
nand U2709 (N_2709,N_1352,N_1765);
or U2710 (N_2710,N_1774,N_1131);
nor U2711 (N_2711,N_1706,N_1656);
xor U2712 (N_2712,N_1419,N_1193);
xor U2713 (N_2713,N_1785,N_1784);
nand U2714 (N_2714,N_1872,N_1752);
nor U2715 (N_2715,N_1762,N_1392);
and U2716 (N_2716,N_1956,N_1511);
nor U2717 (N_2717,N_1514,N_1065);
nand U2718 (N_2718,N_1090,N_1765);
or U2719 (N_2719,N_1981,N_1555);
nand U2720 (N_2720,N_1333,N_1400);
nand U2721 (N_2721,N_1487,N_1380);
nor U2722 (N_2722,N_1722,N_1035);
nor U2723 (N_2723,N_1781,N_1642);
or U2724 (N_2724,N_1101,N_1436);
nor U2725 (N_2725,N_1548,N_1581);
nor U2726 (N_2726,N_1704,N_1926);
xor U2727 (N_2727,N_1443,N_1046);
and U2728 (N_2728,N_1568,N_1270);
and U2729 (N_2729,N_1016,N_1447);
or U2730 (N_2730,N_1270,N_1227);
nor U2731 (N_2731,N_1590,N_1802);
or U2732 (N_2732,N_1957,N_1758);
nand U2733 (N_2733,N_1653,N_1466);
and U2734 (N_2734,N_1594,N_1231);
and U2735 (N_2735,N_1910,N_1749);
nand U2736 (N_2736,N_1350,N_1614);
or U2737 (N_2737,N_1673,N_1343);
or U2738 (N_2738,N_1370,N_1294);
or U2739 (N_2739,N_1796,N_1799);
nand U2740 (N_2740,N_1757,N_1241);
and U2741 (N_2741,N_1093,N_1991);
nor U2742 (N_2742,N_1687,N_1334);
nand U2743 (N_2743,N_1355,N_1487);
nand U2744 (N_2744,N_1211,N_1319);
nor U2745 (N_2745,N_1202,N_1037);
nand U2746 (N_2746,N_1316,N_1420);
nand U2747 (N_2747,N_1826,N_1912);
nor U2748 (N_2748,N_1938,N_1212);
nor U2749 (N_2749,N_1519,N_1777);
nor U2750 (N_2750,N_1629,N_1917);
and U2751 (N_2751,N_1748,N_1742);
nand U2752 (N_2752,N_1245,N_1820);
and U2753 (N_2753,N_1900,N_1462);
nand U2754 (N_2754,N_1306,N_1899);
and U2755 (N_2755,N_1307,N_1660);
nor U2756 (N_2756,N_1940,N_1514);
nor U2757 (N_2757,N_1303,N_1542);
and U2758 (N_2758,N_1967,N_1440);
nor U2759 (N_2759,N_1588,N_1448);
and U2760 (N_2760,N_1166,N_1893);
nand U2761 (N_2761,N_1788,N_1007);
and U2762 (N_2762,N_1110,N_1916);
and U2763 (N_2763,N_1822,N_1609);
nor U2764 (N_2764,N_1637,N_1100);
nand U2765 (N_2765,N_1175,N_1665);
or U2766 (N_2766,N_1946,N_1694);
or U2767 (N_2767,N_1929,N_1266);
nor U2768 (N_2768,N_1479,N_1022);
or U2769 (N_2769,N_1487,N_1614);
nor U2770 (N_2770,N_1057,N_1712);
and U2771 (N_2771,N_1730,N_1469);
xor U2772 (N_2772,N_1711,N_1746);
nand U2773 (N_2773,N_1166,N_1272);
and U2774 (N_2774,N_1135,N_1591);
nand U2775 (N_2775,N_1658,N_1490);
nand U2776 (N_2776,N_1467,N_1190);
and U2777 (N_2777,N_1772,N_1046);
nor U2778 (N_2778,N_1802,N_1963);
and U2779 (N_2779,N_1533,N_1835);
nand U2780 (N_2780,N_1542,N_1798);
and U2781 (N_2781,N_1556,N_1120);
nor U2782 (N_2782,N_1116,N_1934);
nand U2783 (N_2783,N_1139,N_1297);
nor U2784 (N_2784,N_1089,N_1594);
nor U2785 (N_2785,N_1515,N_1821);
nand U2786 (N_2786,N_1761,N_1361);
and U2787 (N_2787,N_1006,N_1399);
nand U2788 (N_2788,N_1951,N_1820);
and U2789 (N_2789,N_1957,N_1048);
nand U2790 (N_2790,N_1360,N_1636);
nor U2791 (N_2791,N_1327,N_1274);
and U2792 (N_2792,N_1997,N_1675);
nand U2793 (N_2793,N_1374,N_1329);
nand U2794 (N_2794,N_1745,N_1438);
or U2795 (N_2795,N_1930,N_1978);
and U2796 (N_2796,N_1211,N_1232);
and U2797 (N_2797,N_1752,N_1461);
and U2798 (N_2798,N_1562,N_1757);
nand U2799 (N_2799,N_1805,N_1050);
nor U2800 (N_2800,N_1814,N_1124);
nand U2801 (N_2801,N_1322,N_1317);
nand U2802 (N_2802,N_1200,N_1449);
nand U2803 (N_2803,N_1213,N_1426);
and U2804 (N_2804,N_1864,N_1664);
or U2805 (N_2805,N_1961,N_1729);
and U2806 (N_2806,N_1452,N_1046);
and U2807 (N_2807,N_1307,N_1321);
and U2808 (N_2808,N_1887,N_1419);
nor U2809 (N_2809,N_1849,N_1820);
or U2810 (N_2810,N_1519,N_1737);
or U2811 (N_2811,N_1553,N_1385);
or U2812 (N_2812,N_1794,N_1352);
nand U2813 (N_2813,N_1331,N_1569);
nand U2814 (N_2814,N_1347,N_1167);
or U2815 (N_2815,N_1012,N_1568);
or U2816 (N_2816,N_1436,N_1807);
and U2817 (N_2817,N_1819,N_1542);
or U2818 (N_2818,N_1520,N_1750);
or U2819 (N_2819,N_1881,N_1534);
nor U2820 (N_2820,N_1593,N_1087);
and U2821 (N_2821,N_1035,N_1894);
and U2822 (N_2822,N_1202,N_1020);
or U2823 (N_2823,N_1402,N_1218);
or U2824 (N_2824,N_1721,N_1029);
or U2825 (N_2825,N_1721,N_1982);
and U2826 (N_2826,N_1531,N_1992);
or U2827 (N_2827,N_1220,N_1322);
or U2828 (N_2828,N_1496,N_1082);
nand U2829 (N_2829,N_1574,N_1734);
nand U2830 (N_2830,N_1112,N_1730);
or U2831 (N_2831,N_1252,N_1510);
and U2832 (N_2832,N_1228,N_1762);
and U2833 (N_2833,N_1008,N_1507);
or U2834 (N_2834,N_1193,N_1724);
or U2835 (N_2835,N_1631,N_1072);
and U2836 (N_2836,N_1827,N_1135);
or U2837 (N_2837,N_1916,N_1593);
nor U2838 (N_2838,N_1527,N_1665);
nand U2839 (N_2839,N_1857,N_1493);
and U2840 (N_2840,N_1637,N_1593);
nand U2841 (N_2841,N_1286,N_1311);
nor U2842 (N_2842,N_1738,N_1109);
nand U2843 (N_2843,N_1658,N_1127);
nand U2844 (N_2844,N_1912,N_1490);
or U2845 (N_2845,N_1032,N_1211);
or U2846 (N_2846,N_1130,N_1948);
nand U2847 (N_2847,N_1913,N_1058);
and U2848 (N_2848,N_1652,N_1211);
nand U2849 (N_2849,N_1554,N_1583);
nor U2850 (N_2850,N_1294,N_1793);
nand U2851 (N_2851,N_1750,N_1547);
nor U2852 (N_2852,N_1931,N_1340);
or U2853 (N_2853,N_1232,N_1005);
xor U2854 (N_2854,N_1397,N_1110);
nand U2855 (N_2855,N_1759,N_1269);
nand U2856 (N_2856,N_1433,N_1933);
and U2857 (N_2857,N_1818,N_1752);
or U2858 (N_2858,N_1860,N_1570);
nand U2859 (N_2859,N_1913,N_1619);
and U2860 (N_2860,N_1103,N_1372);
or U2861 (N_2861,N_1199,N_1020);
or U2862 (N_2862,N_1977,N_1725);
or U2863 (N_2863,N_1502,N_1049);
xnor U2864 (N_2864,N_1558,N_1858);
xnor U2865 (N_2865,N_1091,N_1579);
nand U2866 (N_2866,N_1813,N_1359);
or U2867 (N_2867,N_1613,N_1097);
nand U2868 (N_2868,N_1601,N_1301);
nor U2869 (N_2869,N_1732,N_1186);
or U2870 (N_2870,N_1911,N_1800);
nor U2871 (N_2871,N_1914,N_1838);
or U2872 (N_2872,N_1963,N_1039);
or U2873 (N_2873,N_1887,N_1423);
nand U2874 (N_2874,N_1865,N_1314);
nand U2875 (N_2875,N_1373,N_1118);
or U2876 (N_2876,N_1980,N_1802);
and U2877 (N_2877,N_1577,N_1747);
and U2878 (N_2878,N_1158,N_1906);
nor U2879 (N_2879,N_1784,N_1395);
nand U2880 (N_2880,N_1860,N_1599);
or U2881 (N_2881,N_1568,N_1584);
and U2882 (N_2882,N_1079,N_1984);
and U2883 (N_2883,N_1442,N_1607);
or U2884 (N_2884,N_1763,N_1427);
nor U2885 (N_2885,N_1046,N_1225);
or U2886 (N_2886,N_1219,N_1372);
nand U2887 (N_2887,N_1491,N_1221);
nand U2888 (N_2888,N_1568,N_1622);
nor U2889 (N_2889,N_1828,N_1793);
or U2890 (N_2890,N_1549,N_1629);
and U2891 (N_2891,N_1971,N_1892);
nand U2892 (N_2892,N_1439,N_1817);
nor U2893 (N_2893,N_1124,N_1363);
nand U2894 (N_2894,N_1574,N_1767);
or U2895 (N_2895,N_1531,N_1380);
xor U2896 (N_2896,N_1140,N_1404);
or U2897 (N_2897,N_1658,N_1223);
or U2898 (N_2898,N_1952,N_1325);
nor U2899 (N_2899,N_1443,N_1964);
nand U2900 (N_2900,N_1786,N_1178);
or U2901 (N_2901,N_1741,N_1584);
or U2902 (N_2902,N_1422,N_1328);
and U2903 (N_2903,N_1418,N_1318);
nor U2904 (N_2904,N_1932,N_1204);
nand U2905 (N_2905,N_1068,N_1492);
nand U2906 (N_2906,N_1088,N_1891);
nand U2907 (N_2907,N_1833,N_1760);
and U2908 (N_2908,N_1804,N_1769);
and U2909 (N_2909,N_1757,N_1041);
xnor U2910 (N_2910,N_1974,N_1784);
and U2911 (N_2911,N_1626,N_1966);
or U2912 (N_2912,N_1156,N_1295);
xor U2913 (N_2913,N_1035,N_1257);
or U2914 (N_2914,N_1847,N_1288);
nand U2915 (N_2915,N_1083,N_1215);
nand U2916 (N_2916,N_1906,N_1578);
nor U2917 (N_2917,N_1526,N_1995);
nand U2918 (N_2918,N_1627,N_1580);
or U2919 (N_2919,N_1376,N_1354);
and U2920 (N_2920,N_1424,N_1709);
or U2921 (N_2921,N_1711,N_1186);
nand U2922 (N_2922,N_1423,N_1119);
nor U2923 (N_2923,N_1152,N_1018);
xor U2924 (N_2924,N_1624,N_1088);
or U2925 (N_2925,N_1380,N_1271);
nand U2926 (N_2926,N_1014,N_1766);
nand U2927 (N_2927,N_1679,N_1077);
nor U2928 (N_2928,N_1726,N_1502);
or U2929 (N_2929,N_1235,N_1192);
or U2930 (N_2930,N_1297,N_1290);
nor U2931 (N_2931,N_1851,N_1448);
xnor U2932 (N_2932,N_1150,N_1515);
nand U2933 (N_2933,N_1920,N_1213);
and U2934 (N_2934,N_1870,N_1271);
and U2935 (N_2935,N_1474,N_1124);
and U2936 (N_2936,N_1992,N_1130);
and U2937 (N_2937,N_1482,N_1059);
and U2938 (N_2938,N_1721,N_1143);
nand U2939 (N_2939,N_1747,N_1454);
nor U2940 (N_2940,N_1439,N_1933);
nand U2941 (N_2941,N_1678,N_1551);
nor U2942 (N_2942,N_1500,N_1089);
or U2943 (N_2943,N_1265,N_1025);
or U2944 (N_2944,N_1732,N_1138);
nor U2945 (N_2945,N_1461,N_1201);
nor U2946 (N_2946,N_1136,N_1311);
or U2947 (N_2947,N_1670,N_1791);
and U2948 (N_2948,N_1263,N_1995);
and U2949 (N_2949,N_1646,N_1581);
nand U2950 (N_2950,N_1665,N_1731);
nor U2951 (N_2951,N_1111,N_1839);
and U2952 (N_2952,N_1008,N_1161);
nand U2953 (N_2953,N_1233,N_1857);
nand U2954 (N_2954,N_1076,N_1016);
or U2955 (N_2955,N_1675,N_1200);
or U2956 (N_2956,N_1841,N_1833);
nand U2957 (N_2957,N_1085,N_1240);
and U2958 (N_2958,N_1318,N_1021);
nor U2959 (N_2959,N_1313,N_1742);
nor U2960 (N_2960,N_1875,N_1633);
nor U2961 (N_2961,N_1216,N_1778);
nor U2962 (N_2962,N_1931,N_1080);
or U2963 (N_2963,N_1047,N_1864);
nor U2964 (N_2964,N_1747,N_1355);
nand U2965 (N_2965,N_1425,N_1166);
nand U2966 (N_2966,N_1615,N_1066);
nor U2967 (N_2967,N_1039,N_1835);
or U2968 (N_2968,N_1689,N_1176);
nor U2969 (N_2969,N_1955,N_1807);
or U2970 (N_2970,N_1417,N_1401);
nand U2971 (N_2971,N_1376,N_1727);
nand U2972 (N_2972,N_1705,N_1865);
or U2973 (N_2973,N_1785,N_1919);
xor U2974 (N_2974,N_1242,N_1077);
and U2975 (N_2975,N_1429,N_1840);
and U2976 (N_2976,N_1106,N_1308);
or U2977 (N_2977,N_1731,N_1147);
and U2978 (N_2978,N_1615,N_1856);
nor U2979 (N_2979,N_1310,N_1437);
nand U2980 (N_2980,N_1268,N_1656);
nor U2981 (N_2981,N_1147,N_1909);
xnor U2982 (N_2982,N_1565,N_1729);
nor U2983 (N_2983,N_1384,N_1614);
or U2984 (N_2984,N_1967,N_1711);
nor U2985 (N_2985,N_1880,N_1940);
or U2986 (N_2986,N_1088,N_1361);
nor U2987 (N_2987,N_1088,N_1423);
nand U2988 (N_2988,N_1148,N_1567);
and U2989 (N_2989,N_1037,N_1179);
and U2990 (N_2990,N_1215,N_1843);
nor U2991 (N_2991,N_1523,N_1546);
xnor U2992 (N_2992,N_1024,N_1273);
nor U2993 (N_2993,N_1937,N_1776);
or U2994 (N_2994,N_1303,N_1809);
nor U2995 (N_2995,N_1917,N_1587);
and U2996 (N_2996,N_1302,N_1164);
nor U2997 (N_2997,N_1837,N_1870);
nand U2998 (N_2998,N_1493,N_1461);
or U2999 (N_2999,N_1708,N_1288);
nand UO_0 (O_0,N_2280,N_2385);
nand UO_1 (O_1,N_2861,N_2166);
or UO_2 (O_2,N_2423,N_2155);
nand UO_3 (O_3,N_2800,N_2834);
nand UO_4 (O_4,N_2935,N_2974);
nand UO_5 (O_5,N_2364,N_2424);
and UO_6 (O_6,N_2767,N_2836);
and UO_7 (O_7,N_2776,N_2324);
or UO_8 (O_8,N_2617,N_2810);
nand UO_9 (O_9,N_2415,N_2737);
nor UO_10 (O_10,N_2741,N_2441);
or UO_11 (O_11,N_2140,N_2124);
nor UO_12 (O_12,N_2127,N_2076);
and UO_13 (O_13,N_2173,N_2807);
and UO_14 (O_14,N_2572,N_2125);
nor UO_15 (O_15,N_2611,N_2464);
or UO_16 (O_16,N_2799,N_2506);
and UO_17 (O_17,N_2754,N_2926);
and UO_18 (O_18,N_2349,N_2846);
and UO_19 (O_19,N_2075,N_2882);
nand UO_20 (O_20,N_2784,N_2803);
nand UO_21 (O_21,N_2106,N_2240);
and UO_22 (O_22,N_2956,N_2139);
and UO_23 (O_23,N_2507,N_2779);
nor UO_24 (O_24,N_2516,N_2213);
nand UO_25 (O_25,N_2607,N_2137);
nor UO_26 (O_26,N_2496,N_2413);
and UO_27 (O_27,N_2230,N_2686);
or UO_28 (O_28,N_2063,N_2002);
nor UO_29 (O_29,N_2856,N_2592);
nand UO_30 (O_30,N_2334,N_2520);
or UO_31 (O_31,N_2477,N_2422);
nand UO_32 (O_32,N_2197,N_2820);
and UO_33 (O_33,N_2222,N_2198);
and UO_34 (O_34,N_2255,N_2603);
nor UO_35 (O_35,N_2320,N_2093);
nor UO_36 (O_36,N_2792,N_2388);
nand UO_37 (O_37,N_2463,N_2621);
nand UO_38 (O_38,N_2404,N_2589);
or UO_39 (O_39,N_2838,N_2237);
nand UO_40 (O_40,N_2046,N_2120);
or UO_41 (O_41,N_2628,N_2962);
nand UO_42 (O_42,N_2340,N_2703);
or UO_43 (O_43,N_2157,N_2486);
xnor UO_44 (O_44,N_2937,N_2346);
xnor UO_45 (O_45,N_2262,N_2577);
nand UO_46 (O_46,N_2062,N_2497);
or UO_47 (O_47,N_2397,N_2912);
nor UO_48 (O_48,N_2399,N_2019);
nand UO_49 (O_49,N_2027,N_2499);
nor UO_50 (O_50,N_2566,N_2398);
or UO_51 (O_51,N_2778,N_2406);
or UO_52 (O_52,N_2026,N_2874);
nor UO_53 (O_53,N_2528,N_2259);
nor UO_54 (O_54,N_2261,N_2246);
nor UO_55 (O_55,N_2529,N_2887);
nand UO_56 (O_56,N_2739,N_2037);
or UO_57 (O_57,N_2078,N_2360);
nor UO_58 (O_58,N_2135,N_2475);
nand UO_59 (O_59,N_2457,N_2878);
or UO_60 (O_60,N_2492,N_2450);
nor UO_61 (O_61,N_2050,N_2410);
or UO_62 (O_62,N_2401,N_2546);
and UO_63 (O_63,N_2654,N_2084);
xnor UO_64 (O_64,N_2664,N_2158);
or UO_65 (O_65,N_2941,N_2719);
or UO_66 (O_66,N_2352,N_2122);
nor UO_67 (O_67,N_2631,N_2599);
nor UO_68 (O_68,N_2333,N_2503);
and UO_69 (O_69,N_2227,N_2451);
or UO_70 (O_70,N_2970,N_2430);
and UO_71 (O_71,N_2482,N_2161);
or UO_72 (O_72,N_2001,N_2260);
nand UO_73 (O_73,N_2613,N_2134);
nand UO_74 (O_74,N_2247,N_2278);
nand UO_75 (O_75,N_2304,N_2112);
and UO_76 (O_76,N_2371,N_2618);
nand UO_77 (O_77,N_2688,N_2378);
or UO_78 (O_78,N_2072,N_2403);
nor UO_79 (O_79,N_2321,N_2817);
nand UO_80 (O_80,N_2858,N_2187);
nand UO_81 (O_81,N_2585,N_2829);
or UO_82 (O_82,N_2344,N_2449);
nand UO_83 (O_83,N_2070,N_2625);
and UO_84 (O_84,N_2479,N_2827);
nand UO_85 (O_85,N_2761,N_2927);
or UO_86 (O_86,N_2556,N_2971);
and UO_87 (O_87,N_2272,N_2995);
or UO_88 (O_88,N_2069,N_2024);
nor UO_89 (O_89,N_2752,N_2170);
nand UO_90 (O_90,N_2900,N_2372);
nand UO_91 (O_91,N_2315,N_2409);
or UO_92 (O_92,N_2952,N_2171);
nor UO_93 (O_93,N_2405,N_2115);
or UO_94 (O_94,N_2208,N_2056);
and UO_95 (O_95,N_2215,N_2736);
and UO_96 (O_96,N_2472,N_2593);
or UO_97 (O_97,N_2682,N_2407);
and UO_98 (O_98,N_2203,N_2561);
and UO_99 (O_99,N_2744,N_2299);
and UO_100 (O_100,N_2487,N_2966);
and UO_101 (O_101,N_2563,N_2953);
nor UO_102 (O_102,N_2071,N_2505);
nor UO_103 (O_103,N_2588,N_2092);
nand UO_104 (O_104,N_2281,N_2651);
or UO_105 (O_105,N_2484,N_2708);
nor UO_106 (O_106,N_2055,N_2738);
nor UO_107 (O_107,N_2221,N_2017);
xnor UO_108 (O_108,N_2687,N_2335);
xor UO_109 (O_109,N_2728,N_2411);
nor UO_110 (O_110,N_2036,N_2747);
or UO_111 (O_111,N_2266,N_2250);
nor UO_112 (O_112,N_2057,N_2351);
or UO_113 (O_113,N_2574,N_2059);
or UO_114 (O_114,N_2141,N_2600);
and UO_115 (O_115,N_2949,N_2675);
nor UO_116 (O_116,N_2077,N_2841);
and UO_117 (O_117,N_2855,N_2149);
nand UO_118 (O_118,N_2214,N_2612);
nand UO_119 (O_119,N_2976,N_2053);
or UO_120 (O_120,N_2374,N_2681);
xnor UO_121 (O_121,N_2981,N_2919);
and UO_122 (O_122,N_2323,N_2363);
nor UO_123 (O_123,N_2571,N_2969);
nand UO_124 (O_124,N_2847,N_2853);
and UO_125 (O_125,N_2502,N_2542);
or UO_126 (O_126,N_2726,N_2101);
or UO_127 (O_127,N_2095,N_2504);
nor UO_128 (O_128,N_2151,N_2354);
and UO_129 (O_129,N_2011,N_2753);
and UO_130 (O_130,N_2760,N_2192);
and UO_131 (O_131,N_2515,N_2073);
nor UO_132 (O_132,N_2030,N_2730);
xnor UO_133 (O_133,N_2713,N_2035);
or UO_134 (O_134,N_2996,N_2284);
nor UO_135 (O_135,N_2119,N_2443);
or UO_136 (O_136,N_2945,N_2327);
nor UO_137 (O_137,N_2567,N_2045);
or UO_138 (O_138,N_2328,N_2696);
or UO_139 (O_139,N_2283,N_2832);
and UO_140 (O_140,N_2086,N_2781);
nor UO_141 (O_141,N_2940,N_2025);
and UO_142 (O_142,N_2640,N_2332);
nor UO_143 (O_143,N_2083,N_2908);
nand UO_144 (O_144,N_2559,N_2462);
nand UO_145 (O_145,N_2831,N_2745);
nor UO_146 (O_146,N_2925,N_2645);
nand UO_147 (O_147,N_2153,N_2331);
and UO_148 (O_148,N_2287,N_2749);
nand UO_149 (O_149,N_2438,N_2176);
nor UO_150 (O_150,N_2312,N_2432);
and UO_151 (O_151,N_2903,N_2500);
nand UO_152 (O_152,N_2608,N_2370);
or UO_153 (O_153,N_2715,N_2862);
nor UO_154 (O_154,N_2967,N_2932);
nand UO_155 (O_155,N_2560,N_2032);
and UO_156 (O_156,N_2518,N_2389);
nor UO_157 (O_157,N_2376,N_2110);
nand UO_158 (O_158,N_2793,N_2609);
nor UO_159 (O_159,N_2318,N_2782);
or UO_160 (O_160,N_2308,N_2771);
or UO_161 (O_161,N_2551,N_2126);
and UO_162 (O_162,N_2285,N_2802);
or UO_163 (O_163,N_2590,N_2160);
nand UO_164 (O_164,N_2154,N_2606);
or UO_165 (O_165,N_2762,N_2712);
and UO_166 (O_166,N_2873,N_2750);
nor UO_167 (O_167,N_2938,N_2601);
nor UO_168 (O_168,N_2890,N_2013);
and UO_169 (O_169,N_2074,N_2704);
nor UO_170 (O_170,N_2302,N_2519);
or UO_171 (O_171,N_2523,N_2380);
and UO_172 (O_172,N_2629,N_2954);
or UO_173 (O_173,N_2209,N_2842);
nor UO_174 (O_174,N_2694,N_2396);
nor UO_175 (O_175,N_2860,N_2723);
or UO_176 (O_176,N_2685,N_2196);
or UO_177 (O_177,N_2986,N_2416);
or UO_178 (O_178,N_2564,N_2553);
nand UO_179 (O_179,N_2852,N_2480);
nor UO_180 (O_180,N_2531,N_2489);
and UO_181 (O_181,N_2034,N_2478);
nor UO_182 (O_182,N_2256,N_2991);
nand UO_183 (O_183,N_2768,N_2867);
and UO_184 (O_184,N_2041,N_2298);
xor UO_185 (O_185,N_2907,N_2711);
nand UO_186 (O_186,N_2317,N_2097);
nand UO_187 (O_187,N_2316,N_2658);
nand UO_188 (O_188,N_2641,N_2325);
and UO_189 (O_189,N_2412,N_2337);
xor UO_190 (O_190,N_2647,N_2183);
nand UO_191 (O_191,N_2236,N_2718);
or UO_192 (O_192,N_2948,N_2229);
nand UO_193 (O_193,N_2709,N_2368);
nor UO_194 (O_194,N_2469,N_2445);
nand UO_195 (O_195,N_2845,N_2942);
or UO_196 (O_196,N_2216,N_2452);
and UO_197 (O_197,N_2999,N_2113);
or UO_198 (O_198,N_2624,N_2094);
or UO_199 (O_199,N_2290,N_2693);
nor UO_200 (O_200,N_2476,N_2985);
or UO_201 (O_201,N_2082,N_2047);
and UO_202 (O_202,N_2616,N_2773);
nor UO_203 (O_203,N_2460,N_2899);
nand UO_204 (O_204,N_2795,N_2018);
and UO_205 (O_205,N_2065,N_2205);
nand UO_206 (O_206,N_2883,N_2207);
nand UO_207 (O_207,N_2555,N_2468);
or UO_208 (O_208,N_2079,N_2669);
or UO_209 (O_209,N_2068,N_2794);
nand UO_210 (O_210,N_2843,N_2223);
xnor UO_211 (O_211,N_2929,N_2722);
nor UO_212 (O_212,N_2634,N_2251);
and UO_213 (O_213,N_2851,N_2642);
or UO_214 (O_214,N_2626,N_2978);
or UO_215 (O_215,N_2797,N_2545);
and UO_216 (O_216,N_2764,N_2982);
nand UO_217 (O_217,N_2557,N_2193);
and UO_218 (O_218,N_2393,N_2731);
nand UO_219 (O_219,N_2189,N_2677);
and UO_220 (O_220,N_2454,N_2806);
xor UO_221 (O_221,N_2924,N_2210);
and UO_222 (O_222,N_2444,N_2031);
xnor UO_223 (O_223,N_2185,N_2249);
nand UO_224 (O_224,N_2225,N_2898);
or UO_225 (O_225,N_2200,N_2386);
and UO_226 (O_226,N_2373,N_2228);
and UO_227 (O_227,N_2512,N_2394);
or UO_228 (O_228,N_2253,N_2596);
nor UO_229 (O_229,N_2008,N_2653);
or UO_230 (O_230,N_2267,N_2839);
nand UO_231 (O_231,N_2014,N_2191);
and UO_232 (O_232,N_2530,N_2648);
xor UO_233 (O_233,N_2885,N_2358);
nand UO_234 (O_234,N_2594,N_2038);
and UO_235 (O_235,N_2769,N_2917);
and UO_236 (O_236,N_2180,N_2459);
or UO_237 (O_237,N_2177,N_2786);
or UO_238 (O_238,N_2921,N_2989);
or UO_239 (O_239,N_2421,N_2144);
nand UO_240 (O_240,N_2548,N_2639);
and UO_241 (O_241,N_2695,N_2652);
or UO_242 (O_242,N_2636,N_2414);
and UO_243 (O_243,N_2823,N_2980);
nand UO_244 (O_244,N_2649,N_2785);
or UO_245 (O_245,N_2751,N_2638);
xor UO_246 (O_246,N_2850,N_2714);
or UO_247 (O_247,N_2920,N_2788);
and UO_248 (O_248,N_2022,N_2759);
nor UO_249 (O_249,N_2835,N_2164);
or UO_250 (O_250,N_2345,N_2809);
and UO_251 (O_251,N_2869,N_2252);
and UO_252 (O_252,N_2233,N_2455);
or UO_253 (O_253,N_2911,N_2973);
and UO_254 (O_254,N_2258,N_2665);
nor UO_255 (O_255,N_2264,N_2534);
or UO_256 (O_256,N_2743,N_2000);
or UO_257 (O_257,N_2558,N_2990);
and UO_258 (O_258,N_2620,N_2777);
and UO_259 (O_259,N_2958,N_2182);
nand UO_260 (O_260,N_2081,N_2798);
or UO_261 (O_261,N_2347,N_2959);
nor UO_262 (O_262,N_2586,N_2757);
and UO_263 (O_263,N_2904,N_2089);
or UO_264 (O_264,N_2066,N_2133);
or UO_265 (O_265,N_2550,N_2811);
or UO_266 (O_266,N_2637,N_2175);
nor UO_267 (O_267,N_2003,N_2275);
nand UO_268 (O_268,N_2359,N_2868);
nor UO_269 (O_269,N_2532,N_2871);
nor UO_270 (O_270,N_2309,N_2541);
or UO_271 (O_271,N_2341,N_2150);
nor UO_272 (O_272,N_2968,N_2439);
nor UO_273 (O_273,N_2977,N_2440);
nand UO_274 (O_274,N_2384,N_2698);
nand UO_275 (O_275,N_2067,N_2471);
nand UO_276 (O_276,N_2897,N_2143);
nand UO_277 (O_277,N_2872,N_2395);
nand UO_278 (O_278,N_2565,N_2880);
nand UO_279 (O_279,N_2429,N_2218);
nor UO_280 (O_280,N_2391,N_2543);
and UO_281 (O_281,N_2822,N_2552);
nor UO_282 (O_282,N_2104,N_2544);
or UO_283 (O_283,N_2387,N_2840);
nand UO_284 (O_284,N_2734,N_2453);
nand UO_285 (O_285,N_2268,N_2684);
nor UO_286 (O_286,N_2679,N_2427);
or UO_287 (O_287,N_2951,N_2099);
nor UO_288 (O_288,N_2735,N_2914);
and UO_289 (O_289,N_2501,N_2244);
and UO_290 (O_290,N_2238,N_2123);
nor UO_291 (O_291,N_2655,N_2804);
or UO_292 (O_292,N_2494,N_2549);
nor UO_293 (O_293,N_2576,N_2691);
nand UO_294 (O_294,N_2052,N_2790);
nor UO_295 (O_295,N_2091,N_2188);
nand UO_296 (O_296,N_2051,N_2965);
or UO_297 (O_297,N_2772,N_2305);
and UO_298 (O_298,N_2179,N_2524);
and UO_299 (O_299,N_2231,N_2825);
nand UO_300 (O_300,N_2296,N_2243);
or UO_301 (O_301,N_2998,N_2058);
or UO_302 (O_302,N_2595,N_2306);
or UO_303 (O_303,N_2930,N_2178);
and UO_304 (O_304,N_2659,N_2527);
nand UO_305 (O_305,N_2859,N_2064);
or UO_306 (O_306,N_2526,N_2163);
nor UO_307 (O_307,N_2787,N_2844);
and UO_308 (O_308,N_2756,N_2294);
and UO_309 (O_309,N_2666,N_2049);
or UO_310 (O_310,N_2382,N_2016);
nand UO_311 (O_311,N_2136,N_2604);
or UO_312 (O_312,N_2162,N_2796);
nand UO_313 (O_313,N_2392,N_2905);
or UO_314 (O_314,N_2029,N_2632);
or UO_315 (O_315,N_2879,N_2006);
or UO_316 (O_316,N_2909,N_2533);
or UO_317 (O_317,N_2671,N_2100);
nand UO_318 (O_318,N_2434,N_2495);
nand UO_319 (O_319,N_2291,N_2165);
xor UO_320 (O_320,N_2812,N_2118);
nor UO_321 (O_321,N_2010,N_2428);
or UO_322 (O_322,N_2627,N_2313);
nand UO_323 (O_323,N_2766,N_2437);
and UO_324 (O_324,N_2888,N_2581);
nor UO_325 (O_325,N_2987,N_2511);
and UO_326 (O_326,N_2993,N_2670);
and UO_327 (O_327,N_2934,N_2994);
nand UO_328 (O_328,N_2509,N_2770);
nor UO_329 (O_329,N_2717,N_2538);
nor UO_330 (O_330,N_2270,N_2676);
or UO_331 (O_331,N_2362,N_2383);
nand UO_332 (O_332,N_2348,N_2808);
nor UO_333 (O_333,N_2931,N_2042);
nor UO_334 (O_334,N_2448,N_2891);
nor UO_335 (O_335,N_2828,N_2514);
nand UO_336 (O_336,N_2716,N_2893);
nand UO_337 (O_337,N_2108,N_2245);
nand UO_338 (O_338,N_2473,N_2690);
xor UO_339 (O_339,N_2700,N_2301);
and UO_340 (O_340,N_2521,N_2915);
or UO_341 (O_341,N_2121,N_2366);
and UO_342 (O_342,N_2085,N_2783);
nor UO_343 (O_343,N_2895,N_2537);
nand UO_344 (O_344,N_2818,N_2390);
or UO_345 (O_345,N_2657,N_2184);
and UO_346 (O_346,N_2673,N_2004);
and UO_347 (O_347,N_2864,N_2961);
or UO_348 (O_348,N_2015,N_2582);
nand UO_349 (O_349,N_2224,N_2465);
and UO_350 (O_350,N_2522,N_2918);
and UO_351 (O_351,N_2195,N_2821);
or UO_352 (O_352,N_2303,N_2746);
nor UO_353 (O_353,N_2286,N_2202);
nand UO_354 (O_354,N_2012,N_2780);
nand UO_355 (O_355,N_2343,N_2114);
nor UO_356 (O_356,N_2692,N_2201);
nor UO_357 (O_357,N_2375,N_2663);
or UO_358 (O_358,N_2732,N_2674);
nor UO_359 (O_359,N_2848,N_2950);
or UO_360 (O_360,N_2591,N_2643);
or UO_361 (O_361,N_2960,N_2142);
nor UO_362 (O_362,N_2622,N_2090);
nand UO_363 (O_363,N_2381,N_2367);
or UO_364 (O_364,N_2683,N_2217);
nor UO_365 (O_365,N_2105,N_2147);
nand UO_366 (O_366,N_2039,N_2672);
nand UO_367 (O_367,N_2568,N_2619);
nor UO_368 (O_368,N_2033,N_2656);
nor UO_369 (O_369,N_2630,N_2498);
nor UO_370 (O_370,N_2269,N_2635);
or UO_371 (O_371,N_2801,N_2338);
or UO_372 (O_372,N_2138,N_2466);
or UO_373 (O_373,N_2128,N_2884);
or UO_374 (O_374,N_2254,N_2650);
nor UO_375 (O_375,N_2916,N_2289);
and UO_376 (O_376,N_2854,N_2881);
nor UO_377 (O_377,N_2174,N_2148);
nand UO_378 (O_378,N_2660,N_2436);
nor UO_379 (O_379,N_2152,N_2979);
or UO_380 (O_380,N_2485,N_2540);
and UO_381 (O_381,N_2805,N_2724);
nand UO_382 (O_382,N_2461,N_2234);
and UO_383 (O_383,N_2490,N_2667);
or UO_384 (O_384,N_2172,N_2295);
or UO_385 (O_385,N_2525,N_2866);
nand UO_386 (O_386,N_2865,N_2102);
nand UO_387 (O_387,N_2319,N_2474);
nor UO_388 (O_388,N_2578,N_2307);
and UO_389 (O_389,N_2946,N_2587);
and UO_390 (O_390,N_2539,N_2922);
nor UO_391 (O_391,N_2265,N_2021);
nor UO_392 (O_392,N_2943,N_2156);
or UO_393 (O_393,N_2400,N_2554);
nor UO_394 (O_394,N_2379,N_2763);
nor UO_395 (O_395,N_2181,N_2458);
or UO_396 (O_396,N_2377,N_2116);
or UO_397 (O_397,N_2678,N_2274);
xnor UO_398 (O_398,N_2111,N_2819);
and UO_399 (O_399,N_2293,N_2043);
or UO_400 (O_400,N_2435,N_2662);
nor UO_401 (O_401,N_2562,N_2957);
or UO_402 (O_402,N_2212,N_2194);
nand UO_403 (O_403,N_2889,N_2420);
nand UO_404 (O_404,N_2614,N_2145);
xnor UO_405 (O_405,N_2830,N_2361);
nand UO_406 (O_406,N_2939,N_2984);
or UO_407 (O_407,N_2944,N_2190);
nand UO_408 (O_408,N_2668,N_2199);
and UO_409 (O_409,N_2870,N_2235);
xor UO_410 (O_410,N_2536,N_2837);
and UO_411 (O_411,N_2277,N_2456);
or UO_412 (O_412,N_2239,N_2028);
nor UO_413 (O_413,N_2697,N_2875);
nor UO_414 (O_414,N_2167,N_2356);
and UO_415 (O_415,N_2933,N_2279);
nor UO_416 (O_416,N_2467,N_2727);
or UO_417 (O_417,N_2023,N_2288);
nand UO_418 (O_418,N_2748,N_2992);
or UO_419 (O_419,N_2132,N_2009);
and UO_420 (O_420,N_2758,N_2263);
nand UO_421 (O_421,N_2721,N_2297);
and UO_422 (O_422,N_2007,N_2570);
and UO_423 (O_423,N_2054,N_2680);
or UO_424 (O_424,N_2602,N_2508);
or UO_425 (O_425,N_2876,N_2241);
and UO_426 (O_426,N_2510,N_2044);
or UO_427 (O_427,N_2857,N_2040);
or UO_428 (O_428,N_2775,N_2740);
or UO_429 (O_429,N_2020,N_2913);
or UO_430 (O_430,N_2117,N_2433);
xnor UO_431 (O_431,N_2517,N_2211);
and UO_432 (O_432,N_2339,N_2710);
nor UO_433 (O_433,N_2096,N_2276);
nand UO_434 (O_434,N_2232,N_2964);
nor UO_435 (O_435,N_2923,N_2902);
nand UO_436 (O_436,N_2098,N_2701);
nor UO_437 (O_437,N_2707,N_2610);
nand UO_438 (O_438,N_2605,N_2408);
nor UO_439 (O_439,N_2972,N_2789);
or UO_440 (O_440,N_2080,N_2955);
or UO_441 (O_441,N_2419,N_2271);
and UO_442 (O_442,N_2061,N_2742);
and UO_443 (O_443,N_2633,N_2513);
xnor UO_444 (O_444,N_2579,N_2483);
and UO_445 (O_445,N_2418,N_2720);
and UO_446 (O_446,N_2689,N_2975);
or UO_447 (O_447,N_2547,N_2310);
and UO_448 (O_448,N_2282,N_2330);
nand UO_449 (O_449,N_2575,N_2569);
and UO_450 (O_450,N_2928,N_2623);
and UO_451 (O_451,N_2988,N_2369);
or UO_452 (O_452,N_2292,N_2765);
nand UO_453 (O_453,N_2896,N_2774);
and UO_454 (O_454,N_2906,N_2060);
nand UO_455 (O_455,N_2355,N_2353);
and UO_456 (O_456,N_2877,N_2849);
or UO_457 (O_457,N_2088,N_2242);
and UO_458 (O_458,N_2493,N_2535);
nor UO_459 (O_459,N_2936,N_2107);
nor UO_460 (O_460,N_2580,N_2488);
nand UO_461 (O_461,N_2417,N_2248);
nand UO_462 (O_462,N_2947,N_2357);
nor UO_463 (O_463,N_2431,N_2005);
nand UO_464 (O_464,N_2963,N_2983);
nand UO_465 (O_465,N_2103,N_2109);
nor UO_466 (O_466,N_2257,N_2322);
nand UO_467 (O_467,N_2300,N_2886);
nand UO_468 (O_468,N_2311,N_2426);
and UO_469 (O_469,N_2446,N_2863);
and UO_470 (O_470,N_2597,N_2326);
and UO_471 (O_471,N_2129,N_2273);
or UO_472 (O_472,N_2725,N_2755);
and UO_473 (O_473,N_2470,N_2910);
nor UO_474 (O_474,N_2813,N_2729);
nand UO_475 (O_475,N_2491,N_2442);
or UO_476 (O_476,N_2481,N_2204);
nor UO_477 (O_477,N_2168,N_2336);
and UO_478 (O_478,N_2206,N_2824);
nand UO_479 (O_479,N_2646,N_2699);
or UO_480 (O_480,N_2425,N_2169);
or UO_481 (O_481,N_2314,N_2892);
nand UO_482 (O_482,N_2598,N_2087);
xnor UO_483 (O_483,N_2997,N_2186);
nor UO_484 (O_484,N_2833,N_2146);
or UO_485 (O_485,N_2702,N_2048);
nand UO_486 (O_486,N_2220,N_2615);
nor UO_487 (O_487,N_2573,N_2705);
nand UO_488 (O_488,N_2791,N_2584);
nor UO_489 (O_489,N_2131,N_2219);
nor UO_490 (O_490,N_2226,N_2583);
nor UO_491 (O_491,N_2733,N_2402);
or UO_492 (O_492,N_2901,N_2816);
nand UO_493 (O_493,N_2894,N_2661);
and UO_494 (O_494,N_2447,N_2706);
and UO_495 (O_495,N_2814,N_2644);
and UO_496 (O_496,N_2130,N_2342);
or UO_497 (O_497,N_2159,N_2365);
nand UO_498 (O_498,N_2350,N_2815);
nand UO_499 (O_499,N_2826,N_2329);
endmodule