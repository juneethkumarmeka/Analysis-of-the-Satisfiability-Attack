module basic_3000_30000_3500_15_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_275,In_2613);
nor U1 (N_1,In_1466,In_1853);
and U2 (N_2,In_2473,In_2718);
or U3 (N_3,In_1983,In_38);
nand U4 (N_4,In_2382,In_466);
and U5 (N_5,In_1499,In_2364);
nor U6 (N_6,In_489,In_91);
nor U7 (N_7,In_930,In_727);
xnor U8 (N_8,In_1911,In_2018);
and U9 (N_9,In_2618,In_2808);
or U10 (N_10,In_995,In_2164);
nand U11 (N_11,In_342,In_2506);
nand U12 (N_12,In_2038,In_1559);
or U13 (N_13,In_1461,In_382);
or U14 (N_14,In_1228,In_1120);
and U15 (N_15,In_539,In_532);
nand U16 (N_16,In_1431,In_2475);
and U17 (N_17,In_1832,In_1063);
nand U18 (N_18,In_124,In_343);
and U19 (N_19,In_93,In_1552);
or U20 (N_20,In_1535,In_1523);
nand U21 (N_21,In_2641,In_1369);
nand U22 (N_22,In_2723,In_1644);
nand U23 (N_23,In_156,In_1432);
nand U24 (N_24,In_265,In_2092);
and U25 (N_25,In_2585,In_1414);
xnor U26 (N_26,In_2600,In_242);
xnor U27 (N_27,In_26,In_556);
and U28 (N_28,In_615,In_1815);
nor U29 (N_29,In_1511,In_2591);
xnor U30 (N_30,In_1954,In_2301);
and U31 (N_31,In_731,In_2058);
and U32 (N_32,In_1390,In_2885);
and U33 (N_33,In_1491,In_1699);
and U34 (N_34,In_231,In_1546);
nor U35 (N_35,In_892,In_2537);
nand U36 (N_36,In_243,In_1157);
xnor U37 (N_37,In_1140,In_1805);
nor U38 (N_38,In_168,In_1557);
xnor U39 (N_39,In_2967,In_1870);
or U40 (N_40,In_1335,In_932);
nand U41 (N_41,In_2865,In_898);
and U42 (N_42,In_2539,In_1366);
or U43 (N_43,In_2035,In_1530);
xnor U44 (N_44,In_349,In_2479);
or U45 (N_45,In_1964,In_1517);
xnor U46 (N_46,In_288,In_2961);
nor U47 (N_47,In_625,In_810);
and U48 (N_48,In_1881,In_2330);
xor U49 (N_49,In_1967,In_1018);
nand U50 (N_50,In_1476,In_1939);
or U51 (N_51,In_2208,In_822);
nand U52 (N_52,In_1277,In_1163);
nand U53 (N_53,In_2989,In_1380);
and U54 (N_54,In_1534,In_2448);
or U55 (N_55,In_1438,In_818);
nand U56 (N_56,In_1575,In_1802);
nand U57 (N_57,In_1412,In_1860);
nand U58 (N_58,In_295,In_2528);
or U59 (N_59,In_2168,In_1493);
xor U60 (N_60,In_1705,In_2965);
or U61 (N_61,In_2226,In_618);
and U62 (N_62,In_1444,In_2238);
nor U63 (N_63,In_2548,In_1236);
xor U64 (N_64,In_2428,In_125);
nand U65 (N_65,In_2958,In_1145);
nand U66 (N_66,In_1673,In_209);
and U67 (N_67,In_1314,In_2001);
or U68 (N_68,In_1914,In_1706);
nor U69 (N_69,In_2187,In_184);
or U70 (N_70,In_767,In_2145);
xor U71 (N_71,In_1868,In_505);
or U72 (N_72,In_1008,In_993);
or U73 (N_73,In_198,In_167);
and U74 (N_74,In_2328,In_1113);
and U75 (N_75,In_989,In_1184);
nand U76 (N_76,In_1689,In_2653);
nand U77 (N_77,In_2622,In_2635);
or U78 (N_78,In_494,In_1325);
and U79 (N_79,In_746,In_979);
or U80 (N_80,In_1152,In_481);
nor U81 (N_81,In_2420,In_1264);
or U82 (N_82,In_1251,In_2552);
nor U83 (N_83,In_190,In_2609);
and U84 (N_84,In_2686,In_1115);
and U85 (N_85,In_1410,In_2034);
or U86 (N_86,In_375,In_208);
nand U87 (N_87,In_1179,In_2280);
xnor U88 (N_88,In_109,In_814);
and U89 (N_89,In_2688,In_131);
and U90 (N_90,In_1521,In_204);
xnor U91 (N_91,In_1210,In_1604);
and U92 (N_92,In_35,In_2469);
nand U93 (N_93,In_606,In_1199);
or U94 (N_94,In_1896,In_316);
or U95 (N_95,In_497,In_380);
nand U96 (N_96,In_1985,In_1555);
or U97 (N_97,In_1350,In_1060);
and U98 (N_98,In_74,In_1282);
and U99 (N_99,In_1002,In_1048);
or U100 (N_100,In_94,In_1978);
or U101 (N_101,In_2628,In_2927);
nor U102 (N_102,In_2317,In_703);
nand U103 (N_103,In_122,In_2266);
nor U104 (N_104,In_2336,In_2606);
xor U105 (N_105,In_117,In_2824);
xnor U106 (N_106,In_370,In_2042);
xor U107 (N_107,In_258,In_2495);
nor U108 (N_108,In_1701,In_736);
nand U109 (N_109,In_2302,In_2826);
or U110 (N_110,In_1351,In_1176);
nor U111 (N_111,In_1908,In_2397);
or U112 (N_112,In_1938,In_1255);
nand U113 (N_113,In_2359,In_905);
and U114 (N_114,In_2371,In_2561);
nand U115 (N_115,In_2276,In_2571);
nand U116 (N_116,In_2039,In_1836);
nand U117 (N_117,In_2963,In_2436);
xnor U118 (N_118,In_688,In_2883);
nand U119 (N_119,In_398,In_732);
and U120 (N_120,In_2005,In_127);
xnor U121 (N_121,In_2200,In_2781);
and U122 (N_122,In_2647,In_1993);
or U123 (N_123,In_1769,In_547);
xor U124 (N_124,In_2547,In_1398);
and U125 (N_125,In_1422,In_1258);
nor U126 (N_126,In_613,In_812);
and U127 (N_127,In_1206,In_635);
nand U128 (N_128,In_1666,In_347);
nor U129 (N_129,In_366,In_270);
or U130 (N_130,In_2771,In_2312);
nand U131 (N_131,In_2261,In_3);
nand U132 (N_132,In_813,In_1569);
nand U133 (N_133,In_1791,In_2210);
xor U134 (N_134,In_1672,In_1416);
nor U135 (N_135,In_796,In_1084);
nor U136 (N_136,In_874,In_217);
nor U137 (N_137,In_1065,In_459);
nor U138 (N_138,In_403,In_1471);
and U139 (N_139,In_1687,In_730);
xnor U140 (N_140,In_212,In_2136);
or U141 (N_141,In_619,In_2057);
xor U142 (N_142,In_227,In_571);
and U143 (N_143,In_1167,In_206);
and U144 (N_144,In_25,In_116);
or U145 (N_145,In_1134,In_636);
or U146 (N_146,In_662,In_2017);
xnor U147 (N_147,In_1625,In_901);
and U148 (N_148,In_2942,In_2244);
nor U149 (N_149,In_2480,In_440);
or U150 (N_150,In_684,In_2709);
nor U151 (N_151,In_842,In_58);
nor U152 (N_152,In_2365,In_1252);
and U153 (N_153,In_568,In_2775);
nand U154 (N_154,In_2434,In_1148);
or U155 (N_155,In_2088,In_2912);
nand U156 (N_156,In_1032,In_2992);
nor U157 (N_157,In_737,In_165);
nor U158 (N_158,In_2798,In_724);
nor U159 (N_159,In_1234,In_1405);
and U160 (N_160,In_520,In_2109);
and U161 (N_161,In_423,In_2619);
nand U162 (N_162,In_2309,In_100);
nor U163 (N_163,In_541,In_2268);
and U164 (N_164,In_783,In_542);
nand U165 (N_165,In_1283,In_2075);
nor U166 (N_166,In_789,In_298);
nor U167 (N_167,In_2701,In_1972);
and U168 (N_168,In_2118,In_965);
xnor U169 (N_169,In_2329,In_2660);
nor U170 (N_170,In_988,In_1332);
xor U171 (N_171,In_1391,In_790);
and U172 (N_172,In_279,In_2796);
nor U173 (N_173,In_907,In_1834);
nand U174 (N_174,In_2730,In_560);
xor U175 (N_175,In_2513,In_255);
nor U176 (N_176,In_1962,In_1664);
xor U177 (N_177,In_1987,In_1010);
nor U178 (N_178,In_691,In_2489);
nand U179 (N_179,In_2735,In_2866);
and U180 (N_180,In_960,In_2441);
xnor U181 (N_181,In_1652,In_2300);
xor U182 (N_182,In_2435,In_845);
and U183 (N_183,In_630,In_611);
nor U184 (N_184,In_978,In_2472);
nand U185 (N_185,In_1633,In_154);
and U186 (N_186,In_982,In_2158);
nand U187 (N_187,In_2897,In_1323);
nand U188 (N_188,In_2229,In_1848);
or U189 (N_189,In_340,In_1294);
nand U190 (N_190,In_2380,In_1615);
or U191 (N_191,In_777,In_2454);
or U192 (N_192,In_155,In_1272);
nor U193 (N_193,In_1154,In_2054);
nand U194 (N_194,In_2684,In_2629);
nor U195 (N_195,In_1921,In_2102);
nor U196 (N_196,In_706,In_1551);
and U197 (N_197,In_1957,In_1916);
or U198 (N_198,In_887,In_1614);
and U199 (N_199,In_142,In_453);
or U200 (N_200,In_2283,In_386);
xor U201 (N_201,In_2952,In_1337);
and U202 (N_202,In_163,In_1027);
or U203 (N_203,In_2209,In_2633);
nand U204 (N_204,In_1336,In_1450);
nor U205 (N_205,In_917,In_135);
nor U206 (N_206,In_2199,In_1150);
and U207 (N_207,In_1433,In_402);
or U208 (N_208,In_508,In_2922);
and U209 (N_209,In_1707,In_2886);
and U210 (N_210,In_2903,In_1621);
or U211 (N_211,In_756,In_2127);
and U212 (N_212,In_2758,In_1235);
xor U213 (N_213,In_2322,In_2294);
nor U214 (N_214,In_2937,In_2800);
nand U215 (N_215,In_2707,In_1694);
or U216 (N_216,In_2962,In_387);
nand U217 (N_217,In_2498,In_1315);
and U218 (N_218,In_1822,In_1959);
xor U219 (N_219,In_608,In_19);
or U220 (N_220,In_695,In_792);
or U221 (N_221,In_1028,In_1772);
nor U222 (N_222,In_1188,In_2742);
and U223 (N_223,In_958,In_60);
nor U224 (N_224,In_1801,In_2125);
and U225 (N_225,In_1509,In_871);
and U226 (N_226,In_2426,In_945);
nand U227 (N_227,In_1322,In_1719);
nand U228 (N_228,In_1232,In_772);
and U229 (N_229,In_59,In_660);
nor U230 (N_230,In_2368,In_2066);
nand U231 (N_231,In_1216,In_1500);
xor U232 (N_232,In_2748,In_1117);
nand U233 (N_233,In_1395,In_2504);
xnor U234 (N_234,In_1762,In_563);
xor U235 (N_235,In_604,In_677);
and U236 (N_236,In_798,In_1670);
nand U237 (N_237,In_450,In_2692);
nor U238 (N_238,In_2214,In_322);
and U239 (N_239,In_72,In_1955);
and U240 (N_240,In_1371,In_476);
and U241 (N_241,In_763,In_43);
or U242 (N_242,In_499,In_2047);
nand U243 (N_243,In_1718,In_2750);
nand U244 (N_244,In_856,In_1892);
or U245 (N_245,In_2247,In_944);
or U246 (N_246,In_614,In_1420);
nor U247 (N_247,In_2415,In_880);
nor U248 (N_248,In_913,In_638);
nor U249 (N_249,In_2496,In_236);
nand U250 (N_250,In_2411,In_2588);
xor U251 (N_251,In_729,In_2710);
nand U252 (N_252,In_1217,In_1312);
nand U253 (N_253,In_1190,In_651);
and U254 (N_254,In_1810,In_1947);
or U255 (N_255,In_264,In_2632);
nand U256 (N_256,In_916,In_1483);
nand U257 (N_257,In_2806,In_2011);
nor U258 (N_258,In_2778,In_975);
nand U259 (N_259,In_1160,In_1880);
nand U260 (N_260,In_2273,In_2663);
and U261 (N_261,In_983,In_2315);
and U262 (N_262,In_1442,In_2418);
or U263 (N_263,In_2325,In_2687);
xor U264 (N_264,In_1510,In_1781);
nand U265 (N_265,In_230,In_1934);
or U266 (N_266,In_862,In_362);
and U267 (N_267,In_1992,In_2578);
nand U268 (N_268,In_1948,In_2837);
nor U269 (N_269,In_237,In_2141);
nand U270 (N_270,In_2652,In_1013);
or U271 (N_271,In_866,In_582);
xor U272 (N_272,In_1630,In_238);
and U273 (N_273,In_705,In_1333);
nor U274 (N_274,In_311,In_553);
or U275 (N_275,In_2811,In_1503);
and U276 (N_276,In_2012,In_2427);
and U277 (N_277,In_1421,In_1624);
xnor U278 (N_278,In_115,In_1368);
xor U279 (N_279,In_882,In_2461);
and U280 (N_280,In_1393,In_2049);
or U281 (N_281,In_1164,In_417);
nand U282 (N_282,In_617,In_222);
nand U283 (N_283,In_2178,In_2637);
nand U284 (N_284,In_1982,In_1392);
xor U285 (N_285,In_2417,In_2554);
or U286 (N_286,In_1172,In_2754);
and U287 (N_287,In_782,In_876);
or U288 (N_288,In_1094,In_2706);
nor U289 (N_289,In_2941,In_503);
nor U290 (N_290,In_2094,In_1976);
nand U291 (N_291,In_628,In_1399);
or U292 (N_292,In_2212,In_1838);
nor U293 (N_293,In_1589,In_955);
nand U294 (N_294,In_864,In_1676);
nand U295 (N_295,In_2977,In_2916);
nor U296 (N_296,In_973,In_1149);
and U297 (N_297,In_827,In_2577);
nor U298 (N_298,In_1806,In_2804);
xnor U299 (N_299,In_1564,In_1394);
nand U300 (N_300,In_1794,In_1775);
or U301 (N_301,In_418,In_1161);
or U302 (N_302,In_840,In_2373);
or U303 (N_303,In_2231,In_123);
nand U304 (N_304,In_633,In_2077);
or U305 (N_305,In_2998,In_1946);
or U306 (N_306,In_2825,In_1998);
nand U307 (N_307,In_1891,In_2326);
or U308 (N_308,In_2829,In_2849);
and U309 (N_309,In_1229,In_306);
nand U310 (N_310,In_2101,In_2990);
nor U311 (N_311,In_2589,In_1515);
or U312 (N_312,In_1137,In_1847);
and U313 (N_313,In_1735,In_974);
nor U314 (N_314,In_855,In_1658);
xnor U315 (N_315,In_2953,In_1484);
and U316 (N_316,In_1764,In_2549);
nand U317 (N_317,In_88,In_787);
and U318 (N_318,In_740,In_581);
xnor U319 (N_319,In_1598,In_1403);
and U320 (N_320,In_2003,In_2242);
xnor U321 (N_321,In_1721,In_1606);
xnor U322 (N_322,In_750,In_1078);
or U323 (N_323,In_873,In_1005);
and U324 (N_324,In_332,In_809);
or U325 (N_325,In_171,In_755);
and U326 (N_326,In_574,In_2465);
nand U327 (N_327,In_2911,In_793);
xor U328 (N_328,In_526,In_1133);
or U329 (N_329,In_1844,In_1712);
xnor U330 (N_330,In_1182,In_1003);
and U331 (N_331,In_1423,In_176);
and U332 (N_332,In_90,In_2753);
nand U333 (N_333,In_2521,In_867);
and U334 (N_334,In_788,In_507);
nor U335 (N_335,In_943,In_2031);
nor U336 (N_336,In_2525,In_961);
and U337 (N_337,In_2909,In_779);
nor U338 (N_338,In_1061,In_1873);
xor U339 (N_339,In_98,In_1103);
nand U340 (N_340,In_1994,In_600);
or U341 (N_341,In_2410,In_641);
or U342 (N_342,In_1922,In_1131);
nand U343 (N_343,In_2560,In_111);
or U344 (N_344,In_2651,In_2491);
nand U345 (N_345,In_2982,In_1863);
or U346 (N_346,In_2366,In_971);
nor U347 (N_347,In_1045,In_591);
nand U348 (N_348,In_1024,In_2728);
nand U349 (N_349,In_2112,In_1498);
or U350 (N_350,In_969,In_1726);
xnor U351 (N_351,In_2786,In_406);
or U352 (N_352,In_643,In_513);
and U353 (N_353,In_519,In_2146);
nand U354 (N_354,In_1969,In_1119);
and U355 (N_355,In_1945,In_2000);
xnor U356 (N_356,In_447,In_1330);
nor U357 (N_357,In_336,In_1106);
nand U358 (N_358,In_2345,In_733);
xor U359 (N_359,In_1296,In_420);
xnor U360 (N_360,In_2683,In_2267);
and U361 (N_361,In_592,In_1396);
nand U362 (N_362,In_1226,In_1238);
nor U363 (N_363,In_2216,In_1663);
and U364 (N_364,In_860,In_2111);
nand U365 (N_365,In_1354,In_1617);
xnor U366 (N_366,In_1248,In_1902);
nor U367 (N_367,In_1924,In_2822);
or U368 (N_368,In_2123,In_2691);
and U369 (N_369,In_551,In_2648);
and U370 (N_370,In_1843,In_252);
xor U371 (N_371,In_1588,In_689);
nand U372 (N_372,In_909,In_2955);
nand U373 (N_373,In_1744,In_2139);
and U374 (N_374,In_2620,In_2621);
nor U375 (N_375,In_39,In_1827);
nor U376 (N_376,In_250,In_2021);
nor U377 (N_377,In_931,In_2713);
and U378 (N_378,In_2579,In_2828);
nor U379 (N_379,In_2232,In_835);
xor U380 (N_380,In_1629,In_2788);
and U381 (N_381,In_1619,In_1729);
nor U382 (N_382,In_1977,In_739);
and U383 (N_383,In_259,In_1428);
or U384 (N_384,In_1686,In_1300);
nand U385 (N_385,In_1064,In_2458);
or U386 (N_386,In_2243,In_108);
nand U387 (N_387,In_884,In_2236);
nand U388 (N_388,In_565,In_947);
or U389 (N_389,In_2198,In_1090);
and U390 (N_390,In_990,In_2281);
and U391 (N_391,In_1014,In_2874);
nand U392 (N_392,In_218,In_6);
nor U393 (N_393,In_1109,In_2383);
or U394 (N_394,In_1912,In_2063);
nor U395 (N_395,In_2680,In_698);
xnor U396 (N_396,In_493,In_1372);
nor U397 (N_397,In_324,In_1730);
nand U398 (N_398,In_1571,In_1377);
nand U399 (N_399,In_105,In_2219);
nor U400 (N_400,In_1166,In_2779);
xor U401 (N_401,In_1927,In_1054);
or U402 (N_402,In_1143,In_1849);
nor U403 (N_403,In_2557,In_201);
nor U404 (N_404,In_959,In_500);
and U405 (N_405,In_2037,In_2741);
and U406 (N_406,In_52,In_1752);
and U407 (N_407,In_1773,In_1820);
and U408 (N_408,In_1884,In_1050);
nand U409 (N_409,In_999,In_2274);
xor U410 (N_410,In_310,In_427);
xnor U411 (N_411,In_2801,In_69);
or U412 (N_412,In_1683,In_1577);
nand U413 (N_413,In_2234,In_1807);
and U414 (N_414,In_1518,In_954);
nand U415 (N_415,In_436,In_1460);
nor U416 (N_416,In_197,In_1855);
or U417 (N_417,In_266,In_1488);
and U418 (N_418,In_1841,In_1288);
or U419 (N_419,In_483,In_457);
nor U420 (N_420,In_1244,In_388);
or U421 (N_421,In_2685,In_2681);
xnor U422 (N_422,In_2022,In_1128);
or U423 (N_423,In_2013,In_806);
and U424 (N_424,In_747,In_2869);
or U425 (N_425,In_1837,In_2910);
and U426 (N_426,In_2207,In_2627);
or U427 (N_427,In_1859,In_102);
or U428 (N_428,In_2655,In_583);
and U429 (N_429,In_173,In_2133);
nand U430 (N_430,In_555,In_1803);
nand U431 (N_431,In_1611,In_1426);
nor U432 (N_432,In_369,In_1814);
or U433 (N_433,In_2367,In_1237);
xnor U434 (N_434,In_2477,In_1795);
xnor U435 (N_435,In_1748,In_2716);
nor U436 (N_436,In_2708,In_711);
and U437 (N_437,In_346,In_1742);
and U438 (N_438,In_1130,In_1816);
and U439 (N_439,In_929,In_2898);
or U440 (N_440,In_1440,In_1345);
xnor U441 (N_441,In_2277,In_334);
xnor U442 (N_442,In_1544,In_2605);
nand U443 (N_443,In_535,In_998);
nand U444 (N_444,In_2319,In_1828);
nor U445 (N_445,In_1029,In_2090);
or U446 (N_446,In_1081,In_1451);
and U447 (N_447,In_811,In_1305);
xor U448 (N_448,In_1276,In_649);
nor U449 (N_449,In_1035,In_404);
nand U450 (N_450,In_1638,In_1751);
xor U451 (N_451,In_938,In_421);
or U452 (N_452,In_1623,In_922);
nor U453 (N_453,In_804,In_401);
nor U454 (N_454,In_2803,In_771);
or U455 (N_455,In_2271,In_2926);
nor U456 (N_456,In_2508,In_2442);
nor U457 (N_457,In_199,In_2346);
nor U458 (N_458,In_2356,In_1041);
nand U459 (N_459,In_213,In_2470);
or U460 (N_460,In_1262,In_1684);
xnor U461 (N_461,In_1071,In_1311);
or U462 (N_462,In_1620,In_1733);
and U463 (N_463,In_1558,In_2630);
nand U464 (N_464,In_1317,In_1243);
or U465 (N_465,In_2126,In_1562);
nand U466 (N_466,In_368,In_1334);
xor U467 (N_467,In_1455,In_2205);
xnor U468 (N_468,In_655,In_2340);
nand U469 (N_469,In_2550,In_2440);
and U470 (N_470,In_963,In_1904);
and U471 (N_471,In_1485,In_540);
nor U472 (N_472,In_521,In_348);
xnor U473 (N_473,In_2119,In_2048);
or U474 (N_474,In_87,In_1654);
nor U475 (N_475,In_2726,In_1462);
nand U476 (N_476,In_1383,In_2355);
nand U477 (N_477,In_1241,In_1755);
xor U478 (N_478,In_2339,In_2884);
nand U479 (N_479,In_2201,In_2064);
and U480 (N_480,In_220,In_128);
or U481 (N_481,In_95,In_865);
nor U482 (N_482,In_1636,In_1637);
nor U483 (N_483,In_2848,In_546);
nor U484 (N_484,In_2838,In_99);
and U485 (N_485,In_2695,In_2098);
xnor U486 (N_486,In_1030,In_1640);
xnor U487 (N_487,In_1796,In_2956);
nand U488 (N_488,In_2240,In_354);
nor U489 (N_489,In_699,In_396);
nand U490 (N_490,In_1917,In_632);
xnor U491 (N_491,In_674,In_422);
and U492 (N_492,In_743,In_723);
and U493 (N_493,In_437,In_2156);
or U494 (N_494,In_1533,In_1496);
nor U495 (N_495,In_2531,In_1308);
nand U496 (N_496,In_2757,In_1971);
or U497 (N_497,In_825,In_326);
xor U498 (N_498,In_2752,In_2700);
and U499 (N_499,In_353,In_2004);
and U500 (N_500,In_2640,In_2751);
or U501 (N_501,In_2067,In_407);
nand U502 (N_502,In_2943,In_2740);
and U503 (N_503,In_803,In_203);
nand U504 (N_504,In_1253,In_1622);
nand U505 (N_505,In_1494,In_223);
or U506 (N_506,In_2358,In_2712);
nor U507 (N_507,In_2780,In_690);
or U508 (N_508,In_1215,In_2152);
and U509 (N_509,In_816,In_2791);
and U510 (N_510,In_2639,In_2499);
nor U511 (N_511,In_829,In_1359);
and U512 (N_512,In_676,In_2790);
and U513 (N_513,In_2835,In_1952);
or U514 (N_514,In_2745,In_2792);
and U515 (N_515,In_2905,In_474);
and U516 (N_516,In_430,In_784);
nor U517 (N_517,In_585,In_2009);
nand U518 (N_518,In_2919,In_1220);
or U519 (N_519,In_531,In_2973);
xor U520 (N_520,In_1291,In_725);
xor U521 (N_521,In_1708,In_11);
xnor U522 (N_522,In_2122,In_1039);
nor U523 (N_523,In_27,In_2690);
nand U524 (N_524,In_2643,In_2245);
nand U525 (N_525,In_2512,In_455);
nor U526 (N_526,In_1249,In_1181);
or U527 (N_527,In_1600,In_159);
and U528 (N_528,In_1200,In_103);
and U529 (N_529,In_1845,In_367);
nand U530 (N_530,In_2052,In_1202);
nor U531 (N_531,In_345,In_2888);
xor U532 (N_532,In_2914,In_2467);
nor U533 (N_533,In_672,In_795);
nor U534 (N_534,In_2625,In_644);
nor U535 (N_535,In_1651,In_2762);
nand U536 (N_536,In_160,In_831);
nor U537 (N_537,In_2719,In_1023);
and U538 (N_538,In_1077,In_152);
and U539 (N_539,In_712,In_658);
and U540 (N_540,In_1561,In_1582);
nand U541 (N_541,In_1105,In_2147);
nand U542 (N_542,In_148,In_534);
nand U543 (N_543,In_2527,In_1739);
or U544 (N_544,In_1087,In_1132);
nand U545 (N_545,In_2149,In_2439);
xnor U546 (N_546,In_325,In_1738);
and U547 (N_547,In_463,In_2642);
nand U548 (N_548,In_1866,In_1818);
nor U549 (N_549,In_2036,In_2871);
or U550 (N_550,In_1716,In_926);
nand U551 (N_551,In_1088,In_2015);
or U552 (N_552,In_434,In_1743);
nor U553 (N_553,In_2255,In_1214);
and U554 (N_554,In_1774,In_2517);
xnor U555 (N_555,In_584,In_149);
xor U556 (N_556,In_2065,In_1247);
xnor U557 (N_557,In_2795,In_802);
xor U558 (N_558,In_941,In_1659);
nand U559 (N_559,In_2014,In_1213);
nand U560 (N_560,In_1901,In_2572);
or U561 (N_561,In_2522,In_2068);
nor U562 (N_562,In_673,In_2733);
xor U563 (N_563,In_1990,In_1324);
xnor U564 (N_564,In_2493,In_1445);
and U565 (N_565,In_219,In_2450);
or U566 (N_566,In_384,In_1618);
nand U567 (N_567,In_1108,In_1400);
or U568 (N_568,In_510,In_225);
xor U569 (N_569,In_41,In_465);
xnor U570 (N_570,In_1591,In_107);
nor U571 (N_571,In_214,In_1340);
nor U572 (N_572,In_158,In_888);
and U573 (N_573,In_1903,In_426);
or U574 (N_574,In_1348,In_315);
and U575 (N_575,In_157,In_56);
or U576 (N_576,In_2755,In_2464);
nand U577 (N_577,In_17,In_1168);
nor U578 (N_578,In_1580,In_2756);
xor U579 (N_579,In_2318,In_564);
nor U580 (N_580,In_2586,In_2842);
xnor U581 (N_581,In_664,In_2468);
nand U582 (N_582,In_1825,In_1867);
and U583 (N_583,In_2715,In_2252);
xnor U584 (N_584,In_2290,In_1449);
or U585 (N_585,In_486,In_589);
and U586 (N_586,In_1026,In_2190);
and U587 (N_587,In_282,In_1956);
nor U588 (N_588,In_449,In_281);
and U589 (N_589,In_1812,In_1425);
xor U590 (N_590,In_2293,In_151);
and U591 (N_591,In_2841,In_2964);
xnor U592 (N_592,In_234,In_1920);
or U593 (N_593,In_1069,In_1464);
and U594 (N_594,In_580,In_2096);
nand U595 (N_595,In_694,In_1532);
nor U596 (N_596,In_2502,In_1852);
nor U597 (N_597,In_692,In_847);
nand U598 (N_598,In_1401,In_1800);
and U599 (N_599,In_1536,In_2381);
and U600 (N_600,In_1685,In_2103);
nand U601 (N_601,In_1541,In_2947);
nand U602 (N_602,In_2614,In_329);
nor U603 (N_603,In_861,In_908);
xnor U604 (N_604,In_2163,In_2406);
and U605 (N_605,In_824,In_2348);
xnor U606 (N_606,In_1473,In_966);
xnor U607 (N_607,In_2104,In_896);
xor U608 (N_608,In_957,In_1968);
and U609 (N_609,In_2697,In_1696);
nor U610 (N_610,In_1389,In_2510);
nand U611 (N_611,In_2230,In_2573);
or U612 (N_612,In_2699,In_333);
xnor U613 (N_613,In_1942,In_1126);
or U614 (N_614,In_893,In_1470);
nor U615 (N_615,In_2921,In_1437);
or U616 (N_616,In_2070,In_1646);
and U617 (N_617,In_1224,In_2556);
or U618 (N_618,In_2845,In_719);
and U619 (N_619,In_48,In_1862);
and U620 (N_620,In_169,In_2353);
or U621 (N_621,In_2466,In_2809);
nand U622 (N_622,In_2672,In_1522);
nand U623 (N_623,In_634,In_1116);
xnor U624 (N_624,In_2818,In_671);
nor U625 (N_625,In_523,In_1907);
nor U626 (N_626,In_579,In_621);
xor U627 (N_627,In_2321,In_1502);
or U628 (N_628,In_137,In_853);
nand U629 (N_629,In_1667,In_1665);
nand U630 (N_630,In_2455,In_1655);
nand U631 (N_631,In_2767,In_2433);
nor U632 (N_632,In_2634,In_745);
nand U633 (N_633,In_1413,In_1169);
nand U634 (N_634,In_764,In_2983);
nor U635 (N_635,In_308,In_2567);
nor U636 (N_636,In_588,In_389);
and U637 (N_637,In_287,In_320);
or U638 (N_638,In_1573,In_1760);
or U639 (N_639,In_1319,In_2966);
or U640 (N_640,In_2783,In_987);
and U641 (N_641,In_277,In_376);
nand U642 (N_642,In_2250,In_543);
nor U643 (N_643,In_2285,In_441);
or U644 (N_644,In_2423,In_1427);
nand U645 (N_645,In_1268,In_841);
nor U646 (N_646,In_1819,In_682);
nor U647 (N_647,In_2043,In_1486);
or U648 (N_648,In_445,In_2694);
and U649 (N_649,In_2773,In_716);
or U650 (N_650,In_709,In_2483);
nand U651 (N_651,In_2564,In_832);
and U652 (N_652,In_2725,In_1572);
nor U653 (N_653,In_2046,In_1287);
and U654 (N_654,In_2148,In_2069);
and U655 (N_655,In_2299,In_2060);
nand U656 (N_656,In_312,In_1886);
and U657 (N_657,In_1543,In_1913);
and U658 (N_658,In_2852,In_2463);
nor U659 (N_659,In_2167,In_1177);
or U660 (N_660,In_289,In_710);
nand U661 (N_661,In_828,In_558);
nor U662 (N_662,In_1074,In_1382);
or U663 (N_663,In_2665,In_327);
and U664 (N_664,In_886,In_1292);
xor U665 (N_665,In_2389,In_2303);
nand U666 (N_666,In_2457,In_2860);
nand U667 (N_667,In_2576,In_2253);
nand U668 (N_668,In_1905,In_2763);
and U669 (N_669,In_2867,In_2137);
xnor U670 (N_670,In_2534,In_2565);
and U671 (N_671,In_2378,In_2823);
nand U672 (N_672,In_972,In_33);
nor U673 (N_673,In_2166,In_1271);
nor U674 (N_674,In_2132,In_2656);
xnor U675 (N_675,In_2662,In_900);
xnor U676 (N_676,In_2093,In_2194);
or U677 (N_677,In_1963,In_2970);
nand U678 (N_678,In_1012,In_1443);
or U679 (N_679,In_2186,In_2227);
or U680 (N_680,In_2175,In_1628);
xor U681 (N_681,In_1653,In_936);
and U682 (N_682,In_529,In_2174);
xor U683 (N_683,In_2872,In_928);
xor U684 (N_684,In_1174,In_350);
nor U685 (N_685,In_780,In_2935);
xnor U686 (N_686,In_1941,In_2334);
or U687 (N_687,In_601,In_2581);
or U688 (N_688,In_890,In_390);
or U689 (N_689,In_1467,In_182);
xnor U690 (N_690,In_2887,In_414);
xor U691 (N_691,In_1402,In_549);
or U692 (N_692,In_1704,In_2453);
nor U693 (N_693,In_70,In_1626);
nor U694 (N_694,In_1194,In_1047);
xor U695 (N_695,In_910,In_2541);
xnor U696 (N_696,In_1711,In_1424);
and U697 (N_697,In_1900,In_488);
or U698 (N_698,In_2176,In_303);
or U699 (N_699,In_1227,In_1925);
nand U700 (N_700,In_2583,In_653);
and U701 (N_701,In_680,In_885);
and U702 (N_702,In_1201,In_2129);
or U703 (N_703,In_335,In_2736);
nand U704 (N_704,In_820,In_2235);
xor U705 (N_705,In_2610,In_962);
nor U706 (N_706,In_101,In_2237);
nand U707 (N_707,In_920,In_1608);
nor U708 (N_708,In_2864,In_1096);
or U709 (N_709,In_1329,In_2396);
or U710 (N_710,In_1736,In_1245);
or U711 (N_711,In_1745,In_1700);
or U712 (N_712,In_1720,In_195);
xnor U713 (N_713,In_268,In_1782);
and U714 (N_714,In_595,In_1656);
nand U715 (N_715,In_2193,In_2414);
nor U716 (N_716,In_645,In_456);
and U717 (N_717,In_2677,In_2932);
or U718 (N_718,In_1547,In_781);
or U719 (N_719,In_2189,In_1731);
xnor U720 (N_720,In_371,In_2645);
and U721 (N_721,In_1456,In_1817);
or U722 (N_722,In_2673,In_1597);
or U723 (N_723,In_912,In_1784);
nor U724 (N_724,In_545,In_2333);
or U725 (N_725,In_1098,In_1404);
nor U726 (N_726,In_1887,In_2777);
xor U727 (N_727,In_848,In_1789);
and U728 (N_728,In_2879,In_216);
nor U729 (N_729,In_1811,In_554);
nand U730 (N_730,In_81,In_2337);
nor U731 (N_731,In_836,In_469);
nand U732 (N_732,In_1387,In_2624);
xor U733 (N_733,In_915,In_1890);
xor U734 (N_734,In_262,In_2363);
xnor U735 (N_735,In_1677,In_1376);
and U736 (N_736,In_552,In_1178);
xor U737 (N_737,In_240,In_187);
nand U738 (N_738,In_330,In_2259);
or U739 (N_739,In_1257,In_1974);
or U740 (N_740,In_1527,In_2079);
nand U741 (N_741,In_229,In_610);
xor U742 (N_742,In_2899,In_1919);
and U743 (N_743,In_1568,In_2558);
and U744 (N_744,In_2855,In_1052);
and U745 (N_745,In_749,In_1980);
nand U746 (N_746,In_174,In_2844);
nor U747 (N_747,In_2287,In_2459);
nor U748 (N_748,In_2617,In_323);
xnor U749 (N_749,In_433,In_2987);
nor U750 (N_750,In_2975,In_2814);
nor U751 (N_751,In_1453,In_2304);
nor U752 (N_752,In_86,In_538);
and U753 (N_753,In_2379,In_949);
nor U754 (N_754,In_2344,In_2893);
xor U755 (N_755,In_2915,In_1865);
nor U756 (N_756,In_629,In_761);
xnor U757 (N_757,In_14,In_191);
nand U758 (N_758,In_741,In_1009);
xnor U759 (N_759,In_1218,In_1487);
xnor U760 (N_760,In_294,In_2802);
and U761 (N_761,In_527,In_1639);
nand U762 (N_762,In_2785,In_2968);
nor U763 (N_763,In_1793,In_133);
nor U764 (N_764,In_1,In_2398);
xnor U765 (N_765,In_713,In_2960);
or U766 (N_766,In_717,In_2593);
and U767 (N_767,In_2408,In_2233);
xor U768 (N_768,In_2374,In_2995);
or U769 (N_769,In_1538,In_1930);
nor U770 (N_770,In_2492,In_1407);
or U771 (N_771,In_1070,In_1254);
or U772 (N_772,In_113,In_1507);
nand U773 (N_773,In_192,In_1821);
nand U774 (N_774,In_2760,In_869);
or U775 (N_775,In_2041,In_1349);
or U776 (N_776,In_626,In_55);
xnor U777 (N_777,In_839,In_624);
nor U778 (N_778,In_830,In_490);
xor U779 (N_779,In_405,In_1221);
or U780 (N_780,In_2437,In_2896);
and U781 (N_781,In_859,In_2429);
nand U782 (N_782,In_2292,In_134);
xor U783 (N_783,In_1632,In_1358);
nor U784 (N_784,In_2223,In_1352);
xnor U785 (N_785,In_188,In_2530);
nor U786 (N_786,In_1570,In_1091);
xnor U787 (N_787,In_2296,In_1741);
nor U788 (N_788,In_1187,In_2650);
nor U789 (N_789,In_1940,In_1153);
or U790 (N_790,In_504,In_2646);
xnor U791 (N_791,In_1208,In_251);
nand U792 (N_792,In_515,In_2717);
nand U793 (N_793,In_1767,In_374);
nand U794 (N_794,In_2608,In_2305);
or U795 (N_795,In_964,In_1550);
or U796 (N_796,In_877,In_940);
or U797 (N_797,In_309,In_1780);
nor U798 (N_798,In_1702,In_2386);
nand U799 (N_799,In_1642,In_1100);
xnor U800 (N_800,In_1313,In_71);
nor U801 (N_801,In_2264,In_2769);
nor U802 (N_802,In_2228,In_2907);
nor U803 (N_803,In_919,In_2721);
and U804 (N_804,In_968,In_10);
or U805 (N_805,In_1989,In_1454);
xnor U806 (N_806,In_2615,In_57);
xnor U807 (N_807,In_2485,In_1102);
nand U808 (N_808,In_1233,In_2511);
nand U809 (N_809,In_1492,In_84);
and U810 (N_810,In_1409,In_1339);
or U811 (N_811,In_2091,In_2597);
nand U812 (N_812,In_2851,In_1378);
nand U813 (N_813,In_2759,In_1468);
or U814 (N_814,In_2073,In_2768);
xnor U815 (N_815,In_2574,In_762);
nor U816 (N_816,In_2114,In_2100);
nand U817 (N_817,In_304,In_2611);
xor U818 (N_818,In_1542,In_2850);
xor U819 (N_819,In_977,In_2996);
or U820 (N_820,In_2523,In_1709);
or U821 (N_821,In_2460,In_2890);
nor U822 (N_822,In_1960,In_734);
and U823 (N_823,In_2269,In_952);
nor U824 (N_824,In_1475,In_177);
and U825 (N_825,In_2028,In_1146);
nand U826 (N_826,In_2599,In_2362);
nor U827 (N_827,In_110,In_2197);
nor U828 (N_828,In_2976,In_1321);
and U829 (N_829,In_1275,In_2484);
or U830 (N_830,In_1138,In_1737);
and U831 (N_831,In_1364,In_2424);
and U832 (N_832,In_707,In_1508);
or U833 (N_833,In_1365,In_479);
nor U834 (N_834,In_1171,In_2877);
or U835 (N_835,In_1999,In_1397);
nand U836 (N_836,In_273,In_1036);
nand U837 (N_837,In_443,In_1197);
nor U838 (N_838,In_1599,In_735);
xor U839 (N_839,In_715,In_1770);
xor U840 (N_840,In_1353,In_1660);
nand U841 (N_841,In_1361,In_20);
xor U842 (N_842,In_2350,In_461);
xnor U843 (N_843,In_2392,In_758);
or U844 (N_844,In_1937,In_139);
and U845 (N_845,In_2456,In_757);
and U846 (N_846,In_587,In_2891);
nor U847 (N_847,In_385,In_1265);
nor U848 (N_848,In_145,In_2314);
xnor U849 (N_849,In_708,In_2225);
xnor U850 (N_850,In_400,In_1360);
and U851 (N_851,In_2384,In_1918);
and U852 (N_852,In_2986,In_2980);
and U853 (N_853,In_991,In_603);
nand U854 (N_854,In_1046,In_562);
xor U855 (N_855,In_290,In_2638);
or U856 (N_856,In_2154,In_602);
nand U857 (N_857,In_2270,In_2546);
or U858 (N_858,In_994,In_18);
xnor U859 (N_859,In_902,In_2566);
nand U860 (N_860,In_2405,In_89);
and U861 (N_861,In_28,In_180);
nand U862 (N_862,In_485,In_933);
xor U863 (N_863,In_1877,In_2278);
nor U864 (N_864,In_267,In_2913);
nor U865 (N_865,In_1524,In_720);
nand U866 (N_866,In_1246,In_2857);
nor U867 (N_867,In_146,In_118);
and U868 (N_868,In_2421,In_2138);
nor U869 (N_869,In_2807,In_1043);
and U870 (N_870,In_2529,In_2044);
nor U871 (N_871,In_1273,In_631);
nor U872 (N_872,In_2033,In_2143);
or U873 (N_873,In_2324,In_2744);
nand U874 (N_874,In_1057,In_2376);
nor U875 (N_875,In_2007,In_1357);
nor U876 (N_876,In_881,In_1408);
or U877 (N_877,In_2592,In_1136);
and U878 (N_878,In_1765,In_2949);
or U879 (N_879,In_1062,In_2974);
xor U880 (N_880,In_2602,In_1370);
and U881 (N_881,In_1861,In_1211);
xnor U882 (N_882,In_2575,In_2659);
or U883 (N_883,In_548,In_1162);
or U884 (N_884,In_372,In_844);
xnor U885 (N_885,In_1915,In_1595);
and U886 (N_886,In_1631,In_2939);
nand U887 (N_887,In_697,In_2217);
nand U888 (N_888,In_442,In_1874);
and U889 (N_889,In_1474,In_132);
nand U890 (N_890,In_2476,In_129);
or U891 (N_891,In_640,In_1758);
xor U892 (N_892,In_759,In_1725);
nor U893 (N_893,In_112,In_1033);
nor U894 (N_894,In_1448,In_2516);
or U895 (N_895,In_2732,In_42);
or U896 (N_896,In_578,In_2140);
nor U897 (N_897,In_1727,In_1986);
nor U898 (N_898,In_2930,In_1260);
xnor U899 (N_899,In_516,In_1675);
nand U900 (N_900,In_2682,In_1111);
or U901 (N_901,In_106,In_696);
or U902 (N_902,In_2503,In_302);
nand U903 (N_903,In_2130,In_1223);
and U904 (N_904,In_1165,In_1082);
nor U905 (N_905,In_819,In_314);
and U906 (N_906,In_791,In_2858);
nor U907 (N_907,In_2696,In_2482);
nor U908 (N_908,In_2257,In_296);
and U909 (N_909,In_2040,In_2019);
nand U910 (N_910,In_1482,In_1195);
and U911 (N_911,In_2481,In_1038);
nor U912 (N_912,In_448,In_1031);
and U913 (N_913,In_721,In_924);
or U914 (N_914,In_576,In_1278);
nor U915 (N_915,In_1605,In_1965);
nand U916 (N_916,In_2979,In_2249);
nor U917 (N_917,In_1933,In_32);
nand U918 (N_918,In_1512,In_2150);
nor U919 (N_919,In_2670,In_1222);
nor U920 (N_920,In_2177,In_1574);
xor U921 (N_921,In_1749,In_2875);
nor U922 (N_922,In_2678,In_2446);
and U923 (N_923,In_1452,In_495);
xor U924 (N_924,In_2936,In_271);
and U925 (N_925,In_1280,In_215);
nor U926 (N_926,In_397,In_2128);
nand U927 (N_927,In_1034,In_1850);
nor U928 (N_928,In_904,In_1612);
or U929 (N_929,In_1988,In_2016);
or U930 (N_930,In_1147,In_2819);
nor U931 (N_931,In_623,In_1125);
and U932 (N_932,In_863,In_339);
nand U933 (N_933,In_1501,In_1697);
xor U934 (N_934,In_1124,In_718);
or U935 (N_935,In_1415,In_2416);
xnor U936 (N_936,In_1602,In_260);
nand U937 (N_937,In_393,In_2121);
or U938 (N_938,In_1779,In_2737);
nand U939 (N_939,In_2425,In_2160);
nand U940 (N_940,In_1897,In_1203);
xnor U941 (N_941,In_1531,In_2413);
nor U942 (N_942,In_2862,In_1826);
or U943 (N_943,In_1497,In_2097);
and U944 (N_944,In_2056,In_986);
nand U945 (N_945,In_1750,In_751);
nor U946 (N_946,In_1363,In_1680);
xor U947 (N_947,In_2338,In_1525);
nand U948 (N_948,In_1205,In_2071);
nand U949 (N_949,In_1373,In_2863);
xnor U950 (N_950,In_1436,In_1198);
or U951 (N_951,In_1678,In_996);
nand U952 (N_952,In_2514,In_1417);
or U953 (N_953,In_572,In_1662);
and U954 (N_954,In_1889,In_473);
or U955 (N_955,In_1997,In_726);
and U956 (N_956,In_1936,In_1212);
xor U957 (N_957,In_1754,In_1609);
and U958 (N_958,In_1375,In_261);
nor U959 (N_959,In_2105,In_1384);
and U960 (N_960,In_92,In_153);
xor U961 (N_961,In_189,In_1173);
and U962 (N_962,In_1155,In_2030);
or U963 (N_963,In_2774,In_2159);
xor U964 (N_964,In_2254,In_37);
xor U965 (N_965,In_1469,In_2010);
or U966 (N_966,In_805,In_1016);
xnor U967 (N_967,In_341,In_801);
xor U968 (N_968,In_2518,In_392);
and U969 (N_969,In_394,In_1266);
nand U970 (N_970,In_2906,In_1355);
and U971 (N_971,In_1835,In_491);
xnor U972 (N_972,In_15,In_1086);
nor U973 (N_973,In_49,In_2282);
nor U974 (N_974,In_2307,In_2291);
nor U975 (N_975,In_1189,In_2746);
or U976 (N_976,In_2776,In_2991);
nand U977 (N_977,In_2059,In_1056);
and U978 (N_978,In_286,In_438);
nor U979 (N_979,In_1230,In_411);
and U980 (N_980,In_980,In_2612);
nand U981 (N_981,In_446,In_1872);
xor U982 (N_982,In_2306,In_1753);
and U983 (N_983,In_1560,In_1411);
xnor U984 (N_984,In_2929,In_435);
nand U985 (N_985,In_1059,In_1634);
and U986 (N_986,In_843,In_2739);
and U987 (N_987,In_2388,In_1809);
and U988 (N_988,In_738,In_9);
nor U989 (N_989,In_2053,In_1797);
and U990 (N_990,In_1346,In_2657);
nand U991 (N_991,In_1316,In_1787);
xnor U992 (N_992,In_654,In_2184);
xor U993 (N_993,In_2666,In_906);
nor U994 (N_994,In_2978,In_2051);
and U995 (N_995,In_2868,In_460);
nor U996 (N_996,In_1556,In_1613);
nand U997 (N_997,In_1695,In_12);
nand U998 (N_998,In_693,In_1553);
xnor U999 (N_999,In_2928,In_31);
or U1000 (N_1000,In_2562,In_1763);
xor U1001 (N_1001,In_1196,In_245);
nor U1002 (N_1002,In_1778,In_364);
nand U1003 (N_1003,In_2395,In_1970);
or U1004 (N_1004,In_858,In_166);
xnor U1005 (N_1005,In_2805,In_97);
nor U1006 (N_1006,In_1156,In_1000);
xor U1007 (N_1007,In_2892,In_1768);
or U1008 (N_1008,In_2029,In_193);
xor U1009 (N_1009,In_1519,In_498);
nand U1010 (N_1010,In_1669,In_1643);
or U1011 (N_1011,In_1439,In_1882);
and U1012 (N_1012,In_1732,In_2084);
xor U1013 (N_1013,In_760,In_817);
or U1014 (N_1014,In_607,In_652);
nor U1015 (N_1015,In_2008,In_748);
nand U1016 (N_1016,In_2173,In_46);
xor U1017 (N_1017,In_1225,In_2331);
or U1018 (N_1018,In_1263,In_2993);
xor U1019 (N_1019,In_2540,In_377);
nand U1020 (N_1020,In_1379,In_992);
and U1021 (N_1021,In_1851,In_482);
or U1022 (N_1022,In_895,In_1242);
xor U1023 (N_1023,In_686,In_1089);
and U1024 (N_1024,In_428,In_2729);
and U1025 (N_1025,In_1318,In_879);
xnor U1026 (N_1026,In_1829,In_1645);
xor U1027 (N_1027,In_451,In_2045);
nand U1028 (N_1028,In_834,In_570);
nor U1029 (N_1029,In_13,In_1691);
or U1030 (N_1030,In_415,In_2543);
nor U1031 (N_1031,In_2474,In_2391);
or U1032 (N_1032,In_2820,In_2720);
and U1033 (N_1033,In_2248,In_808);
xnor U1034 (N_1034,In_2981,In_1961);
and U1035 (N_1035,In_2876,In_774);
nor U1036 (N_1036,In_1520,In_76);
nand U1037 (N_1037,In_911,In_2636);
or U1038 (N_1038,In_172,In_2451);
and U1039 (N_1039,In_67,In_2347);
nand U1040 (N_1040,In_2840,In_1495);
xor U1041 (N_1041,In_300,In_2343);
and U1042 (N_1042,In_678,In_2490);
and U1043 (N_1043,In_647,In_2144);
xor U1044 (N_1044,In_2157,In_2352);
or U1045 (N_1045,In_1284,In_2542);
nand U1046 (N_1046,In_2085,In_2239);
nand U1047 (N_1047,In_2675,In_2172);
and U1048 (N_1048,In_1073,In_1671);
or U1049 (N_1049,In_121,In_2295);
or U1050 (N_1050,In_2649,In_2596);
nand U1051 (N_1051,In_2834,In_2526);
or U1052 (N_1052,In_1121,In_769);
xor U1053 (N_1053,In_616,In_2351);
xnor U1054 (N_1054,In_927,In_1883);
nor U1055 (N_1055,In_1526,In_1893);
nand U1056 (N_1056,In_235,In_1949);
or U1057 (N_1057,In_432,In_1447);
and U1058 (N_1058,In_2213,In_2195);
nand U1059 (N_1059,In_605,In_622);
nand U1060 (N_1060,In_609,In_2445);
nand U1061 (N_1061,In_1504,In_1823);
nor U1062 (N_1062,In_2985,In_1489);
or U1063 (N_1063,In_2412,In_670);
nand U1064 (N_1064,In_2743,In_2431);
or U1065 (N_1065,In_1129,In_2357);
or U1066 (N_1066,In_1895,In_1158);
nor U1067 (N_1067,In_2797,In_2452);
or U1068 (N_1068,In_1923,In_1270);
and U1069 (N_1069,In_1979,In_2519);
nand U1070 (N_1070,In_2843,In_2081);
nand U1071 (N_1071,In_1585,In_2086);
and U1072 (N_1072,In_1567,In_852);
or U1073 (N_1073,In_2988,In_2061);
xnor U1074 (N_1074,In_1950,In_637);
nor U1075 (N_1075,In_2889,In_2900);
xnor U1076 (N_1076,In_2394,In_1616);
nand U1077 (N_1077,In_1966,In_205);
xnor U1078 (N_1078,In_143,In_269);
or U1079 (N_1079,In_2568,In_2288);
xnor U1080 (N_1080,In_823,In_0);
nand U1081 (N_1081,In_391,In_247);
and U1082 (N_1082,In_2155,In_34);
nor U1083 (N_1083,In_1191,In_1603);
and U1084 (N_1084,In_1299,In_2764);
nor U1085 (N_1085,In_2153,In_661);
and U1086 (N_1086,In_1592,In_2401);
or U1087 (N_1087,In_1001,In_1290);
or U1088 (N_1088,In_1285,In_1813);
or U1089 (N_1089,In_2587,In_458);
nand U1090 (N_1090,In_179,In_854);
nand U1091 (N_1091,In_2161,In_2667);
nor U1092 (N_1092,In_1261,In_1093);
nand U1093 (N_1093,In_246,In_232);
and U1094 (N_1094,In_1049,In_2626);
or U1095 (N_1095,In_1833,In_1053);
nor U1096 (N_1096,In_1356,In_1301);
xor U1097 (N_1097,In_2812,In_2832);
and U1098 (N_1098,In_1075,In_478);
nand U1099 (N_1099,In_2222,In_254);
xnor U1100 (N_1100,In_2050,In_502);
nand U1101 (N_1101,In_439,In_80);
nand U1102 (N_1102,In_2181,In_1019);
nor U1103 (N_1103,In_1714,In_45);
or U1104 (N_1104,In_903,In_2533);
xor U1105 (N_1105,In_620,In_1710);
nand U1106 (N_1106,In_2595,In_2689);
and U1107 (N_1107,In_1840,In_1771);
xnor U1108 (N_1108,In_1479,In_1688);
or U1109 (N_1109,In_2644,In_239);
nand U1110 (N_1110,In_2419,In_4);
or U1111 (N_1111,In_667,In_1898);
xnor U1112 (N_1112,In_1761,In_2083);
xor U1113 (N_1113,In_138,In_1785);
and U1114 (N_1114,In_1269,In_470);
and U1115 (N_1115,In_1037,In_1151);
or U1116 (N_1116,In_319,In_1864);
and U1117 (N_1117,In_2211,In_1746);
nor U1118 (N_1118,In_2698,In_2430);
and U1119 (N_1119,In_1007,In_83);
and U1120 (N_1120,In_331,In_569);
xnor U1121 (N_1121,In_276,In_665);
and U1122 (N_1122,In_1309,In_590);
xor U1123 (N_1123,In_1250,In_1875);
and U1124 (N_1124,In_1540,In_2224);
nor U1125 (N_1125,In_2487,In_1307);
or U1126 (N_1126,In_186,In_612);
or U1127 (N_1127,In_2462,In_2203);
xnor U1128 (N_1128,In_164,In_1015);
nor U1129 (N_1129,In_2006,In_413);
and U1130 (N_1130,In_1219,In_301);
nor U1131 (N_1131,In_1596,In_2372);
nor U1132 (N_1132,In_1766,In_577);
nand U1133 (N_1133,In_82,In_1777);
nor U1134 (N_1134,In_786,In_2113);
and U1135 (N_1135,In_659,In_1679);
nand U1136 (N_1136,In_1831,In_96);
xor U1137 (N_1137,In_2263,In_2520);
and U1138 (N_1138,In_1703,In_846);
nor U1139 (N_1139,In_1931,In_2948);
and U1140 (N_1140,In_2957,In_2385);
nand U1141 (N_1141,In_768,In_1554);
nand U1142 (N_1142,In_2409,In_1122);
nand U1143 (N_1143,In_1419,In_2279);
xnor U1144 (N_1144,In_2594,In_2918);
nand U1145 (N_1145,In_2738,In_666);
or U1146 (N_1146,In_2747,In_1267);
or U1147 (N_1147,In_2360,In_837);
and U1148 (N_1148,In_951,In_1326);
or U1149 (N_1149,In_2679,In_2062);
nor U1150 (N_1150,In_480,In_525);
nor U1151 (N_1151,In_752,In_1306);
or U1152 (N_1152,In_1516,In_1953);
nor U1153 (N_1153,In_1079,In_1944);
nand U1154 (N_1154,In_1385,In_1022);
nand U1155 (N_1155,In_1548,In_1204);
nor U1156 (N_1156,In_561,In_1581);
or U1157 (N_1157,In_1286,In_2722);
nor U1158 (N_1158,In_2994,In_2215);
nor U1159 (N_1159,In_1118,In_1590);
xor U1160 (N_1160,In_1139,In_487);
and U1161 (N_1161,In_1281,In_2182);
xnor U1162 (N_1162,In_1477,In_284);
and U1163 (N_1163,In_1693,In_821);
or U1164 (N_1164,In_2082,In_1792);
and U1165 (N_1165,In_283,In_2407);
and U1166 (N_1166,In_509,In_1698);
xnor U1167 (N_1167,In_2931,In_359);
xnor U1168 (N_1168,In_2836,In_1097);
nor U1169 (N_1169,In_358,In_373);
or U1170 (N_1170,In_833,In_2933);
nand U1171 (N_1171,In_2917,In_2505);
nor U1172 (N_1172,In_2815,In_2559);
or U1173 (N_1173,In_2313,In_1783);
xnor U1174 (N_1174,In_1274,In_61);
nand U1175 (N_1175,In_2106,In_2555);
and U1176 (N_1176,In_646,In_2859);
and U1177 (N_1177,In_1092,In_1341);
nor U1178 (N_1178,In_2661,In_2323);
nand U1179 (N_1179,In_753,In_2260);
nor U1180 (N_1180,In_1734,In_1858);
and U1181 (N_1181,In_2025,In_24);
and U1182 (N_1182,In_899,In_2945);
or U1183 (N_1183,In_2286,In_872);
nand U1184 (N_1184,In_1641,In_524);
and U1185 (N_1185,In_1418,In_274);
nor U1186 (N_1186,In_2020,In_291);
nand U1187 (N_1187,In_704,In_2604);
xor U1188 (N_1188,In_161,In_1480);
xor U1189 (N_1189,In_2308,In_1441);
nand U1190 (N_1190,In_506,In_1175);
nand U1191 (N_1191,In_307,In_23);
or U1192 (N_1192,In_1040,In_2782);
nand U1193 (N_1193,In_596,In_2188);
xnor U1194 (N_1194,In_889,In_1279);
nand U1195 (N_1195,In_147,In_2623);
or U1196 (N_1196,In_2206,In_2951);
or U1197 (N_1197,In_2494,In_1786);
and U1198 (N_1198,In_181,In_883);
and U1199 (N_1199,In_501,In_875);
or U1200 (N_1200,In_1342,In_2901);
or U1201 (N_1201,In_475,In_472);
or U1202 (N_1202,In_2711,In_292);
or U1203 (N_1203,In_140,In_2089);
xnor U1204 (N_1204,In_656,In_2251);
and U1205 (N_1205,In_2390,In_1209);
or U1206 (N_1206,In_537,In_462);
nand U1207 (N_1207,In_233,In_53);
or U1208 (N_1208,In_2908,In_567);
or U1209 (N_1209,In_241,In_669);
nand U1210 (N_1210,In_1293,In_2072);
and U1211 (N_1211,In_1799,In_2400);
nand U1212 (N_1212,In_2162,In_1338);
xnor U1213 (N_1213,In_2422,In_1025);
or U1214 (N_1214,In_1066,In_2349);
nor U1215 (N_1215,In_1231,In_468);
xnor U1216 (N_1216,In_1958,In_776);
nor U1217 (N_1217,In_51,In_120);
xnor U1218 (N_1218,In_544,In_2563);
xnor U1219 (N_1219,In_1344,In_2196);
xor U1220 (N_1220,In_44,In_352);
nor U1221 (N_1221,In_946,In_1607);
nand U1222 (N_1222,In_78,In_464);
nand U1223 (N_1223,In_2444,In_642);
and U1224 (N_1224,In_2969,In_2761);
and U1225 (N_1225,In_2724,In_2793);
and U1226 (N_1226,In_1975,In_1728);
xnor U1227 (N_1227,In_773,In_1506);
nand U1228 (N_1228,In_1583,In_1932);
and U1229 (N_1229,In_1566,In_2377);
and U1230 (N_1230,In_2925,In_597);
or U1231 (N_1231,In_1928,In_2370);
and U1232 (N_1232,In_1142,In_1006);
nor U1233 (N_1233,In_328,In_939);
and U1234 (N_1234,In_2515,In_338);
nand U1235 (N_1235,In_2507,In_75);
and U1236 (N_1236,In_2856,In_1020);
or U1237 (N_1237,In_30,In_794);
and U1238 (N_1238,In_1899,In_1114);
or U1239 (N_1239,In_857,In_2023);
nor U1240 (N_1240,In_1981,In_64);
nor U1241 (N_1241,In_1722,In_1207);
xor U1242 (N_1242,In_257,In_1127);
nor U1243 (N_1243,In_2218,In_2944);
xor U1244 (N_1244,In_1586,In_1627);
nor U1245 (N_1245,In_2134,In_1240);
and U1246 (N_1246,In_1681,In_2241);
nand U1247 (N_1247,In_2551,In_2272);
or U1248 (N_1248,In_1759,In_2784);
nand U1249 (N_1249,In_1804,In_1565);
or U1250 (N_1250,In_228,In_2169);
nor U1251 (N_1251,In_297,In_1076);
and U1252 (N_1252,In_648,In_144);
nand U1253 (N_1253,In_226,In_2827);
nand U1254 (N_1254,In_2220,In_2488);
or U1255 (N_1255,In_967,In_1472);
nand U1256 (N_1256,In_114,In_381);
nand U1257 (N_1257,In_477,In_679);
xnor U1258 (N_1258,In_1894,In_914);
and U1259 (N_1259,In_2099,In_318);
nor U1260 (N_1260,In_573,In_211);
xor U1261 (N_1261,In_431,In_2658);
and U1262 (N_1262,In_162,In_2972);
or U1263 (N_1263,In_956,In_1068);
xor U1264 (N_1264,In_2880,In_2831);
nand U1265 (N_1265,In_800,In_175);
and U1266 (N_1266,In_785,In_934);
xnor U1267 (N_1267,In_2598,In_1239);
or U1268 (N_1268,In_2787,In_492);
nand U1269 (N_1269,In_1170,In_467);
or U1270 (N_1270,In_2524,In_1302);
and U1271 (N_1271,In_1429,In_1067);
xor U1272 (N_1272,In_2873,In_2882);
or U1273 (N_1273,In_925,In_2954);
nor U1274 (N_1274,In_1909,In_868);
xnor U1275 (N_1275,In_2478,In_2332);
nand U1276 (N_1276,In_683,In_2076);
or U1277 (N_1277,In_2878,In_522);
xnor U1278 (N_1278,In_1083,In_2570);
nor U1279 (N_1279,In_685,In_2830);
nand U1280 (N_1280,In_533,In_1513);
nand U1281 (N_1281,In_918,In_1347);
nand U1282 (N_1282,In_2179,In_1331);
and U1283 (N_1283,In_1996,In_2934);
xnor U1284 (N_1284,In_2170,In_263);
and U1285 (N_1285,In_2142,In_170);
nor U1286 (N_1286,In_2704,In_357);
nor U1287 (N_1287,In_1095,In_1123);
nand U1288 (N_1288,In_2120,In_797);
or U1289 (N_1289,In_280,In_657);
nand U1290 (N_1290,In_2124,In_1692);
or U1291 (N_1291,In_2265,In_2497);
nor U1292 (N_1292,In_775,In_344);
nor U1293 (N_1293,In_1757,In_2335);
xor U1294 (N_1294,In_514,In_2923);
nor U1295 (N_1295,In_714,In_1465);
xnor U1296 (N_1296,In_278,In_444);
or U1297 (N_1297,In_826,In_1650);
nand U1298 (N_1298,In_363,In_1788);
nor U1299 (N_1299,In_950,In_2532);
nor U1300 (N_1300,In_1839,In_1192);
or U1301 (N_1301,In_360,In_1297);
nand U1302 (N_1302,In_429,In_1135);
nor U1303 (N_1303,In_2833,In_2924);
nor U1304 (N_1304,In_1579,In_73);
nand U1305 (N_1305,In_77,In_484);
or U1306 (N_1306,In_1004,In_1505);
or U1307 (N_1307,In_1186,In_104);
nand U1308 (N_1308,In_416,In_1578);
nand U1309 (N_1309,In_1593,In_2603);
and U1310 (N_1310,In_2116,In_1435);
or U1311 (N_1311,In_799,In_410);
nor U1312 (N_1312,In_2676,In_1042);
nor U1313 (N_1313,In_2904,In_1713);
or U1314 (N_1314,In_1798,In_62);
xor U1315 (N_1315,In_79,In_256);
and U1316 (N_1316,In_2765,In_2117);
or U1317 (N_1317,In_47,In_2946);
xnor U1318 (N_1318,In_1085,In_2074);
nor U1319 (N_1319,In_2997,In_1808);
nor U1320 (N_1320,In_2256,In_2115);
or U1321 (N_1321,In_408,In_1185);
xor U1322 (N_1322,In_399,In_2354);
xnor U1323 (N_1323,In_851,In_744);
or U1324 (N_1324,In_29,In_2950);
nor U1325 (N_1325,In_1303,In_2999);
nor U1326 (N_1326,In_50,In_141);
or U1327 (N_1327,In_700,In_2447);
nand U1328 (N_1328,In_1539,In_650);
xor U1329 (N_1329,In_2902,In_1388);
xor U1330 (N_1330,In_2165,In_68);
or U1331 (N_1331,In_1478,In_1463);
and U1332 (N_1332,In_66,In_1104);
or U1333 (N_1333,In_2938,In_361);
xor U1334 (N_1334,In_1430,In_454);
nor U1335 (N_1335,In_2582,In_575);
or U1336 (N_1336,In_1256,In_2693);
xnor U1337 (N_1337,In_518,In_22);
nand U1338 (N_1338,In_2853,In_2703);
nand U1339 (N_1339,In_2375,In_2449);
xnor U1340 (N_1340,In_1674,In_923);
and U1341 (N_1341,In_2,In_8);
nor U1342 (N_1342,In_2438,In_2298);
nand U1343 (N_1343,In_356,In_2607);
and U1344 (N_1344,In_2393,In_183);
or U1345 (N_1345,In_2399,In_1044);
nor U1346 (N_1346,In_2027,In_1842);
nor U1347 (N_1347,In_1991,In_1107);
nand U1348 (N_1348,In_566,In_40);
and U1349 (N_1349,In_2151,In_419);
nand U1350 (N_1350,In_1871,In_668);
nor U1351 (N_1351,In_2202,In_365);
xor U1352 (N_1352,In_1740,In_1776);
xnor U1353 (N_1353,In_2316,In_2569);
nand U1354 (N_1354,In_2275,In_2443);
and U1355 (N_1355,In_1099,In_2471);
and U1356 (N_1356,In_770,In_185);
nor U1357 (N_1357,In_1362,In_2107);
nand U1358 (N_1358,In_2185,In_249);
and U1359 (N_1359,In_512,In_528);
and U1360 (N_1360,In_1367,In_2191);
or U1361 (N_1361,In_2108,In_2538);
and U1362 (N_1362,In_937,In_2714);
nor U1363 (N_1363,In_1830,In_2221);
nor U1364 (N_1364,In_701,In_2971);
or U1365 (N_1365,In_2702,In_1879);
or U1366 (N_1366,In_1289,In_1545);
nor U1367 (N_1367,In_2403,In_1878);
nand U1368 (N_1368,In_1885,In_1406);
xor U1369 (N_1369,In_299,In_355);
nand U1370 (N_1370,In_1576,In_1682);
nor U1371 (N_1371,In_2055,In_953);
nand U1372 (N_1372,In_36,In_379);
nand U1373 (N_1373,In_1295,In_1055);
nor U1374 (N_1374,In_2854,In_1549);
or U1375 (N_1375,In_754,In_2631);
nor U1376 (N_1376,In_200,In_557);
and U1377 (N_1377,In_244,In_2002);
nand U1378 (N_1378,In_2668,In_2799);
xor U1379 (N_1379,In_2289,In_1973);
or U1380 (N_1380,In_2847,In_942);
nor U1381 (N_1381,In_1715,In_1144);
nor U1382 (N_1382,In_305,In_1328);
or U1383 (N_1383,In_2024,In_383);
or U1384 (N_1384,In_1888,In_65);
or U1385 (N_1385,In_2131,In_1869);
xnor U1386 (N_1386,In_409,In_2734);
xor U1387 (N_1387,In_894,In_1529);
xor U1388 (N_1388,In_272,In_1647);
or U1389 (N_1389,In_1854,In_2032);
nor U1390 (N_1390,In_321,In_1141);
nor U1391 (N_1391,In_2404,In_2432);
xnor U1392 (N_1392,In_675,In_1876);
or U1393 (N_1393,In_452,In_1657);
nand U1394 (N_1394,In_2369,In_530);
nor U1395 (N_1395,In_5,In_85);
nor U1396 (N_1396,In_1910,In_2817);
or U1397 (N_1397,In_1101,In_202);
and U1398 (N_1398,In_221,In_2135);
and U1399 (N_1399,In_850,In_1481);
nor U1400 (N_1400,In_870,In_2770);
xnor U1401 (N_1401,In_1584,In_2095);
nor U1402 (N_1402,In_1661,In_2183);
nand U1403 (N_1403,In_2669,In_351);
nor U1404 (N_1404,In_207,In_2940);
and U1405 (N_1405,In_2920,In_976);
xnor U1406 (N_1406,In_2616,In_2262);
nor U1407 (N_1407,In_2861,In_511);
xnor U1408 (N_1408,In_2171,In_550);
nand U1409 (N_1409,In_313,In_2590);
and U1410 (N_1410,In_536,In_878);
xnor U1411 (N_1411,In_639,In_2246);
xnor U1412 (N_1412,In_1072,In_2816);
and U1413 (N_1413,In_2361,In_778);
xor U1414 (N_1414,In_2536,In_2895);
and U1415 (N_1415,In_136,In_2839);
xor U1416 (N_1416,In_1747,In_1310);
or U1417 (N_1417,In_663,In_687);
and U1418 (N_1418,In_1381,In_2654);
or U1419 (N_1419,In_1856,In_2501);
nor U1420 (N_1420,In_1995,In_2749);
nor U1421 (N_1421,In_1717,In_496);
xor U1422 (N_1422,In_2535,In_2789);
and U1423 (N_1423,In_2813,In_1984);
nor U1424 (N_1424,In_2387,In_702);
nand U1425 (N_1425,In_1490,In_424);
xnor U1426 (N_1426,In_1563,In_2341);
nor U1427 (N_1427,In_935,In_1058);
nor U1428 (N_1428,In_2327,In_1587);
nand U1429 (N_1429,In_1386,In_1183);
and U1430 (N_1430,In_2731,In_1951);
and U1431 (N_1431,In_126,In_2509);
nand U1432 (N_1432,In_921,In_2284);
or U1433 (N_1433,In_1180,In_1343);
nor U1434 (N_1434,In_2881,In_2671);
xnor U1435 (N_1435,In_559,In_1649);
nor U1436 (N_1436,In_598,In_1320);
nand U1437 (N_1437,In_948,In_1594);
xnor U1438 (N_1438,In_722,In_2320);
nor U1439 (N_1439,In_2674,In_2959);
nand U1440 (N_1440,In_1514,In_997);
and U1441 (N_1441,In_1668,In_742);
or U1442 (N_1442,In_981,In_1327);
and U1443 (N_1443,In_1926,In_766);
nor U1444 (N_1444,In_2705,In_317);
and U1445 (N_1445,In_985,In_16);
or U1446 (N_1446,In_1756,In_2180);
or U1447 (N_1447,In_1601,In_425);
nor U1448 (N_1448,In_2584,In_2846);
or U1449 (N_1449,In_1193,In_594);
or U1450 (N_1450,In_2500,In_1446);
nand U1451 (N_1451,In_1304,In_1943);
and U1452 (N_1452,In_2311,In_2794);
and U1453 (N_1453,In_517,In_194);
xor U1454 (N_1454,In_1935,In_1723);
or U1455 (N_1455,In_2766,In_2894);
nor U1456 (N_1456,In_21,In_2601);
xnor U1457 (N_1457,In_728,In_2810);
and U1458 (N_1458,In_2078,In_681);
or U1459 (N_1459,In_1259,In_412);
and U1460 (N_1460,In_586,In_970);
nand U1461 (N_1461,In_2544,In_2553);
and U1462 (N_1462,In_1017,In_2821);
nor U1463 (N_1463,In_815,In_395);
xnor U1464 (N_1464,In_1298,In_224);
xnor U1465 (N_1465,In_54,In_1434);
nand U1466 (N_1466,In_2580,In_1011);
nor U1467 (N_1467,In_1610,In_1857);
or U1468 (N_1468,In_1790,In_1528);
nor U1469 (N_1469,In_2297,In_1112);
nor U1470 (N_1470,In_2080,In_130);
and U1471 (N_1471,In_2204,In_293);
nand U1472 (N_1472,In_1374,In_984);
nor U1473 (N_1473,In_178,In_2310);
and U1474 (N_1474,In_2727,In_2342);
or U1475 (N_1475,In_1457,In_2192);
or U1476 (N_1476,In_807,In_765);
and U1477 (N_1477,In_150,In_1021);
nand U1478 (N_1478,In_337,In_2664);
or U1479 (N_1479,In_1846,In_1458);
or U1480 (N_1480,In_2402,In_285);
and U1481 (N_1481,In_1159,In_63);
nor U1482 (N_1482,In_1648,In_849);
xnor U1483 (N_1483,In_891,In_378);
and U1484 (N_1484,In_471,In_196);
nor U1485 (N_1485,In_2486,In_248);
or U1486 (N_1486,In_253,In_593);
nor U1487 (N_1487,In_627,In_1537);
or U1488 (N_1488,In_1459,In_1906);
nand U1489 (N_1489,In_599,In_1724);
xor U1490 (N_1490,In_2545,In_838);
and U1491 (N_1491,In_1110,In_2870);
nor U1492 (N_1492,In_2087,In_897);
xor U1493 (N_1493,In_2772,In_119);
nand U1494 (N_1494,In_1929,In_1824);
and U1495 (N_1495,In_2984,In_1635);
nor U1496 (N_1496,In_1051,In_210);
xnor U1497 (N_1497,In_7,In_2026);
xor U1498 (N_1498,In_1690,In_2110);
xor U1499 (N_1499,In_1080,In_2258);
nor U1500 (N_1500,In_1596,In_1757);
or U1501 (N_1501,In_2654,In_443);
nor U1502 (N_1502,In_2268,In_715);
and U1503 (N_1503,In_2302,In_2472);
nand U1504 (N_1504,In_2336,In_2324);
and U1505 (N_1505,In_2710,In_2799);
xnor U1506 (N_1506,In_2296,In_2392);
or U1507 (N_1507,In_2094,In_1424);
nand U1508 (N_1508,In_1482,In_352);
nand U1509 (N_1509,In_144,In_2325);
xor U1510 (N_1510,In_273,In_2839);
or U1511 (N_1511,In_723,In_2022);
nor U1512 (N_1512,In_1639,In_2567);
nand U1513 (N_1513,In_2271,In_2603);
or U1514 (N_1514,In_1103,In_1448);
nor U1515 (N_1515,In_2006,In_755);
nand U1516 (N_1516,In_2591,In_1150);
xor U1517 (N_1517,In_2154,In_927);
nor U1518 (N_1518,In_2107,In_799);
and U1519 (N_1519,In_1374,In_2630);
and U1520 (N_1520,In_2231,In_2718);
and U1521 (N_1521,In_2445,In_1387);
nand U1522 (N_1522,In_117,In_906);
nand U1523 (N_1523,In_150,In_1938);
nor U1524 (N_1524,In_188,In_1978);
nand U1525 (N_1525,In_1007,In_1149);
xor U1526 (N_1526,In_999,In_887);
or U1527 (N_1527,In_504,In_2671);
and U1528 (N_1528,In_421,In_1126);
nor U1529 (N_1529,In_719,In_27);
nor U1530 (N_1530,In_390,In_1883);
and U1531 (N_1531,In_876,In_2542);
xor U1532 (N_1532,In_2506,In_586);
xnor U1533 (N_1533,In_982,In_1634);
nand U1534 (N_1534,In_2173,In_2921);
nand U1535 (N_1535,In_1801,In_1467);
nand U1536 (N_1536,In_106,In_2961);
nor U1537 (N_1537,In_1426,In_1756);
nor U1538 (N_1538,In_1169,In_1927);
or U1539 (N_1539,In_202,In_2400);
xnor U1540 (N_1540,In_2644,In_2083);
and U1541 (N_1541,In_887,In_1748);
or U1542 (N_1542,In_1947,In_1051);
nand U1543 (N_1543,In_1062,In_1194);
or U1544 (N_1544,In_1180,In_480);
or U1545 (N_1545,In_80,In_1386);
xnor U1546 (N_1546,In_533,In_548);
nor U1547 (N_1547,In_2557,In_1614);
nand U1548 (N_1548,In_2126,In_587);
nor U1549 (N_1549,In_1980,In_398);
nor U1550 (N_1550,In_2556,In_2210);
nand U1551 (N_1551,In_148,In_2738);
nor U1552 (N_1552,In_821,In_2259);
and U1553 (N_1553,In_1358,In_326);
or U1554 (N_1554,In_2604,In_2797);
or U1555 (N_1555,In_2386,In_1818);
nand U1556 (N_1556,In_1315,In_563);
or U1557 (N_1557,In_1256,In_1258);
xnor U1558 (N_1558,In_705,In_1399);
or U1559 (N_1559,In_691,In_1690);
xnor U1560 (N_1560,In_1486,In_622);
or U1561 (N_1561,In_2293,In_517);
nand U1562 (N_1562,In_2956,In_1848);
xor U1563 (N_1563,In_1502,In_1585);
nor U1564 (N_1564,In_1690,In_2472);
and U1565 (N_1565,In_2584,In_1212);
xor U1566 (N_1566,In_767,In_1679);
and U1567 (N_1567,In_1485,In_1235);
nand U1568 (N_1568,In_2963,In_2651);
xor U1569 (N_1569,In_980,In_280);
nand U1570 (N_1570,In_2194,In_1861);
and U1571 (N_1571,In_71,In_2802);
and U1572 (N_1572,In_1497,In_1735);
nand U1573 (N_1573,In_654,In_455);
nand U1574 (N_1574,In_188,In_1367);
nor U1575 (N_1575,In_223,In_1967);
and U1576 (N_1576,In_2211,In_1870);
and U1577 (N_1577,In_1660,In_1130);
and U1578 (N_1578,In_1356,In_1863);
and U1579 (N_1579,In_1668,In_305);
and U1580 (N_1580,In_624,In_1623);
or U1581 (N_1581,In_2764,In_1041);
xor U1582 (N_1582,In_626,In_972);
nand U1583 (N_1583,In_1360,In_2722);
and U1584 (N_1584,In_1409,In_2402);
nor U1585 (N_1585,In_218,In_2101);
xnor U1586 (N_1586,In_1384,In_353);
nand U1587 (N_1587,In_1322,In_2206);
nand U1588 (N_1588,In_1548,In_912);
nor U1589 (N_1589,In_186,In_1784);
and U1590 (N_1590,In_631,In_2043);
nand U1591 (N_1591,In_2233,In_2858);
or U1592 (N_1592,In_749,In_239);
nand U1593 (N_1593,In_899,In_202);
xnor U1594 (N_1594,In_2933,In_694);
and U1595 (N_1595,In_2389,In_181);
and U1596 (N_1596,In_2998,In_273);
or U1597 (N_1597,In_801,In_654);
and U1598 (N_1598,In_363,In_375);
xnor U1599 (N_1599,In_2350,In_2950);
and U1600 (N_1600,In_2778,In_2954);
nand U1601 (N_1601,In_753,In_499);
nand U1602 (N_1602,In_1835,In_1172);
nor U1603 (N_1603,In_2534,In_688);
nand U1604 (N_1604,In_1354,In_1681);
and U1605 (N_1605,In_2750,In_995);
or U1606 (N_1606,In_1669,In_1733);
or U1607 (N_1607,In_1313,In_1280);
nand U1608 (N_1608,In_2580,In_7);
xor U1609 (N_1609,In_1825,In_2334);
nand U1610 (N_1610,In_1008,In_2363);
xor U1611 (N_1611,In_1896,In_2546);
nor U1612 (N_1612,In_2477,In_1296);
nand U1613 (N_1613,In_96,In_848);
nand U1614 (N_1614,In_2207,In_804);
nor U1615 (N_1615,In_560,In_612);
xor U1616 (N_1616,In_1920,In_2692);
xor U1617 (N_1617,In_2929,In_1463);
xnor U1618 (N_1618,In_230,In_1287);
nand U1619 (N_1619,In_291,In_2267);
xor U1620 (N_1620,In_213,In_505);
nor U1621 (N_1621,In_2151,In_1249);
nand U1622 (N_1622,In_1622,In_2158);
and U1623 (N_1623,In_2911,In_455);
xnor U1624 (N_1624,In_637,In_2163);
and U1625 (N_1625,In_1190,In_213);
nand U1626 (N_1626,In_730,In_2819);
nor U1627 (N_1627,In_78,In_680);
or U1628 (N_1628,In_344,In_1145);
nor U1629 (N_1629,In_2818,In_1751);
and U1630 (N_1630,In_1338,In_2599);
nor U1631 (N_1631,In_522,In_1483);
and U1632 (N_1632,In_1741,In_2843);
nand U1633 (N_1633,In_2867,In_2015);
or U1634 (N_1634,In_2543,In_1980);
or U1635 (N_1635,In_554,In_2043);
nor U1636 (N_1636,In_313,In_658);
nor U1637 (N_1637,In_919,In_2683);
and U1638 (N_1638,In_2592,In_703);
xor U1639 (N_1639,In_1822,In_2704);
xor U1640 (N_1640,In_1291,In_2324);
or U1641 (N_1641,In_291,In_845);
nor U1642 (N_1642,In_208,In_2149);
nand U1643 (N_1643,In_290,In_2215);
and U1644 (N_1644,In_197,In_915);
nor U1645 (N_1645,In_1490,In_66);
xor U1646 (N_1646,In_1544,In_282);
xnor U1647 (N_1647,In_612,In_694);
or U1648 (N_1648,In_1354,In_2384);
nor U1649 (N_1649,In_2854,In_2424);
nand U1650 (N_1650,In_2823,In_2861);
nand U1651 (N_1651,In_966,In_2311);
nor U1652 (N_1652,In_57,In_2189);
nor U1653 (N_1653,In_797,In_2202);
nor U1654 (N_1654,In_921,In_2603);
and U1655 (N_1655,In_1674,In_417);
nand U1656 (N_1656,In_124,In_640);
nand U1657 (N_1657,In_1776,In_2678);
or U1658 (N_1658,In_681,In_2586);
and U1659 (N_1659,In_1363,In_2501);
nor U1660 (N_1660,In_490,In_2774);
nor U1661 (N_1661,In_2908,In_2104);
or U1662 (N_1662,In_1049,In_1984);
or U1663 (N_1663,In_1105,In_1174);
or U1664 (N_1664,In_1081,In_622);
nor U1665 (N_1665,In_473,In_1142);
xnor U1666 (N_1666,In_534,In_2611);
nor U1667 (N_1667,In_1256,In_375);
nand U1668 (N_1668,In_2547,In_16);
nor U1669 (N_1669,In_2918,In_1135);
or U1670 (N_1670,In_2305,In_358);
nor U1671 (N_1671,In_1711,In_2513);
or U1672 (N_1672,In_1374,In_1997);
nand U1673 (N_1673,In_2194,In_2905);
nand U1674 (N_1674,In_1418,In_2440);
or U1675 (N_1675,In_2124,In_993);
xor U1676 (N_1676,In_292,In_641);
xnor U1677 (N_1677,In_387,In_1598);
nand U1678 (N_1678,In_25,In_1930);
and U1679 (N_1679,In_2071,In_1426);
xnor U1680 (N_1680,In_2799,In_1321);
nor U1681 (N_1681,In_967,In_1000);
or U1682 (N_1682,In_1050,In_1835);
or U1683 (N_1683,In_1856,In_1392);
nor U1684 (N_1684,In_1393,In_2163);
or U1685 (N_1685,In_268,In_42);
xnor U1686 (N_1686,In_171,In_2374);
or U1687 (N_1687,In_982,In_1278);
nor U1688 (N_1688,In_1054,In_426);
xor U1689 (N_1689,In_1208,In_1951);
xor U1690 (N_1690,In_163,In_861);
or U1691 (N_1691,In_2433,In_2625);
xnor U1692 (N_1692,In_337,In_2927);
and U1693 (N_1693,In_2537,In_1281);
or U1694 (N_1694,In_2321,In_2367);
and U1695 (N_1695,In_1219,In_1896);
xor U1696 (N_1696,In_2746,In_196);
and U1697 (N_1697,In_772,In_62);
nor U1698 (N_1698,In_2277,In_2474);
xor U1699 (N_1699,In_2436,In_2761);
nand U1700 (N_1700,In_1793,In_1309);
xnor U1701 (N_1701,In_1723,In_2534);
nor U1702 (N_1702,In_359,In_1967);
or U1703 (N_1703,In_1977,In_2467);
and U1704 (N_1704,In_545,In_1585);
or U1705 (N_1705,In_1098,In_548);
xor U1706 (N_1706,In_112,In_2562);
nand U1707 (N_1707,In_2714,In_902);
or U1708 (N_1708,In_721,In_1090);
nand U1709 (N_1709,In_2004,In_1140);
xnor U1710 (N_1710,In_809,In_2123);
and U1711 (N_1711,In_63,In_1781);
and U1712 (N_1712,In_1933,In_1115);
nand U1713 (N_1713,In_91,In_1896);
and U1714 (N_1714,In_1302,In_300);
xor U1715 (N_1715,In_724,In_2180);
and U1716 (N_1716,In_460,In_2102);
and U1717 (N_1717,In_1866,In_2693);
and U1718 (N_1718,In_529,In_2867);
or U1719 (N_1719,In_2820,In_2927);
or U1720 (N_1720,In_2836,In_1154);
xor U1721 (N_1721,In_2782,In_2884);
nor U1722 (N_1722,In_239,In_622);
xor U1723 (N_1723,In_2005,In_2031);
or U1724 (N_1724,In_1486,In_2709);
nand U1725 (N_1725,In_725,In_2539);
xnor U1726 (N_1726,In_2809,In_1910);
nor U1727 (N_1727,In_2489,In_1414);
and U1728 (N_1728,In_1476,In_1678);
or U1729 (N_1729,In_2610,In_2627);
xor U1730 (N_1730,In_86,In_1774);
nor U1731 (N_1731,In_1182,In_2139);
and U1732 (N_1732,In_536,In_2522);
or U1733 (N_1733,In_476,In_721);
and U1734 (N_1734,In_2494,In_2024);
or U1735 (N_1735,In_1324,In_1913);
and U1736 (N_1736,In_2059,In_1139);
xor U1737 (N_1737,In_1323,In_814);
nor U1738 (N_1738,In_1436,In_1707);
xnor U1739 (N_1739,In_2157,In_1255);
nand U1740 (N_1740,In_2532,In_150);
or U1741 (N_1741,In_621,In_1968);
or U1742 (N_1742,In_2556,In_1519);
or U1743 (N_1743,In_2095,In_1576);
or U1744 (N_1744,In_2569,In_23);
and U1745 (N_1745,In_2306,In_1974);
and U1746 (N_1746,In_2267,In_2045);
and U1747 (N_1747,In_2713,In_790);
nor U1748 (N_1748,In_438,In_2930);
xnor U1749 (N_1749,In_637,In_2237);
xor U1750 (N_1750,In_43,In_310);
and U1751 (N_1751,In_437,In_2940);
and U1752 (N_1752,In_2355,In_1176);
nand U1753 (N_1753,In_852,In_32);
or U1754 (N_1754,In_936,In_737);
and U1755 (N_1755,In_1494,In_47);
and U1756 (N_1756,In_1538,In_952);
nor U1757 (N_1757,In_1765,In_1111);
nor U1758 (N_1758,In_2068,In_2109);
xnor U1759 (N_1759,In_2869,In_2743);
xnor U1760 (N_1760,In_2719,In_996);
and U1761 (N_1761,In_1149,In_193);
and U1762 (N_1762,In_811,In_1000);
nand U1763 (N_1763,In_2976,In_459);
xnor U1764 (N_1764,In_317,In_1235);
nor U1765 (N_1765,In_1194,In_1356);
xor U1766 (N_1766,In_208,In_191);
xor U1767 (N_1767,In_2555,In_2595);
xnor U1768 (N_1768,In_1152,In_2543);
nand U1769 (N_1769,In_20,In_235);
nor U1770 (N_1770,In_428,In_2534);
and U1771 (N_1771,In_2178,In_1284);
nor U1772 (N_1772,In_2728,In_2810);
nand U1773 (N_1773,In_2590,In_504);
nor U1774 (N_1774,In_461,In_1540);
nand U1775 (N_1775,In_63,In_2834);
or U1776 (N_1776,In_480,In_2769);
or U1777 (N_1777,In_1644,In_213);
or U1778 (N_1778,In_1868,In_2238);
and U1779 (N_1779,In_263,In_2290);
nor U1780 (N_1780,In_1210,In_370);
nand U1781 (N_1781,In_1169,In_1484);
or U1782 (N_1782,In_47,In_1794);
nor U1783 (N_1783,In_2797,In_2250);
and U1784 (N_1784,In_604,In_315);
or U1785 (N_1785,In_271,In_619);
xor U1786 (N_1786,In_1262,In_1580);
or U1787 (N_1787,In_40,In_1225);
or U1788 (N_1788,In_1539,In_252);
nand U1789 (N_1789,In_978,In_2439);
or U1790 (N_1790,In_1918,In_2732);
nor U1791 (N_1791,In_1718,In_1041);
nor U1792 (N_1792,In_2761,In_2253);
nor U1793 (N_1793,In_9,In_486);
nor U1794 (N_1794,In_2193,In_2693);
nand U1795 (N_1795,In_1419,In_1011);
nand U1796 (N_1796,In_431,In_1816);
or U1797 (N_1797,In_2284,In_963);
nor U1798 (N_1798,In_1263,In_2670);
nand U1799 (N_1799,In_2340,In_2447);
nand U1800 (N_1800,In_2421,In_2085);
or U1801 (N_1801,In_647,In_1);
xnor U1802 (N_1802,In_2562,In_2289);
nand U1803 (N_1803,In_2272,In_1794);
nand U1804 (N_1804,In_2469,In_2627);
xor U1805 (N_1805,In_199,In_660);
xnor U1806 (N_1806,In_1737,In_1590);
nand U1807 (N_1807,In_870,In_84);
nand U1808 (N_1808,In_2610,In_2156);
and U1809 (N_1809,In_1724,In_149);
or U1810 (N_1810,In_2402,In_687);
xor U1811 (N_1811,In_2931,In_276);
or U1812 (N_1812,In_196,In_141);
or U1813 (N_1813,In_1882,In_1883);
and U1814 (N_1814,In_415,In_2829);
and U1815 (N_1815,In_210,In_824);
or U1816 (N_1816,In_1209,In_1514);
or U1817 (N_1817,In_2102,In_2291);
and U1818 (N_1818,In_1573,In_1338);
nand U1819 (N_1819,In_799,In_1152);
nand U1820 (N_1820,In_1655,In_2506);
or U1821 (N_1821,In_2730,In_1814);
or U1822 (N_1822,In_2335,In_571);
and U1823 (N_1823,In_1642,In_2825);
nor U1824 (N_1824,In_1013,In_2986);
and U1825 (N_1825,In_93,In_2187);
or U1826 (N_1826,In_2829,In_1671);
and U1827 (N_1827,In_811,In_2017);
and U1828 (N_1828,In_1261,In_2085);
or U1829 (N_1829,In_1104,In_982);
and U1830 (N_1830,In_1993,In_403);
xor U1831 (N_1831,In_2090,In_1618);
and U1832 (N_1832,In_1120,In_1605);
xor U1833 (N_1833,In_906,In_2176);
or U1834 (N_1834,In_2254,In_525);
and U1835 (N_1835,In_2624,In_1437);
xor U1836 (N_1836,In_2738,In_2995);
and U1837 (N_1837,In_513,In_1041);
or U1838 (N_1838,In_877,In_1286);
or U1839 (N_1839,In_2386,In_615);
and U1840 (N_1840,In_2811,In_2946);
xnor U1841 (N_1841,In_1936,In_83);
nand U1842 (N_1842,In_831,In_1711);
xnor U1843 (N_1843,In_2831,In_118);
nand U1844 (N_1844,In_2148,In_1282);
and U1845 (N_1845,In_2478,In_1882);
xor U1846 (N_1846,In_1046,In_132);
nand U1847 (N_1847,In_1178,In_1478);
xnor U1848 (N_1848,In_2519,In_922);
and U1849 (N_1849,In_2903,In_2473);
and U1850 (N_1850,In_2766,In_1163);
nand U1851 (N_1851,In_1040,In_2408);
nand U1852 (N_1852,In_401,In_2466);
nand U1853 (N_1853,In_2438,In_2021);
nand U1854 (N_1854,In_552,In_1447);
or U1855 (N_1855,In_2026,In_1784);
and U1856 (N_1856,In_1383,In_1125);
nor U1857 (N_1857,In_1686,In_1988);
nand U1858 (N_1858,In_2398,In_1121);
nand U1859 (N_1859,In_2140,In_866);
and U1860 (N_1860,In_458,In_2380);
nand U1861 (N_1861,In_981,In_2570);
nor U1862 (N_1862,In_1211,In_1163);
xnor U1863 (N_1863,In_2198,In_963);
or U1864 (N_1864,In_1558,In_263);
nor U1865 (N_1865,In_2476,In_2415);
nor U1866 (N_1866,In_592,In_65);
xor U1867 (N_1867,In_2386,In_2301);
or U1868 (N_1868,In_1085,In_1256);
and U1869 (N_1869,In_90,In_1759);
nand U1870 (N_1870,In_2175,In_1396);
nand U1871 (N_1871,In_2718,In_2604);
or U1872 (N_1872,In_503,In_294);
or U1873 (N_1873,In_1901,In_906);
nand U1874 (N_1874,In_1159,In_2506);
or U1875 (N_1875,In_1349,In_122);
nor U1876 (N_1876,In_2643,In_1055);
xor U1877 (N_1877,In_2576,In_2711);
xnor U1878 (N_1878,In_1518,In_1983);
or U1879 (N_1879,In_400,In_2944);
xor U1880 (N_1880,In_544,In_897);
and U1881 (N_1881,In_1102,In_1510);
nor U1882 (N_1882,In_1767,In_973);
nor U1883 (N_1883,In_989,In_1211);
nand U1884 (N_1884,In_2006,In_1675);
and U1885 (N_1885,In_1753,In_2158);
xnor U1886 (N_1886,In_1168,In_1490);
xnor U1887 (N_1887,In_1253,In_132);
nand U1888 (N_1888,In_1671,In_1607);
nor U1889 (N_1889,In_1940,In_1850);
nor U1890 (N_1890,In_2480,In_2539);
xor U1891 (N_1891,In_2209,In_1104);
and U1892 (N_1892,In_508,In_867);
nor U1893 (N_1893,In_2287,In_617);
or U1894 (N_1894,In_2205,In_2176);
or U1895 (N_1895,In_1367,In_1483);
xor U1896 (N_1896,In_2633,In_2564);
nor U1897 (N_1897,In_100,In_2164);
nand U1898 (N_1898,In_1673,In_2739);
nand U1899 (N_1899,In_1045,In_625);
and U1900 (N_1900,In_2854,In_2517);
nor U1901 (N_1901,In_1813,In_887);
or U1902 (N_1902,In_1856,In_1925);
and U1903 (N_1903,In_1349,In_1379);
nand U1904 (N_1904,In_1284,In_1135);
and U1905 (N_1905,In_2359,In_932);
xor U1906 (N_1906,In_402,In_2740);
xor U1907 (N_1907,In_2446,In_2092);
xor U1908 (N_1908,In_420,In_100);
nand U1909 (N_1909,In_2883,In_2662);
xnor U1910 (N_1910,In_2519,In_1428);
nor U1911 (N_1911,In_702,In_2748);
nor U1912 (N_1912,In_51,In_535);
xnor U1913 (N_1913,In_156,In_1623);
nand U1914 (N_1914,In_1268,In_2328);
and U1915 (N_1915,In_2280,In_2162);
nor U1916 (N_1916,In_1845,In_742);
xnor U1917 (N_1917,In_2718,In_1625);
nor U1918 (N_1918,In_1350,In_48);
nand U1919 (N_1919,In_2504,In_2823);
xor U1920 (N_1920,In_2604,In_2031);
or U1921 (N_1921,In_2637,In_920);
and U1922 (N_1922,In_2526,In_1570);
and U1923 (N_1923,In_396,In_498);
xnor U1924 (N_1924,In_2558,In_2659);
nor U1925 (N_1925,In_1857,In_1517);
nor U1926 (N_1926,In_826,In_2413);
and U1927 (N_1927,In_1481,In_205);
nor U1928 (N_1928,In_414,In_1086);
xor U1929 (N_1929,In_1659,In_1892);
nand U1930 (N_1930,In_2977,In_2551);
and U1931 (N_1931,In_433,In_2536);
xor U1932 (N_1932,In_2788,In_2781);
nand U1933 (N_1933,In_1005,In_2862);
or U1934 (N_1934,In_1408,In_2189);
nor U1935 (N_1935,In_1685,In_2543);
or U1936 (N_1936,In_350,In_2494);
xnor U1937 (N_1937,In_1599,In_695);
xnor U1938 (N_1938,In_1880,In_81);
xor U1939 (N_1939,In_199,In_2973);
nor U1940 (N_1940,In_2450,In_2041);
nor U1941 (N_1941,In_1211,In_206);
or U1942 (N_1942,In_2346,In_2995);
and U1943 (N_1943,In_2354,In_2976);
nand U1944 (N_1944,In_1778,In_170);
nand U1945 (N_1945,In_2524,In_1086);
nor U1946 (N_1946,In_2768,In_2019);
xnor U1947 (N_1947,In_555,In_1773);
xor U1948 (N_1948,In_1759,In_2898);
or U1949 (N_1949,In_1982,In_185);
or U1950 (N_1950,In_2396,In_743);
and U1951 (N_1951,In_48,In_2258);
nand U1952 (N_1952,In_789,In_2612);
nor U1953 (N_1953,In_1278,In_2079);
or U1954 (N_1954,In_2107,In_2934);
nand U1955 (N_1955,In_1988,In_865);
and U1956 (N_1956,In_1841,In_2757);
or U1957 (N_1957,In_140,In_1395);
nand U1958 (N_1958,In_1557,In_2709);
xor U1959 (N_1959,In_1206,In_2483);
and U1960 (N_1960,In_2706,In_335);
or U1961 (N_1961,In_1615,In_1026);
nand U1962 (N_1962,In_1611,In_2474);
nor U1963 (N_1963,In_330,In_2578);
nand U1964 (N_1964,In_2225,In_2337);
and U1965 (N_1965,In_2137,In_2220);
xnor U1966 (N_1966,In_1999,In_1031);
nand U1967 (N_1967,In_837,In_2708);
and U1968 (N_1968,In_2331,In_54);
or U1969 (N_1969,In_2661,In_2939);
nor U1970 (N_1970,In_1842,In_1358);
nand U1971 (N_1971,In_727,In_730);
xor U1972 (N_1972,In_2183,In_267);
or U1973 (N_1973,In_1535,In_459);
and U1974 (N_1974,In_532,In_846);
and U1975 (N_1975,In_1354,In_1985);
xnor U1976 (N_1976,In_2414,In_2624);
and U1977 (N_1977,In_615,In_736);
or U1978 (N_1978,In_1532,In_976);
and U1979 (N_1979,In_2395,In_328);
or U1980 (N_1980,In_2195,In_1816);
nand U1981 (N_1981,In_218,In_2294);
or U1982 (N_1982,In_97,In_578);
nand U1983 (N_1983,In_359,In_2895);
nor U1984 (N_1984,In_1151,In_451);
nor U1985 (N_1985,In_2856,In_1241);
xor U1986 (N_1986,In_786,In_1841);
nor U1987 (N_1987,In_2486,In_2915);
or U1988 (N_1988,In_61,In_721);
or U1989 (N_1989,In_790,In_2369);
nand U1990 (N_1990,In_415,In_182);
nor U1991 (N_1991,In_770,In_2267);
and U1992 (N_1992,In_1545,In_1178);
and U1993 (N_1993,In_480,In_2072);
or U1994 (N_1994,In_756,In_2684);
nand U1995 (N_1995,In_2790,In_1980);
or U1996 (N_1996,In_1622,In_68);
or U1997 (N_1997,In_2699,In_1101);
and U1998 (N_1998,In_2737,In_559);
nor U1999 (N_1999,In_298,In_2266);
and U2000 (N_2000,N_1362,N_167);
and U2001 (N_2001,N_1367,N_1402);
nor U2002 (N_2002,N_1633,N_419);
xnor U2003 (N_2003,N_546,N_1161);
or U2004 (N_2004,N_725,N_604);
xor U2005 (N_2005,N_1037,N_498);
or U2006 (N_2006,N_450,N_635);
nand U2007 (N_2007,N_839,N_1233);
and U2008 (N_2008,N_1414,N_1460);
nor U2009 (N_2009,N_873,N_978);
xor U2010 (N_2010,N_1648,N_1194);
xor U2011 (N_2011,N_732,N_1780);
nand U2012 (N_2012,N_742,N_1966);
or U2013 (N_2013,N_870,N_557);
nand U2014 (N_2014,N_1499,N_1464);
or U2015 (N_2015,N_108,N_503);
xor U2016 (N_2016,N_1897,N_388);
nor U2017 (N_2017,N_356,N_471);
or U2018 (N_2018,N_1811,N_306);
and U2019 (N_2019,N_1721,N_1116);
and U2020 (N_2020,N_1702,N_0);
nor U2021 (N_2021,N_393,N_1436);
and U2022 (N_2022,N_1025,N_1147);
or U2023 (N_2023,N_1355,N_1538);
xnor U2024 (N_2024,N_689,N_355);
and U2025 (N_2025,N_533,N_134);
or U2026 (N_2026,N_1442,N_943);
xor U2027 (N_2027,N_1909,N_1701);
and U2028 (N_2028,N_1497,N_938);
nand U2029 (N_2029,N_1176,N_921);
nand U2030 (N_2030,N_762,N_550);
nand U2031 (N_2031,N_822,N_884);
nor U2032 (N_2032,N_484,N_1934);
xnor U2033 (N_2033,N_1047,N_900);
nand U2034 (N_2034,N_1345,N_705);
nand U2035 (N_2035,N_1220,N_1566);
nand U2036 (N_2036,N_708,N_1576);
and U2037 (N_2037,N_1583,N_432);
xor U2038 (N_2038,N_928,N_109);
nor U2039 (N_2039,N_1311,N_967);
xnor U2040 (N_2040,N_1188,N_200);
nor U2041 (N_2041,N_605,N_723);
nand U2042 (N_2042,N_1670,N_1268);
nor U2043 (N_2043,N_1288,N_1498);
or U2044 (N_2044,N_1554,N_1055);
or U2045 (N_2045,N_767,N_524);
nand U2046 (N_2046,N_495,N_963);
nand U2047 (N_2047,N_1745,N_706);
or U2048 (N_2048,N_1800,N_1927);
or U2049 (N_2049,N_774,N_1998);
xnor U2050 (N_2050,N_422,N_631);
xor U2051 (N_2051,N_1912,N_1654);
xnor U2052 (N_2052,N_1947,N_812);
and U2053 (N_2053,N_1327,N_441);
and U2054 (N_2054,N_407,N_1663);
or U2055 (N_2055,N_1871,N_1712);
and U2056 (N_2056,N_1431,N_1257);
nor U2057 (N_2057,N_1786,N_1420);
nand U2058 (N_2058,N_1724,N_786);
nor U2059 (N_2059,N_1038,N_855);
and U2060 (N_2060,N_1517,N_59);
xnor U2061 (N_2061,N_1335,N_724);
xor U2062 (N_2062,N_1853,N_618);
nor U2063 (N_2063,N_1006,N_1710);
xnor U2064 (N_2064,N_621,N_1491);
nand U2065 (N_2065,N_1103,N_100);
xnor U2066 (N_2066,N_798,N_199);
or U2067 (N_2067,N_1486,N_41);
or U2068 (N_2068,N_1946,N_1060);
and U2069 (N_2069,N_353,N_684);
xor U2070 (N_2070,N_1151,N_1597);
nor U2071 (N_2071,N_212,N_1753);
nor U2072 (N_2072,N_656,N_1155);
nand U2073 (N_2073,N_1048,N_184);
xor U2074 (N_2074,N_1564,N_1412);
or U2075 (N_2075,N_1072,N_61);
or U2076 (N_2076,N_1634,N_1529);
nand U2077 (N_2077,N_1354,N_329);
nor U2078 (N_2078,N_1348,N_114);
nor U2079 (N_2079,N_367,N_747);
nor U2080 (N_2080,N_1146,N_1924);
xnor U2081 (N_2081,N_1477,N_834);
or U2082 (N_2082,N_70,N_647);
or U2083 (N_2083,N_1427,N_517);
nand U2084 (N_2084,N_1352,N_330);
and U2085 (N_2085,N_315,N_1300);
or U2086 (N_2086,N_1870,N_865);
xnor U2087 (N_2087,N_346,N_248);
and U2088 (N_2088,N_1205,N_316);
or U2089 (N_2089,N_1957,N_1678);
xor U2090 (N_2090,N_402,N_1627);
and U2091 (N_2091,N_433,N_719);
nand U2092 (N_2092,N_290,N_587);
nand U2093 (N_2093,N_1112,N_147);
nand U2094 (N_2094,N_1852,N_997);
nand U2095 (N_2095,N_344,N_118);
nor U2096 (N_2096,N_780,N_141);
and U2097 (N_2097,N_1245,N_1942);
or U2098 (N_2098,N_790,N_1388);
or U2099 (N_2099,N_1804,N_673);
xnor U2100 (N_2100,N_1567,N_405);
xor U2101 (N_2101,N_813,N_1299);
xor U2102 (N_2102,N_1138,N_752);
and U2103 (N_2103,N_1131,N_1651);
nor U2104 (N_2104,N_664,N_727);
nand U2105 (N_2105,N_85,N_718);
nor U2106 (N_2106,N_1750,N_321);
nand U2107 (N_2107,N_1244,N_1238);
nor U2108 (N_2108,N_867,N_1900);
nor U2109 (N_2109,N_1172,N_1046);
nor U2110 (N_2110,N_609,N_71);
xor U2111 (N_2111,N_992,N_259);
and U2112 (N_2112,N_166,N_821);
xnor U2113 (N_2113,N_75,N_262);
nor U2114 (N_2114,N_96,N_806);
and U2115 (N_2115,N_815,N_1150);
nand U2116 (N_2116,N_445,N_155);
xnor U2117 (N_2117,N_87,N_1778);
xor U2118 (N_2118,N_714,N_1237);
and U2119 (N_2119,N_1384,N_580);
xor U2120 (N_2120,N_1704,N_734);
or U2121 (N_2121,N_281,N_913);
nor U2122 (N_2122,N_585,N_1630);
or U2123 (N_2123,N_1674,N_1365);
xor U2124 (N_2124,N_894,N_1126);
or U2125 (N_2125,N_304,N_1655);
xor U2126 (N_2126,N_1514,N_1984);
nand U2127 (N_2127,N_804,N_738);
nand U2128 (N_2128,N_983,N_1227);
or U2129 (N_2129,N_1665,N_680);
xor U2130 (N_2130,N_240,N_1313);
and U2131 (N_2131,N_1628,N_532);
or U2132 (N_2132,N_800,N_643);
and U2133 (N_2133,N_567,N_171);
nor U2134 (N_2134,N_982,N_7);
or U2135 (N_2135,N_47,N_1624);
nand U2136 (N_2136,N_1470,N_1504);
and U2137 (N_2137,N_612,N_1242);
nor U2138 (N_2138,N_961,N_444);
nand U2139 (N_2139,N_1179,N_726);
nand U2140 (N_2140,N_1001,N_794);
or U2141 (N_2141,N_364,N_799);
nand U2142 (N_2142,N_335,N_1404);
nor U2143 (N_2143,N_1808,N_1344);
nor U2144 (N_2144,N_1254,N_901);
and U2145 (N_2145,N_1454,N_951);
nor U2146 (N_2146,N_896,N_654);
nor U2147 (N_2147,N_835,N_1203);
or U2148 (N_2148,N_1111,N_1434);
and U2149 (N_2149,N_1209,N_1260);
or U2150 (N_2150,N_373,N_845);
xnor U2151 (N_2151,N_1002,N_1931);
nor U2152 (N_2152,N_1908,N_1976);
nand U2153 (N_2153,N_1988,N_1145);
nor U2154 (N_2154,N_18,N_1773);
and U2155 (N_2155,N_1835,N_1094);
xor U2156 (N_2156,N_516,N_146);
nand U2157 (N_2157,N_831,N_1453);
xor U2158 (N_2158,N_544,N_1088);
xnor U2159 (N_2159,N_1280,N_1895);
xnor U2160 (N_2160,N_236,N_1573);
and U2161 (N_2161,N_970,N_926);
and U2162 (N_2162,N_1973,N_1379);
and U2163 (N_2163,N_431,N_197);
nor U2164 (N_2164,N_1793,N_670);
or U2165 (N_2165,N_1815,N_1789);
or U2166 (N_2166,N_1932,N_552);
xnor U2167 (N_2167,N_424,N_500);
nor U2168 (N_2168,N_1798,N_525);
nor U2169 (N_2169,N_1887,N_1039);
nor U2170 (N_2170,N_1381,N_1500);
and U2171 (N_2171,N_1440,N_1303);
or U2172 (N_2172,N_1547,N_1309);
nand U2173 (N_2173,N_1019,N_230);
and U2174 (N_2174,N_101,N_1940);
xnor U2175 (N_2175,N_1409,N_519);
and U2176 (N_2176,N_1955,N_1078);
nand U2177 (N_2177,N_572,N_404);
and U2178 (N_2178,N_129,N_1671);
xnor U2179 (N_2179,N_269,N_350);
and U2180 (N_2180,N_1575,N_1452);
nor U2181 (N_2181,N_940,N_1021);
and U2182 (N_2182,N_115,N_14);
nand U2183 (N_2183,N_953,N_123);
and U2184 (N_2184,N_1441,N_176);
nor U2185 (N_2185,N_298,N_465);
and U2186 (N_2186,N_1861,N_297);
and U2187 (N_2187,N_1411,N_784);
and U2188 (N_2188,N_1492,N_1247);
or U2189 (N_2189,N_1321,N_1694);
xnor U2190 (N_2190,N_850,N_1034);
xnor U2191 (N_2191,N_887,N_1980);
nand U2192 (N_2192,N_1168,N_1757);
nand U2193 (N_2193,N_1307,N_1368);
nor U2194 (N_2194,N_944,N_79);
nor U2195 (N_2195,N_1264,N_562);
nor U2196 (N_2196,N_1546,N_1765);
and U2197 (N_2197,N_1982,N_861);
or U2198 (N_2198,N_663,N_1814);
and U2199 (N_2199,N_1568,N_1169);
nand U2200 (N_2200,N_1649,N_1532);
and U2201 (N_2201,N_1480,N_158);
xor U2202 (N_2202,N_1974,N_694);
or U2203 (N_2203,N_235,N_1221);
or U2204 (N_2204,N_1278,N_1201);
nand U2205 (N_2205,N_1585,N_229);
or U2206 (N_2206,N_29,N_1621);
nor U2207 (N_2207,N_1347,N_1036);
or U2208 (N_2208,N_1401,N_1403);
nand U2209 (N_2209,N_156,N_1135);
and U2210 (N_2210,N_1999,N_1087);
xnor U2211 (N_2211,N_1228,N_1236);
nor U2212 (N_2212,N_1166,N_1137);
or U2213 (N_2213,N_83,N_310);
or U2214 (N_2214,N_177,N_1139);
xor U2215 (N_2215,N_1050,N_435);
or U2216 (N_2216,N_927,N_384);
xor U2217 (N_2217,N_678,N_1803);
xnor U2218 (N_2218,N_1995,N_905);
xor U2219 (N_2219,N_791,N_261);
nor U2220 (N_2220,N_1259,N_1356);
and U2221 (N_2221,N_716,N_193);
nand U2222 (N_2222,N_1959,N_324);
nand U2223 (N_2223,N_1759,N_763);
xor U2224 (N_2224,N_531,N_276);
nor U2225 (N_2225,N_1856,N_1595);
or U2226 (N_2226,N_897,N_775);
nor U2227 (N_2227,N_1657,N_1462);
xnor U2228 (N_2228,N_860,N_1969);
nand U2229 (N_2229,N_907,N_736);
and U2230 (N_2230,N_1590,N_257);
nand U2231 (N_2231,N_1057,N_1588);
or U2232 (N_2232,N_871,N_617);
or U2233 (N_2233,N_40,N_1734);
nand U2234 (N_2234,N_497,N_929);
and U2235 (N_2235,N_1593,N_1424);
nor U2236 (N_2236,N_1016,N_1467);
nor U2237 (N_2237,N_258,N_614);
xor U2238 (N_2238,N_1574,N_345);
nand U2239 (N_2239,N_106,N_1239);
nand U2240 (N_2240,N_1558,N_999);
nor U2241 (N_2241,N_1693,N_1482);
nor U2242 (N_2242,N_1073,N_1490);
and U2243 (N_2243,N_1519,N_457);
and U2244 (N_2244,N_157,N_296);
nand U2245 (N_2245,N_998,N_1422);
or U2246 (N_2246,N_1026,N_1043);
and U2247 (N_2247,N_299,N_1809);
and U2248 (N_2248,N_1457,N_1881);
nor U2249 (N_2249,N_209,N_893);
and U2250 (N_2250,N_148,N_1761);
nor U2251 (N_2251,N_1539,N_13);
xor U2252 (N_2252,N_1177,N_89);
xnor U2253 (N_2253,N_730,N_1996);
xnor U2254 (N_2254,N_1965,N_172);
or U2255 (N_2255,N_667,N_506);
nor U2256 (N_2256,N_1874,N_1613);
nand U2257 (N_2257,N_1031,N_1680);
or U2258 (N_2258,N_326,N_472);
and U2259 (N_2259,N_162,N_1731);
or U2260 (N_2260,N_1503,N_189);
xor U2261 (N_2261,N_1275,N_826);
and U2262 (N_2262,N_1869,N_877);
and U2263 (N_2263,N_1906,N_1415);
or U2264 (N_2264,N_119,N_17);
and U2265 (N_2265,N_221,N_220);
nand U2266 (N_2266,N_672,N_1698);
nand U2267 (N_2267,N_1611,N_755);
nor U2268 (N_2268,N_607,N_1208);
and U2269 (N_2269,N_841,N_782);
nor U2270 (N_2270,N_263,N_543);
xnor U2271 (N_2271,N_1159,N_246);
or U2272 (N_2272,N_638,N_561);
or U2273 (N_2273,N_1448,N_1069);
nand U2274 (N_2274,N_1173,N_688);
or U2275 (N_2275,N_67,N_1729);
and U2276 (N_2276,N_662,N_76);
nand U2277 (N_2277,N_278,N_869);
nand U2278 (N_2278,N_1056,N_1860);
or U2279 (N_2279,N_1782,N_323);
or U2280 (N_2280,N_1846,N_1748);
nand U2281 (N_2281,N_1580,N_675);
xnor U2282 (N_2282,N_279,N_154);
xor U2283 (N_2283,N_1594,N_187);
and U2284 (N_2284,N_1035,N_912);
nor U2285 (N_2285,N_528,N_611);
nor U2286 (N_2286,N_1825,N_778);
and U2287 (N_2287,N_63,N_753);
and U2288 (N_2288,N_112,N_908);
xor U2289 (N_2289,N_254,N_1127);
nand U2290 (N_2290,N_421,N_1779);
xor U2291 (N_2291,N_1262,N_1143);
xor U2292 (N_2292,N_876,N_682);
and U2293 (N_2293,N_1391,N_590);
and U2294 (N_2294,N_426,N_879);
nor U2295 (N_2295,N_1892,N_1707);
or U2296 (N_2296,N_935,N_216);
xnor U2297 (N_2297,N_1061,N_1374);
nand U2298 (N_2298,N_1185,N_549);
nand U2299 (N_2299,N_1096,N_124);
nand U2300 (N_2300,N_792,N_1224);
xor U2301 (N_2301,N_1746,N_423);
xor U2302 (N_2302,N_1938,N_526);
or U2303 (N_2303,N_1136,N_1322);
xnor U2304 (N_2304,N_286,N_1880);
xnor U2305 (N_2305,N_1487,N_1992);
or U2306 (N_2306,N_624,N_341);
nand U2307 (N_2307,N_1725,N_1534);
or U2308 (N_2308,N_1466,N_681);
and U2309 (N_2309,N_1560,N_43);
nor U2310 (N_2310,N_652,N_1591);
nor U2311 (N_2311,N_251,N_237);
xnor U2312 (N_2312,N_1653,N_899);
nor U2313 (N_2313,N_622,N_513);
or U2314 (N_2314,N_343,N_1925);
xnor U2315 (N_2315,N_1586,N_1720);
nor U2316 (N_2316,N_1733,N_1600);
nor U2317 (N_2317,N_483,N_1785);
nand U2318 (N_2318,N_1225,N_1766);
nor U2319 (N_2319,N_1306,N_50);
and U2320 (N_2320,N_1375,N_1989);
nor U2321 (N_2321,N_1456,N_1783);
nand U2322 (N_2322,N_936,N_11);
nand U2323 (N_2323,N_1181,N_1418);
or U2324 (N_2324,N_842,N_383);
and U2325 (N_2325,N_159,N_1749);
nand U2326 (N_2326,N_186,N_1609);
nand U2327 (N_2327,N_854,N_358);
nor U2328 (N_2328,N_1338,N_1692);
nand U2329 (N_2329,N_922,N_857);
nand U2330 (N_2330,N_173,N_406);
nand U2331 (N_2331,N_1620,N_1637);
nand U2332 (N_2332,N_447,N_1963);
nand U2333 (N_2333,N_989,N_756);
nand U2334 (N_2334,N_1439,N_375);
and U2335 (N_2335,N_1830,N_1937);
xor U2336 (N_2336,N_553,N_440);
or U2337 (N_2337,N_228,N_287);
nand U2338 (N_2338,N_777,N_515);
nor U2339 (N_2339,N_1857,N_213);
nand U2340 (N_2340,N_371,N_1319);
nor U2341 (N_2341,N_16,N_1000);
or U2342 (N_2342,N_1122,N_1059);
nor U2343 (N_2343,N_45,N_1961);
nor U2344 (N_2344,N_518,N_231);
xnor U2345 (N_2345,N_1008,N_19);
xor U2346 (N_2346,N_1396,N_1862);
xnor U2347 (N_2347,N_1863,N_1033);
nor U2348 (N_2348,N_110,N_1183);
nor U2349 (N_2349,N_1935,N_764);
and U2350 (N_2350,N_1582,N_1289);
nand U2351 (N_2351,N_223,N_1258);
nand U2352 (N_2352,N_302,N_1756);
or U2353 (N_2353,N_1304,N_205);
nor U2354 (N_2354,N_874,N_1235);
nor U2355 (N_2355,N_1317,N_1616);
or U2356 (N_2356,N_1618,N_735);
xnor U2357 (N_2357,N_1241,N_1281);
or U2358 (N_2358,N_1521,N_594);
nand U2359 (N_2359,N_277,N_713);
nor U2360 (N_2360,N_847,N_448);
nand U2361 (N_2361,N_981,N_1902);
xnor U2362 (N_2362,N_1629,N_1681);
nor U2363 (N_2363,N_807,N_1661);
and U2364 (N_2364,N_204,N_1430);
nor U2365 (N_2365,N_957,N_1831);
xnor U2366 (N_2366,N_1421,N_895);
and U2367 (N_2367,N_362,N_573);
or U2368 (N_2368,N_66,N_1287);
and U2369 (N_2369,N_1105,N_1858);
xor U2370 (N_2370,N_1787,N_872);
nor U2371 (N_2371,N_1842,N_195);
or U2372 (N_2372,N_245,N_260);
or U2373 (N_2373,N_1876,N_1544);
nand U2374 (N_2374,N_1587,N_1119);
or U2375 (N_2375,N_456,N_1550);
nand U2376 (N_2376,N_389,N_1769);
nand U2377 (N_2377,N_107,N_674);
and U2378 (N_2378,N_458,N_210);
and U2379 (N_2379,N_1124,N_293);
nor U2380 (N_2380,N_1107,N_948);
nand U2381 (N_2381,N_1893,N_1443);
or U2382 (N_2382,N_1271,N_1113);
xor U2383 (N_2383,N_411,N_1751);
nand U2384 (N_2384,N_632,N_1606);
and U2385 (N_2385,N_1141,N_1638);
nor U2386 (N_2386,N_1024,N_1685);
xnor U2387 (N_2387,N_1872,N_1030);
or U2388 (N_2388,N_395,N_1525);
nor U2389 (N_2389,N_428,N_226);
xnor U2390 (N_2390,N_95,N_15);
or U2391 (N_2391,N_491,N_1945);
and U2392 (N_2392,N_394,N_130);
and U2393 (N_2393,N_88,N_1397);
or U2394 (N_2394,N_194,N_593);
nand U2395 (N_2395,N_1747,N_1350);
xnor U2396 (N_2396,N_1070,N_1604);
and U2397 (N_2397,N_127,N_606);
nand U2398 (N_2398,N_1577,N_945);
or U2399 (N_2399,N_280,N_1833);
or U2400 (N_2400,N_1433,N_336);
nand U2401 (N_2401,N_462,N_1919);
xnor U2402 (N_2402,N_771,N_1752);
nand U2403 (N_2403,N_564,N_1913);
and U2404 (N_2404,N_1053,N_904);
nand U2405 (N_2405,N_704,N_1066);
and U2406 (N_2406,N_478,N_1474);
xnor U2407 (N_2407,N_429,N_1154);
nand U2408 (N_2408,N_830,N_868);
nor U2409 (N_2409,N_1417,N_247);
nand U2410 (N_2410,N_1346,N_840);
nor U2411 (N_2411,N_1206,N_1283);
xor U2412 (N_2412,N_542,N_1843);
nor U2413 (N_2413,N_1571,N_1635);
xnor U2414 (N_2414,N_766,N_1435);
xor U2415 (N_2415,N_271,N_668);
nand U2416 (N_2416,N_1719,N_1904);
and U2417 (N_2417,N_192,N_1543);
and U2418 (N_2418,N_642,N_1438);
and U2419 (N_2419,N_1011,N_313);
and U2420 (N_2420,N_1082,N_1512);
nor U2421 (N_2421,N_1741,N_1953);
or U2422 (N_2422,N_1405,N_1885);
or U2423 (N_2423,N_480,N_627);
xnor U2424 (N_2424,N_1496,N_268);
or U2425 (N_2425,N_1389,N_238);
nand U2426 (N_2426,N_748,N_1907);
xnor U2427 (N_2427,N_1475,N_1642);
xor U2428 (N_2428,N_398,N_334);
and U2429 (N_2429,N_97,N_1709);
or U2430 (N_2430,N_1644,N_648);
and U2431 (N_2431,N_952,N_691);
xor U2432 (N_2432,N_1625,N_653);
or U2433 (N_2433,N_849,N_933);
and U2434 (N_2434,N_1723,N_828);
nor U2435 (N_2435,N_274,N_1393);
or U2436 (N_2436,N_303,N_1559);
or U2437 (N_2437,N_1180,N_715);
and U2438 (N_2438,N_529,N_852);
nand U2439 (N_2439,N_434,N_468);
or U2440 (N_2440,N_1607,N_1297);
or U2441 (N_2441,N_486,N_349);
or U2442 (N_2442,N_1518,N_1052);
and U2443 (N_2443,N_1058,N_1357);
and U2444 (N_2444,N_1691,N_150);
nor U2445 (N_2445,N_968,N_733);
or U2446 (N_2446,N_862,N_1358);
nor U2447 (N_2447,N_1555,N_479);
nand U2448 (N_2448,N_102,N_1884);
nor U2449 (N_2449,N_244,N_1832);
nand U2450 (N_2450,N_98,N_520);
and U2451 (N_2451,N_1063,N_82);
and U2452 (N_2452,N_721,N_985);
nor U2453 (N_2453,N_1570,N_233);
nor U2454 (N_2454,N_1549,N_630);
nand U2455 (N_2455,N_490,N_1032);
nor U2456 (N_2456,N_1369,N_53);
and U2457 (N_2457,N_1987,N_939);
xnor U2458 (N_2458,N_1592,N_702);
or U2459 (N_2459,N_1469,N_545);
nand U2460 (N_2460,N_988,N_1584);
xnor U2461 (N_2461,N_320,N_460);
or U2462 (N_2462,N_1410,N_1810);
nand U2463 (N_2463,N_400,N_1398);
xnor U2464 (N_2464,N_750,N_931);
and U2465 (N_2465,N_1643,N_986);
nand U2466 (N_2466,N_234,N_1171);
or U2467 (N_2467,N_1041,N_655);
nand U2468 (N_2468,N_1234,N_991);
xnor U2469 (N_2469,N_1728,N_1153);
nor U2470 (N_2470,N_1372,N_1075);
xor U2471 (N_2471,N_1323,N_1199);
nor U2472 (N_2472,N_796,N_1197);
or U2473 (N_2473,N_1210,N_417);
nand U2474 (N_2474,N_1730,N_496);
nand U2475 (N_2475,N_591,N_1805);
xnor U2476 (N_2476,N_352,N_163);
or U2477 (N_2477,N_401,N_1979);
nand U2478 (N_2478,N_695,N_26);
nor U2479 (N_2479,N_683,N_273);
nor U2480 (N_2480,N_348,N_1950);
or U2481 (N_2481,N_1463,N_788);
or U2482 (N_2482,N_1156,N_161);
xor U2483 (N_2483,N_1949,N_1214);
and U2484 (N_2484,N_1764,N_1615);
xor U2485 (N_2485,N_20,N_709);
nand U2486 (N_2486,N_787,N_1797);
nand U2487 (N_2487,N_720,N_1596);
and U2488 (N_2488,N_722,N_390);
and U2489 (N_2489,N_99,N_1286);
or U2490 (N_2490,N_1777,N_443);
xnor U2491 (N_2491,N_1511,N_144);
nand U2492 (N_2492,N_1461,N_225);
or U2493 (N_2493,N_1478,N_396);
and U2494 (N_2494,N_1376,N_759);
xnor U2495 (N_2495,N_1196,N_308);
or U2496 (N_2496,N_598,N_1978);
xor U2497 (N_2497,N_1636,N_1207);
nand U2498 (N_2498,N_418,N_1695);
nand U2499 (N_2499,N_892,N_937);
nand U2500 (N_2500,N_917,N_1130);
or U2501 (N_2501,N_693,N_789);
xnor U2502 (N_2502,N_1383,N_880);
or U2503 (N_2503,N_578,N_1110);
or U2504 (N_2504,N_744,N_1293);
nand U2505 (N_2505,N_1867,N_427);
and U2506 (N_2506,N_436,N_1922);
xor U2507 (N_2507,N_1144,N_116);
and U2508 (N_2508,N_555,N_536);
or U2509 (N_2509,N_1699,N_601);
and U2510 (N_2510,N_558,N_888);
xor U2511 (N_2511,N_1385,N_252);
nand U2512 (N_2512,N_284,N_960);
or U2513 (N_2513,N_1847,N_1666);
or U2514 (N_2514,N_1152,N_267);
nand U2515 (N_2515,N_333,N_1315);
nand U2516 (N_2516,N_575,N_1109);
nand U2517 (N_2517,N_902,N_838);
xnor U2518 (N_2518,N_10,N_1314);
nand U2519 (N_2519,N_1432,N_690);
nand U2520 (N_2520,N_574,N_474);
and U2521 (N_2521,N_699,N_174);
nor U2522 (N_2522,N_1619,N_21);
nor U2523 (N_2523,N_547,N_534);
nor U2524 (N_2524,N_1971,N_1334);
nor U2525 (N_2525,N_1471,N_844);
nand U2526 (N_2526,N_1958,N_947);
and U2527 (N_2527,N_1090,N_1023);
or U2528 (N_2528,N_1569,N_1123);
nand U2529 (N_2529,N_1530,N_1074);
xor U2530 (N_2530,N_1551,N_23);
nand U2531 (N_2531,N_1711,N_1740);
nand U2532 (N_2532,N_1080,N_1732);
or U2533 (N_2533,N_1284,N_1267);
and U2534 (N_2534,N_1667,N_27);
and U2535 (N_2535,N_1017,N_541);
nor U2536 (N_2536,N_1195,N_1775);
or U2537 (N_2537,N_1437,N_958);
and U2538 (N_2538,N_1563,N_816);
and U2539 (N_2539,N_946,N_1445);
and U2540 (N_2540,N_1515,N_1631);
xnor U2541 (N_2541,N_1255,N_386);
xor U2542 (N_2542,N_1509,N_1784);
nand U2543 (N_2543,N_104,N_1859);
xnor U2544 (N_2544,N_1483,N_291);
nand U2545 (N_2545,N_1994,N_1820);
or U2546 (N_2546,N_1792,N_1817);
and U2547 (N_2547,N_1382,N_1085);
xnor U2548 (N_2548,N_1878,N_1308);
nand U2549 (N_2549,N_743,N_1877);
or U2550 (N_2550,N_145,N_1951);
nand U2551 (N_2551,N_1829,N_363);
or U2552 (N_2552,N_86,N_1873);
nand U2553 (N_2553,N_1968,N_1488);
or U2554 (N_2554,N_941,N_640);
and U2555 (N_2555,N_1602,N_824);
and U2556 (N_2556,N_1706,N_1557);
nand U2557 (N_2557,N_1481,N_382);
nor U2558 (N_2558,N_376,N_42);
nor U2559 (N_2559,N_325,N_1230);
or U2560 (N_2560,N_1472,N_266);
and U2561 (N_2561,N_121,N_739);
nor U2562 (N_2562,N_493,N_1222);
xor U2563 (N_2563,N_208,N_451);
and U2564 (N_2564,N_1249,N_165);
nor U2565 (N_2565,N_1104,N_751);
and U2566 (N_2566,N_1875,N_1589);
or U2567 (N_2567,N_1890,N_476);
or U2568 (N_2568,N_322,N_795);
and U2569 (N_2569,N_46,N_1395);
and U2570 (N_2570,N_1022,N_6);
or U2571 (N_2571,N_360,N_1622);
nor U2572 (N_2572,N_1028,N_911);
nand U2573 (N_2573,N_599,N_760);
xnor U2574 (N_2574,N_1337,N_1077);
or U2575 (N_2575,N_971,N_539);
xnor U2576 (N_2576,N_819,N_1459);
nand U2577 (N_2577,N_1868,N_377);
nand U2578 (N_2578,N_8,N_105);
xor U2579 (N_2579,N_569,N_318);
nand U2580 (N_2580,N_1049,N_4);
and U2581 (N_2581,N_962,N_608);
xor U2582 (N_2582,N_1390,N_188);
or U2583 (N_2583,N_69,N_671);
nor U2584 (N_2584,N_1010,N_1894);
nand U2585 (N_2585,N_381,N_1416);
and U2586 (N_2586,N_214,N_754);
nand U2587 (N_2587,N_1578,N_1495);
nor U2588 (N_2588,N_701,N_1213);
and U2589 (N_2589,N_665,N_1310);
and U2590 (N_2590,N_1605,N_1067);
nand U2591 (N_2591,N_758,N_1330);
nand U2592 (N_2592,N_776,N_919);
nor U2593 (N_2593,N_1541,N_22);
or U2594 (N_2594,N_1363,N_1891);
or U2595 (N_2595,N_1333,N_1167);
and U2596 (N_2596,N_1274,N_1688);
nor U2597 (N_2597,N_201,N_1647);
nand U2598 (N_2598,N_773,N_1943);
xnor U2599 (N_2599,N_9,N_469);
nor U2600 (N_2600,N_1479,N_117);
and U2601 (N_2601,N_697,N_446);
and U2602 (N_2602,N_1342,N_1282);
or U2603 (N_2603,N_626,N_73);
or U2604 (N_2604,N_1505,N_379);
nor U2605 (N_2605,N_1531,N_920);
nor U2606 (N_2606,N_950,N_169);
nor U2607 (N_2607,N_331,N_915);
nand U2608 (N_2608,N_793,N_749);
nor U2609 (N_2609,N_1659,N_805);
xor U2610 (N_2610,N_1926,N_185);
xor U2611 (N_2611,N_783,N_1755);
nor U2612 (N_2612,N_875,N_1668);
xor U2613 (N_2613,N_620,N_1014);
nand U2614 (N_2614,N_1211,N_1447);
and U2615 (N_2615,N_1494,N_576);
nor U2616 (N_2616,N_1834,N_35);
and U2617 (N_2617,N_136,N_1713);
or U2618 (N_2618,N_292,N_634);
or U2619 (N_2619,N_239,N_1331);
nor U2620 (N_2620,N_1776,N_600);
nor U2621 (N_2621,N_918,N_942);
nor U2622 (N_2622,N_582,N_1182);
and U2623 (N_2623,N_1983,N_275);
nand U2624 (N_2624,N_55,N_811);
and U2625 (N_2625,N_1850,N_1425);
nor U2626 (N_2626,N_1009,N_581);
nand U2627 (N_2627,N_1690,N_1295);
and U2628 (N_2628,N_283,N_241);
nand U2629 (N_2629,N_1361,N_1142);
xnor U2630 (N_2630,N_551,N_1990);
or U2631 (N_2631,N_781,N_1276);
xnor U2632 (N_2632,N_1763,N_1535);
nor U2633 (N_2633,N_1682,N_1332);
and U2634 (N_2634,N_589,N_1423);
or U2635 (N_2635,N_1632,N_1336);
and U2636 (N_2636,N_1889,N_975);
nand U2637 (N_2637,N_898,N_470);
nand U2638 (N_2638,N_1370,N_215);
or U2639 (N_2639,N_1537,N_1098);
and U2640 (N_2640,N_499,N_1449);
nand U2641 (N_2641,N_1302,N_803);
nand U2642 (N_2642,N_1045,N_1272);
and U2643 (N_2643,N_60,N_1086);
or U2644 (N_2644,N_1163,N_540);
nor U2645 (N_2645,N_1933,N_1226);
nor U2646 (N_2646,N_645,N_1455);
and U2647 (N_2647,N_1324,N_658);
and U2648 (N_2648,N_1526,N_696);
and U2649 (N_2649,N_437,N_613);
nand U2650 (N_2650,N_916,N_1903);
xor U2651 (N_2651,N_1044,N_282);
or U2652 (N_2652,N_1738,N_1791);
or U2653 (N_2653,N_1216,N_1328);
or U2654 (N_2654,N_442,N_973);
nor U2655 (N_2655,N_837,N_1824);
or U2656 (N_2656,N_1836,N_38);
nand U2657 (N_2657,N_481,N_1528);
nor U2658 (N_2658,N_856,N_1378);
xor U2659 (N_2659,N_1380,N_338);
nor U2660 (N_2660,N_1744,N_1298);
and U2661 (N_2661,N_1837,N_925);
xor U2662 (N_2662,N_387,N_1664);
xor U2663 (N_2663,N_1520,N_1742);
xnor U2664 (N_2664,N_361,N_909);
or U2665 (N_2665,N_1772,N_1914);
and U2666 (N_2666,N_179,N_1818);
or U2667 (N_2667,N_1552,N_1929);
and U2668 (N_2668,N_1641,N_385);
xor U2669 (N_2669,N_833,N_1318);
nand U2670 (N_2670,N_910,N_563);
and U2671 (N_2671,N_138,N_126);
nor U2672 (N_2672,N_464,N_974);
nand U2673 (N_2673,N_615,N_965);
nor U2674 (N_2674,N_1164,N_891);
nand U2675 (N_2675,N_463,N_858);
nand U2676 (N_2676,N_1650,N_1051);
nand U2677 (N_2677,N_1076,N_122);
or U2678 (N_2678,N_1160,N_554);
nand U2679 (N_2679,N_977,N_1465);
nor U2680 (N_2680,N_3,N_1232);
and U2681 (N_2681,N_374,N_1387);
or U2682 (N_2682,N_657,N_242);
nand U2683 (N_2683,N_160,N_808);
nand U2684 (N_2684,N_556,N_1849);
or U2685 (N_2685,N_140,N_37);
xnor U2686 (N_2686,N_1083,N_851);
nor U2687 (N_2687,N_132,N_196);
and U2688 (N_2688,N_1204,N_741);
nand U2689 (N_2689,N_1134,N_1093);
xor U2690 (N_2690,N_596,N_131);
and U2691 (N_2691,N_761,N_906);
nand U2692 (N_2692,N_1265,N_932);
nor U2693 (N_2693,N_319,N_1428);
nor U2694 (N_2694,N_178,N_661);
nand U2695 (N_2695,N_817,N_289);
or U2696 (N_2696,N_1985,N_1012);
nand U2697 (N_2697,N_583,N_452);
nor U2698 (N_2698,N_1855,N_1279);
xor U2699 (N_2699,N_1450,N_1);
and U2700 (N_2700,N_1506,N_164);
nor U2701 (N_2701,N_1918,N_1601);
or U2702 (N_2702,N_1645,N_48);
and U2703 (N_2703,N_1277,N_1610);
and U2704 (N_2704,N_466,N_301);
nor U2705 (N_2705,N_1243,N_1882);
xnor U2706 (N_2706,N_133,N_494);
nor U2707 (N_2707,N_1218,N_505);
nor U2708 (N_2708,N_1071,N_190);
nand U2709 (N_2709,N_1097,N_646);
nand U2710 (N_2710,N_183,N_1320);
and U2711 (N_2711,N_692,N_878);
and U2712 (N_2712,N_625,N_168);
or U2713 (N_2713,N_224,N_1936);
nor U2714 (N_2714,N_328,N_603);
nor U2715 (N_2715,N_1042,N_1928);
nand U2716 (N_2716,N_80,N_300);
nand U2717 (N_2717,N_1305,N_203);
or U2718 (N_2718,N_757,N_1184);
xor U2719 (N_2719,N_1801,N_1770);
nand U2720 (N_2720,N_307,N_1339);
nor U2721 (N_2721,N_1175,N_1905);
and U2722 (N_2722,N_256,N_1954);
or U2723 (N_2723,N_430,N_1312);
nand U2724 (N_2724,N_592,N_669);
xor U2725 (N_2725,N_1091,N_511);
nand U2726 (N_2726,N_1102,N_12);
or U2727 (N_2727,N_1726,N_1451);
nand U2728 (N_2728,N_619,N_537);
nor U2729 (N_2729,N_56,N_1399);
or U2730 (N_2730,N_1827,N_1697);
and U2731 (N_2731,N_1029,N_111);
xor U2732 (N_2732,N_1623,N_410);
xor U2733 (N_2733,N_58,N_425);
and U2734 (N_2734,N_820,N_1256);
nor U2735 (N_2735,N_1930,N_595);
nand U2736 (N_2736,N_1964,N_1005);
and U2737 (N_2737,N_1493,N_34);
nor U2738 (N_2738,N_1991,N_740);
and U2739 (N_2739,N_1677,N_1020);
xnor U2740 (N_2740,N_414,N_1921);
and U2741 (N_2741,N_44,N_560);
nand U2742 (N_2742,N_504,N_1502);
nor U2743 (N_2743,N_1687,N_1148);
nor U2744 (N_2744,N_832,N_628);
and U2745 (N_2745,N_1170,N_135);
or U2746 (N_2746,N_1864,N_1794);
or U2747 (N_2747,N_218,N_964);
or U2748 (N_2748,N_1981,N_801);
and U2749 (N_2749,N_337,N_510);
nand U2750 (N_2750,N_956,N_924);
nand U2751 (N_2751,N_28,N_191);
nor U2752 (N_2752,N_717,N_737);
nor U2753 (N_2753,N_698,N_994);
and U2754 (N_2754,N_182,N_1165);
xor U2755 (N_2755,N_1407,N_616);
xnor U2756 (N_2756,N_993,N_1386);
or U2757 (N_2757,N_1774,N_1522);
xnor U2758 (N_2758,N_354,N_602);
and U2759 (N_2759,N_1353,N_651);
nor U2760 (N_2760,N_885,N_198);
xnor U2761 (N_2761,N_250,N_809);
and U2762 (N_2762,N_1291,N_1215);
or U2763 (N_2763,N_930,N_1292);
nand U2764 (N_2764,N_1246,N_366);
xor U2765 (N_2765,N_1962,N_889);
nand U2766 (N_2766,N_314,N_1117);
or U2767 (N_2767,N_1828,N_151);
nand U2768 (N_2768,N_1948,N_1898);
and U2769 (N_2769,N_170,N_219);
and U2770 (N_2770,N_1696,N_512);
or U2771 (N_2771,N_77,N_1099);
nand U2772 (N_2772,N_5,N_84);
and U2773 (N_2773,N_1108,N_1662);
and U2774 (N_2774,N_488,N_570);
nor U2775 (N_2775,N_1406,N_1917);
and U2776 (N_2776,N_1212,N_1758);
nand U2777 (N_2777,N_68,N_1251);
or U2778 (N_2778,N_1579,N_1736);
and U2779 (N_2779,N_1269,N_955);
and U2780 (N_2780,N_637,N_1198);
or U2781 (N_2781,N_1178,N_1916);
and U2782 (N_2782,N_1684,N_392);
or U2783 (N_2783,N_501,N_728);
nor U2784 (N_2784,N_980,N_24);
or U2785 (N_2785,N_1054,N_1845);
and U2786 (N_2786,N_1250,N_1672);
and U2787 (N_2787,N_1273,N_1366);
and U2788 (N_2788,N_548,N_745);
nor U2789 (N_2789,N_1115,N_636);
and U2790 (N_2790,N_641,N_90);
xnor U2791 (N_2791,N_770,N_568);
nand U2792 (N_2792,N_1866,N_1716);
xnor U2793 (N_2793,N_1767,N_1561);
nor U2794 (N_2794,N_923,N_685);
nor U2795 (N_2795,N_1240,N_1812);
nor U2796 (N_2796,N_1296,N_449);
xor U2797 (N_2797,N_1781,N_1660);
xnor U2798 (N_2798,N_1802,N_507);
nor U2799 (N_2799,N_253,N_829);
and U2800 (N_2800,N_633,N_265);
or U2801 (N_2801,N_814,N_987);
nor U2802 (N_2802,N_1669,N_1266);
nor U2803 (N_2803,N_1737,N_372);
xor U2804 (N_2804,N_914,N_143);
or U2805 (N_2805,N_1508,N_1187);
nand U2806 (N_2806,N_461,N_482);
nor U2807 (N_2807,N_92,N_1540);
nor U2808 (N_2808,N_1760,N_317);
and U2809 (N_2809,N_217,N_1133);
nor U2810 (N_2810,N_1081,N_1548);
and U2811 (N_2811,N_1997,N_103);
xnor U2812 (N_2812,N_863,N_1476);
or U2813 (N_2813,N_934,N_639);
xnor U2814 (N_2814,N_1676,N_351);
nor U2815 (N_2815,N_1658,N_1840);
and U2816 (N_2816,N_1252,N_409);
nand U2817 (N_2817,N_113,N_522);
or U2818 (N_2818,N_31,N_125);
or U2819 (N_2819,N_51,N_1683);
and U2820 (N_2820,N_1879,N_255);
or U2821 (N_2821,N_295,N_1598);
and U2822 (N_2822,N_597,N_1819);
or U2823 (N_2823,N_181,N_883);
xor U2824 (N_2824,N_1114,N_365);
nor U2825 (N_2825,N_1360,N_1326);
and U2826 (N_2826,N_1231,N_1639);
and U2827 (N_2827,N_54,N_65);
xnor U2828 (N_2828,N_32,N_1714);
nor U2829 (N_2829,N_153,N_1768);
and U2830 (N_2830,N_1807,N_467);
nand U2831 (N_2831,N_1162,N_1132);
and U2832 (N_2832,N_660,N_1841);
nor U2833 (N_2833,N_25,N_686);
xor U2834 (N_2834,N_1899,N_769);
and U2835 (N_2835,N_1821,N_1121);
and U2836 (N_2836,N_1565,N_1743);
nor U2837 (N_2837,N_232,N_610);
nand U2838 (N_2838,N_521,N_1656);
xnor U2839 (N_2839,N_1545,N_979);
nor U2840 (N_2840,N_1920,N_36);
and U2841 (N_2841,N_1174,N_846);
or U2842 (N_2842,N_1064,N_1599);
xnor U2843 (N_2843,N_1536,N_1118);
nor U2844 (N_2844,N_454,N_1806);
and U2845 (N_2845,N_1062,N_1343);
xor U2846 (N_2846,N_399,N_1603);
nor U2847 (N_2847,N_1341,N_1040);
xnor U2848 (N_2848,N_453,N_1301);
nor U2849 (N_2849,N_1562,N_1865);
nand U2850 (N_2850,N_1854,N_886);
nor U2851 (N_2851,N_729,N_1484);
or U2852 (N_2852,N_996,N_327);
and U2853 (N_2853,N_959,N_1419);
nand U2854 (N_2854,N_1799,N_332);
nor U2855 (N_2855,N_340,N_1190);
and U2856 (N_2856,N_139,N_1392);
and U2857 (N_2857,N_1727,N_1886);
or U2858 (N_2858,N_1349,N_772);
nor U2859 (N_2859,N_152,N_1722);
xor U2860 (N_2860,N_1956,N_1911);
nor U2861 (N_2861,N_1617,N_644);
xor U2862 (N_2862,N_565,N_1652);
nand U2863 (N_2863,N_1673,N_707);
xnor U2864 (N_2864,N_969,N_514);
and U2865 (N_2865,N_1485,N_1095);
nand U2866 (N_2866,N_1703,N_439);
or U2867 (N_2867,N_475,N_623);
nor U2868 (N_2868,N_1739,N_1351);
nor U2869 (N_2869,N_1542,N_64);
nand U2870 (N_2870,N_1626,N_1189);
nor U2871 (N_2871,N_459,N_1524);
xor U2872 (N_2872,N_711,N_249);
xor U2873 (N_2873,N_1219,N_810);
nor U2874 (N_2874,N_1007,N_1400);
nor U2875 (N_2875,N_966,N_1217);
or U2876 (N_2876,N_882,N_1426);
nand U2877 (N_2877,N_797,N_1762);
xor U2878 (N_2878,N_1458,N_359);
nor U2879 (N_2879,N_972,N_207);
and U2880 (N_2880,N_1364,N_128);
or U2881 (N_2881,N_1608,N_712);
nand U2882 (N_2882,N_1640,N_765);
nand U2883 (N_2883,N_1510,N_1329);
or U2884 (N_2884,N_1202,N_1253);
or U2885 (N_2885,N_1523,N_1125);
nand U2886 (N_2886,N_1004,N_1839);
nand U2887 (N_2887,N_853,N_1715);
and U2888 (N_2888,N_1186,N_1556);
or U2889 (N_2889,N_93,N_309);
or U2890 (N_2890,N_1106,N_1473);
nand U2891 (N_2891,N_577,N_1027);
nor U2892 (N_2892,N_995,N_768);
or U2893 (N_2893,N_1248,N_312);
or U2894 (N_2894,N_378,N_1270);
nand U2895 (N_2895,N_1975,N_1718);
or U2896 (N_2896,N_666,N_1261);
nor U2897 (N_2897,N_1826,N_288);
xnor U2898 (N_2898,N_420,N_416);
and U2899 (N_2899,N_659,N_1823);
nand U2900 (N_2900,N_270,N_984);
nor U2901 (N_2901,N_1084,N_1325);
nor U2902 (N_2902,N_703,N_57);
xnor U2903 (N_2903,N_530,N_1157);
nand U2904 (N_2904,N_222,N_1888);
and U2905 (N_2905,N_180,N_1572);
or U2906 (N_2906,N_380,N_818);
nor U2907 (N_2907,N_74,N_1394);
xor U2908 (N_2908,N_370,N_94);
nand U2909 (N_2909,N_890,N_538);
nor U2910 (N_2910,N_52,N_836);
and U2911 (N_2911,N_1612,N_650);
and U2912 (N_2912,N_62,N_272);
or U2913 (N_2913,N_1675,N_1377);
nor U2914 (N_2914,N_1952,N_1679);
or U2915 (N_2915,N_1100,N_347);
and U2916 (N_2916,N_1285,N_1960);
nor U2917 (N_2917,N_1614,N_566);
xor U2918 (N_2918,N_1089,N_1708);
and U2919 (N_2919,N_120,N_1501);
xor U2920 (N_2920,N_285,N_1068);
nor U2921 (N_2921,N_49,N_1686);
nor U2922 (N_2922,N_1910,N_1813);
xor U2923 (N_2923,N_142,N_1018);
nor U2924 (N_2924,N_1941,N_357);
xnor U2925 (N_2925,N_412,N_1101);
and U2926 (N_2926,N_1468,N_1294);
and U2927 (N_2927,N_369,N_438);
and U2928 (N_2928,N_588,N_731);
nand U2929 (N_2929,N_1489,N_1149);
nor U2930 (N_2930,N_149,N_710);
and U2931 (N_2931,N_629,N_779);
xor U2932 (N_2932,N_990,N_305);
nor U2933 (N_2933,N_485,N_339);
and U2934 (N_2934,N_864,N_976);
xor U2935 (N_2935,N_1796,N_949);
xor U2936 (N_2936,N_527,N_473);
nand U2937 (N_2937,N_30,N_1754);
nor U2938 (N_2938,N_206,N_1646);
nand U2939 (N_2939,N_1970,N_827);
nand U2940 (N_2940,N_843,N_39);
and U2941 (N_2941,N_746,N_1944);
and U2942 (N_2942,N_677,N_586);
nor U2943 (N_2943,N_1516,N_687);
or U2944 (N_2944,N_1158,N_487);
xnor U2945 (N_2945,N_1705,N_1140);
and U2946 (N_2946,N_1788,N_1340);
and U2947 (N_2947,N_1092,N_859);
and U2948 (N_2948,N_571,N_1191);
xor U2949 (N_2949,N_1507,N_1192);
or U2950 (N_2950,N_1263,N_202);
or U2951 (N_2951,N_535,N_502);
or U2952 (N_2952,N_1223,N_1065);
and U2953 (N_2953,N_903,N_72);
and U2954 (N_2954,N_489,N_1915);
and U2955 (N_2955,N_1408,N_1844);
xor U2956 (N_2956,N_1700,N_368);
or U2957 (N_2957,N_1003,N_802);
nand U2958 (N_2958,N_1822,N_1851);
and U2959 (N_2959,N_1015,N_477);
nand U2960 (N_2960,N_825,N_1581);
and U2961 (N_2961,N_881,N_866);
and U2962 (N_2962,N_1553,N_1120);
nand U2963 (N_2963,N_1795,N_81);
xor U2964 (N_2964,N_1444,N_264);
and U2965 (N_2965,N_1939,N_1993);
xor U2966 (N_2966,N_1527,N_342);
and U2967 (N_2967,N_1972,N_2);
nand U2968 (N_2968,N_175,N_211);
xnor U2969 (N_2969,N_391,N_1373);
nor U2970 (N_2970,N_91,N_785);
nand U2971 (N_2971,N_1816,N_1200);
nor U2972 (N_2972,N_1446,N_1128);
or U2973 (N_2973,N_823,N_1533);
nor U2974 (N_2974,N_1735,N_1838);
or U2975 (N_2975,N_584,N_1771);
xnor U2976 (N_2976,N_455,N_1193);
nor U2977 (N_2977,N_408,N_523);
and U2978 (N_2978,N_1790,N_1290);
nand U2979 (N_2979,N_243,N_413);
xor U2980 (N_2980,N_1901,N_1717);
xor U2981 (N_2981,N_509,N_1977);
and U2982 (N_2982,N_1689,N_1316);
or U2983 (N_2983,N_1883,N_1079);
nor U2984 (N_2984,N_227,N_137);
nand U2985 (N_2985,N_700,N_415);
and U2986 (N_2986,N_403,N_649);
xnor U2987 (N_2987,N_1923,N_78);
nand U2988 (N_2988,N_33,N_397);
or U2989 (N_2989,N_579,N_954);
nor U2990 (N_2990,N_1359,N_1413);
nor U2991 (N_2991,N_559,N_1986);
nand U2992 (N_2992,N_492,N_508);
and U2993 (N_2993,N_1967,N_676);
xor U2994 (N_2994,N_679,N_1513);
xor U2995 (N_2995,N_848,N_1129);
and U2996 (N_2996,N_294,N_1896);
or U2997 (N_2997,N_311,N_1013);
xor U2998 (N_2998,N_1848,N_1229);
or U2999 (N_2999,N_1371,N_1429);
nor U3000 (N_3000,N_1484,N_508);
nand U3001 (N_3001,N_1363,N_1127);
or U3002 (N_3002,N_1118,N_1655);
xnor U3003 (N_3003,N_1640,N_740);
and U3004 (N_3004,N_730,N_1071);
nor U3005 (N_3005,N_865,N_477);
nor U3006 (N_3006,N_418,N_1179);
or U3007 (N_3007,N_671,N_1072);
xor U3008 (N_3008,N_851,N_1086);
nand U3009 (N_3009,N_1982,N_1862);
or U3010 (N_3010,N_1898,N_524);
nor U3011 (N_3011,N_760,N_690);
and U3012 (N_3012,N_1702,N_1151);
and U3013 (N_3013,N_45,N_1233);
xnor U3014 (N_3014,N_224,N_1797);
and U3015 (N_3015,N_763,N_1562);
nand U3016 (N_3016,N_348,N_1102);
nand U3017 (N_3017,N_132,N_1797);
xor U3018 (N_3018,N_1480,N_209);
or U3019 (N_3019,N_752,N_1356);
xor U3020 (N_3020,N_1948,N_694);
xor U3021 (N_3021,N_1994,N_234);
xnor U3022 (N_3022,N_1650,N_951);
or U3023 (N_3023,N_60,N_676);
or U3024 (N_3024,N_242,N_696);
xor U3025 (N_3025,N_779,N_1801);
xor U3026 (N_3026,N_1540,N_500);
and U3027 (N_3027,N_1339,N_1073);
nor U3028 (N_3028,N_1742,N_72);
and U3029 (N_3029,N_1110,N_482);
and U3030 (N_3030,N_888,N_531);
xnor U3031 (N_3031,N_1057,N_963);
nor U3032 (N_3032,N_1637,N_486);
nor U3033 (N_3033,N_1251,N_729);
or U3034 (N_3034,N_159,N_662);
xor U3035 (N_3035,N_725,N_1274);
nand U3036 (N_3036,N_654,N_402);
or U3037 (N_3037,N_532,N_1190);
nand U3038 (N_3038,N_1338,N_1588);
nand U3039 (N_3039,N_1006,N_157);
nor U3040 (N_3040,N_1822,N_950);
nand U3041 (N_3041,N_57,N_1876);
nand U3042 (N_3042,N_1718,N_620);
and U3043 (N_3043,N_1383,N_615);
nand U3044 (N_3044,N_1573,N_1724);
nand U3045 (N_3045,N_422,N_1656);
nand U3046 (N_3046,N_1339,N_1369);
nand U3047 (N_3047,N_1665,N_1921);
and U3048 (N_3048,N_1721,N_1260);
or U3049 (N_3049,N_347,N_1514);
nor U3050 (N_3050,N_1601,N_466);
and U3051 (N_3051,N_882,N_1108);
and U3052 (N_3052,N_121,N_410);
and U3053 (N_3053,N_1503,N_613);
and U3054 (N_3054,N_355,N_1995);
nand U3055 (N_3055,N_1458,N_949);
or U3056 (N_3056,N_419,N_992);
nand U3057 (N_3057,N_195,N_406);
and U3058 (N_3058,N_1609,N_1479);
xor U3059 (N_3059,N_531,N_1236);
nor U3060 (N_3060,N_59,N_329);
nand U3061 (N_3061,N_1514,N_212);
nand U3062 (N_3062,N_1548,N_81);
nor U3063 (N_3063,N_226,N_323);
or U3064 (N_3064,N_1072,N_155);
nand U3065 (N_3065,N_1566,N_954);
nand U3066 (N_3066,N_1291,N_70);
nor U3067 (N_3067,N_970,N_1971);
or U3068 (N_3068,N_47,N_1990);
nand U3069 (N_3069,N_90,N_1577);
and U3070 (N_3070,N_1136,N_846);
xor U3071 (N_3071,N_1375,N_410);
and U3072 (N_3072,N_17,N_619);
xor U3073 (N_3073,N_1568,N_561);
nand U3074 (N_3074,N_1226,N_86);
or U3075 (N_3075,N_514,N_1827);
or U3076 (N_3076,N_942,N_1523);
or U3077 (N_3077,N_696,N_1509);
nor U3078 (N_3078,N_1952,N_1621);
nor U3079 (N_3079,N_397,N_1875);
or U3080 (N_3080,N_443,N_762);
or U3081 (N_3081,N_1347,N_622);
nand U3082 (N_3082,N_793,N_1663);
or U3083 (N_3083,N_1967,N_631);
xnor U3084 (N_3084,N_952,N_1411);
nand U3085 (N_3085,N_1300,N_1924);
nand U3086 (N_3086,N_1375,N_20);
nor U3087 (N_3087,N_695,N_1566);
or U3088 (N_3088,N_1941,N_886);
nand U3089 (N_3089,N_83,N_703);
and U3090 (N_3090,N_755,N_744);
nor U3091 (N_3091,N_1293,N_1792);
or U3092 (N_3092,N_989,N_895);
and U3093 (N_3093,N_1253,N_1172);
and U3094 (N_3094,N_706,N_12);
and U3095 (N_3095,N_301,N_1391);
nand U3096 (N_3096,N_1833,N_505);
nor U3097 (N_3097,N_1205,N_485);
or U3098 (N_3098,N_1781,N_1953);
or U3099 (N_3099,N_805,N_1505);
or U3100 (N_3100,N_1914,N_456);
and U3101 (N_3101,N_1106,N_128);
nor U3102 (N_3102,N_1107,N_1264);
or U3103 (N_3103,N_1209,N_1475);
xnor U3104 (N_3104,N_1291,N_1709);
or U3105 (N_3105,N_623,N_1446);
nor U3106 (N_3106,N_648,N_363);
nor U3107 (N_3107,N_1387,N_1545);
and U3108 (N_3108,N_1765,N_350);
nor U3109 (N_3109,N_156,N_1388);
nand U3110 (N_3110,N_98,N_124);
or U3111 (N_3111,N_276,N_1819);
nand U3112 (N_3112,N_1919,N_1455);
and U3113 (N_3113,N_1602,N_1010);
or U3114 (N_3114,N_617,N_651);
or U3115 (N_3115,N_687,N_61);
nor U3116 (N_3116,N_1352,N_506);
nor U3117 (N_3117,N_843,N_387);
xnor U3118 (N_3118,N_467,N_1595);
or U3119 (N_3119,N_1783,N_1379);
xnor U3120 (N_3120,N_1704,N_282);
and U3121 (N_3121,N_898,N_659);
xor U3122 (N_3122,N_640,N_1164);
nor U3123 (N_3123,N_960,N_1231);
and U3124 (N_3124,N_702,N_1467);
nor U3125 (N_3125,N_1641,N_855);
nand U3126 (N_3126,N_453,N_799);
xor U3127 (N_3127,N_798,N_1141);
nor U3128 (N_3128,N_186,N_1588);
and U3129 (N_3129,N_647,N_1926);
and U3130 (N_3130,N_1634,N_153);
nand U3131 (N_3131,N_999,N_1899);
and U3132 (N_3132,N_1165,N_644);
nor U3133 (N_3133,N_1990,N_877);
or U3134 (N_3134,N_635,N_555);
nand U3135 (N_3135,N_1458,N_1703);
or U3136 (N_3136,N_316,N_1567);
xnor U3137 (N_3137,N_1400,N_1452);
nor U3138 (N_3138,N_1600,N_1417);
xnor U3139 (N_3139,N_966,N_188);
xor U3140 (N_3140,N_854,N_927);
and U3141 (N_3141,N_713,N_1774);
xor U3142 (N_3142,N_23,N_558);
nand U3143 (N_3143,N_1195,N_1299);
nor U3144 (N_3144,N_1685,N_481);
nor U3145 (N_3145,N_750,N_181);
nand U3146 (N_3146,N_1912,N_983);
nor U3147 (N_3147,N_45,N_1232);
nand U3148 (N_3148,N_381,N_1568);
xor U3149 (N_3149,N_1149,N_1119);
or U3150 (N_3150,N_1837,N_1288);
xor U3151 (N_3151,N_1406,N_504);
and U3152 (N_3152,N_1731,N_877);
and U3153 (N_3153,N_1716,N_297);
nor U3154 (N_3154,N_1318,N_202);
nor U3155 (N_3155,N_1580,N_1825);
or U3156 (N_3156,N_1060,N_1210);
and U3157 (N_3157,N_1648,N_1493);
nand U3158 (N_3158,N_1747,N_254);
nand U3159 (N_3159,N_241,N_220);
nor U3160 (N_3160,N_636,N_1822);
xor U3161 (N_3161,N_1230,N_1405);
nor U3162 (N_3162,N_1947,N_276);
and U3163 (N_3163,N_532,N_125);
or U3164 (N_3164,N_596,N_1900);
nor U3165 (N_3165,N_403,N_1668);
and U3166 (N_3166,N_563,N_1977);
xnor U3167 (N_3167,N_739,N_649);
or U3168 (N_3168,N_214,N_584);
xnor U3169 (N_3169,N_737,N_621);
xnor U3170 (N_3170,N_388,N_476);
and U3171 (N_3171,N_1886,N_908);
nand U3172 (N_3172,N_1415,N_1292);
nor U3173 (N_3173,N_1648,N_1771);
nand U3174 (N_3174,N_1257,N_1427);
xor U3175 (N_3175,N_1098,N_1941);
and U3176 (N_3176,N_494,N_751);
or U3177 (N_3177,N_1948,N_27);
and U3178 (N_3178,N_159,N_1961);
nand U3179 (N_3179,N_1819,N_301);
nor U3180 (N_3180,N_1132,N_303);
nor U3181 (N_3181,N_1089,N_1857);
or U3182 (N_3182,N_1624,N_1269);
and U3183 (N_3183,N_1910,N_593);
nand U3184 (N_3184,N_1773,N_1469);
or U3185 (N_3185,N_34,N_465);
and U3186 (N_3186,N_395,N_123);
and U3187 (N_3187,N_992,N_1489);
nand U3188 (N_3188,N_289,N_356);
nor U3189 (N_3189,N_651,N_1403);
or U3190 (N_3190,N_1101,N_1515);
xor U3191 (N_3191,N_1772,N_1924);
nor U3192 (N_3192,N_1891,N_3);
nand U3193 (N_3193,N_1350,N_1416);
and U3194 (N_3194,N_1927,N_97);
and U3195 (N_3195,N_1523,N_1931);
xor U3196 (N_3196,N_1524,N_627);
nand U3197 (N_3197,N_1314,N_1107);
nand U3198 (N_3198,N_227,N_1990);
and U3199 (N_3199,N_1690,N_977);
nand U3200 (N_3200,N_844,N_1393);
xnor U3201 (N_3201,N_840,N_1987);
xor U3202 (N_3202,N_1982,N_1461);
xor U3203 (N_3203,N_881,N_724);
nor U3204 (N_3204,N_480,N_1187);
nor U3205 (N_3205,N_1690,N_586);
nand U3206 (N_3206,N_1119,N_1420);
or U3207 (N_3207,N_1078,N_1720);
nor U3208 (N_3208,N_1627,N_1009);
nand U3209 (N_3209,N_975,N_1891);
or U3210 (N_3210,N_1814,N_1149);
and U3211 (N_3211,N_1373,N_610);
or U3212 (N_3212,N_289,N_315);
and U3213 (N_3213,N_721,N_580);
or U3214 (N_3214,N_666,N_267);
xor U3215 (N_3215,N_285,N_1165);
xnor U3216 (N_3216,N_340,N_1236);
nand U3217 (N_3217,N_560,N_456);
nand U3218 (N_3218,N_349,N_1276);
and U3219 (N_3219,N_1583,N_119);
or U3220 (N_3220,N_1926,N_1051);
or U3221 (N_3221,N_172,N_641);
xnor U3222 (N_3222,N_1124,N_1069);
xnor U3223 (N_3223,N_905,N_310);
xor U3224 (N_3224,N_504,N_74);
nand U3225 (N_3225,N_577,N_499);
and U3226 (N_3226,N_615,N_1386);
nand U3227 (N_3227,N_719,N_1895);
and U3228 (N_3228,N_107,N_1403);
nor U3229 (N_3229,N_69,N_926);
and U3230 (N_3230,N_302,N_1694);
or U3231 (N_3231,N_1464,N_11);
xnor U3232 (N_3232,N_377,N_559);
and U3233 (N_3233,N_1557,N_838);
nand U3234 (N_3234,N_373,N_1485);
xor U3235 (N_3235,N_739,N_485);
or U3236 (N_3236,N_1895,N_364);
nor U3237 (N_3237,N_5,N_1106);
and U3238 (N_3238,N_1136,N_1300);
nor U3239 (N_3239,N_64,N_1506);
xnor U3240 (N_3240,N_655,N_1025);
and U3241 (N_3241,N_1757,N_497);
xnor U3242 (N_3242,N_1508,N_60);
nor U3243 (N_3243,N_862,N_718);
xor U3244 (N_3244,N_1269,N_767);
or U3245 (N_3245,N_738,N_132);
nor U3246 (N_3246,N_573,N_25);
nor U3247 (N_3247,N_672,N_210);
xor U3248 (N_3248,N_459,N_1002);
and U3249 (N_3249,N_693,N_1679);
nor U3250 (N_3250,N_263,N_1878);
xor U3251 (N_3251,N_1992,N_592);
nor U3252 (N_3252,N_1496,N_1309);
xnor U3253 (N_3253,N_143,N_50);
and U3254 (N_3254,N_1213,N_1137);
xnor U3255 (N_3255,N_1223,N_684);
or U3256 (N_3256,N_476,N_491);
and U3257 (N_3257,N_1115,N_1874);
nor U3258 (N_3258,N_1669,N_974);
xnor U3259 (N_3259,N_922,N_764);
nand U3260 (N_3260,N_647,N_1972);
nand U3261 (N_3261,N_816,N_729);
xor U3262 (N_3262,N_500,N_1002);
and U3263 (N_3263,N_1514,N_1424);
nand U3264 (N_3264,N_1550,N_285);
nand U3265 (N_3265,N_659,N_1022);
and U3266 (N_3266,N_483,N_635);
or U3267 (N_3267,N_1933,N_1724);
or U3268 (N_3268,N_731,N_1502);
nor U3269 (N_3269,N_1754,N_516);
or U3270 (N_3270,N_1884,N_179);
nand U3271 (N_3271,N_1380,N_436);
and U3272 (N_3272,N_1591,N_1807);
or U3273 (N_3273,N_271,N_83);
xnor U3274 (N_3274,N_1191,N_1678);
xor U3275 (N_3275,N_830,N_840);
or U3276 (N_3276,N_53,N_1048);
nand U3277 (N_3277,N_486,N_1401);
and U3278 (N_3278,N_1888,N_330);
or U3279 (N_3279,N_524,N_641);
or U3280 (N_3280,N_1900,N_897);
nor U3281 (N_3281,N_672,N_641);
xor U3282 (N_3282,N_108,N_1345);
nor U3283 (N_3283,N_461,N_775);
xor U3284 (N_3284,N_1491,N_334);
nand U3285 (N_3285,N_1258,N_466);
or U3286 (N_3286,N_500,N_664);
or U3287 (N_3287,N_623,N_519);
and U3288 (N_3288,N_1671,N_705);
nor U3289 (N_3289,N_805,N_1164);
and U3290 (N_3290,N_1734,N_1244);
or U3291 (N_3291,N_116,N_1878);
nand U3292 (N_3292,N_34,N_1774);
nand U3293 (N_3293,N_377,N_995);
xnor U3294 (N_3294,N_1175,N_1232);
or U3295 (N_3295,N_221,N_1032);
xnor U3296 (N_3296,N_1135,N_122);
and U3297 (N_3297,N_1106,N_1242);
or U3298 (N_3298,N_649,N_301);
nor U3299 (N_3299,N_833,N_1432);
xor U3300 (N_3300,N_1224,N_1860);
nor U3301 (N_3301,N_78,N_511);
or U3302 (N_3302,N_34,N_1603);
nor U3303 (N_3303,N_1332,N_131);
and U3304 (N_3304,N_127,N_106);
xnor U3305 (N_3305,N_893,N_231);
nand U3306 (N_3306,N_631,N_485);
or U3307 (N_3307,N_986,N_959);
xor U3308 (N_3308,N_474,N_1664);
xor U3309 (N_3309,N_1780,N_1915);
xor U3310 (N_3310,N_1233,N_217);
nor U3311 (N_3311,N_105,N_89);
and U3312 (N_3312,N_387,N_1157);
nand U3313 (N_3313,N_972,N_1408);
or U3314 (N_3314,N_1940,N_1016);
nand U3315 (N_3315,N_23,N_203);
or U3316 (N_3316,N_1308,N_282);
xnor U3317 (N_3317,N_1990,N_52);
nand U3318 (N_3318,N_86,N_221);
nor U3319 (N_3319,N_505,N_830);
xor U3320 (N_3320,N_542,N_1280);
or U3321 (N_3321,N_484,N_290);
xnor U3322 (N_3322,N_1342,N_1358);
nand U3323 (N_3323,N_135,N_213);
or U3324 (N_3324,N_1899,N_1659);
nand U3325 (N_3325,N_1386,N_1674);
nor U3326 (N_3326,N_1502,N_932);
nor U3327 (N_3327,N_1673,N_327);
xor U3328 (N_3328,N_1373,N_1867);
nor U3329 (N_3329,N_677,N_121);
or U3330 (N_3330,N_1942,N_1874);
and U3331 (N_3331,N_294,N_1757);
or U3332 (N_3332,N_1061,N_729);
xnor U3333 (N_3333,N_358,N_112);
nor U3334 (N_3334,N_839,N_1927);
nand U3335 (N_3335,N_1390,N_115);
nor U3336 (N_3336,N_108,N_1024);
nand U3337 (N_3337,N_268,N_68);
nor U3338 (N_3338,N_876,N_1695);
or U3339 (N_3339,N_1022,N_660);
or U3340 (N_3340,N_175,N_140);
or U3341 (N_3341,N_435,N_1603);
nor U3342 (N_3342,N_388,N_1419);
nand U3343 (N_3343,N_1392,N_480);
or U3344 (N_3344,N_974,N_1575);
and U3345 (N_3345,N_1499,N_1192);
nand U3346 (N_3346,N_1003,N_1759);
or U3347 (N_3347,N_1099,N_1368);
and U3348 (N_3348,N_1368,N_917);
nand U3349 (N_3349,N_1608,N_1394);
nand U3350 (N_3350,N_1150,N_405);
xor U3351 (N_3351,N_385,N_853);
nor U3352 (N_3352,N_953,N_443);
nor U3353 (N_3353,N_685,N_812);
xnor U3354 (N_3354,N_928,N_958);
and U3355 (N_3355,N_251,N_1812);
and U3356 (N_3356,N_491,N_1788);
nor U3357 (N_3357,N_112,N_1329);
or U3358 (N_3358,N_1408,N_1855);
nor U3359 (N_3359,N_1341,N_402);
xor U3360 (N_3360,N_188,N_1209);
nor U3361 (N_3361,N_335,N_1914);
xnor U3362 (N_3362,N_838,N_816);
and U3363 (N_3363,N_387,N_1566);
nor U3364 (N_3364,N_1485,N_69);
nand U3365 (N_3365,N_288,N_1790);
and U3366 (N_3366,N_1695,N_79);
xor U3367 (N_3367,N_732,N_112);
nor U3368 (N_3368,N_324,N_588);
xor U3369 (N_3369,N_1218,N_997);
xnor U3370 (N_3370,N_1294,N_131);
xnor U3371 (N_3371,N_994,N_1339);
nand U3372 (N_3372,N_811,N_457);
xnor U3373 (N_3373,N_1475,N_1151);
or U3374 (N_3374,N_1069,N_342);
nand U3375 (N_3375,N_455,N_1036);
xor U3376 (N_3376,N_961,N_1572);
xnor U3377 (N_3377,N_606,N_261);
xnor U3378 (N_3378,N_818,N_709);
nand U3379 (N_3379,N_1751,N_1519);
nand U3380 (N_3380,N_1970,N_1134);
xor U3381 (N_3381,N_1300,N_1527);
nand U3382 (N_3382,N_1446,N_1125);
nand U3383 (N_3383,N_549,N_476);
and U3384 (N_3384,N_711,N_1750);
nand U3385 (N_3385,N_814,N_328);
nand U3386 (N_3386,N_577,N_907);
and U3387 (N_3387,N_1089,N_668);
or U3388 (N_3388,N_1000,N_963);
or U3389 (N_3389,N_1523,N_1982);
or U3390 (N_3390,N_740,N_304);
nor U3391 (N_3391,N_1768,N_449);
and U3392 (N_3392,N_175,N_498);
nand U3393 (N_3393,N_1627,N_1901);
or U3394 (N_3394,N_574,N_1699);
xor U3395 (N_3395,N_1193,N_828);
and U3396 (N_3396,N_1442,N_592);
nor U3397 (N_3397,N_932,N_1348);
or U3398 (N_3398,N_838,N_908);
xnor U3399 (N_3399,N_1779,N_1197);
nand U3400 (N_3400,N_1423,N_150);
nand U3401 (N_3401,N_1343,N_1586);
or U3402 (N_3402,N_1733,N_1554);
or U3403 (N_3403,N_5,N_1638);
xor U3404 (N_3404,N_270,N_620);
or U3405 (N_3405,N_1732,N_446);
or U3406 (N_3406,N_851,N_248);
and U3407 (N_3407,N_670,N_757);
or U3408 (N_3408,N_843,N_416);
xnor U3409 (N_3409,N_1873,N_412);
nand U3410 (N_3410,N_1653,N_1745);
and U3411 (N_3411,N_1701,N_1703);
nand U3412 (N_3412,N_121,N_213);
nand U3413 (N_3413,N_1682,N_1440);
nand U3414 (N_3414,N_584,N_693);
or U3415 (N_3415,N_924,N_549);
xnor U3416 (N_3416,N_1966,N_1607);
xnor U3417 (N_3417,N_798,N_340);
xor U3418 (N_3418,N_643,N_1326);
nand U3419 (N_3419,N_1491,N_1472);
nor U3420 (N_3420,N_8,N_558);
and U3421 (N_3421,N_597,N_5);
xor U3422 (N_3422,N_1744,N_961);
nor U3423 (N_3423,N_1468,N_63);
xnor U3424 (N_3424,N_1076,N_1563);
nand U3425 (N_3425,N_1905,N_1186);
xor U3426 (N_3426,N_1090,N_1764);
and U3427 (N_3427,N_863,N_853);
or U3428 (N_3428,N_1673,N_140);
xnor U3429 (N_3429,N_1569,N_1736);
and U3430 (N_3430,N_1415,N_662);
nor U3431 (N_3431,N_771,N_1324);
and U3432 (N_3432,N_1835,N_59);
or U3433 (N_3433,N_966,N_1297);
or U3434 (N_3434,N_1036,N_1797);
or U3435 (N_3435,N_440,N_1320);
nand U3436 (N_3436,N_1544,N_1371);
nor U3437 (N_3437,N_250,N_1479);
nor U3438 (N_3438,N_456,N_1472);
nand U3439 (N_3439,N_95,N_1825);
xnor U3440 (N_3440,N_1738,N_1868);
and U3441 (N_3441,N_889,N_190);
xor U3442 (N_3442,N_66,N_842);
nor U3443 (N_3443,N_1114,N_1145);
nand U3444 (N_3444,N_1672,N_1294);
nor U3445 (N_3445,N_1416,N_1190);
nor U3446 (N_3446,N_1680,N_39);
xor U3447 (N_3447,N_305,N_1076);
nand U3448 (N_3448,N_791,N_1943);
xor U3449 (N_3449,N_163,N_970);
and U3450 (N_3450,N_1799,N_1841);
and U3451 (N_3451,N_1244,N_945);
xor U3452 (N_3452,N_622,N_1569);
nand U3453 (N_3453,N_168,N_1000);
nor U3454 (N_3454,N_1313,N_129);
nor U3455 (N_3455,N_486,N_1185);
nor U3456 (N_3456,N_451,N_1550);
or U3457 (N_3457,N_1140,N_800);
nor U3458 (N_3458,N_1084,N_194);
and U3459 (N_3459,N_1336,N_198);
and U3460 (N_3460,N_752,N_1857);
or U3461 (N_3461,N_121,N_875);
or U3462 (N_3462,N_1052,N_1042);
nor U3463 (N_3463,N_1374,N_1672);
or U3464 (N_3464,N_270,N_87);
nor U3465 (N_3465,N_799,N_1647);
or U3466 (N_3466,N_358,N_744);
xnor U3467 (N_3467,N_1220,N_1727);
or U3468 (N_3468,N_692,N_9);
or U3469 (N_3469,N_1015,N_604);
or U3470 (N_3470,N_1373,N_1414);
nand U3471 (N_3471,N_1276,N_911);
and U3472 (N_3472,N_1304,N_1142);
xnor U3473 (N_3473,N_1558,N_1621);
nor U3474 (N_3474,N_715,N_526);
xor U3475 (N_3475,N_1333,N_374);
nand U3476 (N_3476,N_151,N_515);
or U3477 (N_3477,N_872,N_1430);
nand U3478 (N_3478,N_1207,N_1440);
nand U3479 (N_3479,N_1926,N_989);
or U3480 (N_3480,N_1699,N_1398);
and U3481 (N_3481,N_1144,N_1805);
and U3482 (N_3482,N_1764,N_444);
or U3483 (N_3483,N_1128,N_1340);
and U3484 (N_3484,N_986,N_1611);
or U3485 (N_3485,N_305,N_1038);
xnor U3486 (N_3486,N_1417,N_727);
and U3487 (N_3487,N_1212,N_1440);
nand U3488 (N_3488,N_716,N_886);
and U3489 (N_3489,N_1674,N_928);
nand U3490 (N_3490,N_1408,N_1901);
nand U3491 (N_3491,N_1424,N_1777);
or U3492 (N_3492,N_312,N_1963);
or U3493 (N_3493,N_253,N_804);
or U3494 (N_3494,N_77,N_1653);
xor U3495 (N_3495,N_353,N_1024);
or U3496 (N_3496,N_1171,N_494);
nor U3497 (N_3497,N_436,N_8);
xnor U3498 (N_3498,N_58,N_668);
nand U3499 (N_3499,N_1521,N_86);
and U3500 (N_3500,N_628,N_1825);
xor U3501 (N_3501,N_1745,N_1181);
nand U3502 (N_3502,N_1438,N_751);
and U3503 (N_3503,N_236,N_326);
xnor U3504 (N_3504,N_1619,N_331);
nand U3505 (N_3505,N_1294,N_890);
and U3506 (N_3506,N_1627,N_936);
nor U3507 (N_3507,N_814,N_339);
nand U3508 (N_3508,N_1255,N_1146);
xnor U3509 (N_3509,N_52,N_145);
xor U3510 (N_3510,N_1505,N_169);
nand U3511 (N_3511,N_1211,N_77);
xor U3512 (N_3512,N_356,N_970);
xor U3513 (N_3513,N_394,N_330);
nor U3514 (N_3514,N_1667,N_1090);
nor U3515 (N_3515,N_1573,N_707);
nor U3516 (N_3516,N_317,N_500);
nor U3517 (N_3517,N_1272,N_351);
nand U3518 (N_3518,N_647,N_1528);
or U3519 (N_3519,N_1161,N_1930);
nor U3520 (N_3520,N_783,N_1123);
or U3521 (N_3521,N_561,N_1538);
nand U3522 (N_3522,N_500,N_763);
nor U3523 (N_3523,N_1040,N_1107);
and U3524 (N_3524,N_1195,N_201);
xor U3525 (N_3525,N_1938,N_70);
nand U3526 (N_3526,N_624,N_832);
nand U3527 (N_3527,N_1143,N_292);
xor U3528 (N_3528,N_975,N_677);
xor U3529 (N_3529,N_194,N_905);
nand U3530 (N_3530,N_1477,N_970);
xor U3531 (N_3531,N_1087,N_149);
nand U3532 (N_3532,N_191,N_384);
nor U3533 (N_3533,N_1495,N_413);
xnor U3534 (N_3534,N_1622,N_1979);
and U3535 (N_3535,N_1649,N_233);
xnor U3536 (N_3536,N_1894,N_281);
or U3537 (N_3537,N_1358,N_1778);
or U3538 (N_3538,N_1319,N_787);
nor U3539 (N_3539,N_916,N_76);
xnor U3540 (N_3540,N_1307,N_717);
and U3541 (N_3541,N_815,N_634);
nor U3542 (N_3542,N_1850,N_1289);
nand U3543 (N_3543,N_1156,N_1373);
nor U3544 (N_3544,N_1136,N_1707);
nor U3545 (N_3545,N_1505,N_1839);
and U3546 (N_3546,N_1021,N_1204);
or U3547 (N_3547,N_493,N_301);
nand U3548 (N_3548,N_32,N_36);
xor U3549 (N_3549,N_71,N_870);
or U3550 (N_3550,N_1519,N_1232);
xor U3551 (N_3551,N_258,N_74);
and U3552 (N_3552,N_1106,N_638);
or U3553 (N_3553,N_1685,N_613);
and U3554 (N_3554,N_636,N_132);
nor U3555 (N_3555,N_1980,N_1776);
nand U3556 (N_3556,N_1206,N_1473);
nand U3557 (N_3557,N_1082,N_1147);
or U3558 (N_3558,N_1884,N_709);
xnor U3559 (N_3559,N_638,N_398);
nand U3560 (N_3560,N_1896,N_1659);
nand U3561 (N_3561,N_357,N_1477);
and U3562 (N_3562,N_233,N_136);
or U3563 (N_3563,N_1717,N_865);
nor U3564 (N_3564,N_1672,N_1358);
and U3565 (N_3565,N_1808,N_97);
xor U3566 (N_3566,N_1037,N_780);
nand U3567 (N_3567,N_769,N_1721);
and U3568 (N_3568,N_1677,N_931);
xnor U3569 (N_3569,N_946,N_661);
or U3570 (N_3570,N_729,N_334);
nand U3571 (N_3571,N_1235,N_1090);
xor U3572 (N_3572,N_214,N_199);
xor U3573 (N_3573,N_525,N_571);
nand U3574 (N_3574,N_369,N_1112);
nand U3575 (N_3575,N_311,N_731);
nand U3576 (N_3576,N_1902,N_716);
xnor U3577 (N_3577,N_565,N_1182);
nand U3578 (N_3578,N_1572,N_948);
and U3579 (N_3579,N_1760,N_779);
nor U3580 (N_3580,N_1479,N_121);
nor U3581 (N_3581,N_1321,N_1023);
nor U3582 (N_3582,N_771,N_188);
or U3583 (N_3583,N_924,N_1485);
xnor U3584 (N_3584,N_1616,N_1825);
and U3585 (N_3585,N_254,N_207);
xor U3586 (N_3586,N_1122,N_918);
nand U3587 (N_3587,N_766,N_434);
xnor U3588 (N_3588,N_1087,N_999);
and U3589 (N_3589,N_1506,N_429);
xor U3590 (N_3590,N_633,N_609);
nand U3591 (N_3591,N_1909,N_1603);
nor U3592 (N_3592,N_1209,N_1413);
and U3593 (N_3593,N_173,N_1884);
or U3594 (N_3594,N_1734,N_626);
xnor U3595 (N_3595,N_1240,N_716);
and U3596 (N_3596,N_1934,N_1399);
nand U3597 (N_3597,N_1053,N_889);
or U3598 (N_3598,N_1046,N_1892);
nor U3599 (N_3599,N_654,N_1273);
nand U3600 (N_3600,N_1600,N_835);
nand U3601 (N_3601,N_44,N_1236);
xor U3602 (N_3602,N_905,N_1909);
xnor U3603 (N_3603,N_208,N_150);
nand U3604 (N_3604,N_867,N_1320);
or U3605 (N_3605,N_503,N_1181);
xnor U3606 (N_3606,N_1182,N_9);
and U3607 (N_3607,N_20,N_1283);
nor U3608 (N_3608,N_228,N_661);
or U3609 (N_3609,N_319,N_1004);
xnor U3610 (N_3610,N_972,N_1828);
and U3611 (N_3611,N_1332,N_556);
nor U3612 (N_3612,N_40,N_981);
nor U3613 (N_3613,N_415,N_1552);
nand U3614 (N_3614,N_167,N_391);
xor U3615 (N_3615,N_950,N_438);
and U3616 (N_3616,N_129,N_156);
xor U3617 (N_3617,N_418,N_938);
or U3618 (N_3618,N_1352,N_462);
or U3619 (N_3619,N_516,N_1256);
nand U3620 (N_3620,N_1948,N_889);
xnor U3621 (N_3621,N_1809,N_1043);
or U3622 (N_3622,N_1830,N_363);
nor U3623 (N_3623,N_1218,N_597);
nand U3624 (N_3624,N_1140,N_1428);
nor U3625 (N_3625,N_584,N_585);
or U3626 (N_3626,N_676,N_30);
and U3627 (N_3627,N_1148,N_821);
nand U3628 (N_3628,N_397,N_634);
xor U3629 (N_3629,N_1599,N_1410);
nor U3630 (N_3630,N_1141,N_1921);
nand U3631 (N_3631,N_496,N_1594);
nand U3632 (N_3632,N_835,N_1363);
or U3633 (N_3633,N_1096,N_429);
xnor U3634 (N_3634,N_249,N_182);
or U3635 (N_3635,N_1540,N_545);
or U3636 (N_3636,N_1183,N_1941);
and U3637 (N_3637,N_955,N_707);
nor U3638 (N_3638,N_504,N_352);
nand U3639 (N_3639,N_449,N_207);
nand U3640 (N_3640,N_232,N_1191);
nor U3641 (N_3641,N_1508,N_833);
nand U3642 (N_3642,N_1704,N_1618);
nor U3643 (N_3643,N_365,N_438);
or U3644 (N_3644,N_1712,N_444);
or U3645 (N_3645,N_47,N_635);
nor U3646 (N_3646,N_768,N_480);
xor U3647 (N_3647,N_526,N_1209);
nand U3648 (N_3648,N_1132,N_326);
xnor U3649 (N_3649,N_783,N_1434);
nand U3650 (N_3650,N_1604,N_1965);
nor U3651 (N_3651,N_804,N_1444);
or U3652 (N_3652,N_1180,N_1305);
and U3653 (N_3653,N_866,N_1708);
or U3654 (N_3654,N_1390,N_892);
or U3655 (N_3655,N_54,N_1924);
xor U3656 (N_3656,N_1760,N_1723);
and U3657 (N_3657,N_1033,N_1671);
nor U3658 (N_3658,N_86,N_681);
nor U3659 (N_3659,N_357,N_163);
nand U3660 (N_3660,N_440,N_1083);
or U3661 (N_3661,N_532,N_1431);
xnor U3662 (N_3662,N_471,N_30);
nand U3663 (N_3663,N_928,N_1462);
and U3664 (N_3664,N_529,N_1644);
xor U3665 (N_3665,N_607,N_503);
nor U3666 (N_3666,N_347,N_228);
or U3667 (N_3667,N_520,N_1520);
nand U3668 (N_3668,N_1121,N_1204);
nor U3669 (N_3669,N_1397,N_1794);
and U3670 (N_3670,N_115,N_553);
or U3671 (N_3671,N_134,N_703);
or U3672 (N_3672,N_1933,N_57);
nand U3673 (N_3673,N_1241,N_414);
or U3674 (N_3674,N_1477,N_1259);
xnor U3675 (N_3675,N_1459,N_1308);
and U3676 (N_3676,N_1217,N_1850);
or U3677 (N_3677,N_1343,N_1328);
nor U3678 (N_3678,N_1232,N_1344);
and U3679 (N_3679,N_1566,N_1090);
xor U3680 (N_3680,N_1526,N_326);
nor U3681 (N_3681,N_523,N_1793);
xnor U3682 (N_3682,N_1592,N_530);
nor U3683 (N_3683,N_261,N_850);
nand U3684 (N_3684,N_1299,N_1329);
nor U3685 (N_3685,N_1385,N_1715);
and U3686 (N_3686,N_1075,N_767);
and U3687 (N_3687,N_1594,N_1);
nor U3688 (N_3688,N_727,N_951);
or U3689 (N_3689,N_299,N_1937);
nand U3690 (N_3690,N_1065,N_1392);
nor U3691 (N_3691,N_1644,N_1743);
and U3692 (N_3692,N_1966,N_878);
nor U3693 (N_3693,N_1111,N_1018);
or U3694 (N_3694,N_1178,N_1836);
nand U3695 (N_3695,N_1814,N_1411);
or U3696 (N_3696,N_40,N_801);
and U3697 (N_3697,N_1963,N_1866);
xnor U3698 (N_3698,N_415,N_512);
nand U3699 (N_3699,N_850,N_536);
nand U3700 (N_3700,N_498,N_1278);
nand U3701 (N_3701,N_518,N_1607);
xnor U3702 (N_3702,N_1914,N_695);
or U3703 (N_3703,N_1165,N_761);
or U3704 (N_3704,N_1366,N_1969);
xnor U3705 (N_3705,N_904,N_1245);
or U3706 (N_3706,N_1854,N_714);
and U3707 (N_3707,N_1904,N_391);
xor U3708 (N_3708,N_298,N_1774);
nand U3709 (N_3709,N_675,N_1132);
xnor U3710 (N_3710,N_1388,N_68);
and U3711 (N_3711,N_1603,N_300);
nor U3712 (N_3712,N_730,N_1321);
xor U3713 (N_3713,N_1449,N_684);
nor U3714 (N_3714,N_104,N_1099);
and U3715 (N_3715,N_895,N_969);
xor U3716 (N_3716,N_8,N_1768);
nor U3717 (N_3717,N_5,N_1967);
xnor U3718 (N_3718,N_1082,N_1583);
and U3719 (N_3719,N_833,N_133);
and U3720 (N_3720,N_389,N_1057);
and U3721 (N_3721,N_1373,N_801);
or U3722 (N_3722,N_1081,N_1860);
nand U3723 (N_3723,N_1669,N_675);
and U3724 (N_3724,N_1018,N_350);
nand U3725 (N_3725,N_429,N_1946);
nand U3726 (N_3726,N_94,N_1822);
xnor U3727 (N_3727,N_998,N_1186);
nand U3728 (N_3728,N_142,N_586);
xor U3729 (N_3729,N_950,N_139);
or U3730 (N_3730,N_1980,N_868);
nand U3731 (N_3731,N_1846,N_1197);
xor U3732 (N_3732,N_1202,N_1468);
nand U3733 (N_3733,N_1025,N_264);
or U3734 (N_3734,N_711,N_228);
xor U3735 (N_3735,N_1842,N_1717);
nand U3736 (N_3736,N_1331,N_1142);
or U3737 (N_3737,N_672,N_163);
nor U3738 (N_3738,N_847,N_1292);
xor U3739 (N_3739,N_994,N_1933);
or U3740 (N_3740,N_249,N_1274);
xnor U3741 (N_3741,N_729,N_675);
nand U3742 (N_3742,N_1522,N_1950);
xor U3743 (N_3743,N_610,N_1883);
and U3744 (N_3744,N_1647,N_1701);
nand U3745 (N_3745,N_197,N_646);
xor U3746 (N_3746,N_1008,N_1569);
nor U3747 (N_3747,N_1353,N_899);
and U3748 (N_3748,N_507,N_218);
nor U3749 (N_3749,N_587,N_1374);
nand U3750 (N_3750,N_1971,N_868);
nor U3751 (N_3751,N_1207,N_1773);
xnor U3752 (N_3752,N_900,N_406);
nand U3753 (N_3753,N_739,N_1925);
nor U3754 (N_3754,N_221,N_1318);
nor U3755 (N_3755,N_276,N_502);
or U3756 (N_3756,N_62,N_1955);
nand U3757 (N_3757,N_400,N_1512);
xor U3758 (N_3758,N_15,N_941);
nand U3759 (N_3759,N_1842,N_817);
xor U3760 (N_3760,N_1608,N_1861);
xnor U3761 (N_3761,N_423,N_534);
nor U3762 (N_3762,N_1165,N_434);
xor U3763 (N_3763,N_1660,N_1917);
or U3764 (N_3764,N_1721,N_1150);
xnor U3765 (N_3765,N_546,N_879);
and U3766 (N_3766,N_388,N_1710);
or U3767 (N_3767,N_836,N_523);
nand U3768 (N_3768,N_494,N_231);
or U3769 (N_3769,N_970,N_781);
nand U3770 (N_3770,N_1500,N_1233);
and U3771 (N_3771,N_1282,N_217);
xor U3772 (N_3772,N_672,N_619);
xor U3773 (N_3773,N_83,N_827);
or U3774 (N_3774,N_487,N_1247);
xor U3775 (N_3775,N_1579,N_1911);
xnor U3776 (N_3776,N_368,N_1669);
nor U3777 (N_3777,N_1954,N_523);
nor U3778 (N_3778,N_1069,N_1131);
nor U3779 (N_3779,N_1414,N_19);
xnor U3780 (N_3780,N_915,N_1758);
or U3781 (N_3781,N_1189,N_328);
or U3782 (N_3782,N_1471,N_471);
xor U3783 (N_3783,N_654,N_1119);
or U3784 (N_3784,N_335,N_1769);
nor U3785 (N_3785,N_5,N_713);
xor U3786 (N_3786,N_947,N_1026);
nor U3787 (N_3787,N_993,N_1687);
nor U3788 (N_3788,N_227,N_686);
or U3789 (N_3789,N_1675,N_1708);
or U3790 (N_3790,N_1206,N_1960);
or U3791 (N_3791,N_590,N_735);
xor U3792 (N_3792,N_1351,N_67);
xnor U3793 (N_3793,N_1525,N_985);
and U3794 (N_3794,N_229,N_1902);
and U3795 (N_3795,N_305,N_1221);
nor U3796 (N_3796,N_178,N_149);
nor U3797 (N_3797,N_1547,N_1433);
xor U3798 (N_3798,N_748,N_423);
xor U3799 (N_3799,N_1354,N_995);
or U3800 (N_3800,N_434,N_1917);
and U3801 (N_3801,N_1317,N_1256);
xor U3802 (N_3802,N_503,N_910);
nor U3803 (N_3803,N_471,N_1335);
nand U3804 (N_3804,N_1677,N_1505);
and U3805 (N_3805,N_943,N_529);
nand U3806 (N_3806,N_1631,N_1482);
or U3807 (N_3807,N_1445,N_1381);
and U3808 (N_3808,N_1078,N_1139);
or U3809 (N_3809,N_953,N_1646);
nor U3810 (N_3810,N_813,N_85);
nand U3811 (N_3811,N_1396,N_52);
nand U3812 (N_3812,N_680,N_1478);
nor U3813 (N_3813,N_472,N_454);
nand U3814 (N_3814,N_1754,N_1054);
nand U3815 (N_3815,N_1196,N_1546);
nor U3816 (N_3816,N_1581,N_117);
nor U3817 (N_3817,N_917,N_689);
xnor U3818 (N_3818,N_918,N_17);
nand U3819 (N_3819,N_1798,N_1734);
xnor U3820 (N_3820,N_539,N_358);
and U3821 (N_3821,N_1633,N_356);
and U3822 (N_3822,N_1722,N_789);
nor U3823 (N_3823,N_112,N_1727);
nor U3824 (N_3824,N_1323,N_1154);
nor U3825 (N_3825,N_1211,N_1484);
or U3826 (N_3826,N_1371,N_727);
xnor U3827 (N_3827,N_249,N_772);
nand U3828 (N_3828,N_1499,N_1069);
nor U3829 (N_3829,N_419,N_1363);
nand U3830 (N_3830,N_1961,N_930);
xor U3831 (N_3831,N_1386,N_1560);
and U3832 (N_3832,N_380,N_1120);
or U3833 (N_3833,N_709,N_1875);
or U3834 (N_3834,N_693,N_1641);
and U3835 (N_3835,N_1881,N_923);
xnor U3836 (N_3836,N_522,N_132);
nor U3837 (N_3837,N_135,N_507);
nor U3838 (N_3838,N_730,N_1512);
or U3839 (N_3839,N_592,N_123);
xnor U3840 (N_3840,N_1810,N_233);
xor U3841 (N_3841,N_1347,N_1142);
nor U3842 (N_3842,N_1652,N_1319);
nand U3843 (N_3843,N_1184,N_1070);
nand U3844 (N_3844,N_33,N_661);
nand U3845 (N_3845,N_1979,N_1914);
nand U3846 (N_3846,N_262,N_1502);
and U3847 (N_3847,N_1924,N_1091);
and U3848 (N_3848,N_778,N_70);
and U3849 (N_3849,N_693,N_1849);
nand U3850 (N_3850,N_1428,N_1237);
or U3851 (N_3851,N_766,N_382);
nand U3852 (N_3852,N_1283,N_599);
or U3853 (N_3853,N_563,N_1837);
xnor U3854 (N_3854,N_1091,N_97);
xnor U3855 (N_3855,N_1356,N_1339);
and U3856 (N_3856,N_1648,N_1225);
xnor U3857 (N_3857,N_107,N_1586);
xnor U3858 (N_3858,N_1971,N_618);
xor U3859 (N_3859,N_1971,N_822);
or U3860 (N_3860,N_818,N_1410);
or U3861 (N_3861,N_874,N_317);
or U3862 (N_3862,N_846,N_1508);
xor U3863 (N_3863,N_1606,N_860);
nor U3864 (N_3864,N_1729,N_1451);
nand U3865 (N_3865,N_243,N_1774);
nor U3866 (N_3866,N_817,N_1017);
xor U3867 (N_3867,N_1650,N_1493);
nand U3868 (N_3868,N_1435,N_1785);
and U3869 (N_3869,N_1100,N_1282);
nor U3870 (N_3870,N_204,N_1169);
xor U3871 (N_3871,N_1293,N_436);
and U3872 (N_3872,N_541,N_1998);
and U3873 (N_3873,N_969,N_762);
nor U3874 (N_3874,N_1203,N_1989);
nor U3875 (N_3875,N_685,N_1254);
and U3876 (N_3876,N_140,N_1069);
or U3877 (N_3877,N_685,N_832);
nand U3878 (N_3878,N_1385,N_44);
and U3879 (N_3879,N_1048,N_1303);
xnor U3880 (N_3880,N_793,N_1908);
or U3881 (N_3881,N_1801,N_207);
or U3882 (N_3882,N_753,N_1722);
xor U3883 (N_3883,N_145,N_996);
or U3884 (N_3884,N_699,N_602);
and U3885 (N_3885,N_1325,N_942);
or U3886 (N_3886,N_622,N_694);
xnor U3887 (N_3887,N_74,N_334);
nand U3888 (N_3888,N_1347,N_1094);
and U3889 (N_3889,N_1098,N_48);
and U3890 (N_3890,N_1008,N_1816);
xnor U3891 (N_3891,N_1109,N_1437);
nand U3892 (N_3892,N_1706,N_1439);
nand U3893 (N_3893,N_1566,N_52);
and U3894 (N_3894,N_1198,N_1150);
xnor U3895 (N_3895,N_1231,N_111);
or U3896 (N_3896,N_1953,N_424);
and U3897 (N_3897,N_1007,N_1091);
nand U3898 (N_3898,N_961,N_184);
xnor U3899 (N_3899,N_630,N_1297);
and U3900 (N_3900,N_1631,N_613);
xnor U3901 (N_3901,N_1707,N_564);
and U3902 (N_3902,N_310,N_412);
and U3903 (N_3903,N_1599,N_666);
nand U3904 (N_3904,N_47,N_1181);
nand U3905 (N_3905,N_1298,N_1679);
nor U3906 (N_3906,N_1265,N_311);
xnor U3907 (N_3907,N_362,N_1553);
and U3908 (N_3908,N_373,N_1783);
nand U3909 (N_3909,N_720,N_1277);
nor U3910 (N_3910,N_1209,N_1510);
and U3911 (N_3911,N_1872,N_560);
and U3912 (N_3912,N_179,N_1105);
and U3913 (N_3913,N_587,N_1448);
xnor U3914 (N_3914,N_1306,N_849);
nand U3915 (N_3915,N_1020,N_1516);
nor U3916 (N_3916,N_528,N_999);
nand U3917 (N_3917,N_253,N_1622);
or U3918 (N_3918,N_1101,N_1469);
and U3919 (N_3919,N_1684,N_1333);
and U3920 (N_3920,N_431,N_173);
and U3921 (N_3921,N_354,N_146);
or U3922 (N_3922,N_1250,N_1215);
nand U3923 (N_3923,N_920,N_1893);
nor U3924 (N_3924,N_378,N_516);
xor U3925 (N_3925,N_1737,N_855);
xnor U3926 (N_3926,N_1328,N_1179);
and U3927 (N_3927,N_108,N_1917);
and U3928 (N_3928,N_723,N_769);
and U3929 (N_3929,N_1725,N_49);
nand U3930 (N_3930,N_1627,N_1161);
xnor U3931 (N_3931,N_201,N_1359);
xor U3932 (N_3932,N_890,N_1112);
and U3933 (N_3933,N_1433,N_222);
or U3934 (N_3934,N_1635,N_1210);
nand U3935 (N_3935,N_81,N_1965);
and U3936 (N_3936,N_954,N_1339);
nand U3937 (N_3937,N_861,N_381);
and U3938 (N_3938,N_1965,N_1254);
and U3939 (N_3939,N_533,N_1022);
and U3940 (N_3940,N_1307,N_1179);
and U3941 (N_3941,N_1273,N_684);
xnor U3942 (N_3942,N_84,N_6);
xor U3943 (N_3943,N_604,N_1926);
nor U3944 (N_3944,N_1736,N_1913);
xor U3945 (N_3945,N_847,N_207);
nor U3946 (N_3946,N_302,N_453);
nor U3947 (N_3947,N_1637,N_503);
and U3948 (N_3948,N_779,N_1545);
nand U3949 (N_3949,N_1552,N_636);
nand U3950 (N_3950,N_815,N_710);
and U3951 (N_3951,N_466,N_1073);
nor U3952 (N_3952,N_1811,N_1432);
nor U3953 (N_3953,N_1438,N_461);
nand U3954 (N_3954,N_147,N_1054);
nand U3955 (N_3955,N_63,N_161);
nand U3956 (N_3956,N_1238,N_1681);
nand U3957 (N_3957,N_239,N_358);
or U3958 (N_3958,N_1264,N_926);
nor U3959 (N_3959,N_1976,N_53);
nor U3960 (N_3960,N_544,N_1556);
or U3961 (N_3961,N_904,N_767);
or U3962 (N_3962,N_1821,N_1448);
or U3963 (N_3963,N_929,N_309);
and U3964 (N_3964,N_892,N_421);
xnor U3965 (N_3965,N_1521,N_1734);
nor U3966 (N_3966,N_185,N_189);
and U3967 (N_3967,N_1703,N_889);
xnor U3968 (N_3968,N_1676,N_701);
or U3969 (N_3969,N_18,N_699);
nor U3970 (N_3970,N_1218,N_101);
nor U3971 (N_3971,N_540,N_1255);
nand U3972 (N_3972,N_227,N_1070);
or U3973 (N_3973,N_976,N_500);
xor U3974 (N_3974,N_1601,N_1403);
or U3975 (N_3975,N_1157,N_1937);
and U3976 (N_3976,N_953,N_296);
nor U3977 (N_3977,N_1633,N_402);
nor U3978 (N_3978,N_694,N_376);
nor U3979 (N_3979,N_1409,N_1125);
xnor U3980 (N_3980,N_625,N_1725);
or U3981 (N_3981,N_1947,N_1595);
xor U3982 (N_3982,N_1474,N_1373);
or U3983 (N_3983,N_1410,N_1136);
nand U3984 (N_3984,N_1274,N_274);
nand U3985 (N_3985,N_1734,N_1039);
or U3986 (N_3986,N_832,N_280);
nand U3987 (N_3987,N_311,N_550);
nand U3988 (N_3988,N_123,N_1552);
nor U3989 (N_3989,N_667,N_1973);
and U3990 (N_3990,N_404,N_1126);
xor U3991 (N_3991,N_1921,N_1543);
and U3992 (N_3992,N_354,N_1343);
nand U3993 (N_3993,N_18,N_1646);
xor U3994 (N_3994,N_1826,N_373);
and U3995 (N_3995,N_1414,N_1579);
nor U3996 (N_3996,N_1333,N_1002);
and U3997 (N_3997,N_322,N_135);
nand U3998 (N_3998,N_912,N_248);
or U3999 (N_3999,N_1033,N_697);
and U4000 (N_4000,N_3980,N_2759);
and U4001 (N_4001,N_2775,N_2559);
or U4002 (N_4002,N_2918,N_3383);
or U4003 (N_4003,N_3511,N_3038);
nand U4004 (N_4004,N_2963,N_3378);
and U4005 (N_4005,N_2968,N_3055);
nor U4006 (N_4006,N_3914,N_3426);
xor U4007 (N_4007,N_3606,N_3657);
and U4008 (N_4008,N_2419,N_3146);
nor U4009 (N_4009,N_3185,N_3621);
and U4010 (N_4010,N_2610,N_3842);
nand U4011 (N_4011,N_2232,N_2946);
nand U4012 (N_4012,N_3030,N_3619);
xnor U4013 (N_4013,N_2536,N_3673);
or U4014 (N_4014,N_2062,N_3970);
nor U4015 (N_4015,N_2579,N_2924);
nor U4016 (N_4016,N_3603,N_3044);
nor U4017 (N_4017,N_2582,N_3637);
xor U4018 (N_4018,N_2371,N_3248);
nor U4019 (N_4019,N_2225,N_3157);
xor U4020 (N_4020,N_2233,N_2736);
and U4021 (N_4021,N_2004,N_3547);
nand U4022 (N_4022,N_2838,N_3416);
nor U4023 (N_4023,N_3591,N_3093);
nand U4024 (N_4024,N_2256,N_3481);
and U4025 (N_4025,N_2608,N_3176);
xor U4026 (N_4026,N_3404,N_2278);
or U4027 (N_4027,N_2063,N_3679);
nand U4028 (N_4028,N_2190,N_2722);
or U4029 (N_4029,N_2065,N_2088);
xor U4030 (N_4030,N_2658,N_3908);
or U4031 (N_4031,N_3658,N_3995);
nor U4032 (N_4032,N_2896,N_2200);
and U4033 (N_4033,N_3526,N_3598);
nor U4034 (N_4034,N_2712,N_3401);
xor U4035 (N_4035,N_2217,N_2417);
nand U4036 (N_4036,N_3871,N_3830);
or U4037 (N_4037,N_2038,N_2344);
nor U4038 (N_4038,N_2050,N_3453);
and U4039 (N_4039,N_2377,N_2603);
xor U4040 (N_4040,N_2290,N_2202);
or U4041 (N_4041,N_3990,N_2051);
xnor U4042 (N_4042,N_2273,N_3384);
nor U4043 (N_4043,N_3766,N_3741);
and U4044 (N_4044,N_2335,N_3133);
or U4045 (N_4045,N_2412,N_2984);
nand U4046 (N_4046,N_3262,N_2270);
xnor U4047 (N_4047,N_2828,N_2034);
nand U4048 (N_4048,N_2201,N_2856);
and U4049 (N_4049,N_2053,N_2614);
or U4050 (N_4050,N_2750,N_2823);
nand U4051 (N_4051,N_2199,N_2816);
nand U4052 (N_4052,N_3282,N_2011);
nand U4053 (N_4053,N_2995,N_3186);
and U4054 (N_4054,N_3764,N_3541);
and U4055 (N_4055,N_2863,N_3010);
nand U4056 (N_4056,N_2370,N_2799);
and U4057 (N_4057,N_3145,N_3777);
xnor U4058 (N_4058,N_2134,N_2627);
xor U4059 (N_4059,N_3376,N_3554);
and U4060 (N_4060,N_2133,N_3942);
or U4061 (N_4061,N_2393,N_2709);
nand U4062 (N_4062,N_3045,N_3821);
and U4063 (N_4063,N_2169,N_2840);
nor U4064 (N_4064,N_3791,N_3179);
or U4065 (N_4065,N_3999,N_3004);
nand U4066 (N_4066,N_3775,N_2293);
nor U4067 (N_4067,N_3696,N_2623);
xor U4068 (N_4068,N_2814,N_3820);
xnor U4069 (N_4069,N_3206,N_3706);
nor U4070 (N_4070,N_2472,N_2884);
xor U4071 (N_4071,N_2656,N_3497);
nand U4072 (N_4072,N_2756,N_3704);
nor U4073 (N_4073,N_3827,N_2299);
nor U4074 (N_4074,N_2470,N_2532);
or U4075 (N_4075,N_3243,N_3850);
and U4076 (N_4076,N_2915,N_3337);
or U4077 (N_4077,N_3031,N_2020);
or U4078 (N_4078,N_2301,N_2967);
and U4079 (N_4079,N_3600,N_3237);
and U4080 (N_4080,N_2633,N_3869);
xnor U4081 (N_4081,N_2556,N_3490);
xnor U4082 (N_4082,N_3506,N_3046);
nor U4083 (N_4083,N_3608,N_3252);
or U4084 (N_4084,N_3952,N_3149);
and U4085 (N_4085,N_3319,N_3596);
and U4086 (N_4086,N_3408,N_2499);
or U4087 (N_4087,N_3551,N_3972);
xor U4088 (N_4088,N_3859,N_2731);
or U4089 (N_4089,N_2367,N_2832);
or U4090 (N_4090,N_3000,N_3702);
and U4091 (N_4091,N_3323,N_2643);
or U4092 (N_4092,N_3566,N_3677);
nor U4093 (N_4093,N_3686,N_2860);
and U4094 (N_4094,N_2303,N_3778);
or U4095 (N_4095,N_3504,N_3560);
xor U4096 (N_4096,N_3421,N_3937);
xor U4097 (N_4097,N_3205,N_3641);
nor U4098 (N_4098,N_3138,N_2309);
nor U4099 (N_4099,N_3982,N_2476);
and U4100 (N_4100,N_3835,N_3140);
nand U4101 (N_4101,N_3794,N_3062);
nor U4102 (N_4102,N_2418,N_2404);
xor U4103 (N_4103,N_3544,N_3328);
or U4104 (N_4104,N_3259,N_2167);
nand U4105 (N_4105,N_3348,N_2176);
and U4106 (N_4106,N_3315,N_3210);
xnor U4107 (N_4107,N_3214,N_2017);
and U4108 (N_4108,N_3695,N_2466);
and U4109 (N_4109,N_2369,N_2933);
nor U4110 (N_4110,N_3187,N_3856);
nand U4111 (N_4111,N_2467,N_3082);
nor U4112 (N_4112,N_3690,N_3585);
and U4113 (N_4113,N_2776,N_2526);
or U4114 (N_4114,N_3570,N_3251);
nand U4115 (N_4115,N_2577,N_2573);
nand U4116 (N_4116,N_3838,N_2972);
and U4117 (N_4117,N_2347,N_2649);
xor U4118 (N_4118,N_2315,N_2283);
xor U4119 (N_4119,N_3447,N_2935);
or U4120 (N_4120,N_2405,N_2235);
nor U4121 (N_4121,N_3986,N_3960);
nor U4122 (N_4122,N_2906,N_2005);
nand U4123 (N_4123,N_2937,N_2558);
xor U4124 (N_4124,N_2433,N_3685);
nand U4125 (N_4125,N_3051,N_2626);
xor U4126 (N_4126,N_3022,N_3098);
nor U4127 (N_4127,N_3254,N_2247);
nor U4128 (N_4128,N_3195,N_2879);
nand U4129 (N_4129,N_3762,N_2465);
or U4130 (N_4130,N_3099,N_3088);
and U4131 (N_4131,N_2964,N_3208);
and U4132 (N_4132,N_3671,N_2978);
or U4133 (N_4133,N_2222,N_2187);
and U4134 (N_4134,N_2302,N_2274);
nand U4135 (N_4135,N_2109,N_3819);
or U4136 (N_4136,N_2146,N_3423);
xnor U4137 (N_4137,N_3301,N_2878);
and U4138 (N_4138,N_3634,N_3441);
xor U4139 (N_4139,N_3433,N_2394);
xnor U4140 (N_4140,N_2230,N_3876);
or U4141 (N_4141,N_3825,N_3321);
nand U4142 (N_4142,N_3666,N_2236);
xor U4143 (N_4143,N_3734,N_3979);
xor U4144 (N_4144,N_3412,N_2009);
or U4145 (N_4145,N_3805,N_3998);
nand U4146 (N_4146,N_2920,N_3297);
xor U4147 (N_4147,N_3240,N_2154);
xnor U4148 (N_4148,N_3957,N_3019);
or U4149 (N_4149,N_2031,N_2681);
or U4150 (N_4150,N_2339,N_3236);
or U4151 (N_4151,N_2568,N_3147);
nor U4152 (N_4152,N_2458,N_2027);
and U4153 (N_4153,N_3953,N_3443);
xor U4154 (N_4154,N_3245,N_2834);
or U4155 (N_4155,N_2672,N_2553);
xor U4156 (N_4156,N_2077,N_2368);
or U4157 (N_4157,N_3002,N_3509);
and U4158 (N_4158,N_2671,N_3562);
xor U4159 (N_4159,N_2080,N_2811);
or U4160 (N_4160,N_3875,N_3610);
xnor U4161 (N_4161,N_3189,N_3058);
or U4162 (N_4162,N_3060,N_2748);
or U4163 (N_4163,N_2231,N_2598);
or U4164 (N_4164,N_2121,N_2426);
nand U4165 (N_4165,N_2488,N_2525);
and U4166 (N_4166,N_3811,N_2836);
and U4167 (N_4167,N_2508,N_3561);
xor U4168 (N_4168,N_2818,N_3633);
and U4169 (N_4169,N_3703,N_3933);
nor U4170 (N_4170,N_2351,N_2961);
nand U4171 (N_4171,N_3755,N_3445);
nor U4172 (N_4172,N_2437,N_3353);
or U4173 (N_4173,N_3760,N_2527);
and U4174 (N_4174,N_2079,N_3284);
or U4175 (N_4175,N_3693,N_2300);
nor U4176 (N_4176,N_3689,N_3883);
nor U4177 (N_4177,N_3527,N_2755);
xnor U4178 (N_4178,N_2735,N_3097);
and U4179 (N_4179,N_3091,N_2443);
xor U4180 (N_4180,N_3020,N_2766);
nor U4181 (N_4181,N_3751,N_2903);
or U4182 (N_4182,N_3718,N_2827);
or U4183 (N_4183,N_2621,N_2342);
and U4184 (N_4184,N_2061,N_2664);
xor U4185 (N_4185,N_3951,N_3308);
and U4186 (N_4186,N_3705,N_2260);
nor U4187 (N_4187,N_3122,N_3283);
or U4188 (N_4188,N_3087,N_3723);
or U4189 (N_4189,N_2809,N_3203);
and U4190 (N_4190,N_3799,N_2422);
nand U4191 (N_4191,N_2689,N_2587);
or U4192 (N_4192,N_2846,N_2208);
and U4193 (N_4193,N_3474,N_3041);
and U4194 (N_4194,N_2782,N_3984);
nand U4195 (N_4195,N_3391,N_2126);
nor U4196 (N_4196,N_3161,N_3128);
nor U4197 (N_4197,N_2228,N_2817);
or U4198 (N_4198,N_3272,N_3069);
or U4199 (N_4199,N_2075,N_3491);
xnor U4200 (N_4200,N_3967,N_3246);
nand U4201 (N_4201,N_3430,N_3406);
nand U4202 (N_4202,N_2287,N_3784);
or U4203 (N_4203,N_3191,N_3450);
or U4204 (N_4204,N_3064,N_2153);
and U4205 (N_4205,N_3899,N_3398);
nor U4206 (N_4206,N_2333,N_2789);
or U4207 (N_4207,N_3171,N_3074);
nand U4208 (N_4208,N_3571,N_2956);
or U4209 (N_4209,N_2641,N_3235);
nor U4210 (N_4210,N_2000,N_2498);
xnor U4211 (N_4211,N_3017,N_3556);
nand U4212 (N_4212,N_2446,N_3722);
nand U4213 (N_4213,N_2701,N_2890);
or U4214 (N_4214,N_3878,N_2854);
xnor U4215 (N_4215,N_2706,N_3650);
nor U4216 (N_4216,N_2787,N_2067);
or U4217 (N_4217,N_2866,N_2171);
or U4218 (N_4218,N_3399,N_2459);
nor U4219 (N_4219,N_3977,N_2308);
xnor U4220 (N_4220,N_2557,N_2191);
or U4221 (N_4221,N_2039,N_2486);
nor U4222 (N_4222,N_3867,N_3912);
xor U4223 (N_4223,N_3949,N_3273);
and U4224 (N_4224,N_3873,N_2534);
and U4225 (N_4225,N_2055,N_2469);
or U4226 (N_4226,N_2207,N_2698);
and U4227 (N_4227,N_2742,N_3846);
nand U4228 (N_4228,N_3253,N_2117);
nor U4229 (N_4229,N_2506,N_2630);
nor U4230 (N_4230,N_2489,N_2427);
nand U4231 (N_4231,N_2043,N_2380);
nand U4232 (N_4232,N_2639,N_2304);
xor U4233 (N_4233,N_2733,N_2564);
nand U4234 (N_4234,N_3050,N_3851);
or U4235 (N_4235,N_2364,N_3213);
nor U4236 (N_4236,N_2373,N_3137);
and U4237 (N_4237,N_2528,N_2897);
nor U4238 (N_4238,N_3743,N_3148);
or U4239 (N_4239,N_2276,N_2661);
and U4240 (N_4240,N_2788,N_2562);
or U4241 (N_4241,N_3539,N_3033);
nand U4242 (N_4242,N_3484,N_2849);
nand U4243 (N_4243,N_2583,N_2068);
or U4244 (N_4244,N_3409,N_3455);
and U4245 (N_4245,N_3644,N_3520);
nand U4246 (N_4246,N_3809,N_3864);
nor U4247 (N_4247,N_2830,N_3968);
nand U4248 (N_4248,N_2986,N_3763);
xor U4249 (N_4249,N_2471,N_3535);
nor U4250 (N_4250,N_2275,N_3954);
and U4251 (N_4251,N_3040,N_2606);
nor U4252 (N_4252,N_3394,N_3363);
nand U4253 (N_4253,N_2574,N_3325);
nor U4254 (N_4254,N_3672,N_2994);
nor U4255 (N_4255,N_3215,N_3026);
nor U4256 (N_4256,N_3475,N_3569);
xnor U4257 (N_4257,N_2631,N_2548);
xnor U4258 (N_4258,N_2518,N_3915);
nor U4259 (N_4259,N_2522,N_3260);
and U4260 (N_4260,N_2494,N_2460);
nand U4261 (N_4261,N_3513,N_2353);
nand U4262 (N_4262,N_2271,N_2179);
nand U4263 (N_4263,N_3745,N_3141);
xor U4264 (N_4264,N_3897,N_2045);
and U4265 (N_4265,N_2040,N_3266);
xnor U4266 (N_4266,N_2173,N_3229);
nand U4267 (N_4267,N_3865,N_2195);
and U4268 (N_4268,N_2008,N_3564);
nand U4269 (N_4269,N_2395,N_3126);
or U4270 (N_4270,N_2461,N_2944);
and U4271 (N_4271,N_2957,N_2086);
xnor U4272 (N_4272,N_2729,N_3334);
nor U4273 (N_4273,N_3346,N_3521);
and U4274 (N_4274,N_3369,N_2035);
nor U4275 (N_4275,N_3715,N_2138);
nor U4276 (N_4276,N_2220,N_3293);
and U4277 (N_4277,N_3663,N_2763);
nor U4278 (N_4278,N_2592,N_3837);
or U4279 (N_4279,N_3962,N_3710);
xnor U4280 (N_4280,N_2674,N_3776);
xor U4281 (N_4281,N_3316,N_2769);
nor U4282 (N_4282,N_2640,N_2455);
nand U4283 (N_4283,N_2248,N_2703);
and U4284 (N_4284,N_3936,N_2473);
nand U4285 (N_4285,N_3639,N_2699);
xnor U4286 (N_4286,N_2919,N_3713);
xor U4287 (N_4287,N_3312,N_3559);
nand U4288 (N_4288,N_3437,N_2194);
nand U4289 (N_4289,N_2772,N_2490);
nand U4290 (N_4290,N_3368,N_2747);
nor U4291 (N_4291,N_2148,N_2928);
and U4292 (N_4292,N_2491,N_2997);
nor U4293 (N_4293,N_3701,N_3750);
xnor U4294 (N_4294,N_3540,N_2487);
nand U4295 (N_4295,N_2975,N_2162);
nand U4296 (N_4296,N_3356,N_3172);
and U4297 (N_4297,N_3365,N_2588);
or U4298 (N_4298,N_2873,N_3056);
and U4299 (N_4299,N_2916,N_3893);
xor U4300 (N_4300,N_2687,N_2533);
nor U4301 (N_4301,N_2341,N_3495);
or U4302 (N_4302,N_3861,N_3277);
or U4303 (N_4303,N_3773,N_2001);
xnor U4304 (N_4304,N_2358,N_3855);
nand U4305 (N_4305,N_2032,N_2507);
or U4306 (N_4306,N_3959,N_3920);
nand U4307 (N_4307,N_3467,N_2156);
and U4308 (N_4308,N_3863,N_2815);
and U4309 (N_4309,N_2211,N_2806);
nand U4310 (N_4310,N_2106,N_2773);
nand U4311 (N_4311,N_3971,N_3529);
and U4312 (N_4312,N_2657,N_2645);
xor U4313 (N_4313,N_3158,N_3400);
nor U4314 (N_4314,N_2611,N_2695);
xor U4315 (N_4315,N_3083,N_3654);
or U4316 (N_4316,N_3357,N_2110);
xnor U4317 (N_4317,N_3119,N_2252);
xor U4318 (N_4318,N_2646,N_3395);
nand U4319 (N_4319,N_3815,N_3168);
nand U4320 (N_4320,N_3270,N_3349);
xor U4321 (N_4321,N_2655,N_2165);
xnor U4322 (N_4322,N_3742,N_3879);
nand U4323 (N_4323,N_2145,N_3910);
xor U4324 (N_4324,N_3802,N_2683);
and U4325 (N_4325,N_3358,N_3182);
nand U4326 (N_4326,N_3068,N_3623);
xor U4327 (N_4327,N_2170,N_2740);
xnor U4328 (N_4328,N_3862,N_2399);
nor U4329 (N_4329,N_3813,N_2667);
xor U4330 (N_4330,N_2060,N_2547);
or U4331 (N_4331,N_2496,N_3996);
xor U4332 (N_4332,N_2431,N_2238);
and U4333 (N_4333,N_3785,N_2069);
and U4334 (N_4334,N_2976,N_3525);
and U4335 (N_4335,N_2820,N_2666);
nand U4336 (N_4336,N_3156,N_3110);
or U4337 (N_4337,N_3546,N_2006);
and U4338 (N_4338,N_3220,N_3294);
nor U4339 (N_4339,N_2087,N_2163);
nor U4340 (N_4340,N_3906,N_3003);
nor U4341 (N_4341,N_3482,N_2842);
or U4342 (N_4342,N_2861,N_3303);
xnor U4343 (N_4343,N_3488,N_2240);
or U4344 (N_4344,N_3070,N_3039);
xnor U4345 (N_4345,N_3287,N_2673);
xnor U4346 (N_4346,N_2223,N_2453);
and U4347 (N_4347,N_3162,N_3667);
nand U4348 (N_4348,N_2441,N_2242);
nand U4349 (N_4349,N_2241,N_3190);
xnor U4350 (N_4350,N_3987,N_3749);
xor U4351 (N_4351,N_2929,N_3515);
nand U4352 (N_4352,N_3023,N_3054);
nor U4353 (N_4353,N_2479,N_2572);
xnor U4354 (N_4354,N_2932,N_2285);
or U4355 (N_4355,N_3422,N_2177);
nand U4356 (N_4356,N_2057,N_2795);
xor U4357 (N_4357,N_2883,N_3752);
nor U4358 (N_4358,N_3975,N_2350);
nor U4359 (N_4359,N_3106,N_3001);
nand U4360 (N_4360,N_2119,N_2651);
and U4361 (N_4361,N_2938,N_3940);
nand U4362 (N_4362,N_2741,N_3793);
xor U4363 (N_4363,N_3196,N_3170);
or U4364 (N_4364,N_3613,N_2103);
and U4365 (N_4365,N_3945,N_2048);
nand U4366 (N_4366,N_3903,N_3675);
or U4367 (N_4367,N_3227,N_3913);
nor U4368 (N_4368,N_2375,N_3787);
nor U4369 (N_4369,N_2124,N_2073);
or U4370 (N_4370,N_2922,N_2591);
nor U4371 (N_4371,N_3573,N_2844);
or U4372 (N_4372,N_2286,N_3563);
or U4373 (N_4373,N_3011,N_3670);
nand U4374 (N_4374,N_2804,N_3928);
xnor U4375 (N_4375,N_3981,N_2615);
and U4376 (N_4376,N_2497,N_3923);
xor U4377 (N_4377,N_3514,N_2974);
nor U4378 (N_4378,N_2780,N_2680);
nor U4379 (N_4379,N_3769,N_3456);
nand U4380 (N_4380,N_3342,N_3688);
or U4381 (N_4381,N_2839,N_2737);
nor U4382 (N_4382,N_2535,N_2074);
or U4383 (N_4383,N_2561,N_2540);
nand U4384 (N_4384,N_2677,N_2852);
or U4385 (N_4385,N_2585,N_3275);
or U4386 (N_4386,N_2600,N_3372);
or U4387 (N_4387,N_3052,N_3057);
and U4388 (N_4388,N_2136,N_3592);
xnor U4389 (N_4389,N_2529,N_3405);
nor U4390 (N_4390,N_3567,N_2679);
xnor U4391 (N_4391,N_3896,N_2684);
xor U4392 (N_4392,N_2291,N_2829);
nor U4393 (N_4393,N_3305,N_3084);
xnor U4394 (N_4394,N_3646,N_3717);
xnor U4395 (N_4395,N_3225,N_3343);
xnor U4396 (N_4396,N_3507,N_3605);
nand U4397 (N_4397,N_2337,N_2093);
nor U4398 (N_4398,N_3403,N_3332);
nor U4399 (N_4399,N_2594,N_2140);
or U4400 (N_4400,N_2531,N_2714);
nand U4401 (N_4401,N_3618,N_3034);
or U4402 (N_4402,N_2987,N_3770);
nor U4403 (N_4403,N_3911,N_2098);
nor U4404 (N_4404,N_3310,N_3586);
nand U4405 (N_4405,N_3108,N_3007);
nand U4406 (N_4406,N_2041,N_2962);
and U4407 (N_4407,N_2777,N_3655);
xor U4408 (N_4408,N_3938,N_2143);
nand U4409 (N_4409,N_2357,N_3738);
nand U4410 (N_4410,N_2316,N_2175);
and U4411 (N_4411,N_2253,N_3111);
nand U4412 (N_4412,N_2764,N_2949);
or U4413 (N_4413,N_2127,N_3134);
and U4414 (N_4414,N_2147,N_2930);
xor U4415 (N_4415,N_2663,N_3241);
or U4416 (N_4416,N_2193,N_2477);
or U4417 (N_4417,N_3027,N_2899);
xnor U4418 (N_4418,N_3201,N_2758);
nand U4419 (N_4419,N_2660,N_3796);
xnor U4420 (N_4420,N_3531,N_3988);
and U4421 (N_4421,N_3468,N_2851);
or U4422 (N_4422,N_3373,N_2678);
or U4423 (N_4423,N_2837,N_3891);
or U4424 (N_4424,N_3816,N_2096);
nor U4425 (N_4425,N_2909,N_3402);
xnor U4426 (N_4426,N_2910,N_2255);
nand U4427 (N_4427,N_3744,N_2993);
nor U4428 (N_4428,N_2186,N_2210);
nor U4429 (N_4429,N_2013,N_2421);
nand U4430 (N_4430,N_2317,N_2139);
and U4431 (N_4431,N_3708,N_2181);
xor U4432 (N_4432,N_2189,N_2152);
or U4433 (N_4433,N_3032,N_3609);
xnor U4434 (N_4434,N_3322,N_2372);
nand U4435 (N_4435,N_3188,N_2882);
or U4436 (N_4436,N_3700,N_2708);
xnor U4437 (N_4437,N_3333,N_3800);
nand U4438 (N_4438,N_3094,N_3807);
xor U4439 (N_4439,N_3848,N_3905);
or U4440 (N_4440,N_2894,N_2696);
nor U4441 (N_4441,N_2354,N_3442);
nor U4442 (N_4442,N_2757,N_2575);
nor U4443 (N_4443,N_2590,N_2734);
and U4444 (N_4444,N_2485,N_2454);
and U4445 (N_4445,N_3503,N_2468);
nand U4446 (N_4446,N_3264,N_2841);
nor U4447 (N_4447,N_3089,N_2563);
nand U4448 (N_4448,N_3510,N_2280);
nand U4449 (N_4449,N_2545,N_2745);
and U4450 (N_4450,N_3042,N_2444);
xnor U4451 (N_4451,N_3868,N_3197);
nand U4452 (N_4452,N_2765,N_2346);
xor U4453 (N_4453,N_3828,N_2900);
and U4454 (N_4454,N_3096,N_2613);
nor U4455 (N_4455,N_3462,N_3350);
nand U4456 (N_4456,N_3411,N_3221);
nand U4457 (N_4457,N_2654,N_3486);
xnor U4458 (N_4458,N_2400,N_3013);
or U4459 (N_4459,N_2203,N_2014);
nand U4460 (N_4460,N_3469,N_2898);
xor U4461 (N_4461,N_2693,N_2264);
or U4462 (N_4462,N_3692,N_2783);
or U4463 (N_4463,N_2003,N_2778);
xor U4464 (N_4464,N_2502,N_3651);
xor U4465 (N_4465,N_3530,N_2728);
nor U4466 (N_4466,N_3974,N_2237);
and U4467 (N_4467,N_3247,N_2912);
nand U4468 (N_4468,N_2565,N_3595);
or U4469 (N_4469,N_2505,N_2754);
nand U4470 (N_4470,N_3909,N_3021);
nand U4471 (N_4471,N_2047,N_2616);
nor U4472 (N_4472,N_2249,N_3881);
nand U4473 (N_4473,N_2597,N_3884);
or U4474 (N_4474,N_3662,N_2543);
nand U4475 (N_4475,N_3834,N_2269);
xnor U4476 (N_4476,N_3439,N_3092);
xnor U4477 (N_4477,N_3817,N_2676);
xor U4478 (N_4478,N_2340,N_3839);
and U4479 (N_4479,N_2625,N_3035);
or U4480 (N_4480,N_3077,N_2739);
nor U4481 (N_4481,N_2721,N_2391);
xnor U4482 (N_4482,N_3888,N_3135);
xor U4483 (N_4483,N_3330,N_2101);
nand U4484 (N_4484,N_3360,N_3694);
nand U4485 (N_4485,N_2475,N_2790);
xnor U4486 (N_4486,N_2969,N_3831);
xor U4487 (N_4487,N_3480,N_2212);
nand U4488 (N_4488,N_3582,N_2277);
and U4489 (N_4489,N_2362,N_2807);
nor U4490 (N_4490,N_2746,N_2129);
nand U4491 (N_4491,N_2095,N_2015);
nor U4492 (N_4492,N_3635,N_3028);
or U4493 (N_4493,N_2864,N_2205);
or U4494 (N_4494,N_2917,N_2360);
nand U4495 (N_4495,N_3463,N_3840);
nor U4496 (N_4496,N_3844,N_3757);
or U4497 (N_4497,N_2771,N_3874);
nor U4498 (N_4498,N_3127,N_2125);
nand U4499 (N_4499,N_3533,N_2867);
xnor U4500 (N_4500,N_2180,N_3919);
nand U4501 (N_4501,N_3355,N_3588);
nor U4502 (N_4502,N_2876,N_2516);
nor U4503 (N_4503,N_3025,N_3965);
or U4504 (N_4504,N_2251,N_2066);
and U4505 (N_4505,N_3607,N_3116);
nand U4506 (N_4506,N_2338,N_2719);
nor U4507 (N_4507,N_3917,N_2566);
nor U4508 (N_4508,N_2450,N_2682);
or U4509 (N_4509,N_3120,N_3080);
and U4510 (N_4510,N_2492,N_3081);
xor U4511 (N_4511,N_2183,N_3265);
nor U4512 (N_4512,N_2635,N_3175);
nor U4513 (N_4513,N_3597,N_3173);
and U4514 (N_4514,N_3950,N_2292);
or U4515 (N_4515,N_3900,N_3338);
or U4516 (N_4516,N_2825,N_2523);
xor U4517 (N_4517,N_3076,N_3522);
xnor U4518 (N_4518,N_2297,N_2686);
nand U4519 (N_4519,N_3518,N_3123);
or U4520 (N_4520,N_3307,N_3524);
nor U4521 (N_4521,N_3632,N_2868);
nor U4522 (N_4522,N_3991,N_2311);
nor U4523 (N_4523,N_2442,N_3121);
nand U4524 (N_4524,N_2294,N_3436);
or U4525 (N_4525,N_3396,N_3687);
xnor U4526 (N_4526,N_2348,N_2023);
nand U4527 (N_4527,N_3946,N_3465);
nor U4528 (N_4528,N_2030,N_2911);
xor U4529 (N_4529,N_2859,N_3015);
nand U4530 (N_4530,N_3489,N_3512);
xor U4531 (N_4531,N_3429,N_2213);
and U4532 (N_4532,N_2197,N_2482);
nor U4533 (N_4533,N_3983,N_3494);
nand U4534 (N_4534,N_2174,N_3371);
or U4535 (N_4535,N_2702,N_2717);
xor U4536 (N_4536,N_3024,N_2102);
nor U4537 (N_4537,N_2952,N_3438);
nor U4538 (N_4538,N_2970,N_2797);
nor U4539 (N_4539,N_3709,N_2653);
and U4540 (N_4540,N_2452,N_2259);
xnor U4541 (N_4541,N_2115,N_2385);
nand U4542 (N_4542,N_3499,N_3269);
nand U4543 (N_4543,N_2524,N_3599);
nand U4544 (N_4544,N_3261,N_3166);
or U4545 (N_4545,N_3725,N_2947);
xnor U4546 (N_4546,N_3101,N_2555);
xnor U4547 (N_4547,N_2307,N_3324);
or U4548 (N_4548,N_2150,N_3410);
or U4549 (N_4549,N_3249,N_3178);
nor U4550 (N_4550,N_3647,N_2723);
or U4551 (N_4551,N_3452,N_3801);
nor U4552 (N_4552,N_3558,N_3870);
xor U4553 (N_4553,N_2511,N_2356);
nand U4554 (N_4554,N_3614,N_3545);
xor U4555 (N_4555,N_3483,N_2697);
and U4556 (N_4556,N_3681,N_2111);
nand U4557 (N_4557,N_2435,N_2321);
nor U4558 (N_4558,N_3454,N_3086);
or U4559 (N_4559,N_3318,N_2318);
xnor U4560 (N_4560,N_3579,N_3192);
nor U4561 (N_4561,N_2092,N_2022);
or U4562 (N_4562,N_3072,N_2221);
or U4563 (N_4563,N_2379,N_2891);
xor U4564 (N_4564,N_2082,N_2326);
nor U4565 (N_4565,N_2710,N_3786);
xor U4566 (N_4566,N_3882,N_3291);
nor U4567 (N_4567,N_2243,N_2955);
nor U4568 (N_4568,N_3366,N_2411);
and U4569 (N_4569,N_2659,N_2784);
and U4570 (N_4570,N_3927,N_3783);
and U4571 (N_4571,N_2996,N_2456);
and U4572 (N_4572,N_3841,N_2690);
nor U4573 (N_4573,N_3782,N_3719);
and U4574 (N_4574,N_3103,N_2753);
and U4575 (N_4575,N_2691,N_3218);
and U4576 (N_4576,N_2800,N_3431);
nand U4577 (N_4577,N_2336,N_3219);
nor U4578 (N_4578,N_3823,N_2392);
and U4579 (N_4579,N_2927,N_3994);
or U4580 (N_4580,N_3629,N_2480);
and U4581 (N_4581,N_2361,N_2413);
nand U4582 (N_4582,N_2345,N_3160);
or U4583 (N_4583,N_2512,N_2355);
or U4584 (N_4584,N_3048,N_3552);
and U4585 (N_4585,N_3063,N_2113);
xor U4586 (N_4586,N_2123,N_3362);
nand U4587 (N_4587,N_2546,N_2835);
xor U4588 (N_4588,N_3169,N_2596);
xor U4589 (N_4589,N_2229,N_2711);
nor U4590 (N_4590,N_2282,N_2408);
or U4591 (N_4591,N_3164,N_2382);
nor U4592 (N_4592,N_3890,N_3257);
and U4593 (N_4593,N_2159,N_2390);
xnor U4594 (N_4594,N_3640,N_3536);
xnor U4595 (N_4595,N_3638,N_3313);
nand U4596 (N_4596,N_2637,N_3765);
nand U4597 (N_4597,N_3113,N_3761);
or U4598 (N_4598,N_2327,N_2334);
and U4599 (N_4599,N_2796,N_3887);
xor U4600 (N_4600,N_2137,N_3748);
or U4601 (N_4601,N_2808,N_3726);
nor U4602 (N_4602,N_2705,N_3661);
and U4603 (N_4603,N_2185,N_2449);
xnor U4604 (N_4604,N_2438,N_3012);
or U4605 (N_4605,N_2401,N_2018);
or U4606 (N_4606,N_3387,N_3477);
nor U4607 (N_4607,N_3916,N_2847);
and U4608 (N_4608,N_3964,N_2246);
nor U4609 (N_4609,N_3810,N_3902);
and U4610 (N_4610,N_2936,N_3580);
nand U4611 (N_4611,N_2813,N_3653);
xnor U4612 (N_4612,N_3212,N_2448);
xnor U4613 (N_4613,N_2652,N_2581);
and U4614 (N_4614,N_3630,N_3139);
and U4615 (N_4615,N_2601,N_2451);
nand U4616 (N_4616,N_2245,N_3716);
nand U4617 (N_4617,N_2481,N_2885);
nor U4618 (N_4618,N_3669,N_2064);
nand U4619 (N_4619,N_2052,N_3067);
nand U4620 (N_4620,N_3340,N_3415);
or U4621 (N_4621,N_2415,N_2037);
nand U4622 (N_4622,N_3624,N_2738);
xnor U4623 (N_4623,N_3593,N_3528);
nor U4624 (N_4624,N_2979,N_2644);
nand U4625 (N_4625,N_2990,N_3472);
nand U4626 (N_4626,N_2724,N_2895);
nor U4627 (N_4627,N_2960,N_2387);
or U4628 (N_4628,N_2515,N_3367);
or U4629 (N_4629,N_2732,N_3296);
or U4630 (N_4630,N_3826,N_3627);
or U4631 (N_4631,N_2365,N_3568);
xnor U4632 (N_4632,N_2439,N_2619);
and U4633 (N_4633,N_2054,N_2250);
xnor U4634 (N_4634,N_3549,N_3194);
and U4635 (N_4635,N_3095,N_3652);
nand U4636 (N_4636,N_2389,N_3728);
or U4637 (N_4637,N_2904,N_3471);
xnor U4638 (N_4638,N_3721,N_2056);
xnor U4639 (N_4639,N_2520,N_2794);
and U4640 (N_4640,N_2999,N_2122);
nand U4641 (N_4641,N_2939,N_3458);
and U4642 (N_4642,N_2168,N_3604);
or U4643 (N_4643,N_3130,N_2509);
nor U4644 (N_4644,N_2044,N_3263);
nand U4645 (N_4645,N_2550,N_3379);
or U4646 (N_4646,N_2826,N_3754);
or U4647 (N_4647,N_2114,N_3461);
nor U4648 (N_4648,N_2907,N_2366);
or U4649 (N_4649,N_2406,N_3720);
nor U4650 (N_4650,N_2549,N_2028);
xnor U4651 (N_4651,N_3789,N_2857);
nor U4652 (N_4652,N_3948,N_3601);
nor U4653 (N_4653,N_2227,N_2578);
nand U4654 (N_4654,N_3668,N_3943);
nor U4655 (N_4655,N_3648,N_2091);
nor U4656 (N_4656,N_2801,N_2874);
xor U4657 (N_4657,N_2100,N_3278);
xnor U4658 (N_4658,N_2319,N_3331);
and U4659 (N_4659,N_3466,N_2402);
nor U4660 (N_4660,N_2720,N_2604);
xor U4661 (N_4661,N_2206,N_2284);
and U4662 (N_4662,N_2071,N_3295);
or U4663 (N_4663,N_2239,N_2768);
and U4664 (N_4664,N_3854,N_3798);
nand U4665 (N_4665,N_2848,N_3047);
or U4666 (N_4666,N_3451,N_3124);
xor U4667 (N_4667,N_2538,N_2021);
nand U4668 (N_4668,N_3207,N_3836);
xnor U4669 (N_4669,N_3973,N_3577);
nand U4670 (N_4670,N_3306,N_2036);
and U4671 (N_4671,N_3756,N_2855);
xnor U4672 (N_4672,N_3181,N_2312);
and U4673 (N_4673,N_2108,N_3758);
or U4674 (N_4674,N_2483,N_3853);
or U4675 (N_4675,N_2141,N_3735);
nand U4676 (N_4676,N_3925,N_3341);
and U4677 (N_4677,N_3292,N_2288);
nor U4678 (N_4678,N_2803,N_2514);
nor U4679 (N_4679,N_2716,N_3397);
xor U4680 (N_4680,N_2384,N_2155);
or U4681 (N_4681,N_3699,N_2607);
nor U4682 (N_4682,N_3014,N_2090);
nand U4683 (N_4683,N_2685,N_3018);
xnor U4684 (N_4684,N_2599,N_2893);
nor U4685 (N_4685,N_3361,N_2902);
xnor U4686 (N_4686,N_2634,N_2752);
xor U4687 (N_4687,N_3380,N_3420);
nand U4688 (N_4688,N_3729,N_3885);
or U4689 (N_4689,N_2007,N_2161);
nand U4690 (N_4690,N_3311,N_3947);
and U4691 (N_4691,N_3832,N_2977);
nor U4692 (N_4692,N_2322,N_2992);
nand U4693 (N_4693,N_3818,N_3904);
nor U4694 (N_4694,N_3922,N_2381);
and U4695 (N_4695,N_3385,N_3814);
and U4696 (N_4696,N_3665,N_2078);
nand U4697 (N_4697,N_2810,N_3944);
and U4698 (N_4698,N_3553,N_3643);
nand U4699 (N_4699,N_2012,N_3589);
xnor U4700 (N_4700,N_2668,N_3167);
nor U4701 (N_4701,N_3268,N_2833);
or U4702 (N_4702,N_3419,N_2097);
or U4703 (N_4703,N_3612,N_3392);
xnor U4704 (N_4704,N_3347,N_2870);
nand U4705 (N_4705,N_3872,N_3498);
xor U4706 (N_4706,N_3242,N_2822);
xnor U4707 (N_4707,N_2638,N_2541);
xnor U4708 (N_4708,N_3434,N_3008);
nor U4709 (N_4709,N_2049,N_3731);
xor U4710 (N_4710,N_3500,N_3557);
and U4711 (N_4711,N_2831,N_3388);
nand U4712 (N_4712,N_3425,N_3930);
xor U4713 (N_4713,N_3424,N_2888);
or U4714 (N_4714,N_2002,N_3199);
xnor U4715 (N_4715,N_3550,N_3304);
nand U4716 (N_4716,N_3576,N_3772);
xor U4717 (N_4717,N_3286,N_3781);
xor U4718 (N_4718,N_3642,N_2700);
nor U4719 (N_4719,N_2539,N_3298);
nor U4720 (N_4720,N_2158,N_2942);
and U4721 (N_4721,N_3224,N_3418);
or U4722 (N_4722,N_2058,N_3320);
nand U4723 (N_4723,N_3289,N_3102);
nor U4724 (N_4724,N_2665,N_2586);
nor U4725 (N_4725,N_2116,N_3502);
nor U4726 (N_4726,N_2425,N_3680);
or U4727 (N_4727,N_3963,N_3707);
xnor U4728 (N_4728,N_2554,N_3955);
nand U4729 (N_4729,N_3575,N_3542);
nor U4730 (N_4730,N_2410,N_3895);
or U4731 (N_4731,N_3683,N_3364);
nand U4732 (N_4732,N_3877,N_3314);
nor U4733 (N_4733,N_3117,N_2046);
or U4734 (N_4734,N_3747,N_2845);
and U4735 (N_4735,N_2875,N_2262);
and U4736 (N_4736,N_2802,N_3806);
and U4737 (N_4737,N_3649,N_2692);
xor U4738 (N_4738,N_3714,N_2172);
and U4739 (N_4739,N_3590,N_3232);
nand U4740 (N_4740,N_2537,N_2982);
xnor U4741 (N_4741,N_3656,N_2376);
xnor U4742 (N_4742,N_3691,N_2688);
xor U4743 (N_4743,N_3280,N_2786);
nor U4744 (N_4744,N_3459,N_2104);
or U4745 (N_4745,N_3061,N_2267);
nand U4746 (N_4746,N_2767,N_2343);
nand U4747 (N_4747,N_3339,N_3631);
and U4748 (N_4748,N_3676,N_3843);
or U4749 (N_4749,N_3250,N_2513);
nor U4750 (N_4750,N_3470,N_2219);
and U4751 (N_4751,N_3238,N_3059);
and U4752 (N_4752,N_3543,N_2552);
nand U4753 (N_4753,N_2149,N_3370);
and U4754 (N_4754,N_2430,N_3393);
nand U4755 (N_4755,N_3090,N_3276);
and U4756 (N_4756,N_3460,N_2973);
xnor U4757 (N_4757,N_3594,N_3386);
xor U4758 (N_4758,N_3737,N_3581);
nor U4759 (N_4759,N_3517,N_2266);
and U4760 (N_4760,N_2871,N_3112);
nand U4761 (N_4761,N_2330,N_2407);
and U4762 (N_4762,N_3143,N_2323);
xor U4763 (N_4763,N_3485,N_2295);
or U4764 (N_4764,N_3428,N_3479);
xor U4765 (N_4765,N_2881,N_3724);
nor U4766 (N_4766,N_3931,N_2120);
and U4767 (N_4767,N_3852,N_3628);
and U4768 (N_4768,N_2388,N_2386);
nand U4769 (N_4769,N_3375,N_2484);
nor U4770 (N_4770,N_3359,N_3487);
nor U4771 (N_4771,N_3457,N_2617);
or U4772 (N_4772,N_2966,N_3617);
nand U4773 (N_4773,N_2164,N_2214);
nand U4774 (N_4774,N_3565,N_3966);
or U4775 (N_4775,N_3150,N_2887);
or U4776 (N_4776,N_2718,N_3574);
nand U4777 (N_4777,N_2359,N_2998);
nor U4778 (N_4778,N_3611,N_2542);
or U4779 (N_4779,N_3746,N_3071);
and U4780 (N_4780,N_3660,N_3144);
nand U4781 (N_4781,N_2289,N_2457);
xor U4782 (N_4782,N_2953,N_2628);
nand U4783 (N_4783,N_3142,N_2560);
nand U4784 (N_4784,N_2951,N_3234);
xor U4785 (N_4785,N_3100,N_3105);
nand U4786 (N_4786,N_2029,N_2707);
xnor U4787 (N_4787,N_3523,N_2785);
nand U4788 (N_4788,N_3812,N_2770);
xor U4789 (N_4789,N_2669,N_2862);
nor U4790 (N_4790,N_3740,N_2493);
nor U4791 (N_4791,N_3193,N_3730);
nor U4792 (N_4792,N_3073,N_2132);
xnor U4793 (N_4793,N_3698,N_3163);
xnor U4794 (N_4794,N_2010,N_3374);
or U4795 (N_4795,N_3626,N_3016);
nand U4796 (N_4796,N_3678,N_3389);
xor U4797 (N_4797,N_2019,N_2713);
and U4798 (N_4798,N_2850,N_3104);
xnor U4799 (N_4799,N_2081,N_3898);
or U4800 (N_4800,N_3165,N_2184);
and U4801 (N_4801,N_2072,N_2363);
or U4802 (N_4802,N_3997,N_3941);
nand U4803 (N_4803,N_3244,N_3788);
nor U4804 (N_4804,N_2589,N_2500);
xnor U4805 (N_4805,N_3417,N_3381);
nor U4806 (N_4806,N_3969,N_2216);
and U4807 (N_4807,N_2727,N_2580);
or U4808 (N_4808,N_2504,N_3602);
xnor U4809 (N_4809,N_2821,N_3327);
nor U4810 (N_4810,N_2420,N_3759);
nand U4811 (N_4811,N_3336,N_3448);
and U4812 (N_4812,N_3886,N_2383);
xnor U4813 (N_4813,N_3184,N_2409);
nand U4814 (N_4814,N_2569,N_2901);
nor U4815 (N_4815,N_2258,N_2188);
and U4816 (N_4816,N_3153,N_3053);
nand U4817 (N_4817,N_2478,N_3894);
and U4818 (N_4818,N_2105,N_3377);
nand U4819 (N_4819,N_3697,N_3222);
nand U4820 (N_4820,N_2985,N_2429);
or U4821 (N_4821,N_2016,N_3043);
nor U4822 (N_4822,N_3659,N_2378);
nand U4823 (N_4823,N_3255,N_2436);
xor U4824 (N_4824,N_2779,N_2447);
xnor U4825 (N_4825,N_3845,N_3427);
and U4826 (N_4826,N_2965,N_2445);
xor U4827 (N_4827,N_2934,N_3209);
nor U4828 (N_4828,N_2182,N_2675);
nor U4829 (N_4829,N_2843,N_2877);
nor U4830 (N_4830,N_2196,N_3803);
xnor U4831 (N_4831,N_2314,N_3616);
nor U4832 (N_4832,N_2730,N_2530);
nand U4833 (N_4833,N_3712,N_2923);
and U4834 (N_4834,N_3768,N_3822);
nor U4835 (N_4835,N_3857,N_3493);
xor U4836 (N_4836,N_3733,N_2198);
and U4837 (N_4837,N_2940,N_3345);
xor U4838 (N_4838,N_2070,N_2744);
and U4839 (N_4839,N_2636,N_3258);
nor U4840 (N_4840,N_3078,N_2805);
xor U4841 (N_4841,N_2624,N_2042);
or U4842 (N_4842,N_2567,N_3302);
nand U4843 (N_4843,N_3271,N_3344);
nand U4844 (N_4844,N_2099,N_2296);
xnor U4845 (N_4845,N_3233,N_3152);
nor U4846 (N_4846,N_3792,N_3587);
nand U4847 (N_4847,N_3006,N_3230);
nand U4848 (N_4848,N_3532,N_3935);
nor U4849 (N_4849,N_3636,N_2869);
xnor U4850 (N_4850,N_2593,N_2130);
or U4851 (N_4851,N_2192,N_3674);
nor U4852 (N_4852,N_2076,N_3066);
and U4853 (N_4853,N_3476,N_3989);
xnor U4854 (N_4854,N_3211,N_2749);
or U4855 (N_4855,N_3732,N_2584);
and U4856 (N_4856,N_3274,N_3177);
or U4857 (N_4857,N_2981,N_2157);
nor U4858 (N_4858,N_2905,N_3684);
and U4859 (N_4859,N_3151,N_2298);
and U4860 (N_4860,N_2310,N_2791);
nor U4861 (N_4861,N_2925,N_2760);
xnor U4862 (N_4862,N_2324,N_3352);
and U4863 (N_4863,N_2762,N_2432);
nor U4864 (N_4864,N_2462,N_3464);
nor U4865 (N_4865,N_3354,N_3625);
xor U4866 (N_4866,N_3326,N_2128);
nor U4867 (N_4867,N_2781,N_2135);
nor U4868 (N_4868,N_3584,N_3645);
nor U4869 (N_4869,N_3622,N_3075);
and U4870 (N_4870,N_3932,N_3985);
and U4871 (N_4871,N_2349,N_3125);
or U4872 (N_4872,N_2328,N_3155);
nor U4873 (N_4873,N_3583,N_2166);
xnor U4874 (N_4874,N_3858,N_2650);
nor U4875 (N_4875,N_2872,N_3901);
and U4876 (N_4876,N_3414,N_3281);
nor U4877 (N_4877,N_2503,N_3889);
xnor U4878 (N_4878,N_3407,N_3174);
and U4879 (N_4879,N_2889,N_3309);
xnor U4880 (N_4880,N_2620,N_3516);
xor U4881 (N_4881,N_3880,N_3109);
xnor U4882 (N_4882,N_2254,N_3154);
nor U4883 (N_4883,N_2761,N_3049);
nor U4884 (N_4884,N_2215,N_2495);
nor U4885 (N_4885,N_2218,N_3413);
nor U4886 (N_4886,N_3435,N_2622);
or U4887 (N_4887,N_3711,N_3961);
nand U4888 (N_4888,N_3767,N_2892);
xor U4889 (N_4889,N_2142,N_2544);
and U4890 (N_4890,N_3833,N_2463);
xor U4891 (N_4891,N_2026,N_3390);
xor U4892 (N_4892,N_2519,N_3132);
nand U4893 (N_4893,N_2914,N_3136);
nor U4894 (N_4894,N_2329,N_3065);
xnor U4895 (N_4895,N_2886,N_2948);
nand U4896 (N_4896,N_3519,N_2085);
nor U4897 (N_4897,N_3159,N_3548);
nand U4898 (N_4898,N_3279,N_2988);
and U4899 (N_4899,N_3256,N_3107);
nor U4900 (N_4900,N_2434,N_2858);
xor U4901 (N_4901,N_3615,N_3029);
nor U4902 (N_4902,N_2517,N_2423);
nand U4903 (N_4903,N_2931,N_3824);
xor U4904 (N_4904,N_2725,N_3958);
nor U4905 (N_4905,N_2980,N_2281);
nor U4906 (N_4906,N_3446,N_3180);
nand U4907 (N_4907,N_2824,N_3129);
or U4908 (N_4908,N_2774,N_2083);
or U4909 (N_4909,N_2374,N_2983);
nand U4910 (N_4910,N_2880,N_3795);
or U4911 (N_4911,N_2320,N_3779);
and U4912 (N_4912,N_2397,N_3921);
xnor U4913 (N_4913,N_3079,N_3508);
nand U4914 (N_4914,N_3578,N_3231);
nand U4915 (N_4915,N_2926,N_2853);
xor U4916 (N_4916,N_2024,N_2715);
and U4917 (N_4917,N_3216,N_3939);
and U4918 (N_4918,N_3774,N_3797);
xnor U4919 (N_4919,N_2793,N_3924);
xor U4920 (N_4920,N_3217,N_3496);
or U4921 (N_4921,N_3478,N_2025);
or U4922 (N_4922,N_2261,N_2396);
nor U4923 (N_4923,N_3329,N_2662);
xnor U4924 (N_4924,N_3501,N_3538);
and U4925 (N_4925,N_3866,N_2819);
and U4926 (N_4926,N_2989,N_3860);
xor U4927 (N_4927,N_2325,N_3790);
xor U4928 (N_4928,N_2570,N_3918);
or U4929 (N_4929,N_2313,N_3183);
and U4930 (N_4930,N_2414,N_3440);
and U4931 (N_4931,N_2670,N_3537);
and U4932 (N_4932,N_2424,N_2059);
xnor U4933 (N_4933,N_3808,N_3664);
nand U4934 (N_4934,N_2428,N_3009);
xnor U4935 (N_4935,N_2118,N_2244);
xnor U4936 (N_4936,N_3929,N_2551);
xor U4937 (N_4937,N_3572,N_3449);
and U4938 (N_4938,N_3085,N_2609);
nor U4939 (N_4939,N_2160,N_2151);
and U4940 (N_4940,N_3005,N_3382);
or U4941 (N_4941,N_3226,N_2204);
xor U4942 (N_4942,N_2474,N_2107);
nor U4943 (N_4943,N_2954,N_3267);
or U4944 (N_4944,N_3727,N_2632);
nor U4945 (N_4945,N_2226,N_3907);
nor U4946 (N_4946,N_2440,N_2812);
or U4947 (N_4947,N_3036,N_2331);
or U4948 (N_4948,N_3335,N_2908);
nand U4949 (N_4949,N_3223,N_3829);
and U4950 (N_4950,N_2921,N_2751);
or U4951 (N_4951,N_2268,N_2618);
and U4952 (N_4952,N_3771,N_2224);
and U4953 (N_4953,N_2991,N_3037);
xnor U4954 (N_4954,N_2112,N_3317);
xor U4955 (N_4955,N_2971,N_2398);
and U4956 (N_4956,N_2306,N_3202);
or U4957 (N_4957,N_2959,N_3351);
and U4958 (N_4958,N_2571,N_3198);
or U4959 (N_4959,N_3739,N_2416);
or U4960 (N_4960,N_2265,N_2178);
or U4961 (N_4961,N_2642,N_3492);
nand U4962 (N_4962,N_3992,N_3753);
or U4963 (N_4963,N_3849,N_3682);
xnor U4964 (N_4964,N_2913,N_2865);
nand U4965 (N_4965,N_3200,N_3473);
nand U4966 (N_4966,N_2595,N_2279);
or U4967 (N_4967,N_2958,N_3780);
nand U4968 (N_4968,N_3505,N_3976);
nor U4969 (N_4969,N_3432,N_2209);
or U4970 (N_4970,N_3204,N_2501);
or U4971 (N_4971,N_3290,N_2629);
nor U4972 (N_4972,N_3118,N_2305);
and U4973 (N_4973,N_2332,N_3288);
nand U4974 (N_4974,N_2694,N_3847);
xor U4975 (N_4975,N_3114,N_2234);
or U4976 (N_4976,N_3736,N_3620);
xnor U4977 (N_4977,N_2945,N_2605);
nand U4978 (N_4978,N_2033,N_2084);
nand U4979 (N_4979,N_3299,N_2352);
and U4980 (N_4980,N_3978,N_2089);
xor U4981 (N_4981,N_3956,N_2094);
xor U4982 (N_4982,N_2272,N_2950);
nand U4983 (N_4983,N_3131,N_3534);
or U4984 (N_4984,N_3444,N_2798);
nand U4985 (N_4985,N_2602,N_2576);
or U4986 (N_4986,N_2647,N_2792);
nor U4987 (N_4987,N_2648,N_2131);
or U4988 (N_4988,N_3239,N_2743);
nor U4989 (N_4989,N_3892,N_3228);
or U4990 (N_4990,N_2612,N_2403);
or U4991 (N_4991,N_2510,N_2521);
and U4992 (N_4992,N_3285,N_3804);
nand U4993 (N_4993,N_2144,N_2263);
or U4994 (N_4994,N_2941,N_3555);
xnor U4995 (N_4995,N_3300,N_2726);
or U4996 (N_4996,N_3926,N_3934);
xnor U4997 (N_4997,N_3993,N_2943);
or U4998 (N_4998,N_2704,N_2464);
nand U4999 (N_4999,N_2257,N_3115);
nand U5000 (N_5000,N_2954,N_3001);
nor U5001 (N_5001,N_3356,N_2118);
nand U5002 (N_5002,N_3719,N_3448);
nor U5003 (N_5003,N_2964,N_2711);
nor U5004 (N_5004,N_3392,N_3029);
nand U5005 (N_5005,N_3038,N_3133);
xor U5006 (N_5006,N_2408,N_3675);
nor U5007 (N_5007,N_3842,N_3830);
nor U5008 (N_5008,N_2525,N_2902);
nand U5009 (N_5009,N_3430,N_2283);
nor U5010 (N_5010,N_2500,N_2786);
nor U5011 (N_5011,N_3668,N_2343);
xnor U5012 (N_5012,N_2925,N_2911);
nor U5013 (N_5013,N_2198,N_3592);
nand U5014 (N_5014,N_2762,N_3332);
or U5015 (N_5015,N_2201,N_3755);
xor U5016 (N_5016,N_3662,N_3409);
xor U5017 (N_5017,N_2601,N_2084);
or U5018 (N_5018,N_2375,N_3839);
nor U5019 (N_5019,N_3445,N_3418);
and U5020 (N_5020,N_2999,N_3163);
nand U5021 (N_5021,N_3815,N_2542);
and U5022 (N_5022,N_3388,N_2530);
xnor U5023 (N_5023,N_2178,N_2116);
xor U5024 (N_5024,N_3566,N_3269);
and U5025 (N_5025,N_2453,N_3345);
or U5026 (N_5026,N_2324,N_2262);
or U5027 (N_5027,N_2478,N_2800);
and U5028 (N_5028,N_2147,N_3768);
and U5029 (N_5029,N_3548,N_3296);
nand U5030 (N_5030,N_3654,N_3481);
nor U5031 (N_5031,N_2095,N_2093);
nand U5032 (N_5032,N_3310,N_2958);
and U5033 (N_5033,N_3845,N_2858);
and U5034 (N_5034,N_2637,N_2493);
nor U5035 (N_5035,N_3592,N_3239);
xnor U5036 (N_5036,N_2385,N_2397);
or U5037 (N_5037,N_3435,N_2306);
nand U5038 (N_5038,N_2254,N_2305);
nor U5039 (N_5039,N_2263,N_3493);
or U5040 (N_5040,N_3307,N_2050);
nand U5041 (N_5041,N_3925,N_3060);
nor U5042 (N_5042,N_2896,N_3956);
and U5043 (N_5043,N_2604,N_2612);
nand U5044 (N_5044,N_2417,N_2592);
and U5045 (N_5045,N_2937,N_2610);
or U5046 (N_5046,N_2895,N_2328);
nor U5047 (N_5047,N_2160,N_2066);
nand U5048 (N_5048,N_2598,N_3621);
and U5049 (N_5049,N_3744,N_2154);
or U5050 (N_5050,N_3064,N_3045);
xnor U5051 (N_5051,N_3343,N_2396);
nand U5052 (N_5052,N_3701,N_2664);
or U5053 (N_5053,N_2990,N_3694);
nor U5054 (N_5054,N_3816,N_2638);
or U5055 (N_5055,N_3874,N_2519);
or U5056 (N_5056,N_2374,N_3662);
nand U5057 (N_5057,N_2308,N_3487);
nor U5058 (N_5058,N_2523,N_2187);
nor U5059 (N_5059,N_3425,N_2423);
xor U5060 (N_5060,N_3543,N_2273);
and U5061 (N_5061,N_3141,N_2120);
nand U5062 (N_5062,N_3308,N_3366);
nand U5063 (N_5063,N_2441,N_3363);
xor U5064 (N_5064,N_3086,N_3682);
and U5065 (N_5065,N_2334,N_3446);
xor U5066 (N_5066,N_2759,N_3939);
xnor U5067 (N_5067,N_2300,N_3471);
or U5068 (N_5068,N_2218,N_2269);
nand U5069 (N_5069,N_2170,N_3122);
xnor U5070 (N_5070,N_2867,N_2705);
xor U5071 (N_5071,N_3522,N_3494);
xnor U5072 (N_5072,N_2586,N_3748);
nand U5073 (N_5073,N_3897,N_2009);
xnor U5074 (N_5074,N_3783,N_2886);
xnor U5075 (N_5075,N_2991,N_3401);
or U5076 (N_5076,N_3703,N_3057);
nand U5077 (N_5077,N_3320,N_3670);
nor U5078 (N_5078,N_3637,N_2116);
nand U5079 (N_5079,N_2472,N_2091);
and U5080 (N_5080,N_2279,N_2678);
and U5081 (N_5081,N_3964,N_3954);
and U5082 (N_5082,N_3433,N_2725);
nor U5083 (N_5083,N_3216,N_3215);
xor U5084 (N_5084,N_3999,N_3825);
and U5085 (N_5085,N_2177,N_2690);
or U5086 (N_5086,N_3697,N_3207);
or U5087 (N_5087,N_3862,N_2943);
xor U5088 (N_5088,N_2155,N_3818);
nor U5089 (N_5089,N_3134,N_3452);
and U5090 (N_5090,N_3037,N_2795);
xor U5091 (N_5091,N_3246,N_3860);
or U5092 (N_5092,N_2229,N_3906);
xnor U5093 (N_5093,N_3315,N_3651);
xor U5094 (N_5094,N_2358,N_3486);
and U5095 (N_5095,N_3831,N_3867);
xnor U5096 (N_5096,N_2418,N_3843);
nor U5097 (N_5097,N_2229,N_2243);
nor U5098 (N_5098,N_2465,N_2653);
xnor U5099 (N_5099,N_3386,N_3866);
and U5100 (N_5100,N_3720,N_2866);
xnor U5101 (N_5101,N_3389,N_3029);
nor U5102 (N_5102,N_2016,N_2627);
nor U5103 (N_5103,N_3001,N_3163);
and U5104 (N_5104,N_3121,N_3393);
nor U5105 (N_5105,N_2515,N_2184);
or U5106 (N_5106,N_2153,N_3937);
nand U5107 (N_5107,N_3657,N_3076);
and U5108 (N_5108,N_3501,N_3719);
and U5109 (N_5109,N_2743,N_2697);
and U5110 (N_5110,N_3940,N_3827);
or U5111 (N_5111,N_3437,N_3032);
or U5112 (N_5112,N_3448,N_3378);
xor U5113 (N_5113,N_2652,N_2210);
xor U5114 (N_5114,N_3747,N_3998);
nand U5115 (N_5115,N_2718,N_2509);
and U5116 (N_5116,N_2092,N_3424);
or U5117 (N_5117,N_2954,N_2261);
xnor U5118 (N_5118,N_2280,N_2106);
and U5119 (N_5119,N_3260,N_2108);
nand U5120 (N_5120,N_3094,N_3146);
or U5121 (N_5121,N_3361,N_2012);
and U5122 (N_5122,N_2261,N_3851);
or U5123 (N_5123,N_3022,N_2533);
xor U5124 (N_5124,N_2420,N_3502);
xnor U5125 (N_5125,N_2773,N_3393);
and U5126 (N_5126,N_3260,N_2198);
nor U5127 (N_5127,N_2153,N_3271);
nor U5128 (N_5128,N_2709,N_3838);
nor U5129 (N_5129,N_3404,N_2589);
and U5130 (N_5130,N_2750,N_3536);
nor U5131 (N_5131,N_2485,N_2292);
xnor U5132 (N_5132,N_3132,N_2727);
and U5133 (N_5133,N_2671,N_2611);
and U5134 (N_5134,N_3382,N_2709);
nand U5135 (N_5135,N_2841,N_3126);
nand U5136 (N_5136,N_3285,N_2532);
and U5137 (N_5137,N_3458,N_2743);
xnor U5138 (N_5138,N_3621,N_2181);
or U5139 (N_5139,N_2879,N_2401);
or U5140 (N_5140,N_3435,N_2751);
and U5141 (N_5141,N_3754,N_3823);
or U5142 (N_5142,N_3513,N_2970);
and U5143 (N_5143,N_3828,N_2096);
or U5144 (N_5144,N_2269,N_2976);
or U5145 (N_5145,N_2583,N_3259);
nand U5146 (N_5146,N_3324,N_2411);
or U5147 (N_5147,N_3965,N_3697);
nand U5148 (N_5148,N_2175,N_2111);
or U5149 (N_5149,N_3338,N_3253);
or U5150 (N_5150,N_2418,N_2919);
xnor U5151 (N_5151,N_2057,N_2025);
or U5152 (N_5152,N_3661,N_2420);
and U5153 (N_5153,N_3500,N_3009);
and U5154 (N_5154,N_3190,N_3196);
or U5155 (N_5155,N_2894,N_2344);
and U5156 (N_5156,N_2878,N_2034);
xor U5157 (N_5157,N_3865,N_3346);
xor U5158 (N_5158,N_2274,N_2992);
or U5159 (N_5159,N_2769,N_3799);
xnor U5160 (N_5160,N_2356,N_2850);
nor U5161 (N_5161,N_3048,N_2586);
and U5162 (N_5162,N_2920,N_3527);
nand U5163 (N_5163,N_2688,N_2194);
nor U5164 (N_5164,N_3044,N_3106);
xor U5165 (N_5165,N_2003,N_3302);
nand U5166 (N_5166,N_2470,N_3612);
xnor U5167 (N_5167,N_2150,N_3660);
xnor U5168 (N_5168,N_3607,N_3049);
nand U5169 (N_5169,N_3277,N_2342);
or U5170 (N_5170,N_3037,N_3951);
nor U5171 (N_5171,N_3253,N_2839);
or U5172 (N_5172,N_3732,N_3710);
nor U5173 (N_5173,N_2783,N_2452);
and U5174 (N_5174,N_2789,N_2668);
or U5175 (N_5175,N_2859,N_3740);
nand U5176 (N_5176,N_2389,N_3589);
and U5177 (N_5177,N_2758,N_2727);
xnor U5178 (N_5178,N_3390,N_3553);
nor U5179 (N_5179,N_3556,N_2837);
and U5180 (N_5180,N_3686,N_3777);
or U5181 (N_5181,N_3660,N_3366);
xor U5182 (N_5182,N_2248,N_2695);
nor U5183 (N_5183,N_2054,N_3169);
xor U5184 (N_5184,N_2616,N_2814);
nand U5185 (N_5185,N_3571,N_2897);
nor U5186 (N_5186,N_2060,N_3274);
or U5187 (N_5187,N_2420,N_3006);
or U5188 (N_5188,N_3897,N_3382);
nand U5189 (N_5189,N_2428,N_3649);
nand U5190 (N_5190,N_3562,N_2742);
nor U5191 (N_5191,N_3195,N_2016);
nand U5192 (N_5192,N_2503,N_2917);
or U5193 (N_5193,N_2641,N_3020);
nand U5194 (N_5194,N_3647,N_3451);
nand U5195 (N_5195,N_3115,N_3698);
xnor U5196 (N_5196,N_3709,N_2034);
nand U5197 (N_5197,N_3573,N_2763);
nand U5198 (N_5198,N_2333,N_2898);
and U5199 (N_5199,N_3551,N_3043);
or U5200 (N_5200,N_3862,N_3647);
nor U5201 (N_5201,N_2664,N_2146);
or U5202 (N_5202,N_2542,N_3499);
or U5203 (N_5203,N_3158,N_2560);
xnor U5204 (N_5204,N_2900,N_3073);
nand U5205 (N_5205,N_3098,N_2726);
nand U5206 (N_5206,N_2147,N_2155);
or U5207 (N_5207,N_2629,N_3990);
nor U5208 (N_5208,N_2419,N_3106);
and U5209 (N_5209,N_3820,N_3340);
nor U5210 (N_5210,N_3974,N_3730);
nand U5211 (N_5211,N_2636,N_3917);
nand U5212 (N_5212,N_3146,N_3922);
and U5213 (N_5213,N_3711,N_2994);
nand U5214 (N_5214,N_3062,N_2548);
or U5215 (N_5215,N_2951,N_2737);
nor U5216 (N_5216,N_3577,N_2109);
nand U5217 (N_5217,N_3267,N_3569);
nor U5218 (N_5218,N_2756,N_3625);
and U5219 (N_5219,N_2748,N_2754);
nand U5220 (N_5220,N_2046,N_3743);
nor U5221 (N_5221,N_3360,N_3181);
and U5222 (N_5222,N_2922,N_2622);
nor U5223 (N_5223,N_2438,N_2914);
or U5224 (N_5224,N_2292,N_3063);
xnor U5225 (N_5225,N_3895,N_3281);
or U5226 (N_5226,N_3283,N_3836);
nand U5227 (N_5227,N_3883,N_2437);
or U5228 (N_5228,N_3558,N_2747);
nand U5229 (N_5229,N_3368,N_2675);
and U5230 (N_5230,N_3656,N_2065);
nand U5231 (N_5231,N_3875,N_2863);
nand U5232 (N_5232,N_3192,N_2199);
and U5233 (N_5233,N_3483,N_3385);
nor U5234 (N_5234,N_3769,N_2846);
and U5235 (N_5235,N_2919,N_3612);
nand U5236 (N_5236,N_2936,N_2002);
or U5237 (N_5237,N_3314,N_3550);
and U5238 (N_5238,N_2472,N_3376);
nor U5239 (N_5239,N_2617,N_3299);
nand U5240 (N_5240,N_3010,N_2630);
or U5241 (N_5241,N_2079,N_3805);
nor U5242 (N_5242,N_2426,N_2122);
nor U5243 (N_5243,N_2138,N_3133);
and U5244 (N_5244,N_2691,N_3942);
or U5245 (N_5245,N_3058,N_3966);
and U5246 (N_5246,N_2366,N_3801);
and U5247 (N_5247,N_3473,N_2995);
xor U5248 (N_5248,N_3080,N_3104);
nand U5249 (N_5249,N_3078,N_3295);
and U5250 (N_5250,N_3246,N_2330);
or U5251 (N_5251,N_3572,N_3483);
xor U5252 (N_5252,N_2887,N_3254);
or U5253 (N_5253,N_3763,N_3699);
or U5254 (N_5254,N_2899,N_3555);
xor U5255 (N_5255,N_2968,N_2984);
and U5256 (N_5256,N_3041,N_2743);
xor U5257 (N_5257,N_3860,N_3445);
nor U5258 (N_5258,N_3393,N_2447);
xor U5259 (N_5259,N_2771,N_2250);
and U5260 (N_5260,N_3478,N_3510);
xnor U5261 (N_5261,N_3504,N_2244);
nor U5262 (N_5262,N_3552,N_2847);
nand U5263 (N_5263,N_2564,N_3385);
and U5264 (N_5264,N_2265,N_3003);
or U5265 (N_5265,N_2266,N_3423);
nor U5266 (N_5266,N_3630,N_3414);
nor U5267 (N_5267,N_2506,N_3943);
and U5268 (N_5268,N_3949,N_2767);
and U5269 (N_5269,N_3069,N_3625);
xor U5270 (N_5270,N_3763,N_2181);
and U5271 (N_5271,N_2441,N_3381);
nor U5272 (N_5272,N_2886,N_3313);
nand U5273 (N_5273,N_2832,N_2966);
xnor U5274 (N_5274,N_2406,N_2271);
xor U5275 (N_5275,N_2696,N_2234);
and U5276 (N_5276,N_3616,N_3218);
and U5277 (N_5277,N_2614,N_2686);
nor U5278 (N_5278,N_2381,N_2220);
nor U5279 (N_5279,N_2434,N_3139);
or U5280 (N_5280,N_2248,N_3775);
nand U5281 (N_5281,N_2618,N_3989);
or U5282 (N_5282,N_3951,N_3076);
and U5283 (N_5283,N_2374,N_3229);
and U5284 (N_5284,N_3996,N_2118);
nor U5285 (N_5285,N_3187,N_2884);
or U5286 (N_5286,N_3465,N_3431);
nor U5287 (N_5287,N_3466,N_3952);
xnor U5288 (N_5288,N_2071,N_2594);
nor U5289 (N_5289,N_3149,N_2073);
nor U5290 (N_5290,N_2770,N_3714);
nor U5291 (N_5291,N_2014,N_2904);
and U5292 (N_5292,N_2149,N_3308);
and U5293 (N_5293,N_3030,N_3789);
xnor U5294 (N_5294,N_3849,N_3857);
xnor U5295 (N_5295,N_3261,N_2118);
or U5296 (N_5296,N_2775,N_2509);
xnor U5297 (N_5297,N_2623,N_3950);
and U5298 (N_5298,N_3394,N_3828);
nor U5299 (N_5299,N_3375,N_2653);
xor U5300 (N_5300,N_3485,N_3351);
nand U5301 (N_5301,N_3402,N_3028);
and U5302 (N_5302,N_2482,N_2878);
nor U5303 (N_5303,N_2413,N_3085);
nand U5304 (N_5304,N_2337,N_2302);
nor U5305 (N_5305,N_3451,N_3515);
and U5306 (N_5306,N_3485,N_2227);
nand U5307 (N_5307,N_2518,N_3947);
nor U5308 (N_5308,N_3120,N_3917);
nor U5309 (N_5309,N_2172,N_2449);
nand U5310 (N_5310,N_3811,N_3595);
nor U5311 (N_5311,N_3060,N_3246);
and U5312 (N_5312,N_2517,N_3893);
nand U5313 (N_5313,N_2053,N_2417);
xor U5314 (N_5314,N_2607,N_2180);
or U5315 (N_5315,N_2838,N_2280);
nor U5316 (N_5316,N_2768,N_3212);
and U5317 (N_5317,N_3938,N_3367);
or U5318 (N_5318,N_3142,N_2889);
nand U5319 (N_5319,N_2811,N_3214);
nor U5320 (N_5320,N_3421,N_3828);
xnor U5321 (N_5321,N_3657,N_2808);
and U5322 (N_5322,N_2028,N_3534);
and U5323 (N_5323,N_3781,N_2174);
and U5324 (N_5324,N_3562,N_3958);
nand U5325 (N_5325,N_2241,N_2951);
xnor U5326 (N_5326,N_3260,N_3687);
or U5327 (N_5327,N_3604,N_3187);
xor U5328 (N_5328,N_3436,N_3629);
nand U5329 (N_5329,N_3569,N_3819);
nand U5330 (N_5330,N_3231,N_2880);
nand U5331 (N_5331,N_2930,N_2795);
xor U5332 (N_5332,N_3591,N_3273);
nand U5333 (N_5333,N_3098,N_3967);
or U5334 (N_5334,N_2424,N_2154);
and U5335 (N_5335,N_3886,N_2267);
or U5336 (N_5336,N_2574,N_2149);
nor U5337 (N_5337,N_3425,N_2127);
nand U5338 (N_5338,N_3587,N_3647);
or U5339 (N_5339,N_3118,N_3495);
xnor U5340 (N_5340,N_2697,N_2479);
nand U5341 (N_5341,N_3564,N_2945);
nor U5342 (N_5342,N_3191,N_2211);
nor U5343 (N_5343,N_2732,N_2341);
xor U5344 (N_5344,N_2948,N_2063);
nor U5345 (N_5345,N_2678,N_3518);
and U5346 (N_5346,N_2062,N_2833);
nand U5347 (N_5347,N_3590,N_2637);
xnor U5348 (N_5348,N_3899,N_2188);
and U5349 (N_5349,N_2759,N_2596);
xnor U5350 (N_5350,N_2857,N_2889);
nand U5351 (N_5351,N_3648,N_3493);
nand U5352 (N_5352,N_3094,N_3997);
xor U5353 (N_5353,N_3128,N_3239);
xnor U5354 (N_5354,N_2878,N_3147);
or U5355 (N_5355,N_3160,N_3443);
and U5356 (N_5356,N_2664,N_3080);
xor U5357 (N_5357,N_2135,N_3589);
xnor U5358 (N_5358,N_2254,N_2623);
and U5359 (N_5359,N_2205,N_2677);
xor U5360 (N_5360,N_2562,N_3540);
xor U5361 (N_5361,N_2764,N_3685);
and U5362 (N_5362,N_2183,N_2663);
and U5363 (N_5363,N_2655,N_3154);
and U5364 (N_5364,N_2185,N_3457);
nor U5365 (N_5365,N_3212,N_2290);
xnor U5366 (N_5366,N_3472,N_3458);
nor U5367 (N_5367,N_3923,N_2363);
and U5368 (N_5368,N_2367,N_3639);
or U5369 (N_5369,N_3267,N_2070);
or U5370 (N_5370,N_3710,N_2221);
nand U5371 (N_5371,N_3232,N_3995);
nor U5372 (N_5372,N_3437,N_2856);
and U5373 (N_5373,N_2729,N_2356);
xor U5374 (N_5374,N_2774,N_2576);
nand U5375 (N_5375,N_2634,N_2067);
xnor U5376 (N_5376,N_3390,N_2580);
xnor U5377 (N_5377,N_2366,N_2690);
or U5378 (N_5378,N_3021,N_2867);
or U5379 (N_5379,N_2688,N_2877);
and U5380 (N_5380,N_3222,N_3811);
xor U5381 (N_5381,N_3461,N_3939);
and U5382 (N_5382,N_2870,N_3767);
and U5383 (N_5383,N_2984,N_2988);
nand U5384 (N_5384,N_3292,N_3013);
xor U5385 (N_5385,N_3660,N_3047);
xor U5386 (N_5386,N_3326,N_3510);
nand U5387 (N_5387,N_3104,N_3085);
or U5388 (N_5388,N_2804,N_3592);
nor U5389 (N_5389,N_3547,N_2153);
nor U5390 (N_5390,N_3102,N_3069);
nand U5391 (N_5391,N_2465,N_2244);
xnor U5392 (N_5392,N_3550,N_2037);
nor U5393 (N_5393,N_2148,N_3611);
or U5394 (N_5394,N_3925,N_3251);
and U5395 (N_5395,N_3278,N_3509);
xor U5396 (N_5396,N_3905,N_3058);
nand U5397 (N_5397,N_2923,N_3154);
nor U5398 (N_5398,N_3908,N_2577);
xor U5399 (N_5399,N_2079,N_2394);
nor U5400 (N_5400,N_3571,N_3570);
or U5401 (N_5401,N_2140,N_3496);
nand U5402 (N_5402,N_3691,N_3500);
xnor U5403 (N_5403,N_3223,N_3641);
and U5404 (N_5404,N_2292,N_2762);
and U5405 (N_5405,N_3409,N_2445);
and U5406 (N_5406,N_3930,N_2289);
nor U5407 (N_5407,N_3953,N_2225);
or U5408 (N_5408,N_2984,N_2431);
xor U5409 (N_5409,N_3103,N_2109);
and U5410 (N_5410,N_3542,N_2002);
and U5411 (N_5411,N_2544,N_3679);
nor U5412 (N_5412,N_2732,N_2991);
nor U5413 (N_5413,N_3305,N_2840);
or U5414 (N_5414,N_3889,N_3024);
and U5415 (N_5415,N_2590,N_2880);
xor U5416 (N_5416,N_2650,N_3365);
nor U5417 (N_5417,N_3834,N_2997);
xnor U5418 (N_5418,N_3436,N_3694);
and U5419 (N_5419,N_3634,N_2805);
and U5420 (N_5420,N_2478,N_2050);
and U5421 (N_5421,N_3599,N_2798);
nor U5422 (N_5422,N_3301,N_2046);
xnor U5423 (N_5423,N_3557,N_3525);
and U5424 (N_5424,N_2044,N_3255);
and U5425 (N_5425,N_2303,N_2389);
and U5426 (N_5426,N_2079,N_3057);
nor U5427 (N_5427,N_2523,N_3400);
xor U5428 (N_5428,N_2852,N_3490);
nor U5429 (N_5429,N_3002,N_2771);
nor U5430 (N_5430,N_3733,N_2350);
xnor U5431 (N_5431,N_2046,N_2258);
nor U5432 (N_5432,N_2423,N_3618);
nand U5433 (N_5433,N_3054,N_3865);
nor U5434 (N_5434,N_3519,N_2087);
nor U5435 (N_5435,N_3234,N_3698);
nand U5436 (N_5436,N_3317,N_3127);
nor U5437 (N_5437,N_3435,N_3459);
nand U5438 (N_5438,N_2122,N_3697);
nor U5439 (N_5439,N_3259,N_2315);
and U5440 (N_5440,N_2056,N_2108);
or U5441 (N_5441,N_2569,N_3368);
and U5442 (N_5442,N_3405,N_3675);
nand U5443 (N_5443,N_3550,N_3213);
or U5444 (N_5444,N_3257,N_2019);
or U5445 (N_5445,N_3098,N_3200);
xor U5446 (N_5446,N_3069,N_3071);
or U5447 (N_5447,N_3618,N_2349);
xor U5448 (N_5448,N_3656,N_3360);
or U5449 (N_5449,N_2420,N_2882);
or U5450 (N_5450,N_2723,N_2398);
xor U5451 (N_5451,N_2423,N_3121);
or U5452 (N_5452,N_2839,N_3704);
and U5453 (N_5453,N_3889,N_2725);
nand U5454 (N_5454,N_2558,N_3626);
or U5455 (N_5455,N_2778,N_2891);
xor U5456 (N_5456,N_2755,N_3121);
or U5457 (N_5457,N_3821,N_3565);
or U5458 (N_5458,N_2664,N_2749);
and U5459 (N_5459,N_2266,N_3553);
nand U5460 (N_5460,N_2718,N_2850);
or U5461 (N_5461,N_3049,N_2442);
nor U5462 (N_5462,N_3899,N_3719);
or U5463 (N_5463,N_3748,N_2930);
or U5464 (N_5464,N_3905,N_2351);
nor U5465 (N_5465,N_2697,N_2500);
and U5466 (N_5466,N_3556,N_3587);
nor U5467 (N_5467,N_3041,N_3900);
xnor U5468 (N_5468,N_3274,N_2961);
and U5469 (N_5469,N_3561,N_2401);
xor U5470 (N_5470,N_2787,N_3402);
or U5471 (N_5471,N_2120,N_2132);
nand U5472 (N_5472,N_2743,N_2606);
or U5473 (N_5473,N_3626,N_2013);
and U5474 (N_5474,N_3858,N_3090);
nand U5475 (N_5475,N_3799,N_2388);
or U5476 (N_5476,N_3649,N_2621);
nor U5477 (N_5477,N_3701,N_2212);
nor U5478 (N_5478,N_2428,N_3428);
xnor U5479 (N_5479,N_2093,N_2672);
nand U5480 (N_5480,N_3131,N_2917);
nand U5481 (N_5481,N_3759,N_3461);
nand U5482 (N_5482,N_2519,N_2720);
nor U5483 (N_5483,N_3620,N_2789);
and U5484 (N_5484,N_3990,N_2389);
xor U5485 (N_5485,N_2074,N_2277);
nand U5486 (N_5486,N_2793,N_3419);
xnor U5487 (N_5487,N_2938,N_2839);
or U5488 (N_5488,N_2562,N_2423);
xor U5489 (N_5489,N_2834,N_2811);
nor U5490 (N_5490,N_2537,N_2052);
and U5491 (N_5491,N_3270,N_2693);
and U5492 (N_5492,N_3204,N_2781);
nand U5493 (N_5493,N_2023,N_3056);
and U5494 (N_5494,N_3425,N_2017);
and U5495 (N_5495,N_2854,N_2308);
nor U5496 (N_5496,N_3283,N_2769);
or U5497 (N_5497,N_3342,N_2604);
and U5498 (N_5498,N_3168,N_2388);
or U5499 (N_5499,N_2492,N_2710);
or U5500 (N_5500,N_2634,N_2156);
nand U5501 (N_5501,N_2897,N_2665);
or U5502 (N_5502,N_2879,N_2750);
xnor U5503 (N_5503,N_3115,N_3081);
nand U5504 (N_5504,N_3247,N_2750);
and U5505 (N_5505,N_3637,N_2205);
nand U5506 (N_5506,N_3221,N_2305);
nor U5507 (N_5507,N_2651,N_2141);
nor U5508 (N_5508,N_2504,N_3676);
and U5509 (N_5509,N_2585,N_2078);
and U5510 (N_5510,N_3254,N_2029);
nor U5511 (N_5511,N_3037,N_3610);
or U5512 (N_5512,N_2615,N_3660);
and U5513 (N_5513,N_2929,N_3159);
xor U5514 (N_5514,N_2227,N_3065);
xor U5515 (N_5515,N_2484,N_2993);
nand U5516 (N_5516,N_3140,N_2112);
nor U5517 (N_5517,N_2398,N_3676);
xnor U5518 (N_5518,N_2610,N_3166);
nand U5519 (N_5519,N_2641,N_2484);
nand U5520 (N_5520,N_3576,N_2352);
or U5521 (N_5521,N_3931,N_3593);
and U5522 (N_5522,N_2856,N_3340);
nand U5523 (N_5523,N_3470,N_3716);
xor U5524 (N_5524,N_3428,N_2393);
or U5525 (N_5525,N_3509,N_3988);
or U5526 (N_5526,N_2921,N_2569);
or U5527 (N_5527,N_2880,N_2938);
nor U5528 (N_5528,N_3832,N_2875);
xor U5529 (N_5529,N_3952,N_3174);
or U5530 (N_5530,N_3154,N_3746);
or U5531 (N_5531,N_3529,N_2932);
or U5532 (N_5532,N_3884,N_3631);
nand U5533 (N_5533,N_3629,N_3382);
xnor U5534 (N_5534,N_2413,N_2275);
xor U5535 (N_5535,N_2585,N_2835);
nor U5536 (N_5536,N_2057,N_3938);
xor U5537 (N_5537,N_3560,N_3107);
nor U5538 (N_5538,N_3572,N_3593);
or U5539 (N_5539,N_2554,N_3239);
xnor U5540 (N_5540,N_2927,N_3901);
nand U5541 (N_5541,N_2821,N_2314);
nor U5542 (N_5542,N_2411,N_3037);
xnor U5543 (N_5543,N_3941,N_3090);
and U5544 (N_5544,N_2417,N_2015);
xor U5545 (N_5545,N_2217,N_3060);
or U5546 (N_5546,N_2870,N_3615);
nand U5547 (N_5547,N_2496,N_2664);
xnor U5548 (N_5548,N_3885,N_3954);
and U5549 (N_5549,N_2098,N_2575);
and U5550 (N_5550,N_2968,N_2541);
nor U5551 (N_5551,N_2532,N_2212);
xor U5552 (N_5552,N_2372,N_3959);
xor U5553 (N_5553,N_2868,N_3565);
xor U5554 (N_5554,N_2601,N_2826);
xor U5555 (N_5555,N_2836,N_3752);
nand U5556 (N_5556,N_2020,N_3791);
xnor U5557 (N_5557,N_2474,N_2458);
nor U5558 (N_5558,N_3310,N_2108);
or U5559 (N_5559,N_2059,N_2109);
and U5560 (N_5560,N_2841,N_3505);
nor U5561 (N_5561,N_3549,N_3405);
and U5562 (N_5562,N_3438,N_2580);
xor U5563 (N_5563,N_2890,N_2004);
and U5564 (N_5564,N_2284,N_3687);
nand U5565 (N_5565,N_3875,N_2277);
nand U5566 (N_5566,N_2364,N_3468);
and U5567 (N_5567,N_3512,N_3443);
nor U5568 (N_5568,N_2224,N_3226);
nor U5569 (N_5569,N_2522,N_3410);
nand U5570 (N_5570,N_2643,N_2727);
and U5571 (N_5571,N_3253,N_2130);
or U5572 (N_5572,N_3807,N_3594);
nor U5573 (N_5573,N_3196,N_3033);
or U5574 (N_5574,N_2913,N_3802);
and U5575 (N_5575,N_3128,N_2627);
or U5576 (N_5576,N_3153,N_2828);
or U5577 (N_5577,N_2452,N_2976);
nor U5578 (N_5578,N_3563,N_2357);
xnor U5579 (N_5579,N_3905,N_3628);
xor U5580 (N_5580,N_2307,N_2430);
and U5581 (N_5581,N_3003,N_3076);
and U5582 (N_5582,N_3530,N_2081);
xnor U5583 (N_5583,N_3072,N_2593);
nor U5584 (N_5584,N_2595,N_3668);
or U5585 (N_5585,N_2316,N_2429);
xnor U5586 (N_5586,N_2021,N_2413);
nand U5587 (N_5587,N_2531,N_2041);
nand U5588 (N_5588,N_2178,N_2248);
nor U5589 (N_5589,N_2034,N_3017);
nor U5590 (N_5590,N_2376,N_2940);
xnor U5591 (N_5591,N_3635,N_3728);
nand U5592 (N_5592,N_2119,N_2812);
and U5593 (N_5593,N_3270,N_3648);
or U5594 (N_5594,N_2162,N_3107);
nand U5595 (N_5595,N_2720,N_3894);
nand U5596 (N_5596,N_3667,N_2513);
xnor U5597 (N_5597,N_2849,N_3030);
or U5598 (N_5598,N_3991,N_3228);
and U5599 (N_5599,N_2617,N_3675);
nand U5600 (N_5600,N_2541,N_2745);
nor U5601 (N_5601,N_2837,N_2455);
or U5602 (N_5602,N_2892,N_2777);
nand U5603 (N_5603,N_3697,N_2314);
and U5604 (N_5604,N_3224,N_2026);
nor U5605 (N_5605,N_3896,N_2095);
nor U5606 (N_5606,N_3078,N_3622);
and U5607 (N_5607,N_2487,N_2871);
or U5608 (N_5608,N_2049,N_3740);
or U5609 (N_5609,N_3935,N_2327);
and U5610 (N_5610,N_3079,N_2645);
nand U5611 (N_5611,N_2321,N_2903);
xor U5612 (N_5612,N_3025,N_2898);
nor U5613 (N_5613,N_3831,N_3578);
or U5614 (N_5614,N_3021,N_2549);
xor U5615 (N_5615,N_2226,N_3689);
or U5616 (N_5616,N_3102,N_2579);
or U5617 (N_5617,N_3873,N_2857);
nor U5618 (N_5618,N_3001,N_3677);
nor U5619 (N_5619,N_2513,N_3136);
or U5620 (N_5620,N_2790,N_2558);
or U5621 (N_5621,N_2133,N_3075);
nand U5622 (N_5622,N_3762,N_3052);
and U5623 (N_5623,N_2819,N_2224);
xor U5624 (N_5624,N_2278,N_3612);
and U5625 (N_5625,N_2105,N_2098);
and U5626 (N_5626,N_3411,N_3715);
xnor U5627 (N_5627,N_2046,N_3943);
and U5628 (N_5628,N_3981,N_2804);
and U5629 (N_5629,N_2152,N_3521);
nand U5630 (N_5630,N_2433,N_3108);
or U5631 (N_5631,N_3441,N_3436);
nand U5632 (N_5632,N_2669,N_3248);
and U5633 (N_5633,N_2266,N_2480);
and U5634 (N_5634,N_3151,N_3560);
or U5635 (N_5635,N_3169,N_2286);
nor U5636 (N_5636,N_2645,N_3744);
xor U5637 (N_5637,N_2032,N_2683);
and U5638 (N_5638,N_3192,N_3341);
nand U5639 (N_5639,N_3711,N_3851);
or U5640 (N_5640,N_2868,N_3095);
or U5641 (N_5641,N_3757,N_2695);
or U5642 (N_5642,N_3593,N_2946);
or U5643 (N_5643,N_3948,N_2071);
xnor U5644 (N_5644,N_3960,N_2252);
nand U5645 (N_5645,N_3586,N_2427);
nand U5646 (N_5646,N_3435,N_2359);
xor U5647 (N_5647,N_3878,N_2843);
xnor U5648 (N_5648,N_2540,N_3538);
xnor U5649 (N_5649,N_3350,N_2793);
and U5650 (N_5650,N_2484,N_2076);
and U5651 (N_5651,N_2921,N_3008);
nor U5652 (N_5652,N_2287,N_3874);
or U5653 (N_5653,N_2106,N_3744);
or U5654 (N_5654,N_2409,N_2349);
and U5655 (N_5655,N_3279,N_2220);
xnor U5656 (N_5656,N_3551,N_3523);
and U5657 (N_5657,N_2004,N_2754);
nand U5658 (N_5658,N_3573,N_3029);
xor U5659 (N_5659,N_2858,N_2716);
or U5660 (N_5660,N_2038,N_3067);
or U5661 (N_5661,N_2456,N_2600);
nand U5662 (N_5662,N_3148,N_2643);
nor U5663 (N_5663,N_2595,N_2937);
xor U5664 (N_5664,N_3946,N_3905);
or U5665 (N_5665,N_3497,N_2204);
xor U5666 (N_5666,N_3287,N_3967);
nand U5667 (N_5667,N_2502,N_2151);
xnor U5668 (N_5668,N_3735,N_2597);
or U5669 (N_5669,N_2374,N_2717);
and U5670 (N_5670,N_3945,N_3044);
and U5671 (N_5671,N_2570,N_3242);
nor U5672 (N_5672,N_3257,N_3277);
and U5673 (N_5673,N_3909,N_2676);
nor U5674 (N_5674,N_3107,N_2223);
nand U5675 (N_5675,N_2508,N_3475);
nand U5676 (N_5676,N_2760,N_2709);
and U5677 (N_5677,N_2498,N_2975);
xnor U5678 (N_5678,N_2533,N_2738);
and U5679 (N_5679,N_3135,N_2301);
nor U5680 (N_5680,N_3595,N_2707);
nand U5681 (N_5681,N_2411,N_2082);
nand U5682 (N_5682,N_2716,N_3375);
or U5683 (N_5683,N_3972,N_3315);
nand U5684 (N_5684,N_2563,N_3968);
and U5685 (N_5685,N_3040,N_3310);
or U5686 (N_5686,N_3301,N_3046);
or U5687 (N_5687,N_3795,N_3238);
xor U5688 (N_5688,N_3846,N_2073);
or U5689 (N_5689,N_2501,N_2036);
xor U5690 (N_5690,N_3688,N_3800);
xor U5691 (N_5691,N_2679,N_2878);
xor U5692 (N_5692,N_2496,N_3296);
nand U5693 (N_5693,N_2255,N_2331);
or U5694 (N_5694,N_3064,N_2000);
and U5695 (N_5695,N_3008,N_3099);
and U5696 (N_5696,N_2410,N_2854);
nand U5697 (N_5697,N_3076,N_2593);
and U5698 (N_5698,N_2511,N_3100);
nand U5699 (N_5699,N_3842,N_3281);
and U5700 (N_5700,N_2736,N_2182);
nand U5701 (N_5701,N_3349,N_2972);
nand U5702 (N_5702,N_2660,N_3203);
nor U5703 (N_5703,N_3913,N_3325);
nor U5704 (N_5704,N_3104,N_2664);
and U5705 (N_5705,N_3861,N_2005);
xnor U5706 (N_5706,N_2492,N_3485);
and U5707 (N_5707,N_2674,N_2205);
xor U5708 (N_5708,N_2951,N_2972);
nor U5709 (N_5709,N_2397,N_3527);
nor U5710 (N_5710,N_2446,N_2220);
and U5711 (N_5711,N_3996,N_3881);
nand U5712 (N_5712,N_2699,N_2320);
or U5713 (N_5713,N_3009,N_2758);
and U5714 (N_5714,N_2425,N_2171);
or U5715 (N_5715,N_3245,N_2275);
xnor U5716 (N_5716,N_3447,N_2364);
nor U5717 (N_5717,N_2653,N_2902);
xnor U5718 (N_5718,N_2381,N_3635);
or U5719 (N_5719,N_3326,N_3673);
and U5720 (N_5720,N_3197,N_2151);
nor U5721 (N_5721,N_3980,N_3867);
nor U5722 (N_5722,N_3470,N_2596);
xor U5723 (N_5723,N_3586,N_2945);
xor U5724 (N_5724,N_3088,N_3387);
xor U5725 (N_5725,N_3086,N_2017);
nor U5726 (N_5726,N_2326,N_3035);
xor U5727 (N_5727,N_2579,N_2135);
or U5728 (N_5728,N_3176,N_3414);
and U5729 (N_5729,N_3748,N_2891);
nand U5730 (N_5730,N_3410,N_3901);
nand U5731 (N_5731,N_3413,N_3934);
nor U5732 (N_5732,N_3136,N_2705);
xor U5733 (N_5733,N_2497,N_2511);
and U5734 (N_5734,N_3327,N_3264);
xnor U5735 (N_5735,N_3772,N_3231);
and U5736 (N_5736,N_2223,N_2795);
nand U5737 (N_5737,N_2570,N_2760);
nor U5738 (N_5738,N_3590,N_2117);
nand U5739 (N_5739,N_2702,N_2758);
nor U5740 (N_5740,N_3002,N_2400);
and U5741 (N_5741,N_3487,N_3263);
nand U5742 (N_5742,N_3789,N_2186);
and U5743 (N_5743,N_3159,N_3204);
or U5744 (N_5744,N_3684,N_3329);
and U5745 (N_5745,N_3226,N_2501);
or U5746 (N_5746,N_3259,N_2050);
nand U5747 (N_5747,N_3334,N_2385);
nand U5748 (N_5748,N_3527,N_3961);
and U5749 (N_5749,N_3837,N_2405);
or U5750 (N_5750,N_3836,N_2247);
nor U5751 (N_5751,N_3429,N_3227);
and U5752 (N_5752,N_2154,N_3063);
nand U5753 (N_5753,N_3007,N_2685);
nand U5754 (N_5754,N_2854,N_2251);
nand U5755 (N_5755,N_2815,N_3361);
and U5756 (N_5756,N_2820,N_3319);
xor U5757 (N_5757,N_2650,N_3498);
xor U5758 (N_5758,N_3679,N_3749);
nand U5759 (N_5759,N_3444,N_2687);
nand U5760 (N_5760,N_2155,N_3633);
xor U5761 (N_5761,N_3154,N_3247);
and U5762 (N_5762,N_2327,N_3834);
nand U5763 (N_5763,N_2324,N_2293);
nor U5764 (N_5764,N_3015,N_3550);
nor U5765 (N_5765,N_3340,N_3879);
nand U5766 (N_5766,N_3681,N_2554);
or U5767 (N_5767,N_3126,N_3542);
and U5768 (N_5768,N_2097,N_3505);
and U5769 (N_5769,N_2841,N_3496);
nor U5770 (N_5770,N_2291,N_3965);
and U5771 (N_5771,N_2953,N_2733);
and U5772 (N_5772,N_3860,N_3194);
nor U5773 (N_5773,N_2745,N_2635);
and U5774 (N_5774,N_2801,N_2909);
xor U5775 (N_5775,N_3937,N_3119);
and U5776 (N_5776,N_3120,N_3375);
and U5777 (N_5777,N_2306,N_3399);
xnor U5778 (N_5778,N_2239,N_3693);
or U5779 (N_5779,N_3758,N_2592);
or U5780 (N_5780,N_2067,N_2313);
nor U5781 (N_5781,N_2324,N_2463);
and U5782 (N_5782,N_2827,N_2217);
nand U5783 (N_5783,N_2011,N_3189);
nand U5784 (N_5784,N_2887,N_2466);
nand U5785 (N_5785,N_3592,N_3504);
nor U5786 (N_5786,N_3972,N_2195);
and U5787 (N_5787,N_2574,N_2366);
nand U5788 (N_5788,N_3153,N_2930);
nor U5789 (N_5789,N_2352,N_3569);
nor U5790 (N_5790,N_3603,N_3818);
or U5791 (N_5791,N_3573,N_3931);
nand U5792 (N_5792,N_2657,N_3266);
xnor U5793 (N_5793,N_3290,N_3729);
xnor U5794 (N_5794,N_3009,N_3168);
nand U5795 (N_5795,N_3116,N_3499);
nand U5796 (N_5796,N_2588,N_3481);
and U5797 (N_5797,N_2208,N_2844);
or U5798 (N_5798,N_3998,N_3613);
nor U5799 (N_5799,N_2256,N_2566);
nand U5800 (N_5800,N_2631,N_3939);
xor U5801 (N_5801,N_2273,N_3046);
nor U5802 (N_5802,N_3692,N_3286);
nor U5803 (N_5803,N_3074,N_3971);
nor U5804 (N_5804,N_3291,N_3151);
nand U5805 (N_5805,N_3676,N_3768);
and U5806 (N_5806,N_2188,N_2401);
or U5807 (N_5807,N_3716,N_2806);
nor U5808 (N_5808,N_3362,N_3101);
xor U5809 (N_5809,N_2379,N_3646);
xor U5810 (N_5810,N_3100,N_2453);
xor U5811 (N_5811,N_3214,N_2091);
nor U5812 (N_5812,N_3513,N_3974);
nor U5813 (N_5813,N_3352,N_2506);
nor U5814 (N_5814,N_3622,N_3947);
and U5815 (N_5815,N_3193,N_3003);
or U5816 (N_5816,N_3028,N_2689);
nor U5817 (N_5817,N_3258,N_3668);
xor U5818 (N_5818,N_3044,N_3561);
xnor U5819 (N_5819,N_2973,N_3751);
nand U5820 (N_5820,N_3857,N_3606);
and U5821 (N_5821,N_3015,N_3242);
xnor U5822 (N_5822,N_3037,N_3308);
nor U5823 (N_5823,N_3607,N_3179);
and U5824 (N_5824,N_3222,N_2467);
and U5825 (N_5825,N_2231,N_3934);
xnor U5826 (N_5826,N_2992,N_3394);
and U5827 (N_5827,N_2874,N_2036);
nor U5828 (N_5828,N_2701,N_3171);
xnor U5829 (N_5829,N_3876,N_2177);
nand U5830 (N_5830,N_3841,N_2023);
nor U5831 (N_5831,N_3917,N_3540);
or U5832 (N_5832,N_2763,N_2573);
nor U5833 (N_5833,N_2288,N_2887);
and U5834 (N_5834,N_3361,N_2422);
and U5835 (N_5835,N_2464,N_2319);
and U5836 (N_5836,N_2865,N_2130);
nor U5837 (N_5837,N_2295,N_2221);
or U5838 (N_5838,N_3190,N_2551);
nor U5839 (N_5839,N_2653,N_2347);
nand U5840 (N_5840,N_2690,N_2261);
and U5841 (N_5841,N_2134,N_3697);
xnor U5842 (N_5842,N_3617,N_2284);
and U5843 (N_5843,N_2986,N_2190);
nand U5844 (N_5844,N_3334,N_3328);
nand U5845 (N_5845,N_3257,N_3653);
xor U5846 (N_5846,N_2389,N_2627);
nand U5847 (N_5847,N_3258,N_3889);
and U5848 (N_5848,N_3455,N_2562);
and U5849 (N_5849,N_2541,N_3653);
nor U5850 (N_5850,N_3235,N_3877);
nand U5851 (N_5851,N_2403,N_2483);
or U5852 (N_5852,N_3693,N_3170);
nand U5853 (N_5853,N_3926,N_3852);
xnor U5854 (N_5854,N_3930,N_2825);
nand U5855 (N_5855,N_3523,N_2783);
or U5856 (N_5856,N_3730,N_2180);
nor U5857 (N_5857,N_2269,N_2112);
nor U5858 (N_5858,N_2391,N_2821);
nor U5859 (N_5859,N_3450,N_3885);
and U5860 (N_5860,N_2686,N_3727);
or U5861 (N_5861,N_2352,N_2506);
nor U5862 (N_5862,N_2244,N_2995);
nor U5863 (N_5863,N_2845,N_2348);
xor U5864 (N_5864,N_2370,N_3124);
nand U5865 (N_5865,N_3921,N_3511);
and U5866 (N_5866,N_3610,N_2080);
and U5867 (N_5867,N_3134,N_2002);
or U5868 (N_5868,N_2312,N_2636);
and U5869 (N_5869,N_3658,N_2699);
nand U5870 (N_5870,N_2137,N_2576);
xor U5871 (N_5871,N_3575,N_2560);
and U5872 (N_5872,N_3203,N_2001);
nand U5873 (N_5873,N_3299,N_3384);
or U5874 (N_5874,N_2506,N_2478);
nor U5875 (N_5875,N_3525,N_2313);
nand U5876 (N_5876,N_2900,N_3146);
xor U5877 (N_5877,N_3065,N_2742);
or U5878 (N_5878,N_3320,N_3098);
or U5879 (N_5879,N_3656,N_3685);
xor U5880 (N_5880,N_2722,N_3136);
and U5881 (N_5881,N_2323,N_2024);
nor U5882 (N_5882,N_2784,N_3363);
and U5883 (N_5883,N_2762,N_3484);
and U5884 (N_5884,N_2087,N_2422);
nand U5885 (N_5885,N_2176,N_3173);
xnor U5886 (N_5886,N_3434,N_2275);
nor U5887 (N_5887,N_2158,N_2511);
or U5888 (N_5888,N_3195,N_2476);
nand U5889 (N_5889,N_3127,N_3251);
and U5890 (N_5890,N_3845,N_3501);
or U5891 (N_5891,N_3958,N_2142);
xnor U5892 (N_5892,N_3769,N_2703);
or U5893 (N_5893,N_2538,N_2272);
or U5894 (N_5894,N_3278,N_2825);
xor U5895 (N_5895,N_3459,N_2504);
xor U5896 (N_5896,N_2325,N_3233);
and U5897 (N_5897,N_2822,N_2986);
and U5898 (N_5898,N_3534,N_3875);
xor U5899 (N_5899,N_3197,N_2101);
nor U5900 (N_5900,N_3032,N_2823);
nor U5901 (N_5901,N_2171,N_3062);
nand U5902 (N_5902,N_3074,N_2929);
xnor U5903 (N_5903,N_3141,N_3270);
xor U5904 (N_5904,N_2515,N_2246);
nor U5905 (N_5905,N_2151,N_2096);
nor U5906 (N_5906,N_3678,N_2186);
nand U5907 (N_5907,N_2360,N_2340);
xor U5908 (N_5908,N_3971,N_3635);
nor U5909 (N_5909,N_2144,N_2352);
and U5910 (N_5910,N_2601,N_3336);
nor U5911 (N_5911,N_2894,N_2335);
nand U5912 (N_5912,N_3898,N_2722);
nor U5913 (N_5913,N_3962,N_3882);
nand U5914 (N_5914,N_3485,N_2661);
nor U5915 (N_5915,N_2847,N_3868);
nand U5916 (N_5916,N_2801,N_2084);
nor U5917 (N_5917,N_2961,N_3584);
xor U5918 (N_5918,N_3248,N_3386);
xor U5919 (N_5919,N_2880,N_2249);
and U5920 (N_5920,N_2923,N_3459);
nor U5921 (N_5921,N_3418,N_3102);
nand U5922 (N_5922,N_2477,N_2184);
or U5923 (N_5923,N_2629,N_2226);
nand U5924 (N_5924,N_2289,N_2646);
nor U5925 (N_5925,N_2251,N_3345);
nor U5926 (N_5926,N_2197,N_3766);
and U5927 (N_5927,N_3742,N_3053);
or U5928 (N_5928,N_3193,N_2370);
nand U5929 (N_5929,N_2367,N_3819);
and U5930 (N_5930,N_3932,N_2644);
and U5931 (N_5931,N_3418,N_2233);
nor U5932 (N_5932,N_2039,N_3892);
and U5933 (N_5933,N_2380,N_3050);
or U5934 (N_5934,N_3297,N_3790);
xor U5935 (N_5935,N_3386,N_2661);
or U5936 (N_5936,N_3242,N_2588);
nand U5937 (N_5937,N_2594,N_2245);
xor U5938 (N_5938,N_2534,N_2630);
nor U5939 (N_5939,N_3678,N_2345);
xor U5940 (N_5940,N_3706,N_3966);
and U5941 (N_5941,N_2549,N_2310);
or U5942 (N_5942,N_2416,N_3053);
xor U5943 (N_5943,N_3921,N_2403);
nand U5944 (N_5944,N_3871,N_2353);
xor U5945 (N_5945,N_2083,N_2457);
or U5946 (N_5946,N_2649,N_2459);
and U5947 (N_5947,N_2175,N_3209);
nand U5948 (N_5948,N_3929,N_2811);
xnor U5949 (N_5949,N_3190,N_2211);
or U5950 (N_5950,N_2662,N_2680);
and U5951 (N_5951,N_2176,N_2270);
nand U5952 (N_5952,N_3451,N_3690);
nor U5953 (N_5953,N_3129,N_2135);
xnor U5954 (N_5954,N_2924,N_2539);
nand U5955 (N_5955,N_2429,N_2742);
xor U5956 (N_5956,N_3247,N_3219);
and U5957 (N_5957,N_3708,N_3342);
nand U5958 (N_5958,N_3565,N_3726);
nor U5959 (N_5959,N_2127,N_2790);
nand U5960 (N_5960,N_3684,N_2437);
or U5961 (N_5961,N_2729,N_2280);
nor U5962 (N_5962,N_3030,N_3924);
or U5963 (N_5963,N_2366,N_3894);
nor U5964 (N_5964,N_3011,N_2019);
nand U5965 (N_5965,N_2172,N_3691);
and U5966 (N_5966,N_2352,N_3698);
and U5967 (N_5967,N_3386,N_3276);
nor U5968 (N_5968,N_2487,N_2941);
or U5969 (N_5969,N_3039,N_3508);
and U5970 (N_5970,N_3673,N_3710);
and U5971 (N_5971,N_3351,N_3563);
nor U5972 (N_5972,N_3075,N_3561);
or U5973 (N_5973,N_2888,N_3055);
and U5974 (N_5974,N_2101,N_3202);
nand U5975 (N_5975,N_3002,N_3731);
or U5976 (N_5976,N_3604,N_3184);
nand U5977 (N_5977,N_3601,N_2106);
xor U5978 (N_5978,N_2971,N_2661);
xnor U5979 (N_5979,N_3821,N_3624);
or U5980 (N_5980,N_3229,N_3170);
and U5981 (N_5981,N_3285,N_3130);
or U5982 (N_5982,N_3827,N_2938);
or U5983 (N_5983,N_3651,N_3370);
and U5984 (N_5984,N_2795,N_2286);
xnor U5985 (N_5985,N_2150,N_3067);
or U5986 (N_5986,N_2415,N_2184);
nor U5987 (N_5987,N_2179,N_3848);
xnor U5988 (N_5988,N_2688,N_3804);
xor U5989 (N_5989,N_2457,N_2568);
or U5990 (N_5990,N_3955,N_2220);
nor U5991 (N_5991,N_3239,N_2254);
or U5992 (N_5992,N_2986,N_2205);
and U5993 (N_5993,N_2386,N_2926);
xnor U5994 (N_5994,N_2154,N_2851);
nor U5995 (N_5995,N_2337,N_3229);
nor U5996 (N_5996,N_3794,N_2512);
and U5997 (N_5997,N_2380,N_3250);
nand U5998 (N_5998,N_3935,N_3895);
or U5999 (N_5999,N_2509,N_3874);
nand U6000 (N_6000,N_4799,N_4738);
xnor U6001 (N_6001,N_4004,N_5158);
nor U6002 (N_6002,N_5223,N_4448);
nand U6003 (N_6003,N_5848,N_5486);
nand U6004 (N_6004,N_4119,N_4968);
and U6005 (N_6005,N_5658,N_5881);
and U6006 (N_6006,N_4519,N_5795);
and U6007 (N_6007,N_4274,N_4449);
xor U6008 (N_6008,N_5650,N_4992);
or U6009 (N_6009,N_4813,N_4275);
and U6010 (N_6010,N_5363,N_5275);
xnor U6011 (N_6011,N_5443,N_4722);
nor U6012 (N_6012,N_4701,N_4697);
xor U6013 (N_6013,N_4835,N_4467);
xor U6014 (N_6014,N_5273,N_4524);
xor U6015 (N_6015,N_4852,N_5195);
xnor U6016 (N_6016,N_4312,N_5062);
and U6017 (N_6017,N_4198,N_4262);
nand U6018 (N_6018,N_5709,N_5822);
nand U6019 (N_6019,N_5430,N_4452);
and U6020 (N_6020,N_4908,N_4193);
xnor U6021 (N_6021,N_5447,N_5362);
nor U6022 (N_6022,N_4313,N_5396);
xnor U6023 (N_6023,N_5990,N_5775);
or U6024 (N_6024,N_5526,N_4610);
xnor U6025 (N_6025,N_4357,N_5873);
nand U6026 (N_6026,N_4389,N_4911);
or U6027 (N_6027,N_4522,N_5786);
nand U6028 (N_6028,N_5064,N_4732);
xnor U6029 (N_6029,N_5318,N_5514);
and U6030 (N_6030,N_5225,N_4696);
nand U6031 (N_6031,N_5520,N_4816);
nor U6032 (N_6032,N_4535,N_5259);
and U6033 (N_6033,N_5431,N_5993);
nand U6034 (N_6034,N_5006,N_4571);
nand U6035 (N_6035,N_5596,N_4343);
xor U6036 (N_6036,N_5071,N_5503);
xnor U6037 (N_6037,N_4954,N_4322);
or U6038 (N_6038,N_4867,N_5513);
or U6039 (N_6039,N_5459,N_4241);
nor U6040 (N_6040,N_4095,N_4488);
xor U6041 (N_6041,N_5785,N_4367);
nand U6042 (N_6042,N_5246,N_5367);
and U6043 (N_6043,N_4024,N_5221);
or U6044 (N_6044,N_4286,N_4092);
nand U6045 (N_6045,N_4960,N_5497);
nor U6046 (N_6046,N_5945,N_4784);
and U6047 (N_6047,N_5949,N_5585);
nand U6048 (N_6048,N_5402,N_5304);
nor U6049 (N_6049,N_4144,N_4397);
xnor U6050 (N_6050,N_4675,N_5380);
nor U6051 (N_6051,N_4721,N_4113);
or U6052 (N_6052,N_4555,N_5673);
nor U6053 (N_6053,N_5537,N_5583);
nand U6054 (N_6054,N_4366,N_5724);
xor U6055 (N_6055,N_4001,N_4189);
nand U6056 (N_6056,N_4962,N_5688);
nand U6057 (N_6057,N_4026,N_5791);
nand U6058 (N_6058,N_5052,N_5611);
and U6059 (N_6059,N_4007,N_4282);
nand U6060 (N_6060,N_5959,N_4763);
nand U6061 (N_6061,N_4231,N_4705);
nand U6062 (N_6062,N_5025,N_5900);
nand U6063 (N_6063,N_5712,N_5297);
xnor U6064 (N_6064,N_5435,N_4768);
nor U6065 (N_6065,N_4063,N_4009);
nand U6066 (N_6066,N_5908,N_5125);
xor U6067 (N_6067,N_5080,N_5828);
and U6068 (N_6068,N_5613,N_4444);
nor U6069 (N_6069,N_4377,N_4743);
and U6070 (N_6070,N_4091,N_4659);
or U6071 (N_6071,N_4183,N_4082);
or U6072 (N_6072,N_5935,N_5999);
xnor U6073 (N_6073,N_5130,N_5150);
xnor U6074 (N_6074,N_5948,N_5352);
nand U6075 (N_6075,N_5835,N_5399);
nor U6076 (N_6076,N_5189,N_4994);
nand U6077 (N_6077,N_4808,N_5970);
and U6078 (N_6078,N_5457,N_5824);
nand U6079 (N_6079,N_5143,N_4711);
or U6080 (N_6080,N_5111,N_4577);
or U6081 (N_6081,N_5651,N_4351);
nor U6082 (N_6082,N_4409,N_4761);
and U6083 (N_6083,N_4718,N_4551);
and U6084 (N_6084,N_5663,N_5621);
or U6085 (N_6085,N_4131,N_4170);
xor U6086 (N_6086,N_5722,N_5748);
nor U6087 (N_6087,N_4773,N_5705);
and U6088 (N_6088,N_4319,N_5743);
nor U6089 (N_6089,N_5851,N_5810);
and U6090 (N_6090,N_4174,N_4217);
or U6091 (N_6091,N_5700,N_4036);
or U6092 (N_6092,N_4056,N_4990);
or U6093 (N_6093,N_4010,N_5799);
nor U6094 (N_6094,N_5423,N_4491);
or U6095 (N_6095,N_4267,N_5206);
nand U6096 (N_6096,N_4611,N_4388);
nand U6097 (N_6097,N_4450,N_5733);
xnor U6098 (N_6098,N_4942,N_5161);
and U6099 (N_6099,N_4515,N_4633);
and U6100 (N_6100,N_4729,N_5030);
nor U6101 (N_6101,N_5445,N_5233);
xor U6102 (N_6102,N_5355,N_5026);
and U6103 (N_6103,N_4583,N_4569);
nand U6104 (N_6104,N_4544,N_5617);
nand U6105 (N_6105,N_5668,N_4049);
and U6106 (N_6106,N_4014,N_5293);
and U6107 (N_6107,N_5797,N_4489);
and U6108 (N_6108,N_5226,N_4106);
xor U6109 (N_6109,N_4127,N_4023);
nand U6110 (N_6110,N_4074,N_4061);
nor U6111 (N_6111,N_5863,N_5042);
nand U6112 (N_6112,N_5112,N_4907);
and U6113 (N_6113,N_5922,N_4318);
or U6114 (N_6114,N_4655,N_4900);
xnor U6115 (N_6115,N_4406,N_4054);
nand U6116 (N_6116,N_5814,N_4477);
xnor U6117 (N_6117,N_5910,N_4547);
and U6118 (N_6118,N_5315,N_5886);
nor U6119 (N_6119,N_4600,N_5008);
nor U6120 (N_6120,N_5333,N_4593);
nand U6121 (N_6121,N_5172,N_5971);
or U6122 (N_6122,N_4109,N_5731);
xnor U6123 (N_6123,N_4956,N_5119);
or U6124 (N_6124,N_5204,N_5427);
and U6125 (N_6125,N_4093,N_5888);
nor U6126 (N_6126,N_5449,N_4629);
nor U6127 (N_6127,N_5612,N_5793);
xor U6128 (N_6128,N_4775,N_5710);
xor U6129 (N_6129,N_4788,N_4324);
nand U6130 (N_6130,N_5882,N_5539);
nor U6131 (N_6131,N_5313,N_5483);
nor U6132 (N_6132,N_5110,N_4381);
or U6133 (N_6133,N_5385,N_5693);
or U6134 (N_6134,N_5269,N_4211);
nand U6135 (N_6135,N_4264,N_5361);
nor U6136 (N_6136,N_4430,N_4462);
xor U6137 (N_6137,N_5105,N_5992);
nor U6138 (N_6138,N_4358,N_5856);
and U6139 (N_6139,N_4133,N_4046);
nand U6140 (N_6140,N_5813,N_4589);
xnor U6141 (N_6141,N_4832,N_5199);
or U6142 (N_6142,N_4951,N_4809);
and U6143 (N_6143,N_4871,N_5581);
or U6144 (N_6144,N_5151,N_5577);
nor U6145 (N_6145,N_4003,N_5051);
nand U6146 (N_6146,N_5788,N_5662);
and U6147 (N_6147,N_4215,N_5419);
xnor U6148 (N_6148,N_5562,N_5565);
xnor U6149 (N_6149,N_4958,N_5805);
nand U6150 (N_6150,N_4631,N_4212);
nand U6151 (N_6151,N_4303,N_4151);
or U6152 (N_6152,N_4427,N_4426);
nor U6153 (N_6153,N_5395,N_4993);
and U6154 (N_6154,N_5345,N_4260);
and U6155 (N_6155,N_4889,N_4099);
nor U6156 (N_6156,N_5601,N_5640);
and U6157 (N_6157,N_4829,N_4419);
nand U6158 (N_6158,N_4019,N_4626);
nand U6159 (N_6159,N_4320,N_5939);
and U6160 (N_6160,N_5806,N_4636);
nor U6161 (N_6161,N_4529,N_5260);
xnor U6162 (N_6162,N_4929,N_4309);
xnor U6163 (N_6163,N_4186,N_5919);
or U6164 (N_6164,N_4135,N_4114);
or U6165 (N_6165,N_4390,N_4602);
or U6166 (N_6166,N_5392,N_4691);
or U6167 (N_6167,N_4272,N_5850);
and U6168 (N_6168,N_4130,N_5923);
xor U6169 (N_6169,N_5292,N_4155);
and U6170 (N_6170,N_4790,N_5069);
or U6171 (N_6171,N_4253,N_4485);
xnor U6172 (N_6172,N_4029,N_5239);
nor U6173 (N_6173,N_4361,N_4123);
nand U6174 (N_6174,N_4739,N_5406);
nand U6175 (N_6175,N_4734,N_4306);
or U6176 (N_6176,N_4086,N_5515);
xor U6177 (N_6177,N_4985,N_5815);
xor U6178 (N_6178,N_4826,N_4285);
and U6179 (N_6179,N_4684,N_5120);
xor U6180 (N_6180,N_5780,N_4665);
nand U6181 (N_6181,N_4256,N_4468);
nor U6182 (N_6182,N_4208,N_5506);
nand U6183 (N_6183,N_4818,N_4380);
or U6184 (N_6184,N_4201,N_5364);
or U6185 (N_6185,N_4481,N_5568);
xnor U6186 (N_6186,N_4724,N_5021);
and U6187 (N_6187,N_5698,N_4574);
nor U6188 (N_6188,N_5017,N_4534);
and U6189 (N_6189,N_5542,N_4483);
nand U6190 (N_6190,N_4949,N_4982);
and U6191 (N_6191,N_4273,N_4899);
xor U6192 (N_6192,N_4719,N_4165);
and U6193 (N_6193,N_4585,N_5618);
and U6194 (N_6194,N_4421,N_4578);
and U6195 (N_6195,N_5794,N_4647);
nand U6196 (N_6196,N_4048,N_4128);
nand U6197 (N_6197,N_4674,N_4403);
or U6198 (N_6198,N_5998,N_5867);
nor U6199 (N_6199,N_5580,N_5963);
xnor U6200 (N_6200,N_4823,N_4059);
xor U6201 (N_6201,N_5912,N_5827);
nand U6202 (N_6202,N_4500,N_5774);
or U6203 (N_6203,N_5418,N_4905);
xnor U6204 (N_6204,N_5126,N_4791);
and U6205 (N_6205,N_4974,N_4821);
nand U6206 (N_6206,N_4008,N_5525);
or U6207 (N_6207,N_5560,N_4297);
xor U6208 (N_6208,N_4336,N_5634);
or U6209 (N_6209,N_5609,N_4033);
or U6210 (N_6210,N_5365,N_4162);
xor U6211 (N_6211,N_4707,N_4461);
and U6212 (N_6212,N_5598,N_4382);
and U6213 (N_6213,N_5257,N_5523);
nor U6214 (N_6214,N_5737,N_5277);
nand U6215 (N_6215,N_4460,N_5301);
and U6216 (N_6216,N_4439,N_4373);
nand U6217 (N_6217,N_5216,N_4681);
xnor U6218 (N_6218,N_4735,N_4786);
or U6219 (N_6219,N_5348,N_5687);
or U6220 (N_6220,N_4979,N_5653);
nand U6221 (N_6221,N_5615,N_5723);
nor U6222 (N_6222,N_4362,N_4516);
xnor U6223 (N_6223,N_4752,N_4759);
or U6224 (N_6224,N_4769,N_5123);
xnor U6225 (N_6225,N_5013,N_4552);
or U6226 (N_6226,N_4070,N_5494);
xor U6227 (N_6227,N_5370,N_4065);
xor U6228 (N_6228,N_5747,N_5517);
or U6229 (N_6229,N_4032,N_5770);
and U6230 (N_6230,N_5652,N_4153);
nor U6231 (N_6231,N_4041,N_4614);
or U6232 (N_6232,N_4726,N_4172);
nand U6233 (N_6233,N_5768,N_4694);
and U6234 (N_6234,N_4970,N_4570);
or U6235 (N_6235,N_4693,N_5274);
or U6236 (N_6236,N_4042,N_5891);
nor U6237 (N_6237,N_4470,N_4802);
xor U6238 (N_6238,N_5933,N_5758);
xnor U6239 (N_6239,N_5060,N_5102);
nor U6240 (N_6240,N_5820,N_5579);
nand U6241 (N_6241,N_5325,N_4058);
nor U6242 (N_6242,N_5298,N_5323);
nand U6243 (N_6243,N_4234,N_5592);
and U6244 (N_6244,N_5976,N_5371);
nor U6245 (N_6245,N_4510,N_5101);
or U6246 (N_6246,N_4582,N_4706);
nor U6247 (N_6247,N_5819,N_5282);
or U6248 (N_6248,N_4598,N_5256);
xor U6249 (N_6249,N_5512,N_4085);
nor U6250 (N_6250,N_4429,N_4538);
xnor U6251 (N_6251,N_4011,N_4148);
xor U6252 (N_6252,N_4801,N_5033);
xor U6253 (N_6253,N_4353,N_5475);
and U6254 (N_6254,N_4747,N_5839);
xnor U6255 (N_6255,N_4930,N_5179);
nor U6256 (N_6256,N_5812,N_4414);
nor U6257 (N_6257,N_4505,N_4034);
nor U6258 (N_6258,N_4475,N_4828);
or U6259 (N_6259,N_4337,N_4836);
or U6260 (N_6260,N_5883,N_4271);
xnor U6261 (N_6261,N_5398,N_5242);
nand U6262 (N_6262,N_5296,N_4575);
nor U6263 (N_6263,N_4640,N_5789);
and U6264 (N_6264,N_4064,N_5741);
nor U6265 (N_6265,N_4599,N_4700);
xnor U6266 (N_6266,N_4129,N_4758);
xor U6267 (N_6267,N_5674,N_5118);
xor U6268 (N_6268,N_5295,N_4044);
nor U6269 (N_6269,N_5884,N_4134);
or U6270 (N_6270,N_4347,N_5196);
xor U6271 (N_6271,N_5203,N_5059);
nand U6272 (N_6272,N_4977,N_4643);
and U6273 (N_6273,N_5376,N_5584);
nand U6274 (N_6274,N_4031,N_5214);
xor U6275 (N_6275,N_5053,N_5659);
xor U6276 (N_6276,N_5453,N_4022);
and U6277 (N_6277,N_4825,N_5755);
xnor U6278 (N_6278,N_5997,N_4392);
nand U6279 (N_6279,N_4713,N_4730);
nor U6280 (N_6280,N_5155,N_4553);
and U6281 (N_6281,N_5833,N_5067);
and U6282 (N_6282,N_5682,N_4459);
or U6283 (N_6283,N_5248,N_4683);
and U6284 (N_6284,N_5879,N_5340);
nand U6285 (N_6285,N_4232,N_4712);
or U6286 (N_6286,N_4557,N_5076);
xnor U6287 (N_6287,N_5134,N_4290);
nand U6288 (N_6288,N_5969,N_4338);
xor U6289 (N_6289,N_4422,N_5776);
nand U6290 (N_6290,N_5684,N_5750);
nor U6291 (N_6291,N_5564,N_5465);
nand U6292 (N_6292,N_5078,N_5994);
nand U6293 (N_6293,N_4848,N_4433);
nand U6294 (N_6294,N_5916,N_5738);
nor U6295 (N_6295,N_5007,N_4616);
or U6296 (N_6296,N_5009,N_4948);
and U6297 (N_6297,N_5522,N_5178);
or U6298 (N_6298,N_4307,N_5336);
or U6299 (N_6299,N_4559,N_4531);
nand U6300 (N_6300,N_4893,N_4294);
nor U6301 (N_6301,N_5896,N_5029);
nor U6302 (N_6302,N_4843,N_4774);
and U6303 (N_6303,N_5661,N_4096);
nand U6304 (N_6304,N_4445,N_4898);
xnor U6305 (N_6305,N_5639,N_5046);
and U6306 (N_6306,N_5310,N_4143);
and U6307 (N_6307,N_5582,N_5907);
nand U6308 (N_6308,N_4150,N_4118);
or U6309 (N_6309,N_4443,N_4139);
and U6310 (N_6310,N_4071,N_4226);
and U6311 (N_6311,N_5114,N_5200);
and U6312 (N_6312,N_5803,N_5428);
xor U6313 (N_6313,N_5589,N_4762);
or U6314 (N_6314,N_5625,N_5644);
and U6315 (N_6315,N_4975,N_4101);
and U6316 (N_6316,N_5086,N_5034);
xnor U6317 (N_6317,N_5670,N_5610);
nor U6318 (N_6318,N_5420,N_4654);
nand U6319 (N_6319,N_5469,N_4863);
or U6320 (N_6320,N_4910,N_4918);
and U6321 (N_6321,N_4239,N_4770);
nor U6322 (N_6322,N_4645,N_4878);
nor U6323 (N_6323,N_4989,N_4230);
nor U6324 (N_6324,N_5587,N_4933);
nand U6325 (N_6325,N_4685,N_4870);
nand U6326 (N_6326,N_4913,N_5594);
xor U6327 (N_6327,N_5779,N_5887);
nand U6328 (N_6328,N_5057,N_5759);
and U6329 (N_6329,N_4431,N_5965);
nor U6330 (N_6330,N_4947,N_5100);
nand U6331 (N_6331,N_5308,N_4660);
xnor U6332 (N_6332,N_5981,N_5180);
and U6333 (N_6333,N_5656,N_4767);
or U6334 (N_6334,N_5458,N_4157);
xnor U6335 (N_6335,N_4545,N_5329);
nor U6336 (N_6336,N_4400,N_4238);
nand U6337 (N_6337,N_4120,N_5771);
nor U6338 (N_6338,N_4455,N_4125);
nand U6339 (N_6339,N_5544,N_4780);
xnor U6340 (N_6340,N_4012,N_5142);
or U6341 (N_6341,N_4943,N_5518);
nor U6342 (N_6342,N_5527,N_4378);
xnor U6343 (N_6343,N_5268,N_4744);
and U6344 (N_6344,N_5231,N_4334);
xor U6345 (N_6345,N_5765,N_4269);
and U6346 (N_6346,N_5253,N_4717);
and U6347 (N_6347,N_5356,N_4904);
or U6348 (N_6348,N_4486,N_5980);
nor U6349 (N_6349,N_4349,N_5466);
or U6350 (N_6350,N_4617,N_4728);
nor U6351 (N_6351,N_4259,N_5946);
xnor U6352 (N_6352,N_5600,N_5605);
nor U6353 (N_6353,N_5556,N_4384);
and U6354 (N_6354,N_4881,N_5084);
or U6355 (N_6355,N_5147,N_4687);
and U6356 (N_6356,N_4772,N_5689);
nand U6357 (N_6357,N_4757,N_4677);
nor U6358 (N_6358,N_4210,N_4509);
or U6359 (N_6359,N_4699,N_5400);
nor U6360 (N_6360,N_5866,N_4754);
nor U6361 (N_6361,N_4368,N_5711);
and U6362 (N_6362,N_5085,N_4702);
xor U6363 (N_6363,N_5728,N_5243);
or U6364 (N_6364,N_4973,N_4850);
and U6365 (N_6365,N_5591,N_4953);
or U6366 (N_6366,N_5319,N_4180);
and U6367 (N_6367,N_4903,N_5697);
xor U6368 (N_6368,N_5679,N_4147);
nor U6369 (N_6369,N_5186,N_5626);
nand U6370 (N_6370,N_4496,N_4976);
and U6371 (N_6371,N_5553,N_4592);
or U6372 (N_6372,N_4698,N_4163);
xor U6373 (N_6373,N_4849,N_4209);
nand U6374 (N_6374,N_5426,N_4216);
nand U6375 (N_6375,N_5262,N_4110);
and U6376 (N_6376,N_5138,N_4880);
or U6377 (N_6377,N_5389,N_5010);
nor U6378 (N_6378,N_5182,N_4177);
xor U6379 (N_6379,N_5885,N_4391);
or U6380 (N_6380,N_4595,N_5417);
or U6381 (N_6381,N_4891,N_5245);
and U6382 (N_6382,N_5903,N_5250);
nand U6383 (N_6383,N_4401,N_5769);
nand U6384 (N_6384,N_5860,N_4420);
xor U6385 (N_6385,N_5720,N_4229);
xor U6386 (N_6386,N_4709,N_5849);
nor U6387 (N_6387,N_4961,N_5359);
and U6388 (N_6388,N_4190,N_5092);
nand U6389 (N_6389,N_4466,N_4619);
and U6390 (N_6390,N_5316,N_5409);
nand U6391 (N_6391,N_4844,N_5505);
nand U6392 (N_6392,N_4199,N_4890);
and U6393 (N_6393,N_4025,N_5079);
nand U6394 (N_6394,N_4983,N_4090);
and U6395 (N_6395,N_4244,N_5022);
and U6396 (N_6396,N_5058,N_5533);
nand U6397 (N_6397,N_4417,N_5590);
nand U6398 (N_6398,N_4142,N_4805);
xor U6399 (N_6399,N_4122,N_5635);
or U6400 (N_6400,N_4300,N_5487);
xor U6401 (N_6401,N_5460,N_5211);
or U6402 (N_6402,N_4884,N_5039);
and U6403 (N_6403,N_4243,N_5349);
xor U6404 (N_6404,N_4376,N_5902);
nand U6405 (N_6405,N_4221,N_5063);
nor U6406 (N_6406,N_4865,N_4872);
nor U6407 (N_6407,N_4432,N_4579);
xnor U6408 (N_6408,N_5176,N_4356);
or U6409 (N_6409,N_5499,N_4237);
or U6410 (N_6410,N_5121,N_5838);
xnor U6411 (N_6411,N_5930,N_5864);
or U6412 (N_6412,N_4167,N_5403);
and U6413 (N_6413,N_4815,N_5001);
and U6414 (N_6414,N_5975,N_4955);
nor U6415 (N_6415,N_5408,N_4746);
xor U6416 (N_6416,N_5045,N_5578);
nand U6417 (N_6417,N_5957,N_5501);
nand U6418 (N_6418,N_5772,N_4673);
and U6419 (N_6419,N_5287,N_5072);
and U6420 (N_6420,N_4176,N_4332);
and U6421 (N_6421,N_4957,N_4441);
or U6422 (N_6422,N_4532,N_5906);
nand U6423 (N_6423,N_5853,N_4517);
and U6424 (N_6424,N_4442,N_5649);
xor U6425 (N_6425,N_4723,N_4882);
xnor U6426 (N_6426,N_4539,N_4493);
xor U6427 (N_6427,N_5703,N_4803);
or U6428 (N_6428,N_4415,N_5561);
and U6429 (N_6429,N_4081,N_4440);
and U6430 (N_6430,N_4576,N_4006);
and U6431 (N_6431,N_5918,N_5869);
nand U6432 (N_6432,N_4301,N_4037);
nand U6433 (N_6433,N_4437,N_4169);
or U6434 (N_6434,N_4246,N_4644);
nand U6435 (N_6435,N_5066,N_5538);
or U6436 (N_6436,N_4627,N_4395);
and U6437 (N_6437,N_5841,N_5847);
nand U6438 (N_6438,N_4076,N_5492);
nand U6439 (N_6439,N_5832,N_4051);
nand U6440 (N_6440,N_5068,N_5425);
and U6441 (N_6441,N_4520,N_4158);
nor U6442 (N_6442,N_4457,N_4895);
or U6443 (N_6443,N_5153,N_4959);
nor U6444 (N_6444,N_4714,N_4354);
and U6445 (N_6445,N_5163,N_4187);
nand U6446 (N_6446,N_5169,N_4811);
and U6447 (N_6447,N_5279,N_4372);
and U6448 (N_6448,N_4972,N_4197);
nor U6449 (N_6449,N_5681,N_4628);
xor U6450 (N_6450,N_5437,N_4804);
and U6451 (N_6451,N_5777,N_4078);
nor U6452 (N_6452,N_4068,N_4017);
nor U6453 (N_6453,N_4479,N_4787);
and U6454 (N_6454,N_4482,N_4922);
xor U6455 (N_6455,N_5146,N_4411);
xnor U6456 (N_6456,N_5122,N_5895);
and U6457 (N_6457,N_5441,N_5899);
or U6458 (N_6458,N_5929,N_4521);
nand U6459 (N_6459,N_5093,N_5521);
nand U6460 (N_6460,N_5436,N_5339);
or U6461 (N_6461,N_5572,N_4249);
nor U6462 (N_6462,N_5773,N_4277);
nand U6463 (N_6463,N_4478,N_5602);
or U6464 (N_6464,N_5136,N_4727);
nand U6465 (N_6465,N_5149,N_4100);
nor U6466 (N_6466,N_5476,N_4926);
and U6467 (N_6467,N_4506,N_4149);
or U6468 (N_6468,N_5749,N_5341);
nand U6469 (N_6469,N_4689,N_5987);
xnor U6470 (N_6470,N_4344,N_5185);
or U6471 (N_6471,N_5116,N_4383);
or U6472 (N_6472,N_4289,N_4857);
nand U6473 (N_6473,N_4112,N_5942);
nor U6474 (N_6474,N_4639,N_4305);
and U6475 (N_6475,N_5870,N_4225);
xnor U6476 (N_6476,N_4369,N_4015);
nor U6477 (N_6477,N_5889,N_5893);
nor U6478 (N_6478,N_4995,N_4326);
and U6479 (N_6479,N_4073,N_4618);
and U6480 (N_6480,N_4137,N_5157);
nor U6481 (N_6481,N_5950,N_5931);
nand U6482 (N_6482,N_5450,N_5781);
xnor U6483 (N_6483,N_4967,N_4472);
nor U6484 (N_6484,N_4340,N_5224);
and U6485 (N_6485,N_5690,N_5227);
xor U6486 (N_6486,N_4393,N_5914);
nor U6487 (N_6487,N_5088,N_4751);
nand U6488 (N_6488,N_4346,N_4615);
xor U6489 (N_6489,N_4554,N_4480);
or U6490 (N_6490,N_5381,N_5638);
and U6491 (N_6491,N_4055,N_5383);
and U6492 (N_6492,N_5686,N_4281);
nand U6493 (N_6493,N_5174,N_4495);
nor U6494 (N_6494,N_4839,N_5548);
nand U6495 (N_6495,N_5035,N_4288);
xor U6496 (N_6496,N_5011,N_4254);
xnor U6497 (N_6497,N_4292,N_4588);
and U6498 (N_6498,N_4625,N_4733);
nand U6499 (N_6499,N_4605,N_5135);
xnor U6500 (N_6500,N_4310,N_5019);
nor U6501 (N_6501,N_4080,N_5377);
nand U6502 (N_6502,N_5081,N_5766);
xnor U6503 (N_6503,N_4508,N_5936);
and U6504 (N_6504,N_4792,N_4311);
xor U6505 (N_6505,N_4407,N_4885);
or U6506 (N_6506,N_5397,N_5463);
nor U6507 (N_6507,N_4653,N_4258);
or U6508 (N_6508,N_4845,N_5666);
xor U6509 (N_6509,N_5831,N_5541);
or U6510 (N_6510,N_4423,N_4161);
or U6511 (N_6511,N_4664,N_5124);
or U6512 (N_6512,N_5306,N_4630);
nand U6513 (N_6513,N_4748,N_4612);
nor U6514 (N_6514,N_4590,N_5655);
nor U6515 (N_6515,N_4869,N_4206);
or U6516 (N_6516,N_5220,N_5438);
xnor U6517 (N_6517,N_5825,N_4020);
nand U6518 (N_6518,N_5551,N_5240);
nand U6519 (N_6519,N_5286,N_5843);
nand U6520 (N_6520,N_4072,N_5107);
xnor U6521 (N_6521,N_4035,N_4196);
xnor U6522 (N_6522,N_5790,N_5171);
nor U6523 (N_6523,N_4657,N_5654);
nor U6524 (N_6524,N_5165,N_5432);
xor U6525 (N_6525,N_4121,N_4079);
nand U6526 (N_6526,N_4146,N_5159);
or U6527 (N_6527,N_4950,N_5816);
nand U6528 (N_6528,N_4132,N_5455);
nand U6529 (N_6529,N_5353,N_4451);
and U6530 (N_6530,N_5616,N_4668);
or U6531 (N_6531,N_5543,N_5128);
and U6532 (N_6532,N_5859,N_4536);
nand U6533 (N_6533,N_4325,N_4996);
nand U6534 (N_6534,N_5620,N_4404);
nor U6535 (N_6535,N_5778,N_5290);
or U6536 (N_6536,N_4965,N_5865);
nor U6537 (N_6537,N_4789,N_4641);
and U6538 (N_6538,N_5586,N_5559);
and U6539 (N_6539,N_4278,N_4560);
nor U6540 (N_6540,N_4386,N_5576);
xor U6541 (N_6541,N_4370,N_4240);
and U6542 (N_6542,N_4919,N_4862);
xnor U6543 (N_6543,N_5558,N_5020);
and U6544 (N_6544,N_5056,N_5549);
nand U6545 (N_6545,N_5872,N_4141);
nand U6546 (N_6546,N_5484,N_5236);
nor U6547 (N_6547,N_4827,N_4750);
nand U6548 (N_6548,N_4573,N_5491);
xor U6549 (N_6549,N_4991,N_5575);
and U6550 (N_6550,N_4710,N_5982);
nor U6551 (N_6551,N_5382,N_4425);
or U6552 (N_6552,N_5804,N_5960);
xor U6553 (N_6553,N_4476,N_5244);
or U6554 (N_6554,N_4335,N_5739);
xor U6555 (N_6555,N_5255,N_4266);
nor U6556 (N_6556,N_4126,N_4888);
and U6557 (N_6557,N_5258,N_5630);
nor U6558 (N_6558,N_5588,N_4255);
or U6559 (N_6559,N_5628,N_5861);
nand U6560 (N_6560,N_5489,N_5809);
and U6561 (N_6561,N_5041,N_4923);
nor U6562 (N_6562,N_4901,N_4077);
and U6563 (N_6563,N_4124,N_4667);
and U6564 (N_6564,N_4464,N_4105);
or U6565 (N_6565,N_4766,N_5347);
and U6566 (N_6566,N_5495,N_5545);
nor U6567 (N_6567,N_5173,N_5229);
xnor U6568 (N_6568,N_5368,N_4501);
nand U6569 (N_6569,N_5730,N_5456);
nand U6570 (N_6570,N_5852,N_5593);
xor U6571 (N_6571,N_4834,N_5452);
and U6572 (N_6572,N_5995,N_5909);
nand U6573 (N_6573,N_5955,N_5000);
nor U6574 (N_6574,N_4291,N_5351);
or U6575 (N_6575,N_5753,N_5877);
nor U6576 (N_6576,N_5097,N_5346);
and U6577 (N_6577,N_5194,N_5956);
xnor U6578 (N_6578,N_4650,N_4649);
and U6579 (N_6579,N_4672,N_4765);
or U6580 (N_6580,N_4159,N_5552);
xor U6581 (N_6581,N_5327,N_5717);
nor U6582 (N_6582,N_5660,N_5665);
nand U6583 (N_6583,N_4107,N_5528);
and U6584 (N_6584,N_4469,N_5191);
xnor U6585 (N_6585,N_4178,N_5137);
nand U6586 (N_6586,N_5106,N_4964);
or U6587 (N_6587,N_5500,N_5217);
xor U6588 (N_6588,N_4543,N_4117);
and U6589 (N_6589,N_5307,N_5958);
nand U6590 (N_6590,N_4028,N_4398);
nor U6591 (N_6591,N_4587,N_5272);
or U6592 (N_6592,N_5451,N_4601);
xor U6593 (N_6593,N_5181,N_5490);
nand U6594 (N_6594,N_4864,N_5386);
nand U6595 (N_6595,N_5429,N_5488);
xor U6596 (N_6596,N_5312,N_5837);
nor U6597 (N_6597,N_4140,N_5818);
nand U6598 (N_6598,N_4083,N_4638);
or U6599 (N_6599,N_4315,N_4855);
and U6600 (N_6600,N_5675,N_4005);
nand U6601 (N_6601,N_5937,N_4195);
nor U6602 (N_6602,N_5844,N_4963);
or U6603 (N_6603,N_4695,N_4830);
xor U6604 (N_6604,N_4795,N_4116);
xnor U6605 (N_6605,N_5314,N_5354);
nor U6606 (N_6606,N_4798,N_5387);
xor U6607 (N_6607,N_5028,N_4971);
and U6608 (N_6608,N_4875,N_4027);
nand U6609 (N_6609,N_5413,N_4749);
and U6610 (N_6610,N_5842,N_4102);
nand U6611 (N_6611,N_5573,N_5834);
xor U6612 (N_6612,N_4250,N_4669);
nand U6613 (N_6613,N_5144,N_5800);
or U6614 (N_6614,N_5251,N_5075);
xor U6615 (N_6615,N_4348,N_5201);
nor U6616 (N_6616,N_5751,N_5115);
nor U6617 (N_6617,N_4295,N_4235);
nor U6618 (N_6618,N_5732,N_5954);
nor U6619 (N_6619,N_4652,N_4637);
nand U6620 (N_6620,N_4374,N_5725);
nor U6621 (N_6621,N_4435,N_5978);
and U6622 (N_6622,N_5696,N_5407);
nand U6623 (N_6623,N_4854,N_5205);
and U6624 (N_6624,N_4263,N_4530);
and U6625 (N_6625,N_4715,N_5875);
or U6626 (N_6626,N_4634,N_4257);
nor U6627 (N_6627,N_4219,N_5024);
xor U6628 (N_6628,N_4666,N_4567);
or U6629 (N_6629,N_4045,N_5924);
and U6630 (N_6630,N_4050,N_5261);
nand U6631 (N_6631,N_5444,N_4245);
nand U6632 (N_6632,N_4581,N_4632);
nor U6633 (N_6633,N_4341,N_4548);
or U6634 (N_6634,N_5324,N_5715);
or U6635 (N_6635,N_5234,N_5133);
nor U6636 (N_6636,N_4586,N_5154);
nor U6637 (N_6637,N_4793,N_4981);
nor U6638 (N_6638,N_5421,N_4188);
xnor U6639 (N_6639,N_5464,N_5643);
and U6640 (N_6640,N_5740,N_4566);
xnor U6641 (N_6641,N_5692,N_4528);
nand U6642 (N_6642,N_4473,N_5405);
nand U6643 (N_6643,N_4690,N_5038);
xnor U6644 (N_6644,N_4270,N_4662);
and U6645 (N_6645,N_4861,N_5817);
and U6646 (N_6646,N_4218,N_4860);
and U6647 (N_6647,N_4352,N_4359);
nand U6648 (N_6648,N_5332,N_4446);
or U6649 (N_6649,N_5162,N_4998);
nor U6650 (N_6650,N_4293,N_4363);
and U6651 (N_6651,N_5073,N_4944);
xor U6652 (N_6652,N_4945,N_5676);
nor U6653 (N_6653,N_5317,N_5707);
and U6654 (N_6654,N_4642,N_4814);
and U6655 (N_6655,N_4806,N_5055);
nor U6656 (N_6656,N_4868,N_5566);
and U6657 (N_6657,N_4220,N_5311);
and U6658 (N_6658,N_5934,N_5004);
nand U6659 (N_6659,N_5254,N_5905);
nand U6660 (N_6660,N_4859,N_4527);
and U6661 (N_6661,N_4164,N_4207);
nand U6662 (N_6662,N_4447,N_5480);
or U6663 (N_6663,N_4252,N_4651);
and U6664 (N_6664,N_5358,N_4931);
nor U6665 (N_6665,N_4000,N_5299);
or U6666 (N_6666,N_5546,N_5271);
xnor U6667 (N_6667,N_4021,N_4883);
or U6668 (N_6668,N_5247,N_4379);
and U6669 (N_6669,N_5015,N_4075);
nor U6670 (N_6670,N_4564,N_4405);
or U6671 (N_6671,N_5641,N_4138);
and U6672 (N_6672,N_5267,N_5477);
nor U6673 (N_6673,N_4345,N_5003);
nand U6674 (N_6674,N_4456,N_4168);
and U6675 (N_6675,N_5595,N_5904);
xor U6676 (N_6676,N_5979,N_5798);
nand U6677 (N_6677,N_5393,N_4261);
nor U6678 (N_6678,N_4304,N_4565);
nor U6679 (N_6679,N_4676,N_4987);
or U6680 (N_6680,N_4454,N_4502);
nor U6681 (N_6681,N_5369,N_4997);
nor U6682 (N_6682,N_4498,N_5599);
and U6683 (N_6683,N_4783,N_5694);
nand U6684 (N_6684,N_4499,N_5871);
or U6685 (N_6685,N_5984,N_4540);
or U6686 (N_6686,N_4200,N_4194);
or U6687 (N_6687,N_5614,N_5603);
and U6688 (N_6688,N_5270,N_5091);
xor U6689 (N_6689,N_4686,N_4233);
and U6690 (N_6690,N_4541,N_4413);
xor U6691 (N_6691,N_4542,N_4604);
and U6692 (N_6692,N_5284,N_4002);
xnor U6693 (N_6693,N_4396,N_5023);
and U6694 (N_6694,N_4621,N_4333);
xnor U6695 (N_6695,N_5141,N_5187);
or U6696 (N_6696,N_5734,N_5760);
xnor U6697 (N_6697,N_5757,N_4912);
xnor U6698 (N_6698,N_4284,N_5840);
nand U6699 (N_6699,N_4978,N_4866);
or U6700 (N_6700,N_5947,N_4166);
xor U6701 (N_6701,N_5534,N_4785);
and U6702 (N_6702,N_4103,N_5334);
nand U6703 (N_6703,N_4394,N_5952);
nor U6704 (N_6704,N_5898,N_4661);
and U6705 (N_6705,N_5763,N_5303);
nor U6706 (N_6706,N_5782,N_5736);
or U6707 (N_6707,N_4779,N_5964);
xor U6708 (N_6708,N_4833,N_4192);
nand U6709 (N_6709,N_5478,N_4914);
or U6710 (N_6710,N_5830,N_4287);
or U6711 (N_6711,N_5504,N_4966);
or U6712 (N_6712,N_4399,N_5913);
xnor U6713 (N_6713,N_5854,N_4778);
or U6714 (N_6714,N_4607,N_5519);
nor U6715 (N_6715,N_5228,N_5378);
xnor U6716 (N_6716,N_4682,N_4526);
and U6717 (N_6717,N_5198,N_5230);
nand U6718 (N_6718,N_5482,N_5754);
xnor U6719 (N_6719,N_5471,N_5467);
and U6720 (N_6720,N_5631,N_4523);
nand U6721 (N_6721,N_4892,N_4606);
or U6722 (N_6722,N_4902,N_4794);
nor U6723 (N_6723,N_5448,N_5481);
xor U6724 (N_6724,N_4594,N_4283);
nand U6725 (N_6725,N_4663,N_4928);
nor U6726 (N_6726,N_4512,N_5322);
or U6727 (N_6727,N_5410,N_5606);
nor U6728 (N_6728,N_4563,N_5440);
xor U6729 (N_6729,N_4355,N_4136);
and U6730 (N_6730,N_4412,N_5212);
nor U6731 (N_6731,N_5373,N_5264);
or U6732 (N_6732,N_4060,N_4946);
nand U6733 (N_6733,N_4438,N_4807);
or U6734 (N_6734,N_5433,N_5090);
or U6735 (N_6735,N_5192,N_4365);
nor U6736 (N_6736,N_4596,N_4518);
nand U6737 (N_6737,N_5632,N_5977);
and U6738 (N_6738,N_5232,N_5953);
and U6739 (N_6739,N_4402,N_5972);
xor U6740 (N_6740,N_4646,N_4203);
xor U6741 (N_6741,N_5714,N_4648);
nor U6742 (N_6742,N_5170,N_4688);
nor U6743 (N_6743,N_5764,N_4191);
nand U6744 (N_6744,N_5473,N_5695);
or U6745 (N_6745,N_4537,N_4920);
nand U6746 (N_6746,N_4731,N_5507);
or U6747 (N_6747,N_4331,N_5555);
and U6748 (N_6748,N_5252,N_5951);
xor U6749 (N_6749,N_5829,N_4474);
nor U6750 (N_6750,N_5160,N_5394);
nor U6751 (N_6751,N_5411,N_4624);
or U6752 (N_6752,N_4492,N_4436);
xnor U6753 (N_6753,N_4387,N_5350);
nor U6754 (N_6754,N_4487,N_5563);
or U6755 (N_6755,N_4434,N_4182);
xor U6756 (N_6756,N_5985,N_5607);
xnor U6757 (N_6757,N_5077,N_5862);
and U6758 (N_6758,N_4952,N_4782);
or U6759 (N_6759,N_4416,N_4222);
and U6760 (N_6760,N_5932,N_4317);
nor U6761 (N_6761,N_4716,N_4819);
xor U6762 (N_6762,N_4704,N_4316);
and U6763 (N_6763,N_4841,N_5082);
nand U6764 (N_6764,N_5372,N_5745);
or U6765 (N_6765,N_5140,N_5801);
nand U6766 (N_6766,N_5569,N_5219);
nand U6767 (N_6767,N_5095,N_5925);
nor U6768 (N_6768,N_4087,N_5040);
nor U6769 (N_6769,N_5657,N_4013);
xnor U6770 (N_6770,N_5043,N_4896);
or U6771 (N_6771,N_5288,N_4251);
nor U6772 (N_6772,N_4658,N_4236);
nand U6773 (N_6773,N_5014,N_4737);
nand U6774 (N_6774,N_5103,N_5917);
or U6775 (N_6775,N_4927,N_5968);
or U6776 (N_6776,N_5721,N_4609);
nor U6777 (N_6777,N_5388,N_4680);
nor U6778 (N_6778,N_5177,N_5266);
and U6779 (N_6779,N_5479,N_4760);
xnor U6780 (N_6780,N_4154,N_4504);
nand U6781 (N_6781,N_4184,N_5604);
nand U6782 (N_6782,N_5646,N_4066);
xor U6783 (N_6783,N_5087,N_5719);
nand U6784 (N_6784,N_5498,N_4308);
or U6785 (N_6785,N_5099,N_4810);
or U6786 (N_6786,N_5027,N_5235);
nand U6787 (N_6787,N_4796,N_5624);
and U6788 (N_6788,N_5375,N_4736);
nor U6789 (N_6789,N_4465,N_5222);
xnor U6790 (N_6790,N_5018,N_4580);
nor U6791 (N_6791,N_5516,N_5190);
nor U6792 (N_6792,N_5281,N_5928);
xnor U6793 (N_6793,N_5280,N_5424);
and U6794 (N_6794,N_5127,N_4067);
nand U6795 (N_6795,N_4094,N_4753);
and U6796 (N_6796,N_4781,N_4204);
nor U6797 (N_6797,N_5716,N_4507);
nor U6798 (N_6798,N_4988,N_4463);
xor U6799 (N_6799,N_5249,N_4740);
and U6800 (N_6800,N_5648,N_4069);
xor U6801 (N_6801,N_4556,N_5152);
or U6802 (N_6802,N_4838,N_4935);
and U6803 (N_6803,N_5320,N_4776);
xnor U6804 (N_6804,N_5070,N_5802);
nor U6805 (N_6805,N_4925,N_4679);
xor U6806 (N_6806,N_4016,N_5213);
and U6807 (N_6807,N_5197,N_5404);
and U6808 (N_6808,N_5164,N_5671);
or U6809 (N_6809,N_5744,N_4938);
xnor U6810 (N_6810,N_4296,N_5996);
nand U6811 (N_6811,N_5472,N_5167);
nand U6812 (N_6812,N_4549,N_4104);
and U6813 (N_6813,N_4375,N_5961);
and U6814 (N_6814,N_5032,N_5422);
xor U6815 (N_6815,N_5047,N_4088);
or U6816 (N_6816,N_4228,N_4703);
and U6817 (N_6817,N_5622,N_5927);
or U6818 (N_6818,N_4185,N_5857);
nor U6819 (N_6819,N_5890,N_4608);
or U6820 (N_6820,N_4410,N_4916);
nand U6821 (N_6821,N_5300,N_5729);
or U6822 (N_6822,N_5704,N_4550);
nor U6823 (N_6823,N_5535,N_5302);
nor U6824 (N_6824,N_4858,N_5983);
xnor U6825 (N_6825,N_4503,N_4145);
and U6826 (N_6826,N_4418,N_4214);
and U6827 (N_6827,N_5874,N_5708);
xor U6828 (N_6828,N_5608,N_4108);
xor U6829 (N_6829,N_4525,N_5074);
nand U6830 (N_6830,N_4428,N_5357);
or U6831 (N_6831,N_4494,N_5701);
nand U6832 (N_6832,N_4777,N_5184);
nand U6833 (N_6833,N_4745,N_5678);
nand U6834 (N_6834,N_4853,N_5485);
or U6835 (N_6835,N_4932,N_4817);
xnor U6836 (N_6836,N_5148,N_4800);
xnor U6837 (N_6837,N_4298,N_4268);
nand U6838 (N_6838,N_5826,N_5098);
xnor U6839 (N_6839,N_5132,N_5343);
nor U6840 (N_6840,N_5104,N_4160);
and U6841 (N_6841,N_5108,N_5237);
nor U6842 (N_6842,N_5944,N_5263);
xor U6843 (N_6843,N_4453,N_4350);
or U6844 (N_6844,N_4847,N_4248);
nor U6845 (N_6845,N_5366,N_5215);
or U6846 (N_6846,N_5294,N_5002);
and U6847 (N_6847,N_5291,N_5335);
xnor U6848 (N_6848,N_4840,N_5031);
nand U6849 (N_6849,N_5880,N_5054);
nor U6850 (N_6850,N_5360,N_5742);
xor U6851 (N_6851,N_4924,N_5811);
and U6852 (N_6852,N_4678,N_5379);
xor U6853 (N_6853,N_5633,N_5065);
nor U6854 (N_6854,N_5557,N_5208);
nand U6855 (N_6855,N_4156,N_4897);
xnor U6856 (N_6856,N_4279,N_5331);
and U6857 (N_6857,N_5496,N_5642);
and U6858 (N_6858,N_4591,N_5337);
nand U6859 (N_6859,N_5973,N_5321);
nand U6860 (N_6860,N_5005,N_5188);
and U6861 (N_6861,N_4040,N_5858);
and U6862 (N_6862,N_5636,N_4906);
nor U6863 (N_6863,N_5109,N_5718);
nand U6864 (N_6864,N_5474,N_4755);
xnor U6865 (N_6865,N_5702,N_4242);
xor U6866 (N_6866,N_5532,N_4057);
xor U6867 (N_6867,N_5344,N_4635);
nand U6868 (N_6868,N_4558,N_5746);
and U6869 (N_6869,N_5061,N_4039);
or U6870 (N_6870,N_4327,N_5283);
nor U6871 (N_6871,N_4111,N_5943);
nor U6872 (N_6872,N_5597,N_5988);
or U6873 (N_6873,N_4314,N_5278);
nor U6874 (N_6874,N_4342,N_5752);
and U6875 (N_6875,N_4328,N_5415);
or U6876 (N_6876,N_5524,N_5823);
xnor U6877 (N_6877,N_5637,N_5048);
or U6878 (N_6878,N_5412,N_5326);
or U6879 (N_6879,N_5209,N_4276);
nand U6880 (N_6880,N_5049,N_4364);
nand U6881 (N_6881,N_4873,N_5462);
nand U6882 (N_6882,N_5089,N_5113);
and U6883 (N_6883,N_4053,N_4089);
and U6884 (N_6884,N_5567,N_5685);
nand U6885 (N_6885,N_5767,N_4597);
nand U6886 (N_6886,N_5166,N_4062);
xnor U6887 (N_6887,N_5012,N_5442);
nor U6888 (N_6888,N_4179,N_4205);
or U6889 (N_6889,N_4708,N_5974);
or U6890 (N_6890,N_4572,N_4886);
nand U6891 (N_6891,N_4603,N_4038);
nand U6892 (N_6892,N_5878,N_5962);
xor U6893 (N_6893,N_4561,N_5416);
nand U6894 (N_6894,N_4941,N_4584);
nand U6895 (N_6895,N_4692,N_4671);
xor U6896 (N_6896,N_4371,N_4385);
xnor U6897 (N_6897,N_4323,N_5285);
xor U6898 (N_6898,N_5894,N_4856);
or U6899 (N_6899,N_5667,N_4052);
or U6900 (N_6900,N_4842,N_4822);
nand U6901 (N_6901,N_5915,N_5706);
or U6902 (N_6902,N_4513,N_5664);
nor U6903 (N_6903,N_4490,N_5783);
nand U6904 (N_6904,N_5726,N_5342);
xor U6905 (N_6905,N_5554,N_5966);
and U6906 (N_6906,N_5784,N_4360);
nor U6907 (N_6907,N_5309,N_5761);
nor U6908 (N_6908,N_4181,N_4224);
and U6909 (N_6909,N_4984,N_5083);
nor U6910 (N_6910,N_5168,N_4047);
xnor U6911 (N_6911,N_4175,N_5911);
or U6912 (N_6912,N_4874,N_4670);
or U6913 (N_6913,N_4934,N_5530);
nand U6914 (N_6914,N_4831,N_5876);
or U6915 (N_6915,N_4742,N_5627);
nand U6916 (N_6916,N_4546,N_4299);
nor U6917 (N_6917,N_4986,N_5808);
nor U6918 (N_6918,N_4720,N_5183);
and U6919 (N_6919,N_4458,N_5139);
or U6920 (N_6920,N_4741,N_4321);
nor U6921 (N_6921,N_5623,N_4152);
or U6922 (N_6922,N_5210,N_5338);
or U6923 (N_6923,N_5175,N_4620);
nand U6924 (N_6924,N_5677,N_5401);
xnor U6925 (N_6925,N_4018,N_5647);
or U6926 (N_6926,N_5238,N_5855);
nor U6927 (N_6927,N_4030,N_5629);
and U6928 (N_6928,N_5796,N_5938);
xnor U6929 (N_6929,N_4894,N_4471);
nand U6930 (N_6930,N_5713,N_4562);
nand U6931 (N_6931,N_5384,N_4568);
and U6932 (N_6932,N_5672,N_4497);
xor U6933 (N_6933,N_5454,N_5305);
nor U6934 (N_6934,N_4173,N_5967);
xor U6935 (N_6935,N_4837,N_5756);
and U6936 (N_6936,N_5330,N_4223);
and U6937 (N_6937,N_5921,N_5193);
xor U6938 (N_6938,N_4812,N_4247);
xnor U6939 (N_6939,N_5461,N_5683);
nand U6940 (N_6940,N_4820,N_5845);
and U6941 (N_6941,N_5531,N_5691);
xnor U6942 (N_6942,N_5989,N_4408);
or U6943 (N_6943,N_4909,N_4876);
or U6944 (N_6944,N_4171,N_5156);
or U6945 (N_6945,N_4514,N_5036);
or U6946 (N_6946,N_4887,N_5414);
or U6947 (N_6947,N_4280,N_4424);
or U6948 (N_6948,N_5940,N_4329);
xnor U6949 (N_6949,N_5762,N_5570);
and U6950 (N_6950,N_5207,N_5131);
and U6951 (N_6951,N_4940,N_4115);
xnor U6952 (N_6952,N_5434,N_5669);
and U6953 (N_6953,N_4879,N_5509);
or U6954 (N_6954,N_4877,N_4656);
xnor U6955 (N_6955,N_5547,N_5470);
nor U6956 (N_6956,N_4797,N_5735);
nor U6957 (N_6957,N_4725,N_5792);
nand U6958 (N_6958,N_4227,N_5096);
nor U6959 (N_6959,N_4265,N_4824);
xnor U6960 (N_6960,N_5390,N_5807);
nor U6961 (N_6961,N_4936,N_4756);
nor U6962 (N_6962,N_4937,N_5117);
nor U6963 (N_6963,N_4511,N_5536);
and U6964 (N_6964,N_5493,N_5901);
nand U6965 (N_6965,N_4098,N_4764);
nand U6966 (N_6966,N_4097,N_5508);
and U6967 (N_6967,N_5446,N_5289);
and U6968 (N_6968,N_4846,N_5926);
nor U6969 (N_6969,N_5846,N_4980);
or U6970 (N_6970,N_4213,N_4622);
nor U6971 (N_6971,N_4613,N_5391);
or U6972 (N_6972,N_5145,N_5094);
nand U6973 (N_6973,N_5571,N_4999);
nand U6974 (N_6974,N_5328,N_5218);
and U6975 (N_6975,N_5016,N_5241);
or U6976 (N_6976,N_5920,N_5202);
and U6977 (N_6977,N_5511,N_5468);
xnor U6978 (N_6978,N_4302,N_4969);
or U6979 (N_6979,N_4084,N_5037);
nor U6980 (N_6980,N_4771,N_5645);
nand U6981 (N_6981,N_4043,N_5439);
xor U6982 (N_6982,N_5276,N_5529);
and U6983 (N_6983,N_5550,N_4623);
nor U6984 (N_6984,N_5897,N_4330);
and U6985 (N_6985,N_5986,N_5727);
or U6986 (N_6986,N_4851,N_4917);
or U6987 (N_6987,N_5044,N_5265);
or U6988 (N_6988,N_5129,N_5374);
and U6989 (N_6989,N_4533,N_4939);
xnor U6990 (N_6990,N_5868,N_5619);
nor U6991 (N_6991,N_5991,N_5699);
xnor U6992 (N_6992,N_5680,N_5510);
nand U6993 (N_6993,N_5540,N_5941);
nand U6994 (N_6994,N_4921,N_5574);
or U6995 (N_6995,N_5836,N_5502);
nor U6996 (N_6996,N_5892,N_5821);
nor U6997 (N_6997,N_5787,N_5050);
and U6998 (N_6998,N_4915,N_4484);
nand U6999 (N_6999,N_4339,N_4202);
nor U7000 (N_7000,N_4283,N_5888);
or U7001 (N_7001,N_5790,N_4686);
nor U7002 (N_7002,N_4070,N_4794);
nor U7003 (N_7003,N_4881,N_5709);
or U7004 (N_7004,N_4972,N_4685);
nor U7005 (N_7005,N_5835,N_5266);
nor U7006 (N_7006,N_5384,N_5610);
nand U7007 (N_7007,N_4750,N_4570);
nor U7008 (N_7008,N_5442,N_4627);
xnor U7009 (N_7009,N_4780,N_5711);
nand U7010 (N_7010,N_5912,N_4011);
xnor U7011 (N_7011,N_4083,N_5235);
nand U7012 (N_7012,N_5408,N_5046);
and U7013 (N_7013,N_4956,N_5135);
xnor U7014 (N_7014,N_4461,N_5450);
xnor U7015 (N_7015,N_5684,N_4920);
nand U7016 (N_7016,N_5281,N_5871);
nor U7017 (N_7017,N_5731,N_4301);
nor U7018 (N_7018,N_4478,N_4851);
xor U7019 (N_7019,N_4903,N_4783);
nand U7020 (N_7020,N_4936,N_4097);
and U7021 (N_7021,N_5505,N_5759);
nor U7022 (N_7022,N_4275,N_5681);
nand U7023 (N_7023,N_5757,N_4168);
nor U7024 (N_7024,N_4524,N_5626);
and U7025 (N_7025,N_5577,N_4355);
and U7026 (N_7026,N_4294,N_4961);
and U7027 (N_7027,N_4018,N_4983);
nor U7028 (N_7028,N_5073,N_5685);
or U7029 (N_7029,N_4457,N_5648);
nor U7030 (N_7030,N_5930,N_4753);
nand U7031 (N_7031,N_5222,N_4749);
nand U7032 (N_7032,N_4297,N_5201);
or U7033 (N_7033,N_5690,N_5390);
and U7034 (N_7034,N_4157,N_4081);
nor U7035 (N_7035,N_5145,N_4621);
xor U7036 (N_7036,N_4096,N_5036);
nand U7037 (N_7037,N_4211,N_4231);
or U7038 (N_7038,N_5489,N_5099);
nand U7039 (N_7039,N_4102,N_4195);
nor U7040 (N_7040,N_4210,N_5733);
or U7041 (N_7041,N_5175,N_4265);
nor U7042 (N_7042,N_5047,N_5021);
nor U7043 (N_7043,N_4691,N_5908);
xnor U7044 (N_7044,N_4689,N_4914);
nor U7045 (N_7045,N_5103,N_5087);
xnor U7046 (N_7046,N_5926,N_5144);
nor U7047 (N_7047,N_4286,N_5620);
and U7048 (N_7048,N_4568,N_5423);
and U7049 (N_7049,N_5829,N_4687);
nor U7050 (N_7050,N_4384,N_5202);
or U7051 (N_7051,N_5758,N_5545);
nand U7052 (N_7052,N_5124,N_5273);
xnor U7053 (N_7053,N_5056,N_4546);
nor U7054 (N_7054,N_5302,N_4832);
or U7055 (N_7055,N_5618,N_4494);
and U7056 (N_7056,N_4357,N_5356);
nor U7057 (N_7057,N_4975,N_4504);
and U7058 (N_7058,N_5660,N_5947);
and U7059 (N_7059,N_5042,N_5544);
xor U7060 (N_7060,N_5691,N_5484);
nand U7061 (N_7061,N_4895,N_5176);
xor U7062 (N_7062,N_4256,N_5451);
or U7063 (N_7063,N_5475,N_4048);
or U7064 (N_7064,N_4163,N_4034);
nor U7065 (N_7065,N_4184,N_5220);
nor U7066 (N_7066,N_5277,N_4825);
nand U7067 (N_7067,N_5790,N_4661);
xnor U7068 (N_7068,N_4429,N_5288);
nand U7069 (N_7069,N_4455,N_5383);
nand U7070 (N_7070,N_5759,N_4634);
and U7071 (N_7071,N_4324,N_4916);
nand U7072 (N_7072,N_5318,N_4898);
nor U7073 (N_7073,N_4279,N_4050);
nor U7074 (N_7074,N_4307,N_5544);
nor U7075 (N_7075,N_4537,N_5588);
or U7076 (N_7076,N_4730,N_4686);
xor U7077 (N_7077,N_5750,N_4232);
or U7078 (N_7078,N_4001,N_4325);
or U7079 (N_7079,N_5908,N_5066);
xor U7080 (N_7080,N_5588,N_4645);
nand U7081 (N_7081,N_4739,N_4678);
nor U7082 (N_7082,N_5644,N_4959);
or U7083 (N_7083,N_5810,N_4609);
or U7084 (N_7084,N_4945,N_5192);
nor U7085 (N_7085,N_4515,N_4348);
or U7086 (N_7086,N_5872,N_4775);
nor U7087 (N_7087,N_4309,N_5730);
xor U7088 (N_7088,N_4067,N_5419);
nor U7089 (N_7089,N_5876,N_4373);
xor U7090 (N_7090,N_4961,N_5587);
and U7091 (N_7091,N_5853,N_5660);
or U7092 (N_7092,N_5665,N_5930);
xnor U7093 (N_7093,N_5011,N_5119);
nand U7094 (N_7094,N_5373,N_5219);
and U7095 (N_7095,N_4035,N_4188);
nand U7096 (N_7096,N_4891,N_4515);
nand U7097 (N_7097,N_5396,N_4019);
nand U7098 (N_7098,N_5231,N_4901);
xor U7099 (N_7099,N_4299,N_5569);
nand U7100 (N_7100,N_5707,N_5984);
xor U7101 (N_7101,N_4363,N_5465);
xor U7102 (N_7102,N_4470,N_4369);
nand U7103 (N_7103,N_4755,N_5062);
and U7104 (N_7104,N_4433,N_5304);
and U7105 (N_7105,N_4289,N_4413);
nor U7106 (N_7106,N_4923,N_4039);
nor U7107 (N_7107,N_5104,N_4841);
nor U7108 (N_7108,N_4628,N_4433);
nand U7109 (N_7109,N_5403,N_5577);
or U7110 (N_7110,N_4970,N_5575);
nand U7111 (N_7111,N_4147,N_5631);
xnor U7112 (N_7112,N_4057,N_5175);
and U7113 (N_7113,N_5430,N_4321);
or U7114 (N_7114,N_4873,N_4875);
nor U7115 (N_7115,N_5354,N_5957);
nand U7116 (N_7116,N_5022,N_5442);
nor U7117 (N_7117,N_5332,N_5324);
nor U7118 (N_7118,N_5543,N_4246);
nor U7119 (N_7119,N_5119,N_5591);
or U7120 (N_7120,N_4350,N_5523);
nand U7121 (N_7121,N_4117,N_4631);
or U7122 (N_7122,N_5818,N_5729);
or U7123 (N_7123,N_4890,N_4907);
or U7124 (N_7124,N_5724,N_5715);
nand U7125 (N_7125,N_5089,N_5357);
nor U7126 (N_7126,N_4737,N_5798);
xnor U7127 (N_7127,N_5759,N_4703);
nor U7128 (N_7128,N_4599,N_5855);
xnor U7129 (N_7129,N_4914,N_4246);
xnor U7130 (N_7130,N_4630,N_4748);
nor U7131 (N_7131,N_5782,N_5295);
and U7132 (N_7132,N_5734,N_5559);
and U7133 (N_7133,N_5890,N_4421);
nor U7134 (N_7134,N_4975,N_5018);
nor U7135 (N_7135,N_4107,N_5037);
nand U7136 (N_7136,N_5146,N_5251);
and U7137 (N_7137,N_5753,N_5910);
nand U7138 (N_7138,N_4686,N_4030);
nand U7139 (N_7139,N_5557,N_5290);
nand U7140 (N_7140,N_4314,N_4303);
and U7141 (N_7141,N_5422,N_4396);
nand U7142 (N_7142,N_5996,N_5755);
xor U7143 (N_7143,N_5779,N_4594);
and U7144 (N_7144,N_4033,N_5157);
or U7145 (N_7145,N_5537,N_5943);
nor U7146 (N_7146,N_5080,N_5712);
and U7147 (N_7147,N_5075,N_4880);
nor U7148 (N_7148,N_5765,N_5256);
nor U7149 (N_7149,N_4418,N_5516);
and U7150 (N_7150,N_5961,N_5742);
nand U7151 (N_7151,N_4996,N_5494);
nand U7152 (N_7152,N_5568,N_5218);
and U7153 (N_7153,N_4550,N_5930);
or U7154 (N_7154,N_5626,N_5393);
or U7155 (N_7155,N_4436,N_5868);
nand U7156 (N_7156,N_5964,N_5757);
and U7157 (N_7157,N_5335,N_4024);
xor U7158 (N_7158,N_5465,N_5174);
or U7159 (N_7159,N_4624,N_5690);
xor U7160 (N_7160,N_5678,N_4294);
nand U7161 (N_7161,N_5155,N_5510);
nor U7162 (N_7162,N_5265,N_4992);
nor U7163 (N_7163,N_5594,N_4376);
xnor U7164 (N_7164,N_4692,N_4125);
xnor U7165 (N_7165,N_5148,N_4725);
and U7166 (N_7166,N_5569,N_5886);
xnor U7167 (N_7167,N_5526,N_5513);
nor U7168 (N_7168,N_4392,N_5843);
or U7169 (N_7169,N_5989,N_4076);
xnor U7170 (N_7170,N_4536,N_5520);
xor U7171 (N_7171,N_4229,N_4658);
or U7172 (N_7172,N_5170,N_4928);
and U7173 (N_7173,N_4394,N_5497);
or U7174 (N_7174,N_4090,N_4277);
or U7175 (N_7175,N_5130,N_5767);
and U7176 (N_7176,N_4062,N_5880);
nand U7177 (N_7177,N_5453,N_4001);
or U7178 (N_7178,N_4566,N_4265);
nor U7179 (N_7179,N_4739,N_4851);
or U7180 (N_7180,N_5742,N_4329);
nor U7181 (N_7181,N_4184,N_5655);
or U7182 (N_7182,N_5737,N_5490);
xor U7183 (N_7183,N_4246,N_4188);
nor U7184 (N_7184,N_4768,N_5832);
nor U7185 (N_7185,N_4233,N_5819);
and U7186 (N_7186,N_5616,N_5015);
xnor U7187 (N_7187,N_4683,N_5182);
nor U7188 (N_7188,N_4799,N_4820);
and U7189 (N_7189,N_4596,N_4853);
nand U7190 (N_7190,N_5523,N_5233);
nor U7191 (N_7191,N_5620,N_4161);
and U7192 (N_7192,N_5805,N_4866);
and U7193 (N_7193,N_4578,N_5888);
and U7194 (N_7194,N_5945,N_5604);
xnor U7195 (N_7195,N_4340,N_4242);
nor U7196 (N_7196,N_4054,N_5101);
nand U7197 (N_7197,N_5696,N_5572);
and U7198 (N_7198,N_5269,N_5663);
nand U7199 (N_7199,N_5876,N_5889);
xnor U7200 (N_7200,N_4047,N_4895);
and U7201 (N_7201,N_4367,N_4149);
or U7202 (N_7202,N_5291,N_4002);
nand U7203 (N_7203,N_5017,N_5061);
nand U7204 (N_7204,N_5906,N_5195);
nor U7205 (N_7205,N_4380,N_4443);
nand U7206 (N_7206,N_4254,N_4601);
or U7207 (N_7207,N_4558,N_5676);
nand U7208 (N_7208,N_5285,N_5093);
nor U7209 (N_7209,N_5313,N_4796);
nor U7210 (N_7210,N_5779,N_5732);
nand U7211 (N_7211,N_4509,N_5571);
xnor U7212 (N_7212,N_5630,N_5342);
nor U7213 (N_7213,N_4211,N_5592);
nand U7214 (N_7214,N_4850,N_5734);
xnor U7215 (N_7215,N_5702,N_5558);
or U7216 (N_7216,N_4532,N_4366);
and U7217 (N_7217,N_5927,N_5683);
and U7218 (N_7218,N_4840,N_4360);
and U7219 (N_7219,N_4707,N_4757);
or U7220 (N_7220,N_5046,N_5737);
or U7221 (N_7221,N_5740,N_5066);
and U7222 (N_7222,N_4970,N_5117);
nand U7223 (N_7223,N_4464,N_5010);
or U7224 (N_7224,N_5699,N_4108);
nor U7225 (N_7225,N_4923,N_4209);
nand U7226 (N_7226,N_5340,N_5561);
nand U7227 (N_7227,N_4150,N_5887);
xnor U7228 (N_7228,N_4274,N_5310);
or U7229 (N_7229,N_5628,N_4949);
or U7230 (N_7230,N_4981,N_5220);
nand U7231 (N_7231,N_4557,N_4781);
xor U7232 (N_7232,N_4892,N_5085);
nor U7233 (N_7233,N_4004,N_4616);
or U7234 (N_7234,N_5406,N_4636);
nor U7235 (N_7235,N_5401,N_4738);
or U7236 (N_7236,N_4851,N_4686);
or U7237 (N_7237,N_5103,N_5881);
or U7238 (N_7238,N_5179,N_5037);
and U7239 (N_7239,N_5073,N_4223);
nor U7240 (N_7240,N_5247,N_5761);
or U7241 (N_7241,N_4046,N_4816);
xnor U7242 (N_7242,N_5642,N_4583);
or U7243 (N_7243,N_5812,N_4859);
xnor U7244 (N_7244,N_4535,N_5986);
and U7245 (N_7245,N_4772,N_4484);
and U7246 (N_7246,N_4674,N_4261);
or U7247 (N_7247,N_5562,N_4993);
or U7248 (N_7248,N_4278,N_5882);
and U7249 (N_7249,N_4317,N_5873);
and U7250 (N_7250,N_5076,N_4081);
nand U7251 (N_7251,N_4735,N_4334);
nor U7252 (N_7252,N_4329,N_5227);
nor U7253 (N_7253,N_5870,N_4723);
and U7254 (N_7254,N_5171,N_4388);
xnor U7255 (N_7255,N_5614,N_5021);
and U7256 (N_7256,N_4849,N_5663);
or U7257 (N_7257,N_4639,N_5149);
nor U7258 (N_7258,N_4316,N_4476);
or U7259 (N_7259,N_5640,N_5528);
xnor U7260 (N_7260,N_5568,N_5619);
and U7261 (N_7261,N_4551,N_5838);
or U7262 (N_7262,N_5753,N_4983);
nand U7263 (N_7263,N_4322,N_5144);
and U7264 (N_7264,N_5678,N_5194);
and U7265 (N_7265,N_4244,N_4994);
nor U7266 (N_7266,N_5231,N_5452);
nor U7267 (N_7267,N_4923,N_5470);
and U7268 (N_7268,N_5970,N_4370);
nor U7269 (N_7269,N_4287,N_4149);
xor U7270 (N_7270,N_5787,N_5023);
nand U7271 (N_7271,N_4572,N_4228);
nor U7272 (N_7272,N_4052,N_5805);
nand U7273 (N_7273,N_4302,N_5647);
or U7274 (N_7274,N_4733,N_5875);
nor U7275 (N_7275,N_5552,N_4517);
and U7276 (N_7276,N_4833,N_5967);
nor U7277 (N_7277,N_5330,N_5242);
nand U7278 (N_7278,N_5872,N_5448);
or U7279 (N_7279,N_4785,N_5833);
xnor U7280 (N_7280,N_5264,N_4929);
xnor U7281 (N_7281,N_5819,N_4393);
nor U7282 (N_7282,N_4871,N_4765);
or U7283 (N_7283,N_5097,N_4173);
xnor U7284 (N_7284,N_5586,N_4137);
xnor U7285 (N_7285,N_4712,N_4436);
and U7286 (N_7286,N_5954,N_5081);
or U7287 (N_7287,N_4467,N_4962);
or U7288 (N_7288,N_4567,N_4723);
or U7289 (N_7289,N_4858,N_5319);
or U7290 (N_7290,N_4732,N_4641);
nor U7291 (N_7291,N_5230,N_4240);
nor U7292 (N_7292,N_4210,N_4356);
nor U7293 (N_7293,N_5918,N_4867);
xnor U7294 (N_7294,N_5760,N_5639);
xnor U7295 (N_7295,N_4118,N_4480);
and U7296 (N_7296,N_4557,N_4075);
nor U7297 (N_7297,N_4917,N_4280);
and U7298 (N_7298,N_4797,N_4922);
and U7299 (N_7299,N_4233,N_4092);
and U7300 (N_7300,N_4214,N_5353);
nor U7301 (N_7301,N_4267,N_5633);
and U7302 (N_7302,N_4050,N_4441);
xnor U7303 (N_7303,N_4156,N_5600);
or U7304 (N_7304,N_5608,N_5246);
xnor U7305 (N_7305,N_4735,N_4375);
or U7306 (N_7306,N_5765,N_5779);
and U7307 (N_7307,N_5504,N_5220);
and U7308 (N_7308,N_4566,N_4814);
nand U7309 (N_7309,N_5259,N_4755);
nor U7310 (N_7310,N_4035,N_5127);
nand U7311 (N_7311,N_5287,N_4537);
and U7312 (N_7312,N_4400,N_4456);
and U7313 (N_7313,N_4466,N_4438);
nor U7314 (N_7314,N_4986,N_5951);
or U7315 (N_7315,N_5574,N_5994);
xnor U7316 (N_7316,N_5612,N_4816);
nand U7317 (N_7317,N_4958,N_4352);
nand U7318 (N_7318,N_4165,N_4679);
nor U7319 (N_7319,N_4218,N_4704);
nand U7320 (N_7320,N_4042,N_5516);
nor U7321 (N_7321,N_4115,N_4167);
or U7322 (N_7322,N_5224,N_4991);
nor U7323 (N_7323,N_5918,N_5240);
or U7324 (N_7324,N_4362,N_5202);
and U7325 (N_7325,N_4460,N_4691);
or U7326 (N_7326,N_5497,N_4361);
xnor U7327 (N_7327,N_5345,N_4235);
nand U7328 (N_7328,N_5246,N_4601);
or U7329 (N_7329,N_5668,N_5777);
nor U7330 (N_7330,N_5734,N_5971);
xnor U7331 (N_7331,N_5240,N_4232);
nand U7332 (N_7332,N_5000,N_4548);
or U7333 (N_7333,N_4451,N_4020);
nand U7334 (N_7334,N_5943,N_4659);
nor U7335 (N_7335,N_5057,N_5294);
nand U7336 (N_7336,N_5701,N_4934);
or U7337 (N_7337,N_4460,N_4188);
or U7338 (N_7338,N_5994,N_4947);
and U7339 (N_7339,N_5849,N_4559);
or U7340 (N_7340,N_5987,N_4981);
nand U7341 (N_7341,N_4838,N_4928);
nand U7342 (N_7342,N_5339,N_4394);
nand U7343 (N_7343,N_4608,N_4690);
nor U7344 (N_7344,N_5886,N_5783);
or U7345 (N_7345,N_5017,N_5026);
xor U7346 (N_7346,N_5534,N_5600);
or U7347 (N_7347,N_5555,N_4819);
nor U7348 (N_7348,N_4754,N_5542);
and U7349 (N_7349,N_4212,N_4607);
or U7350 (N_7350,N_4714,N_4060);
and U7351 (N_7351,N_4835,N_4318);
nor U7352 (N_7352,N_4394,N_5658);
nor U7353 (N_7353,N_5890,N_4118);
nor U7354 (N_7354,N_5719,N_5763);
nor U7355 (N_7355,N_5994,N_5645);
or U7356 (N_7356,N_4904,N_5822);
or U7357 (N_7357,N_5294,N_4829);
nand U7358 (N_7358,N_5258,N_4708);
and U7359 (N_7359,N_4068,N_5777);
xor U7360 (N_7360,N_5009,N_5830);
and U7361 (N_7361,N_4646,N_4340);
or U7362 (N_7362,N_5118,N_4999);
nor U7363 (N_7363,N_4168,N_5868);
xnor U7364 (N_7364,N_5429,N_4772);
nor U7365 (N_7365,N_4650,N_4299);
nor U7366 (N_7366,N_4497,N_5586);
nand U7367 (N_7367,N_4063,N_5640);
nand U7368 (N_7368,N_5662,N_5359);
or U7369 (N_7369,N_5996,N_5690);
xor U7370 (N_7370,N_4280,N_4154);
and U7371 (N_7371,N_4602,N_5760);
nand U7372 (N_7372,N_4018,N_5089);
nor U7373 (N_7373,N_4265,N_4595);
xor U7374 (N_7374,N_4811,N_4064);
and U7375 (N_7375,N_5723,N_4625);
nand U7376 (N_7376,N_5262,N_4766);
or U7377 (N_7377,N_5133,N_5151);
nand U7378 (N_7378,N_5580,N_5916);
nor U7379 (N_7379,N_4952,N_5157);
or U7380 (N_7380,N_4465,N_5216);
or U7381 (N_7381,N_5421,N_5733);
or U7382 (N_7382,N_5253,N_4377);
or U7383 (N_7383,N_5299,N_5522);
xor U7384 (N_7384,N_4140,N_5028);
and U7385 (N_7385,N_4234,N_4105);
or U7386 (N_7386,N_5475,N_5650);
or U7387 (N_7387,N_5779,N_5609);
or U7388 (N_7388,N_4163,N_5666);
or U7389 (N_7389,N_5706,N_4792);
nand U7390 (N_7390,N_4317,N_4368);
nor U7391 (N_7391,N_4999,N_4064);
nor U7392 (N_7392,N_4451,N_5491);
nand U7393 (N_7393,N_4529,N_4762);
nand U7394 (N_7394,N_5522,N_5880);
nand U7395 (N_7395,N_5976,N_5326);
and U7396 (N_7396,N_5907,N_4463);
nor U7397 (N_7397,N_5817,N_5331);
and U7398 (N_7398,N_4696,N_5982);
xnor U7399 (N_7399,N_4937,N_4262);
nand U7400 (N_7400,N_5938,N_4883);
nor U7401 (N_7401,N_5997,N_5195);
nand U7402 (N_7402,N_5557,N_4449);
and U7403 (N_7403,N_4669,N_4833);
nand U7404 (N_7404,N_5042,N_4586);
and U7405 (N_7405,N_4754,N_5952);
and U7406 (N_7406,N_4117,N_5780);
xor U7407 (N_7407,N_5487,N_5896);
xor U7408 (N_7408,N_5195,N_5308);
or U7409 (N_7409,N_4577,N_4191);
nor U7410 (N_7410,N_5718,N_5807);
nor U7411 (N_7411,N_4642,N_4274);
nor U7412 (N_7412,N_5483,N_5330);
nand U7413 (N_7413,N_5875,N_4606);
or U7414 (N_7414,N_4245,N_5569);
or U7415 (N_7415,N_4636,N_4510);
nor U7416 (N_7416,N_4579,N_5008);
xnor U7417 (N_7417,N_5201,N_5250);
nand U7418 (N_7418,N_4065,N_4384);
or U7419 (N_7419,N_5846,N_4270);
nand U7420 (N_7420,N_5576,N_4041);
xnor U7421 (N_7421,N_4580,N_5556);
or U7422 (N_7422,N_5485,N_4595);
xor U7423 (N_7423,N_5817,N_4177);
nand U7424 (N_7424,N_4992,N_4074);
xnor U7425 (N_7425,N_4830,N_5213);
nor U7426 (N_7426,N_4341,N_5420);
nor U7427 (N_7427,N_5348,N_4426);
nor U7428 (N_7428,N_5217,N_4556);
xor U7429 (N_7429,N_4569,N_4566);
and U7430 (N_7430,N_4141,N_4102);
nand U7431 (N_7431,N_4783,N_4309);
xor U7432 (N_7432,N_4732,N_5872);
or U7433 (N_7433,N_5058,N_4906);
and U7434 (N_7434,N_5956,N_5569);
and U7435 (N_7435,N_5686,N_5160);
and U7436 (N_7436,N_4710,N_4983);
nand U7437 (N_7437,N_5898,N_4584);
nand U7438 (N_7438,N_4773,N_4543);
or U7439 (N_7439,N_5040,N_5037);
xnor U7440 (N_7440,N_4916,N_4954);
and U7441 (N_7441,N_5129,N_5840);
nor U7442 (N_7442,N_4304,N_4584);
or U7443 (N_7443,N_4528,N_5402);
xnor U7444 (N_7444,N_4601,N_4524);
or U7445 (N_7445,N_4837,N_5076);
nor U7446 (N_7446,N_5628,N_4665);
xnor U7447 (N_7447,N_4671,N_4180);
and U7448 (N_7448,N_5111,N_5221);
xnor U7449 (N_7449,N_5312,N_5074);
or U7450 (N_7450,N_4767,N_4977);
nor U7451 (N_7451,N_4055,N_4535);
nand U7452 (N_7452,N_5436,N_5323);
xor U7453 (N_7453,N_4356,N_4824);
and U7454 (N_7454,N_4130,N_4989);
xnor U7455 (N_7455,N_4329,N_5928);
nand U7456 (N_7456,N_4353,N_4996);
and U7457 (N_7457,N_5255,N_4409);
or U7458 (N_7458,N_4433,N_4662);
or U7459 (N_7459,N_5948,N_4057);
xnor U7460 (N_7460,N_4842,N_4542);
or U7461 (N_7461,N_4672,N_5537);
nand U7462 (N_7462,N_5467,N_5052);
xor U7463 (N_7463,N_5858,N_4391);
and U7464 (N_7464,N_4744,N_5551);
xnor U7465 (N_7465,N_5326,N_5403);
and U7466 (N_7466,N_4980,N_4156);
or U7467 (N_7467,N_5994,N_4049);
nor U7468 (N_7468,N_4534,N_4049);
xnor U7469 (N_7469,N_5214,N_5593);
nand U7470 (N_7470,N_4312,N_5005);
or U7471 (N_7471,N_5466,N_5035);
nand U7472 (N_7472,N_4297,N_5554);
and U7473 (N_7473,N_5689,N_4661);
nor U7474 (N_7474,N_5699,N_4540);
nand U7475 (N_7475,N_4295,N_5482);
nand U7476 (N_7476,N_5818,N_4821);
or U7477 (N_7477,N_5721,N_4885);
nor U7478 (N_7478,N_5870,N_4138);
nor U7479 (N_7479,N_4047,N_4814);
or U7480 (N_7480,N_4098,N_5439);
xor U7481 (N_7481,N_4357,N_5979);
nand U7482 (N_7482,N_4753,N_5859);
nor U7483 (N_7483,N_5440,N_5627);
xor U7484 (N_7484,N_4933,N_4154);
and U7485 (N_7485,N_5828,N_5356);
or U7486 (N_7486,N_4798,N_4406);
xnor U7487 (N_7487,N_4845,N_4815);
and U7488 (N_7488,N_4511,N_5637);
or U7489 (N_7489,N_4126,N_4349);
xnor U7490 (N_7490,N_5585,N_4735);
or U7491 (N_7491,N_4625,N_4274);
nand U7492 (N_7492,N_5655,N_5843);
nor U7493 (N_7493,N_5213,N_4543);
nand U7494 (N_7494,N_4840,N_5024);
nor U7495 (N_7495,N_4973,N_5611);
xnor U7496 (N_7496,N_5862,N_5428);
or U7497 (N_7497,N_4851,N_4810);
xor U7498 (N_7498,N_4533,N_4575);
xnor U7499 (N_7499,N_5430,N_4847);
xor U7500 (N_7500,N_4151,N_4503);
or U7501 (N_7501,N_4146,N_5911);
xor U7502 (N_7502,N_5401,N_5440);
xor U7503 (N_7503,N_4505,N_4628);
xnor U7504 (N_7504,N_4406,N_5597);
and U7505 (N_7505,N_5397,N_4062);
and U7506 (N_7506,N_4548,N_5818);
and U7507 (N_7507,N_4338,N_4688);
or U7508 (N_7508,N_5490,N_5356);
xnor U7509 (N_7509,N_4291,N_5105);
nand U7510 (N_7510,N_4634,N_4033);
xor U7511 (N_7511,N_5218,N_4482);
xnor U7512 (N_7512,N_4918,N_4668);
nand U7513 (N_7513,N_5482,N_4464);
xnor U7514 (N_7514,N_4812,N_5164);
or U7515 (N_7515,N_4648,N_5930);
and U7516 (N_7516,N_4799,N_5903);
nand U7517 (N_7517,N_5638,N_4201);
and U7518 (N_7518,N_4042,N_5329);
xor U7519 (N_7519,N_4199,N_4373);
xor U7520 (N_7520,N_5003,N_5109);
and U7521 (N_7521,N_4313,N_5122);
nand U7522 (N_7522,N_4002,N_5774);
and U7523 (N_7523,N_5195,N_4466);
or U7524 (N_7524,N_5298,N_5609);
or U7525 (N_7525,N_4263,N_4855);
nor U7526 (N_7526,N_4894,N_5255);
or U7527 (N_7527,N_4257,N_4041);
xnor U7528 (N_7528,N_4230,N_5338);
xor U7529 (N_7529,N_5838,N_4064);
nor U7530 (N_7530,N_5115,N_5759);
xor U7531 (N_7531,N_4023,N_5888);
nand U7532 (N_7532,N_5433,N_4569);
nand U7533 (N_7533,N_4420,N_5651);
and U7534 (N_7534,N_5639,N_5202);
and U7535 (N_7535,N_5262,N_5908);
and U7536 (N_7536,N_5292,N_5141);
nor U7537 (N_7537,N_4822,N_4747);
nand U7538 (N_7538,N_5218,N_5494);
or U7539 (N_7539,N_5727,N_4716);
or U7540 (N_7540,N_5879,N_4723);
nand U7541 (N_7541,N_4945,N_4836);
nor U7542 (N_7542,N_5365,N_5526);
or U7543 (N_7543,N_5483,N_5305);
nor U7544 (N_7544,N_5334,N_4233);
nand U7545 (N_7545,N_5226,N_4894);
nand U7546 (N_7546,N_5980,N_5060);
or U7547 (N_7547,N_4147,N_4668);
xnor U7548 (N_7548,N_4907,N_5070);
or U7549 (N_7549,N_4868,N_5689);
nand U7550 (N_7550,N_5824,N_5678);
and U7551 (N_7551,N_4109,N_4634);
nor U7552 (N_7552,N_4229,N_5290);
xor U7553 (N_7553,N_5741,N_4251);
and U7554 (N_7554,N_4526,N_4480);
nand U7555 (N_7555,N_5916,N_5185);
nor U7556 (N_7556,N_4578,N_5143);
xor U7557 (N_7557,N_4467,N_5278);
nor U7558 (N_7558,N_5900,N_5106);
nand U7559 (N_7559,N_4785,N_4412);
nand U7560 (N_7560,N_5168,N_4654);
xor U7561 (N_7561,N_5047,N_4519);
xnor U7562 (N_7562,N_4291,N_4509);
xnor U7563 (N_7563,N_5663,N_5041);
xnor U7564 (N_7564,N_4137,N_5727);
xor U7565 (N_7565,N_5174,N_4016);
nor U7566 (N_7566,N_4208,N_5791);
or U7567 (N_7567,N_5136,N_5039);
xor U7568 (N_7568,N_4250,N_5254);
nor U7569 (N_7569,N_5477,N_5629);
xnor U7570 (N_7570,N_4868,N_5824);
xor U7571 (N_7571,N_4114,N_5556);
or U7572 (N_7572,N_4161,N_5669);
or U7573 (N_7573,N_5419,N_4664);
nand U7574 (N_7574,N_5571,N_5301);
xor U7575 (N_7575,N_5487,N_5454);
xnor U7576 (N_7576,N_5613,N_4183);
nor U7577 (N_7577,N_5564,N_5215);
or U7578 (N_7578,N_5273,N_4082);
nor U7579 (N_7579,N_4808,N_5721);
nand U7580 (N_7580,N_4607,N_4170);
or U7581 (N_7581,N_4759,N_5663);
and U7582 (N_7582,N_5727,N_5264);
xnor U7583 (N_7583,N_5828,N_4427);
and U7584 (N_7584,N_5428,N_4968);
and U7585 (N_7585,N_4021,N_5005);
nor U7586 (N_7586,N_5758,N_4149);
xor U7587 (N_7587,N_5505,N_5891);
and U7588 (N_7588,N_4937,N_4585);
and U7589 (N_7589,N_5416,N_4619);
and U7590 (N_7590,N_5937,N_4988);
and U7591 (N_7591,N_4972,N_5792);
nor U7592 (N_7592,N_4142,N_4051);
xnor U7593 (N_7593,N_5647,N_4948);
nand U7594 (N_7594,N_4123,N_4607);
nor U7595 (N_7595,N_5322,N_5287);
and U7596 (N_7596,N_4550,N_4887);
and U7597 (N_7597,N_4610,N_5653);
xnor U7598 (N_7598,N_5330,N_4388);
or U7599 (N_7599,N_5498,N_5454);
and U7600 (N_7600,N_5642,N_5537);
xor U7601 (N_7601,N_5548,N_4220);
nor U7602 (N_7602,N_5705,N_4409);
xnor U7603 (N_7603,N_4152,N_4558);
nor U7604 (N_7604,N_5960,N_5151);
xor U7605 (N_7605,N_5111,N_4726);
nand U7606 (N_7606,N_5271,N_5845);
xor U7607 (N_7607,N_5320,N_4911);
xnor U7608 (N_7608,N_4729,N_5546);
and U7609 (N_7609,N_4622,N_5850);
and U7610 (N_7610,N_4128,N_4455);
nand U7611 (N_7611,N_5472,N_5099);
or U7612 (N_7612,N_5023,N_5045);
and U7613 (N_7613,N_4103,N_5920);
nor U7614 (N_7614,N_5417,N_4467);
nand U7615 (N_7615,N_4915,N_4181);
and U7616 (N_7616,N_4153,N_4085);
nand U7617 (N_7617,N_4776,N_4401);
nor U7618 (N_7618,N_4930,N_5304);
and U7619 (N_7619,N_5366,N_5920);
nor U7620 (N_7620,N_4757,N_4175);
and U7621 (N_7621,N_4901,N_4110);
nand U7622 (N_7622,N_5420,N_5757);
nor U7623 (N_7623,N_5532,N_5874);
nand U7624 (N_7624,N_5397,N_4465);
or U7625 (N_7625,N_5409,N_4660);
nor U7626 (N_7626,N_5142,N_4556);
and U7627 (N_7627,N_4020,N_4370);
or U7628 (N_7628,N_4837,N_5353);
and U7629 (N_7629,N_5439,N_5437);
xor U7630 (N_7630,N_4098,N_4944);
nand U7631 (N_7631,N_5173,N_4851);
or U7632 (N_7632,N_5367,N_4131);
or U7633 (N_7633,N_5230,N_5048);
xnor U7634 (N_7634,N_4289,N_4075);
xnor U7635 (N_7635,N_4199,N_5000);
nand U7636 (N_7636,N_5738,N_4106);
or U7637 (N_7637,N_4920,N_4184);
nand U7638 (N_7638,N_5842,N_5538);
or U7639 (N_7639,N_4734,N_5526);
or U7640 (N_7640,N_5981,N_4248);
nor U7641 (N_7641,N_5305,N_5633);
nor U7642 (N_7642,N_5900,N_4252);
nor U7643 (N_7643,N_5353,N_4015);
nand U7644 (N_7644,N_4901,N_5355);
nand U7645 (N_7645,N_5472,N_5249);
xor U7646 (N_7646,N_4514,N_4311);
and U7647 (N_7647,N_5569,N_5481);
or U7648 (N_7648,N_5872,N_5020);
nand U7649 (N_7649,N_4307,N_4562);
xor U7650 (N_7650,N_5152,N_5839);
or U7651 (N_7651,N_4204,N_4293);
xor U7652 (N_7652,N_5434,N_5684);
xnor U7653 (N_7653,N_4547,N_4166);
or U7654 (N_7654,N_5954,N_4975);
and U7655 (N_7655,N_4874,N_5509);
nor U7656 (N_7656,N_5841,N_5286);
nand U7657 (N_7657,N_5870,N_4557);
nor U7658 (N_7658,N_4130,N_5088);
and U7659 (N_7659,N_4098,N_5655);
and U7660 (N_7660,N_4714,N_5372);
nor U7661 (N_7661,N_4440,N_5399);
or U7662 (N_7662,N_4824,N_5916);
nor U7663 (N_7663,N_5493,N_5479);
nand U7664 (N_7664,N_4874,N_5304);
nand U7665 (N_7665,N_5987,N_5017);
nor U7666 (N_7666,N_5377,N_5307);
and U7667 (N_7667,N_5149,N_4666);
nand U7668 (N_7668,N_4565,N_5426);
and U7669 (N_7669,N_4948,N_4189);
nand U7670 (N_7670,N_4915,N_4795);
nor U7671 (N_7671,N_5152,N_5465);
or U7672 (N_7672,N_5665,N_4468);
and U7673 (N_7673,N_4710,N_4868);
nand U7674 (N_7674,N_4721,N_5189);
nand U7675 (N_7675,N_4021,N_5017);
nand U7676 (N_7676,N_5199,N_4163);
and U7677 (N_7677,N_5070,N_5882);
nor U7678 (N_7678,N_5600,N_5652);
nor U7679 (N_7679,N_5353,N_4039);
nand U7680 (N_7680,N_5114,N_5696);
nor U7681 (N_7681,N_4659,N_5312);
nand U7682 (N_7682,N_5830,N_5488);
and U7683 (N_7683,N_4196,N_4994);
and U7684 (N_7684,N_5955,N_4295);
nor U7685 (N_7685,N_4979,N_5037);
nand U7686 (N_7686,N_4081,N_5503);
and U7687 (N_7687,N_5709,N_5116);
nor U7688 (N_7688,N_5194,N_4780);
nand U7689 (N_7689,N_5066,N_4390);
and U7690 (N_7690,N_4638,N_5295);
nor U7691 (N_7691,N_5885,N_5210);
xor U7692 (N_7692,N_5358,N_5045);
and U7693 (N_7693,N_5911,N_5450);
xnor U7694 (N_7694,N_4406,N_5517);
or U7695 (N_7695,N_4866,N_4692);
nor U7696 (N_7696,N_4236,N_4550);
or U7697 (N_7697,N_5487,N_4503);
and U7698 (N_7698,N_4738,N_4744);
or U7699 (N_7699,N_5367,N_5318);
nor U7700 (N_7700,N_5230,N_4074);
xnor U7701 (N_7701,N_5473,N_4213);
or U7702 (N_7702,N_5577,N_5098);
nor U7703 (N_7703,N_4735,N_5713);
nor U7704 (N_7704,N_4988,N_4499);
nand U7705 (N_7705,N_4183,N_4407);
nor U7706 (N_7706,N_4215,N_5166);
or U7707 (N_7707,N_4223,N_5763);
or U7708 (N_7708,N_4330,N_5439);
nand U7709 (N_7709,N_5541,N_5093);
xnor U7710 (N_7710,N_4241,N_5186);
nor U7711 (N_7711,N_4019,N_4976);
nor U7712 (N_7712,N_5071,N_4404);
and U7713 (N_7713,N_4775,N_5581);
and U7714 (N_7714,N_4015,N_4029);
or U7715 (N_7715,N_5242,N_4032);
nor U7716 (N_7716,N_4560,N_4063);
nand U7717 (N_7717,N_4075,N_4711);
xnor U7718 (N_7718,N_4871,N_4669);
nor U7719 (N_7719,N_4538,N_4356);
xnor U7720 (N_7720,N_4149,N_5308);
nor U7721 (N_7721,N_4968,N_5836);
nand U7722 (N_7722,N_5210,N_4687);
or U7723 (N_7723,N_5469,N_5047);
nor U7724 (N_7724,N_4360,N_4764);
nor U7725 (N_7725,N_4705,N_4750);
and U7726 (N_7726,N_4822,N_5902);
nand U7727 (N_7727,N_5350,N_5214);
xor U7728 (N_7728,N_5823,N_4557);
nor U7729 (N_7729,N_4905,N_5412);
xor U7730 (N_7730,N_5090,N_5571);
or U7731 (N_7731,N_5175,N_4539);
nor U7732 (N_7732,N_5579,N_4029);
nand U7733 (N_7733,N_4034,N_4922);
xnor U7734 (N_7734,N_5826,N_5971);
or U7735 (N_7735,N_5134,N_4309);
xnor U7736 (N_7736,N_5604,N_5636);
nor U7737 (N_7737,N_4130,N_5390);
and U7738 (N_7738,N_5357,N_5076);
and U7739 (N_7739,N_5388,N_4368);
xor U7740 (N_7740,N_4530,N_5227);
and U7741 (N_7741,N_4467,N_4830);
or U7742 (N_7742,N_4589,N_4290);
nor U7743 (N_7743,N_4996,N_5678);
xnor U7744 (N_7744,N_5343,N_4199);
nand U7745 (N_7745,N_5826,N_4988);
xnor U7746 (N_7746,N_4168,N_5361);
nor U7747 (N_7747,N_4045,N_4088);
xnor U7748 (N_7748,N_5561,N_5959);
nand U7749 (N_7749,N_5313,N_5828);
nand U7750 (N_7750,N_4288,N_5386);
or U7751 (N_7751,N_4454,N_5407);
xnor U7752 (N_7752,N_5816,N_5198);
nand U7753 (N_7753,N_5840,N_4467);
nand U7754 (N_7754,N_5252,N_5089);
and U7755 (N_7755,N_5392,N_5889);
nand U7756 (N_7756,N_5004,N_5228);
or U7757 (N_7757,N_5594,N_5059);
and U7758 (N_7758,N_4589,N_4289);
nor U7759 (N_7759,N_5097,N_5081);
nand U7760 (N_7760,N_4506,N_4318);
or U7761 (N_7761,N_4677,N_4494);
or U7762 (N_7762,N_5061,N_4084);
xnor U7763 (N_7763,N_5775,N_5357);
xor U7764 (N_7764,N_5738,N_4834);
xor U7765 (N_7765,N_4414,N_4719);
xor U7766 (N_7766,N_4971,N_5745);
and U7767 (N_7767,N_5589,N_5848);
nor U7768 (N_7768,N_5003,N_4557);
nor U7769 (N_7769,N_5634,N_4523);
or U7770 (N_7770,N_5032,N_5449);
and U7771 (N_7771,N_4025,N_5518);
or U7772 (N_7772,N_4451,N_4998);
xor U7773 (N_7773,N_4789,N_4423);
nand U7774 (N_7774,N_5333,N_5282);
xnor U7775 (N_7775,N_4973,N_4693);
and U7776 (N_7776,N_5563,N_4462);
and U7777 (N_7777,N_4805,N_4188);
nor U7778 (N_7778,N_4167,N_4170);
nor U7779 (N_7779,N_5880,N_4336);
xor U7780 (N_7780,N_4708,N_5324);
or U7781 (N_7781,N_5132,N_4056);
nor U7782 (N_7782,N_5790,N_4257);
or U7783 (N_7783,N_4978,N_4346);
or U7784 (N_7784,N_4577,N_5059);
nor U7785 (N_7785,N_5386,N_5499);
nand U7786 (N_7786,N_5621,N_4142);
nor U7787 (N_7787,N_5093,N_5515);
and U7788 (N_7788,N_4363,N_5044);
xor U7789 (N_7789,N_5322,N_4387);
xor U7790 (N_7790,N_5014,N_5332);
or U7791 (N_7791,N_4938,N_4320);
xor U7792 (N_7792,N_4320,N_4458);
or U7793 (N_7793,N_4022,N_5485);
xnor U7794 (N_7794,N_4803,N_4496);
and U7795 (N_7795,N_5479,N_4757);
nor U7796 (N_7796,N_5203,N_5062);
nor U7797 (N_7797,N_5647,N_5869);
nand U7798 (N_7798,N_4716,N_4871);
or U7799 (N_7799,N_4718,N_4213);
and U7800 (N_7800,N_5922,N_5520);
and U7801 (N_7801,N_4342,N_4932);
nor U7802 (N_7802,N_4366,N_4695);
xor U7803 (N_7803,N_5267,N_4517);
and U7804 (N_7804,N_4012,N_4475);
xnor U7805 (N_7805,N_4231,N_5952);
and U7806 (N_7806,N_4327,N_5124);
xor U7807 (N_7807,N_4284,N_5778);
and U7808 (N_7808,N_4186,N_4820);
and U7809 (N_7809,N_4635,N_4142);
xnor U7810 (N_7810,N_4261,N_4270);
xnor U7811 (N_7811,N_4426,N_5702);
xor U7812 (N_7812,N_4578,N_5262);
nor U7813 (N_7813,N_5710,N_5276);
nand U7814 (N_7814,N_5724,N_5266);
nand U7815 (N_7815,N_5539,N_5480);
or U7816 (N_7816,N_4129,N_4907);
nand U7817 (N_7817,N_5975,N_5192);
or U7818 (N_7818,N_4730,N_4189);
nand U7819 (N_7819,N_5604,N_5950);
xor U7820 (N_7820,N_4248,N_4394);
and U7821 (N_7821,N_4880,N_5259);
or U7822 (N_7822,N_4711,N_4823);
and U7823 (N_7823,N_5267,N_5904);
and U7824 (N_7824,N_5424,N_5061);
nand U7825 (N_7825,N_4830,N_4565);
nor U7826 (N_7826,N_4366,N_5705);
nor U7827 (N_7827,N_4655,N_5636);
nor U7828 (N_7828,N_4113,N_5538);
or U7829 (N_7829,N_4914,N_4160);
and U7830 (N_7830,N_5366,N_5865);
nand U7831 (N_7831,N_4833,N_4229);
and U7832 (N_7832,N_5755,N_4059);
or U7833 (N_7833,N_5681,N_4777);
or U7834 (N_7834,N_4761,N_4604);
nor U7835 (N_7835,N_4058,N_5006);
nor U7836 (N_7836,N_5064,N_5065);
xor U7837 (N_7837,N_4964,N_4030);
nor U7838 (N_7838,N_5535,N_5811);
and U7839 (N_7839,N_4050,N_5991);
nand U7840 (N_7840,N_4543,N_4059);
nand U7841 (N_7841,N_4870,N_5627);
and U7842 (N_7842,N_4758,N_4654);
and U7843 (N_7843,N_4576,N_4467);
or U7844 (N_7844,N_5859,N_5221);
xnor U7845 (N_7845,N_5360,N_4821);
xnor U7846 (N_7846,N_4474,N_4343);
xor U7847 (N_7847,N_5899,N_5229);
nor U7848 (N_7848,N_4858,N_4426);
or U7849 (N_7849,N_4855,N_4822);
nand U7850 (N_7850,N_5194,N_5228);
and U7851 (N_7851,N_5626,N_5164);
or U7852 (N_7852,N_5172,N_4834);
nand U7853 (N_7853,N_4524,N_4829);
xnor U7854 (N_7854,N_4529,N_5679);
nand U7855 (N_7855,N_4418,N_4192);
and U7856 (N_7856,N_5087,N_4646);
or U7857 (N_7857,N_4895,N_5318);
or U7858 (N_7858,N_4439,N_4099);
nor U7859 (N_7859,N_5563,N_4942);
and U7860 (N_7860,N_4727,N_4290);
nand U7861 (N_7861,N_5649,N_4278);
and U7862 (N_7862,N_5982,N_4004);
nand U7863 (N_7863,N_5478,N_4647);
nand U7864 (N_7864,N_4396,N_4968);
nor U7865 (N_7865,N_5611,N_5826);
or U7866 (N_7866,N_5933,N_4070);
xor U7867 (N_7867,N_5487,N_4060);
or U7868 (N_7868,N_5275,N_4454);
or U7869 (N_7869,N_4429,N_4376);
nor U7870 (N_7870,N_4940,N_4140);
xnor U7871 (N_7871,N_4683,N_5615);
xor U7872 (N_7872,N_5858,N_5341);
xor U7873 (N_7873,N_5947,N_4173);
nand U7874 (N_7874,N_5400,N_4390);
xnor U7875 (N_7875,N_4168,N_4299);
xnor U7876 (N_7876,N_4606,N_5946);
and U7877 (N_7877,N_5811,N_5965);
xnor U7878 (N_7878,N_4982,N_5273);
and U7879 (N_7879,N_5898,N_4866);
and U7880 (N_7880,N_4888,N_4265);
xor U7881 (N_7881,N_5582,N_4017);
xor U7882 (N_7882,N_5184,N_5346);
nor U7883 (N_7883,N_4651,N_5625);
nand U7884 (N_7884,N_5871,N_4452);
xnor U7885 (N_7885,N_5206,N_5400);
xnor U7886 (N_7886,N_4192,N_5147);
nor U7887 (N_7887,N_5592,N_4457);
xor U7888 (N_7888,N_4131,N_4028);
and U7889 (N_7889,N_4956,N_4553);
nand U7890 (N_7890,N_4643,N_4494);
or U7891 (N_7891,N_4919,N_4242);
xnor U7892 (N_7892,N_5418,N_5479);
and U7893 (N_7893,N_5999,N_5729);
nand U7894 (N_7894,N_5211,N_4888);
xnor U7895 (N_7895,N_5770,N_4383);
or U7896 (N_7896,N_5531,N_4417);
nand U7897 (N_7897,N_4338,N_4751);
nor U7898 (N_7898,N_4372,N_4352);
nor U7899 (N_7899,N_5445,N_5611);
nor U7900 (N_7900,N_5531,N_4242);
or U7901 (N_7901,N_4356,N_4404);
and U7902 (N_7902,N_4827,N_4364);
xnor U7903 (N_7903,N_4595,N_4239);
nand U7904 (N_7904,N_5307,N_5921);
or U7905 (N_7905,N_4648,N_5985);
xnor U7906 (N_7906,N_5233,N_4630);
or U7907 (N_7907,N_5501,N_5568);
nor U7908 (N_7908,N_5257,N_5170);
nand U7909 (N_7909,N_5627,N_5316);
or U7910 (N_7910,N_4555,N_4758);
xor U7911 (N_7911,N_5693,N_5278);
nand U7912 (N_7912,N_5229,N_4285);
and U7913 (N_7913,N_4438,N_4995);
or U7914 (N_7914,N_4408,N_5782);
nand U7915 (N_7915,N_4739,N_4694);
nand U7916 (N_7916,N_5681,N_4226);
and U7917 (N_7917,N_4352,N_5414);
or U7918 (N_7918,N_4245,N_5026);
nor U7919 (N_7919,N_5930,N_4910);
or U7920 (N_7920,N_5909,N_5641);
nand U7921 (N_7921,N_4466,N_5627);
nor U7922 (N_7922,N_5309,N_5489);
and U7923 (N_7923,N_4097,N_4107);
nand U7924 (N_7924,N_4871,N_5183);
or U7925 (N_7925,N_5168,N_5985);
nand U7926 (N_7926,N_5091,N_4174);
or U7927 (N_7927,N_5554,N_4877);
and U7928 (N_7928,N_4972,N_5912);
and U7929 (N_7929,N_5821,N_5119);
and U7930 (N_7930,N_4197,N_5150);
or U7931 (N_7931,N_4045,N_4806);
nand U7932 (N_7932,N_4140,N_5306);
or U7933 (N_7933,N_4950,N_5702);
xnor U7934 (N_7934,N_5140,N_5677);
nand U7935 (N_7935,N_4404,N_5946);
xnor U7936 (N_7936,N_5346,N_5917);
nand U7937 (N_7937,N_5630,N_4165);
and U7938 (N_7938,N_5111,N_5263);
or U7939 (N_7939,N_4418,N_5297);
or U7940 (N_7940,N_4982,N_5616);
nor U7941 (N_7941,N_5420,N_5847);
nand U7942 (N_7942,N_5591,N_4428);
xor U7943 (N_7943,N_5951,N_5148);
xor U7944 (N_7944,N_5842,N_4490);
nor U7945 (N_7945,N_5258,N_4803);
nand U7946 (N_7946,N_4150,N_5552);
and U7947 (N_7947,N_4600,N_4604);
nor U7948 (N_7948,N_5558,N_5105);
xnor U7949 (N_7949,N_5449,N_5787);
xor U7950 (N_7950,N_4882,N_4690);
nand U7951 (N_7951,N_4137,N_4962);
xnor U7952 (N_7952,N_5412,N_5971);
and U7953 (N_7953,N_5694,N_4089);
nor U7954 (N_7954,N_4242,N_5161);
xnor U7955 (N_7955,N_5827,N_4531);
or U7956 (N_7956,N_5187,N_5206);
and U7957 (N_7957,N_5555,N_4466);
nor U7958 (N_7958,N_4289,N_5332);
nor U7959 (N_7959,N_5913,N_4569);
nor U7960 (N_7960,N_4581,N_4101);
or U7961 (N_7961,N_4948,N_5073);
xnor U7962 (N_7962,N_4151,N_5742);
xor U7963 (N_7963,N_5234,N_4653);
and U7964 (N_7964,N_5288,N_5368);
xnor U7965 (N_7965,N_5469,N_4314);
nand U7966 (N_7966,N_4458,N_4797);
xor U7967 (N_7967,N_4838,N_5868);
nor U7968 (N_7968,N_5905,N_4777);
nand U7969 (N_7969,N_5652,N_5746);
nor U7970 (N_7970,N_4011,N_5435);
xnor U7971 (N_7971,N_5942,N_4734);
and U7972 (N_7972,N_4777,N_5281);
nand U7973 (N_7973,N_4566,N_5129);
nor U7974 (N_7974,N_4850,N_5536);
and U7975 (N_7975,N_4819,N_5289);
and U7976 (N_7976,N_5687,N_5849);
nor U7977 (N_7977,N_4136,N_5590);
and U7978 (N_7978,N_5982,N_4497);
nor U7979 (N_7979,N_4257,N_4311);
and U7980 (N_7980,N_5860,N_5306);
and U7981 (N_7981,N_5006,N_4924);
and U7982 (N_7982,N_4838,N_5085);
xor U7983 (N_7983,N_4974,N_4274);
nand U7984 (N_7984,N_4082,N_5388);
or U7985 (N_7985,N_5232,N_4256);
nor U7986 (N_7986,N_4801,N_5037);
nor U7987 (N_7987,N_5539,N_4889);
nor U7988 (N_7988,N_4864,N_5732);
and U7989 (N_7989,N_5553,N_5917);
nand U7990 (N_7990,N_4830,N_5601);
xor U7991 (N_7991,N_5525,N_5791);
and U7992 (N_7992,N_5915,N_4451);
nand U7993 (N_7993,N_4135,N_4142);
xnor U7994 (N_7994,N_4178,N_4684);
xnor U7995 (N_7995,N_4066,N_5998);
or U7996 (N_7996,N_5143,N_4182);
or U7997 (N_7997,N_5427,N_5622);
nand U7998 (N_7998,N_5133,N_5381);
xor U7999 (N_7999,N_4615,N_5710);
or U8000 (N_8000,N_7780,N_7846);
nand U8001 (N_8001,N_7096,N_6988);
nand U8002 (N_8002,N_7759,N_6210);
or U8003 (N_8003,N_6712,N_6923);
nand U8004 (N_8004,N_7136,N_6498);
nor U8005 (N_8005,N_7376,N_7040);
xor U8006 (N_8006,N_7983,N_6907);
or U8007 (N_8007,N_6910,N_7716);
or U8008 (N_8008,N_7927,N_7124);
and U8009 (N_8009,N_6025,N_7169);
nor U8010 (N_8010,N_7192,N_7229);
or U8011 (N_8011,N_6483,N_6062);
xnor U8012 (N_8012,N_6359,N_6790);
xor U8013 (N_8013,N_6200,N_7517);
nand U8014 (N_8014,N_6517,N_7670);
xnor U8015 (N_8015,N_6085,N_6233);
nor U8016 (N_8016,N_7313,N_6129);
nor U8017 (N_8017,N_6920,N_7285);
or U8018 (N_8018,N_7159,N_6100);
xnor U8019 (N_8019,N_7340,N_7348);
nor U8020 (N_8020,N_6348,N_6662);
and U8021 (N_8021,N_7978,N_6575);
or U8022 (N_8022,N_7492,N_7940);
nor U8023 (N_8023,N_6049,N_7583);
and U8024 (N_8024,N_6482,N_7312);
or U8025 (N_8025,N_6061,N_6165);
or U8026 (N_8026,N_7037,N_7370);
xnor U8027 (N_8027,N_7950,N_7710);
xor U8028 (N_8028,N_6340,N_6629);
and U8029 (N_8029,N_7178,N_7156);
nand U8030 (N_8030,N_7976,N_6029);
nand U8031 (N_8031,N_7856,N_6206);
nand U8032 (N_8032,N_6695,N_6779);
and U8033 (N_8033,N_7924,N_6802);
and U8034 (N_8034,N_6286,N_6812);
xor U8035 (N_8035,N_6432,N_7416);
nand U8036 (N_8036,N_6037,N_7424);
nor U8037 (N_8037,N_6202,N_7081);
or U8038 (N_8038,N_6684,N_6282);
nand U8039 (N_8039,N_7938,N_7436);
xnor U8040 (N_8040,N_6831,N_6195);
and U8041 (N_8041,N_6814,N_7961);
or U8042 (N_8042,N_6637,N_7822);
nand U8043 (N_8043,N_6591,N_6589);
and U8044 (N_8044,N_6746,N_7250);
xnor U8045 (N_8045,N_6614,N_7000);
nand U8046 (N_8046,N_6410,N_7540);
nor U8047 (N_8047,N_7617,N_7199);
and U8048 (N_8048,N_6978,N_6368);
or U8049 (N_8049,N_6048,N_7164);
or U8050 (N_8050,N_7672,N_6848);
nand U8051 (N_8051,N_7724,N_6000);
or U8052 (N_8052,N_6357,N_6440);
and U8053 (N_8053,N_6504,N_6745);
nand U8054 (N_8054,N_6305,N_6413);
nand U8055 (N_8055,N_7048,N_7733);
nor U8056 (N_8056,N_7981,N_7032);
nor U8057 (N_8057,N_7440,N_7914);
or U8058 (N_8058,N_7262,N_6411);
nand U8059 (N_8059,N_6423,N_7879);
xor U8060 (N_8060,N_7612,N_7105);
nand U8061 (N_8061,N_7460,N_6058);
and U8062 (N_8062,N_7082,N_6832);
nand U8063 (N_8063,N_7462,N_6307);
nand U8064 (N_8064,N_6968,N_6647);
or U8065 (N_8065,N_7108,N_6811);
nor U8066 (N_8066,N_7461,N_6215);
nand U8067 (N_8067,N_6162,N_7012);
nand U8068 (N_8068,N_7236,N_7015);
or U8069 (N_8069,N_7381,N_7499);
xnor U8070 (N_8070,N_7358,N_6260);
nor U8071 (N_8071,N_7067,N_7147);
nor U8072 (N_8072,N_7613,N_7541);
nand U8073 (N_8073,N_7784,N_7548);
or U8074 (N_8074,N_6751,N_7330);
nor U8075 (N_8075,N_7212,N_7937);
xnor U8076 (N_8076,N_7553,N_6807);
and U8077 (N_8077,N_6399,N_6648);
or U8078 (N_8078,N_6677,N_6219);
or U8079 (N_8079,N_7252,N_7438);
xnor U8080 (N_8080,N_6117,N_6913);
nand U8081 (N_8081,N_7463,N_6038);
nor U8082 (N_8082,N_6388,N_7152);
and U8083 (N_8083,N_7409,N_6155);
and U8084 (N_8084,N_6073,N_7668);
nand U8085 (N_8085,N_7042,N_6919);
nand U8086 (N_8086,N_7293,N_7790);
nor U8087 (N_8087,N_6886,N_6378);
nand U8088 (N_8088,N_7133,N_7238);
nor U8089 (N_8089,N_7132,N_7335);
nor U8090 (N_8090,N_6633,N_6864);
nor U8091 (N_8091,N_7812,N_7507);
and U8092 (N_8092,N_6014,N_6229);
and U8093 (N_8093,N_6001,N_6557);
nor U8094 (N_8094,N_6764,N_6606);
nor U8095 (N_8095,N_7624,N_6326);
nor U8096 (N_8096,N_6698,N_6820);
xnor U8097 (N_8097,N_7743,N_6881);
or U8098 (N_8098,N_6412,N_6642);
nand U8099 (N_8099,N_6005,N_6990);
nor U8100 (N_8100,N_7401,N_6559);
nand U8101 (N_8101,N_6216,N_7529);
and U8102 (N_8102,N_6435,N_7194);
or U8103 (N_8103,N_7899,N_6600);
nor U8104 (N_8104,N_7992,N_7008);
and U8105 (N_8105,N_7479,N_6341);
or U8106 (N_8106,N_6555,N_6707);
and U8107 (N_8107,N_6320,N_6580);
nand U8108 (N_8108,N_6276,N_7411);
or U8109 (N_8109,N_6173,N_6394);
and U8110 (N_8110,N_7649,N_7653);
nand U8111 (N_8111,N_6475,N_7390);
xor U8112 (N_8112,N_6460,N_7766);
nand U8113 (N_8113,N_7117,N_7570);
and U8114 (N_8114,N_7395,N_7841);
and U8115 (N_8115,N_7607,N_7647);
and U8116 (N_8116,N_7234,N_6094);
nand U8117 (N_8117,N_7066,N_6592);
or U8118 (N_8118,N_7665,N_7657);
nand U8119 (N_8119,N_7973,N_7405);
or U8120 (N_8120,N_7767,N_7003);
and U8121 (N_8121,N_6433,N_7974);
xnor U8122 (N_8122,N_7104,N_7053);
or U8123 (N_8123,N_6946,N_6963);
or U8124 (N_8124,N_7369,N_6187);
xor U8125 (N_8125,N_7443,N_7889);
xnor U8126 (N_8126,N_7208,N_7071);
or U8127 (N_8127,N_6955,N_7623);
xnor U8128 (N_8128,N_6650,N_7038);
xor U8129 (N_8129,N_6901,N_7457);
and U8130 (N_8130,N_6414,N_7235);
nor U8131 (N_8131,N_7611,N_7368);
nor U8132 (N_8132,N_7887,N_7594);
xnor U8133 (N_8133,N_7906,N_6644);
xor U8134 (N_8134,N_7793,N_7145);
and U8135 (N_8135,N_7820,N_6776);
nor U8136 (N_8136,N_7866,N_6488);
nor U8137 (N_8137,N_6740,N_6500);
and U8138 (N_8138,N_7636,N_6581);
xnor U8139 (N_8139,N_6290,N_6209);
nor U8140 (N_8140,N_6965,N_6631);
xnor U8141 (N_8141,N_6113,N_6363);
nand U8142 (N_8142,N_7771,N_7838);
nor U8143 (N_8143,N_6860,N_6291);
or U8144 (N_8144,N_6981,N_6911);
nor U8145 (N_8145,N_7600,N_6622);
nor U8146 (N_8146,N_6053,N_7249);
and U8147 (N_8147,N_6529,N_7651);
xor U8148 (N_8148,N_7497,N_7228);
nand U8149 (N_8149,N_7847,N_7685);
nor U8150 (N_8150,N_7469,N_7472);
nor U8151 (N_8151,N_7593,N_7315);
nor U8152 (N_8152,N_7997,N_7569);
xnor U8153 (N_8153,N_6103,N_6755);
nand U8154 (N_8154,N_6838,N_6241);
nand U8155 (N_8155,N_6610,N_7799);
and U8156 (N_8156,N_6739,N_6514);
and U8157 (N_8157,N_7239,N_7814);
nor U8158 (N_8158,N_6510,N_7379);
or U8159 (N_8159,N_7107,N_6834);
nor U8160 (N_8160,N_6128,N_7935);
or U8161 (N_8161,N_7149,N_7317);
or U8162 (N_8162,N_7397,N_6143);
xor U8163 (N_8163,N_6759,N_6952);
nor U8164 (N_8164,N_7183,N_6780);
or U8165 (N_8165,N_6930,N_7699);
nor U8166 (N_8166,N_7833,N_7445);
and U8167 (N_8167,N_6914,N_7709);
nor U8168 (N_8168,N_6771,N_7148);
nor U8169 (N_8169,N_6294,N_7732);
xor U8170 (N_8170,N_7546,N_7224);
or U8171 (N_8171,N_6894,N_6883);
nor U8172 (N_8172,N_7488,N_6833);
or U8173 (N_8173,N_6661,N_6194);
xor U8174 (N_8174,N_6844,N_7708);
and U8175 (N_8175,N_6004,N_7962);
nor U8176 (N_8176,N_6731,N_7007);
xnor U8177 (N_8177,N_7635,N_7151);
xor U8178 (N_8178,N_6039,N_6304);
xnor U8179 (N_8179,N_7230,N_6322);
or U8180 (N_8180,N_7614,N_6651);
and U8181 (N_8181,N_6567,N_6758);
nand U8182 (N_8182,N_6835,N_6705);
and U8183 (N_8183,N_7726,N_7022);
nand U8184 (N_8184,N_7723,N_7321);
xor U8185 (N_8185,N_6578,N_7802);
xor U8186 (N_8186,N_6799,N_7747);
and U8187 (N_8187,N_7214,N_7456);
nand U8188 (N_8188,N_7939,N_7915);
and U8189 (N_8189,N_7933,N_6816);
nor U8190 (N_8190,N_7103,N_6463);
or U8191 (N_8191,N_7310,N_6601);
xor U8192 (N_8192,N_6688,N_6392);
nor U8193 (N_8193,N_7917,N_7426);
xor U8194 (N_8194,N_7674,N_6337);
xnor U8195 (N_8195,N_6034,N_6605);
xnor U8196 (N_8196,N_7265,N_7832);
and U8197 (N_8197,N_6694,N_6521);
nor U8198 (N_8198,N_7043,N_6762);
nor U8199 (N_8199,N_7301,N_7632);
and U8200 (N_8200,N_7789,N_6047);
xnor U8201 (N_8201,N_7894,N_7084);
nor U8202 (N_8202,N_6728,N_7909);
or U8203 (N_8203,N_7074,N_7433);
xor U8204 (N_8204,N_7761,N_7057);
or U8205 (N_8205,N_6172,N_7324);
nand U8206 (N_8206,N_6754,N_7299);
xnor U8207 (N_8207,N_7587,N_6214);
or U8208 (N_8208,N_6537,N_7157);
or U8209 (N_8209,N_7524,N_7957);
and U8210 (N_8210,N_7953,N_7059);
nor U8211 (N_8211,N_6499,N_6525);
nor U8212 (N_8212,N_6686,N_6123);
nor U8213 (N_8213,N_6800,N_6493);
xnor U8214 (N_8214,N_6088,N_6130);
nor U8215 (N_8215,N_7967,N_7464);
nor U8216 (N_8216,N_6408,N_6634);
nand U8217 (N_8217,N_6108,N_6057);
nor U8218 (N_8218,N_7470,N_6896);
or U8219 (N_8219,N_7020,N_6636);
or U8220 (N_8220,N_6271,N_7535);
nor U8221 (N_8221,N_7858,N_7389);
nand U8222 (N_8222,N_6097,N_7558);
and U8223 (N_8223,N_6075,N_6213);
or U8224 (N_8224,N_6249,N_6718);
and U8225 (N_8225,N_7028,N_7890);
nand U8226 (N_8226,N_7396,N_6274);
nor U8227 (N_8227,N_6957,N_7075);
xnor U8228 (N_8228,N_6670,N_7511);
or U8229 (N_8229,N_6397,N_7220);
nand U8230 (N_8230,N_7680,N_6372);
or U8231 (N_8231,N_6809,N_6288);
nor U8232 (N_8232,N_7804,N_6984);
xnor U8233 (N_8233,N_7884,N_7063);
or U8234 (N_8234,N_7621,N_7948);
and U8235 (N_8235,N_7615,N_7567);
nor U8236 (N_8236,N_6954,N_7362);
and U8237 (N_8237,N_7618,N_7807);
xnor U8238 (N_8238,N_7878,N_7153);
nor U8239 (N_8239,N_6046,N_6389);
and U8240 (N_8240,N_6616,N_7865);
and U8241 (N_8241,N_6658,N_7191);
nand U8242 (N_8242,N_7231,N_7393);
nor U8243 (N_8243,N_7947,N_7956);
or U8244 (N_8244,N_6178,N_7682);
nor U8245 (N_8245,N_7552,N_6856);
nand U8246 (N_8246,N_6766,N_7141);
nor U8247 (N_8247,N_7805,N_6285);
and U8248 (N_8248,N_7627,N_6361);
xor U8249 (N_8249,N_7854,N_7083);
and U8250 (N_8250,N_7165,N_6077);
nor U8251 (N_8251,N_6474,N_6302);
xor U8252 (N_8252,N_6464,N_7429);
nand U8253 (N_8253,N_7345,N_7065);
and U8254 (N_8254,N_6664,N_7683);
xnor U8255 (N_8255,N_7778,N_6553);
and U8256 (N_8256,N_6657,N_7064);
and U8257 (N_8257,N_6570,N_6931);
and U8258 (N_8258,N_7316,N_6084);
and U8259 (N_8259,N_7661,N_7205);
and U8260 (N_8260,N_7131,N_7322);
nor U8261 (N_8261,N_6470,N_7744);
or U8262 (N_8262,N_6163,N_6681);
xnor U8263 (N_8263,N_7213,N_6347);
or U8264 (N_8264,N_7987,N_7885);
nand U8265 (N_8265,N_6671,N_7167);
nor U8266 (N_8266,N_6089,N_6607);
xnor U8267 (N_8267,N_6763,N_6749);
nand U8268 (N_8268,N_6246,N_7910);
nor U8269 (N_8269,N_6752,N_7837);
and U8270 (N_8270,N_6479,N_6859);
nand U8271 (N_8271,N_6157,N_7590);
nor U8272 (N_8272,N_7266,N_6110);
nor U8273 (N_8273,N_7097,N_6767);
nor U8274 (N_8274,N_6218,N_6197);
and U8275 (N_8275,N_6016,N_6055);
or U8276 (N_8276,N_6243,N_6724);
and U8277 (N_8277,N_7702,N_6709);
or U8278 (N_8278,N_7563,N_7863);
nor U8279 (N_8279,N_6821,N_6942);
xor U8280 (N_8280,N_6925,N_6769);
nand U8281 (N_8281,N_6452,N_6114);
and U8282 (N_8282,N_6893,N_7707);
nor U8283 (N_8283,N_7993,N_7338);
or U8284 (N_8284,N_6852,N_7525);
or U8285 (N_8285,N_7571,N_7694);
nand U8286 (N_8286,N_7811,N_6438);
and U8287 (N_8287,N_6120,N_7977);
xor U8288 (N_8288,N_6808,N_6737);
nand U8289 (N_8289,N_7639,N_7127);
nor U8290 (N_8290,N_6104,N_7382);
nand U8291 (N_8291,N_6238,N_6937);
nor U8292 (N_8292,N_6270,N_6723);
and U8293 (N_8293,N_6405,N_6107);
nor U8294 (N_8294,N_6006,N_7551);
or U8295 (N_8295,N_7496,N_6993);
and U8296 (N_8296,N_7343,N_7144);
xnor U8297 (N_8297,N_7990,N_6519);
nand U8298 (N_8298,N_7966,N_7645);
and U8299 (N_8299,N_7999,N_7877);
or U8300 (N_8300,N_6144,N_6619);
nand U8301 (N_8301,N_6092,N_6335);
nor U8302 (N_8302,N_7970,N_6943);
xor U8303 (N_8303,N_7264,N_6311);
nor U8304 (N_8304,N_7673,N_6355);
or U8305 (N_8305,N_7364,N_7675);
nor U8306 (N_8306,N_6180,N_7971);
nand U8307 (N_8307,N_6188,N_7658);
nor U8308 (N_8308,N_7484,N_6393);
nand U8309 (N_8309,N_6170,N_7308);
and U8310 (N_8310,N_7773,N_6126);
nor U8311 (N_8311,N_6490,N_7475);
nor U8312 (N_8312,N_7454,N_6649);
or U8313 (N_8313,N_6836,N_6122);
nor U8314 (N_8314,N_6242,N_6970);
xor U8315 (N_8315,N_7800,N_7662);
or U8316 (N_8316,N_6445,N_6316);
nor U8317 (N_8317,N_6639,N_7297);
nand U8318 (N_8318,N_7388,N_7319);
and U8319 (N_8319,N_7045,N_7829);
nor U8320 (N_8320,N_6778,N_6185);
nand U8321 (N_8321,N_6146,N_7209);
nor U8322 (N_8322,N_6549,N_6720);
or U8323 (N_8323,N_7663,N_6703);
and U8324 (N_8324,N_6186,N_6823);
nand U8325 (N_8325,N_6839,N_7643);
xor U8326 (N_8326,N_6171,N_6880);
nand U8327 (N_8327,N_7994,N_6511);
and U8328 (N_8328,N_7347,N_7787);
or U8329 (N_8329,N_7217,N_7143);
nor U8330 (N_8330,N_6045,N_7786);
and U8331 (N_8331,N_7677,N_7543);
nand U8332 (N_8332,N_6421,N_6467);
nand U8333 (N_8333,N_7334,N_6689);
and U8334 (N_8334,N_7835,N_6627);
or U8335 (N_8335,N_6220,N_6736);
and U8336 (N_8336,N_7809,N_6051);
nand U8337 (N_8337,N_6871,N_6635);
xnor U8338 (N_8338,N_7748,N_6468);
nand U8339 (N_8339,N_6456,N_6334);
or U8340 (N_8340,N_7155,N_6091);
xnor U8341 (N_8341,N_6673,N_6572);
or U8342 (N_8342,N_7242,N_6266);
and U8343 (N_8343,N_7089,N_7428);
nand U8344 (N_8344,N_7925,N_7574);
xor U8345 (N_8345,N_7085,N_6403);
xor U8346 (N_8346,N_7500,N_7849);
and U8347 (N_8347,N_6147,N_7985);
xnor U8348 (N_8348,N_6794,N_6283);
or U8349 (N_8349,N_7712,N_7951);
xor U8350 (N_8350,N_6227,N_6785);
or U8351 (N_8351,N_6679,N_6454);
and U8352 (N_8352,N_7098,N_7969);
and U8353 (N_8353,N_6028,N_7339);
nand U8354 (N_8354,N_6314,N_7542);
nor U8355 (N_8355,N_6429,N_7882);
xnor U8356 (N_8356,N_7911,N_6135);
xor U8357 (N_8357,N_7295,N_6278);
nand U8358 (N_8358,N_6083,N_7620);
or U8359 (N_8359,N_6628,N_6632);
nand U8360 (N_8360,N_6193,N_7046);
and U8361 (N_8361,N_7537,N_7051);
or U8362 (N_8362,N_7049,N_7115);
xor U8363 (N_8363,N_6507,N_7751);
nand U8364 (N_8364,N_7233,N_6583);
nand U8365 (N_8365,N_6448,N_6858);
xnor U8366 (N_8366,N_7554,N_7871);
nand U8367 (N_8367,N_7932,N_6874);
xnor U8368 (N_8368,N_7803,N_6124);
and U8369 (N_8369,N_7420,N_7373);
nand U8370 (N_8370,N_6546,N_7502);
nand U8371 (N_8371,N_6528,N_6887);
and U8372 (N_8372,N_7130,N_7311);
or U8373 (N_8373,N_7810,N_7286);
or U8374 (N_8374,N_6574,N_6682);
xor U8375 (N_8375,N_6941,N_7325);
nor U8376 (N_8376,N_6338,N_6899);
or U8377 (N_8377,N_7047,N_6356);
nor U8378 (N_8378,N_7504,N_7629);
nor U8379 (N_8379,N_6604,N_7202);
xor U8380 (N_8380,N_6112,N_6160);
or U8381 (N_8381,N_6228,N_7834);
xnor U8382 (N_8382,N_6599,N_6577);
xnor U8383 (N_8383,N_7414,N_7585);
nor U8384 (N_8384,N_7770,N_7934);
and U8385 (N_8385,N_7146,N_6863);
nand U8386 (N_8386,N_7795,N_6306);
xnor U8387 (N_8387,N_6564,N_7891);
nor U8388 (N_8388,N_7407,N_6395);
and U8389 (N_8389,N_6732,N_7298);
nor U8390 (N_8390,N_7431,N_7959);
and U8391 (N_8391,N_6030,N_7073);
xor U8392 (N_8392,N_6867,N_6462);
nand U8393 (N_8393,N_6608,N_7459);
xnor U8394 (N_8394,N_6164,N_7385);
nor U8395 (N_8395,N_6258,N_6653);
or U8396 (N_8396,N_6722,N_6585);
or U8397 (N_8397,N_6022,N_6152);
or U8398 (N_8398,N_6875,N_7588);
nor U8399 (N_8399,N_6977,N_7516);
nand U8400 (N_8400,N_6207,N_6358);
xor U8401 (N_8401,N_7122,N_7446);
xor U8402 (N_8402,N_7873,N_6441);
nor U8403 (N_8403,N_6985,N_7642);
xor U8404 (N_8404,N_6313,N_6862);
xnor U8405 (N_8405,N_6956,N_7077);
and U8406 (N_8406,N_7907,N_6344);
nor U8407 (N_8407,N_7101,N_7099);
xor U8408 (N_8408,N_6548,N_6437);
nand U8409 (N_8409,N_7869,N_6101);
nand U8410 (N_8410,N_7112,N_7606);
or U8411 (N_8411,N_6131,N_7188);
or U8412 (N_8412,N_7700,N_6487);
and U8413 (N_8413,N_6327,N_7988);
nor U8414 (N_8414,N_6044,N_6853);
or U8415 (N_8415,N_6926,N_6383);
nor U8416 (N_8416,N_6588,N_7825);
nand U8417 (N_8417,N_7931,N_7300);
nand U8418 (N_8418,N_7260,N_7268);
nand U8419 (N_8419,N_7696,N_7764);
nor U8420 (N_8420,N_6527,N_7134);
xnor U8421 (N_8421,N_7275,N_7468);
and U8422 (N_8422,N_7855,N_6096);
nand U8423 (N_8423,N_6786,N_6263);
and U8424 (N_8424,N_6222,N_6828);
and U8425 (N_8425,N_7912,N_7986);
xor U8426 (N_8426,N_6530,N_6903);
and U8427 (N_8427,N_7881,N_6950);
nor U8428 (N_8428,N_7061,N_6640);
nor U8429 (N_8429,N_6909,N_6247);
or U8430 (N_8430,N_7333,N_6168);
xnor U8431 (N_8431,N_7527,N_7023);
nand U8432 (N_8432,N_7534,N_6806);
or U8433 (N_8433,N_6331,N_7128);
nand U8434 (N_8434,N_6175,N_7692);
nor U8435 (N_8435,N_6565,N_6265);
nand U8436 (N_8436,N_7892,N_6804);
nor U8437 (N_8437,N_6960,N_7539);
nor U8438 (N_8438,N_6211,N_7086);
or U8439 (N_8439,N_7383,N_6885);
and U8440 (N_8440,N_6465,N_7307);
nand U8441 (N_8441,N_6774,N_7030);
and U8442 (N_8442,N_7344,N_7850);
and U8443 (N_8443,N_6992,N_6757);
nor U8444 (N_8444,N_6609,N_6715);
nor U8445 (N_8445,N_6547,N_6167);
and U8446 (N_8446,N_7626,N_7952);
xnor U8447 (N_8447,N_7745,N_7113);
or U8448 (N_8448,N_7519,N_7356);
nor U8449 (N_8449,N_7331,N_6568);
nor U8450 (N_8450,N_7905,N_6318);
xnor U8451 (N_8451,N_6424,N_7261);
nor U8452 (N_8452,N_6332,N_7671);
or U8453 (N_8453,N_6753,N_6976);
and U8454 (N_8454,N_7058,N_7450);
xor U8455 (N_8455,N_7886,N_6773);
or U8456 (N_8456,N_6391,N_6775);
and U8457 (N_8457,N_6156,N_6127);
and U8458 (N_8458,N_6250,N_7565);
or U8459 (N_8459,N_7681,N_7365);
xnor U8460 (N_8460,N_6351,N_7138);
xor U8461 (N_8461,N_6336,N_6259);
or U8462 (N_8462,N_6281,N_7399);
xnor U8463 (N_8463,N_7523,N_7868);
or U8464 (N_8464,N_7092,N_6018);
nand U8465 (N_8465,N_6293,N_7291);
nand U8466 (N_8466,N_6665,N_6617);
nor U8467 (N_8467,N_7875,N_7547);
nor U8468 (N_8468,N_7272,N_7964);
and U8469 (N_8469,N_7170,N_7314);
and U8470 (N_8470,N_6532,N_7444);
xor U8471 (N_8471,N_6052,N_6287);
nor U8472 (N_8472,N_6491,N_7544);
nand U8473 (N_8473,N_6534,N_6561);
or U8474 (N_8474,N_6400,N_6011);
or U8475 (N_8475,N_7410,N_7140);
xnor U8476 (N_8476,N_7175,N_7660);
or U8477 (N_8477,N_6573,N_7510);
and U8478 (N_8478,N_7550,N_7403);
nor U8479 (N_8479,N_7664,N_6154);
and U8480 (N_8480,N_6742,N_7177);
nor U8481 (N_8481,N_7110,N_6721);
or U8482 (N_8482,N_6176,N_7018);
and U8483 (N_8483,N_7304,N_7597);
xor U8484 (N_8484,N_7292,N_7963);
nor U8485 (N_8485,N_7512,N_7686);
xnor U8486 (N_8486,N_7184,N_7698);
and U8487 (N_8487,N_7509,N_6596);
xnor U8488 (N_8488,N_6457,N_7474);
nand U8489 (N_8489,N_7287,N_7305);
and U8490 (N_8490,N_7619,N_6367);
or U8491 (N_8491,N_7650,N_6230);
and U8492 (N_8492,N_6912,N_7185);
or U8493 (N_8493,N_7477,N_7102);
and U8494 (N_8494,N_7240,N_7486);
xnor U8495 (N_8495,N_6822,N_6109);
and U8496 (N_8496,N_7792,N_6623);
xnor U8497 (N_8497,N_6319,N_6535);
or U8498 (N_8498,N_6918,N_7853);
and U8499 (N_8499,N_7921,N_7734);
xor U8500 (N_8500,N_7387,N_6234);
nand U8501 (N_8501,N_6508,N_6478);
and U8502 (N_8502,N_6842,N_6221);
nand U8503 (N_8503,N_7069,N_6396);
and U8504 (N_8504,N_6485,N_6643);
nand U8505 (N_8505,N_6272,N_7025);
xor U8506 (N_8506,N_7729,N_7274);
nand U8507 (N_8507,N_6652,N_7087);
nand U8508 (N_8508,N_7655,N_6569);
xor U8509 (N_8509,N_7481,N_7284);
or U8510 (N_8510,N_6339,N_7276);
nand U8511 (N_8511,N_6343,N_6268);
xnor U8512 (N_8512,N_7035,N_7050);
or U8513 (N_8513,N_7027,N_7372);
nor U8514 (N_8514,N_6480,N_7193);
or U8515 (N_8515,N_6387,N_6079);
xnor U8516 (N_8516,N_7946,N_7100);
nor U8517 (N_8517,N_6315,N_6416);
and U8518 (N_8518,N_7599,N_6184);
nand U8519 (N_8519,N_7813,N_6932);
or U8520 (N_8520,N_7843,N_7688);
nor U8521 (N_8521,N_6974,N_6450);
nor U8522 (N_8522,N_7466,N_6455);
and U8523 (N_8523,N_7201,N_7419);
and U8524 (N_8524,N_6239,N_7336);
or U8525 (N_8525,N_6615,N_7190);
xnor U8526 (N_8526,N_7631,N_6819);
nor U8527 (N_8527,N_7377,N_7836);
or U8528 (N_8528,N_6076,N_7306);
or U8529 (N_8529,N_6477,N_7715);
nor U8530 (N_8530,N_6384,N_6801);
or U8531 (N_8531,N_6915,N_6846);
or U8532 (N_8532,N_6725,N_7095);
nand U8533 (N_8533,N_6513,N_6253);
or U8534 (N_8534,N_6861,N_7898);
xor U8535 (N_8535,N_6054,N_7968);
xor U8536 (N_8536,N_6098,N_7648);
xor U8537 (N_8537,N_6563,N_6983);
or U8538 (N_8538,N_7806,N_6295);
nor U8539 (N_8539,N_6224,N_6916);
or U8540 (N_8540,N_6093,N_6713);
or U8541 (N_8541,N_6503,N_7378);
nor U8542 (N_8542,N_6518,N_7706);
nor U8543 (N_8543,N_7019,N_6382);
nand U8544 (N_8544,N_6869,N_6542);
nand U8545 (N_8545,N_7954,N_6524);
xnor U8546 (N_8546,N_7255,N_6865);
and U8547 (N_8547,N_7638,N_7736);
and U8548 (N_8548,N_6626,N_7161);
xor U8549 (N_8549,N_7289,N_7052);
nor U8550 (N_8550,N_7772,N_6476);
nor U8551 (N_8551,N_6791,N_6308);
nand U8552 (N_8552,N_6562,N_6081);
nor U8553 (N_8553,N_7458,N_6191);
xor U8554 (N_8554,N_7738,N_7913);
nor U8555 (N_8555,N_7536,N_6473);
xor U8556 (N_8556,N_6036,N_6060);
nand U8557 (N_8557,N_7029,N_6940);
and U8558 (N_8558,N_7602,N_6404);
xnor U8559 (N_8559,N_6667,N_7204);
xnor U8560 (N_8560,N_7485,N_7503);
nor U8561 (N_8561,N_7109,N_7269);
nor U8562 (N_8562,N_6010,N_7622);
and U8563 (N_8563,N_6374,N_6134);
and U8564 (N_8564,N_7776,N_7088);
and U8565 (N_8565,N_6136,N_6360);
or U8566 (N_8566,N_7271,N_6849);
or U8567 (N_8567,N_7918,N_7896);
and U8568 (N_8568,N_6364,N_6882);
and U8569 (N_8569,N_7596,N_6002);
nor U8570 (N_8570,N_7021,N_6189);
nand U8571 (N_8571,N_6065,N_6254);
xor U8572 (N_8572,N_7839,N_6678);
nor U8573 (N_8573,N_7118,N_7120);
nand U8574 (N_8574,N_7163,N_7294);
nand U8575 (N_8575,N_6533,N_6021);
xor U8576 (N_8576,N_6453,N_6299);
nand U8577 (N_8577,N_6967,N_7575);
nor U8578 (N_8578,N_6362,N_7353);
and U8579 (N_8579,N_6872,N_6969);
nand U8580 (N_8580,N_7779,N_6795);
nand U8581 (N_8581,N_7979,N_7452);
and U8582 (N_8582,N_6945,N_7232);
nand U8583 (N_8583,N_7801,N_6947);
and U8584 (N_8584,N_7320,N_6813);
nand U8585 (N_8585,N_6980,N_6516);
or U8586 (N_8586,N_6826,N_7568);
and U8587 (N_8587,N_7538,N_7137);
and U8588 (N_8588,N_6927,N_6444);
nand U8589 (N_8589,N_7874,N_7280);
xor U8590 (N_8590,N_6489,N_6428);
xnor U8591 (N_8591,N_6070,N_6119);
nor U8592 (N_8592,N_7010,N_7666);
xor U8593 (N_8593,N_7592,N_7253);
nand U8594 (N_8594,N_7827,N_6252);
or U8595 (N_8595,N_7350,N_7421);
nand U8596 (N_8596,N_6866,N_7756);
nand U8597 (N_8597,N_6182,N_6042);
xnor U8598 (N_8598,N_7408,N_6105);
or U8599 (N_8599,N_7644,N_7366);
nor U8600 (N_8600,N_6830,N_7697);
xnor U8601 (N_8601,N_7174,N_6892);
and U8602 (N_8602,N_7323,N_7139);
nand U8603 (N_8603,N_6373,N_6929);
nand U8604 (N_8604,N_6099,N_7900);
nor U8605 (N_8605,N_7768,N_6409);
nand U8606 (N_8606,N_6630,N_6422);
nor U8607 (N_8607,N_7125,N_7168);
xnor U8608 (N_8608,N_7060,N_6118);
xor U8609 (N_8609,N_6935,N_6466);
nor U8610 (N_8610,N_6890,N_7342);
and U8611 (N_8611,N_7173,N_7728);
or U8612 (N_8612,N_6370,N_6257);
or U8613 (N_8613,N_6675,N_6255);
nor U8614 (N_8614,N_7689,N_7785);
nor U8615 (N_8615,N_6708,N_6289);
nor U8616 (N_8616,N_7758,N_6012);
and U8617 (N_8617,N_7417,N_7186);
and U8618 (N_8618,N_6020,N_7425);
and U8619 (N_8619,N_7374,N_6797);
xnor U8620 (N_8620,N_6035,N_6431);
nand U8621 (N_8621,N_7093,N_6273);
nor U8622 (N_8622,N_6434,N_6556);
or U8623 (N_8623,N_7011,N_7926);
nand U8624 (N_8624,N_7490,N_6687);
nor U8625 (N_8625,N_6087,N_6072);
or U8626 (N_8626,N_7589,N_6019);
nand U8627 (N_8627,N_6704,N_6953);
or U8628 (N_8628,N_7902,N_7637);
nor U8629 (N_8629,N_7888,N_7782);
nor U8630 (N_8630,N_6621,N_7549);
and U8631 (N_8631,N_6904,N_6324);
xor U8632 (N_8632,N_7625,N_7998);
xnor U8633 (N_8633,N_7564,N_6256);
nor U8634 (N_8634,N_7561,N_7415);
nor U8635 (N_8635,N_7828,N_6906);
or U8636 (N_8636,N_6248,N_7412);
nor U8637 (N_8637,N_6818,N_7363);
xor U8638 (N_8638,N_6280,N_7755);
xnor U8639 (N_8639,N_6380,N_6121);
and U8640 (N_8640,N_6069,N_6033);
and U8641 (N_8641,N_7687,N_6743);
nand U8642 (N_8642,N_6727,N_7989);
or U8643 (N_8643,N_6843,N_7975);
xor U8644 (N_8644,N_7727,N_6354);
or U8645 (N_8645,N_6279,N_7494);
nand U8646 (N_8646,N_6868,N_6663);
and U8647 (N_8647,N_6618,N_7150);
and U8648 (N_8648,N_6139,N_7434);
and U8649 (N_8649,N_7996,N_7222);
nor U8650 (N_8650,N_6515,N_7652);
or U8651 (N_8651,N_7072,N_6597);
nor U8652 (N_8652,N_6669,N_7659);
or U8653 (N_8653,N_6245,N_7302);
xnor U8654 (N_8654,N_6151,N_7106);
nand U8655 (N_8655,N_6590,N_6223);
or U8656 (N_8656,N_7941,N_6659);
and U8657 (N_8657,N_6310,N_7815);
and U8658 (N_8658,N_6461,N_6979);
nor U8659 (N_8659,N_6192,N_7080);
nor U8660 (N_8660,N_6401,N_6566);
nand U8661 (N_8661,N_6958,N_7219);
and U8662 (N_8662,N_6402,N_7676);
nor U8663 (N_8663,N_6032,N_7944);
nor U8664 (N_8664,N_6997,N_7277);
nand U8665 (N_8665,N_6439,N_6654);
and U8666 (N_8666,N_6710,N_6158);
nand U8667 (N_8667,N_7493,N_7903);
xor U8668 (N_8668,N_7965,N_6040);
or U8669 (N_8669,N_7641,N_6680);
nor U8670 (N_8670,N_7482,N_6426);
and U8671 (N_8671,N_7530,N_7701);
nand U8672 (N_8672,N_7923,N_6505);
or U8673 (N_8673,N_7851,N_7326);
nor U8674 (N_8674,N_7942,N_6975);
xnor U8675 (N_8675,N_7521,N_7346);
and U8676 (N_8676,N_6169,N_6734);
and U8677 (N_8677,N_7719,N_7752);
nand U8678 (N_8678,N_7400,N_6323);
and U8679 (N_8679,N_7371,N_7526);
nor U8680 (N_8680,N_6905,N_7016);
nand U8681 (N_8681,N_6442,N_6352);
and U8682 (N_8682,N_6777,N_7718);
nand U8683 (N_8683,N_6013,N_7187);
nor U8684 (N_8684,N_6959,N_7465);
xnor U8685 (N_8685,N_6697,N_7009);
nor U8686 (N_8686,N_6551,N_6484);
or U8687 (N_8687,N_7505,N_6277);
and U8688 (N_8688,N_7922,N_7960);
nand U8689 (N_8689,N_7427,N_7406);
or U8690 (N_8690,N_7256,N_7172);
nor U8691 (N_8691,N_6458,N_6026);
xor U8692 (N_8692,N_6190,N_6692);
nand U8693 (N_8693,N_7380,N_7288);
xor U8694 (N_8694,N_6153,N_6345);
and U8695 (N_8695,N_6624,N_6150);
nor U8696 (N_8696,N_7203,N_7578);
and U8697 (N_8697,N_7002,N_7327);
nor U8698 (N_8698,N_7777,N_7870);
nand U8699 (N_8699,N_6674,N_7223);
and U8700 (N_8700,N_6744,N_7211);
or U8701 (N_8701,N_6330,N_6558);
nand U8702 (N_8702,N_7991,N_6090);
xnor U8703 (N_8703,N_6620,N_7984);
nand U8704 (N_8704,N_6655,N_7586);
nor U8705 (N_8705,N_6066,N_7721);
nor U8706 (N_8706,N_6879,N_7189);
nor U8707 (N_8707,N_6870,N_7341);
nand U8708 (N_8708,N_7423,N_7669);
nor U8709 (N_8709,N_7355,N_6994);
nor U8710 (N_8710,N_7577,N_7263);
and U8711 (N_8711,N_6798,N_6668);
nand U8712 (N_8712,N_6691,N_6840);
nand U8713 (N_8713,N_6196,N_6803);
xor U8714 (N_8714,N_7560,N_6586);
nand U8715 (N_8715,N_7982,N_6082);
and U8716 (N_8716,N_7044,N_6349);
and U8717 (N_8717,N_6827,N_6520);
nor U8718 (N_8718,N_7557,N_7197);
nand U8719 (N_8719,N_7876,N_7283);
nor U8720 (N_8720,N_6982,N_7522);
nor U8721 (N_8721,N_7533,N_7439);
or U8722 (N_8722,N_6594,N_7735);
nand U8723 (N_8723,N_6201,N_6264);
nand U8724 (N_8724,N_6041,N_7861);
nor U8725 (N_8725,N_7840,N_7754);
xor U8726 (N_8726,N_6877,N_7972);
and U8727 (N_8727,N_7357,N_6922);
xnor U8728 (N_8728,N_7026,N_6159);
or U8729 (N_8729,N_6086,N_7225);
and U8730 (N_8730,N_6571,N_7830);
nand U8731 (N_8731,N_7704,N_7483);
xnor U8732 (N_8732,N_7413,N_7904);
xnor U8733 (N_8733,N_7824,N_6999);
xor U8734 (N_8734,N_7603,N_7605);
nor U8735 (N_8735,N_7532,N_6699);
xor U8736 (N_8736,N_7678,N_6350);
and U8737 (N_8737,N_7359,N_6756);
nor U8738 (N_8738,N_7111,N_7135);
or U8739 (N_8739,N_6179,N_7775);
xor U8740 (N_8740,N_6398,N_7818);
nand U8741 (N_8741,N_7955,N_7742);
and U8742 (N_8742,N_6995,N_6231);
and U8743 (N_8743,N_6951,N_6973);
nand U8744 (N_8744,N_6540,N_7608);
and U8745 (N_8745,N_7769,N_6921);
nand U8746 (N_8746,N_6140,N_6067);
and U8747 (N_8747,N_6235,N_7750);
nor U8748 (N_8748,N_6837,N_7337);
nor U8749 (N_8749,N_7241,N_7279);
nor U8750 (N_8750,N_6284,N_6436);
nor U8751 (N_8751,N_6481,N_6502);
nand U8752 (N_8752,N_6613,N_6902);
xor U8753 (N_8753,N_6204,N_7309);
and U8754 (N_8754,N_6765,N_7783);
and U8755 (N_8755,N_6888,N_7154);
or U8756 (N_8756,N_6625,N_7004);
or U8757 (N_8757,N_6693,N_6471);
or U8758 (N_8758,N_7404,N_6430);
nand U8759 (N_8759,N_6787,N_6102);
or U8760 (N_8760,N_7245,N_6296);
nor U8761 (N_8761,N_6495,N_7816);
nor U8762 (N_8762,N_6784,N_6638);
xnor U8763 (N_8763,N_7254,N_6847);
nor U8764 (N_8764,N_6593,N_6878);
or U8765 (N_8765,N_7014,N_6972);
nand U8766 (N_8766,N_7566,N_7725);
nand U8767 (N_8767,N_6074,N_7079);
nand U8768 (N_8768,N_6845,N_7226);
and U8769 (N_8769,N_7259,N_7062);
or U8770 (N_8770,N_6702,N_6181);
nor U8771 (N_8771,N_7765,N_7604);
xnor U8772 (N_8772,N_7006,N_6137);
nor U8773 (N_8773,N_6897,N_6125);
nor U8774 (N_8774,N_7693,N_6560);
xnor U8775 (N_8775,N_6895,N_6138);
nand U8776 (N_8776,N_7281,N_7763);
xor U8777 (N_8777,N_6741,N_6690);
xor U8778 (N_8778,N_6805,N_6796);
or U8779 (N_8779,N_6418,N_6469);
and U8780 (N_8780,N_7555,N_7731);
or U8781 (N_8781,N_6446,N_6321);
and U8782 (N_8782,N_6161,N_7746);
nor U8783 (N_8783,N_6050,N_6768);
nand U8784 (N_8784,N_7572,N_7491);
and U8785 (N_8785,N_6017,N_7872);
or U8786 (N_8786,N_7394,N_6961);
or U8787 (N_8787,N_7595,N_6177);
or U8788 (N_8788,N_6928,N_6825);
nand U8789 (N_8789,N_7703,N_7796);
and U8790 (N_8790,N_7121,N_7930);
nor U8791 (N_8791,N_7897,N_7584);
nor U8792 (N_8792,N_7730,N_6174);
nor U8793 (N_8793,N_7506,N_6068);
nor U8794 (N_8794,N_7920,N_6003);
xnor U8795 (N_8795,N_7498,N_6509);
nand U8796 (N_8796,N_7844,N_7826);
and U8797 (N_8797,N_7119,N_6711);
nand U8798 (N_8798,N_6996,N_6325);
xor U8799 (N_8799,N_7257,N_7760);
nor U8800 (N_8800,N_7518,N_6407);
and U8801 (N_8801,N_6415,N_6964);
nand U8802 (N_8802,N_7936,N_7684);
xnor U8803 (N_8803,N_7349,N_7031);
or U8804 (N_8804,N_6933,N_6523);
xnor U8805 (N_8805,N_6526,N_7303);
nor U8806 (N_8806,N_6936,N_7545);
nand U8807 (N_8807,N_7068,N_6576);
nand U8808 (N_8808,N_6217,N_7740);
xor U8809 (N_8809,N_7774,N_7332);
nor U8810 (N_8810,N_6015,N_7360);
and U8811 (N_8811,N_6810,N_6494);
nand U8812 (N_8812,N_7514,N_7630);
nand U8813 (N_8813,N_6376,N_6660);
nand U8814 (N_8814,N_7949,N_6717);
and U8815 (N_8815,N_6726,N_7513);
or U8816 (N_8816,N_6934,N_7781);
nand U8817 (N_8817,N_6366,N_7195);
xor U8818 (N_8818,N_7958,N_7860);
and U8819 (N_8819,N_6854,N_7221);
nand U8820 (N_8820,N_7114,N_6917);
xor U8821 (N_8821,N_6949,N_6782);
nand U8822 (N_8822,N_7005,N_6598);
nor U8823 (N_8823,N_6080,N_7508);
and U8824 (N_8824,N_6237,N_7476);
nor U8825 (N_8825,N_6582,N_7453);
and U8826 (N_8826,N_6716,N_7601);
nand U8827 (N_8827,N_6251,N_7609);
nand U8828 (N_8828,N_6225,N_7034);
xnor U8829 (N_8829,N_7573,N_7916);
or U8830 (N_8830,N_6522,N_7024);
and U8831 (N_8831,N_6781,N_6346);
and U8832 (N_8832,N_7392,N_6998);
xor U8833 (N_8833,N_7893,N_7591);
nand U8834 (N_8834,N_6148,N_6554);
or U8835 (N_8835,N_6550,N_6579);
nand U8836 (N_8836,N_7580,N_6208);
and U8837 (N_8837,N_6390,N_7176);
xnor U8838 (N_8838,N_7248,N_6656);
and U8839 (N_8839,N_6133,N_6317);
xor U8840 (N_8840,N_7654,N_6261);
nand U8841 (N_8841,N_7480,N_7995);
and U8842 (N_8842,N_6027,N_7036);
or U8843 (N_8843,N_6236,N_7640);
and U8844 (N_8844,N_7070,N_6447);
nor U8845 (N_8845,N_7753,N_6031);
and U8846 (N_8846,N_6748,N_7367);
nand U8847 (N_8847,N_6884,N_6141);
nand U8848 (N_8848,N_6506,N_7207);
and U8849 (N_8849,N_7056,N_6329);
nand U8850 (N_8850,N_6730,N_7447);
nand U8851 (N_8851,N_6706,N_7857);
xnor U8852 (N_8852,N_7928,N_7908);
xor U8853 (N_8853,N_7258,N_6924);
and U8854 (N_8854,N_6672,N_7762);
xnor U8855 (N_8855,N_7182,N_6783);
and U8856 (N_8856,N_7842,N_7244);
nor U8857 (N_8857,N_7646,N_7039);
nand U8858 (N_8858,N_6719,N_6512);
and U8859 (N_8859,N_6043,N_7864);
xnor U8860 (N_8860,N_7487,N_6989);
nand U8861 (N_8861,N_6541,N_7788);
or U8862 (N_8862,N_7581,N_7160);
nand U8863 (N_8863,N_7033,N_6232);
xnor U8864 (N_8864,N_6427,N_7435);
nand U8865 (N_8865,N_6106,N_7218);
and U8866 (N_8866,N_7817,N_7739);
and U8867 (N_8867,N_7290,N_7200);
and U8868 (N_8868,N_6451,N_6064);
nor U8869 (N_8869,N_7610,N_7180);
xnor U8870 (N_8870,N_6183,N_6666);
and U8871 (N_8871,N_7562,N_6889);
xor U8872 (N_8872,N_7848,N_7328);
and U8873 (N_8873,N_7442,N_6948);
nor U8874 (N_8874,N_6966,N_6851);
nor U8875 (N_8875,N_6760,N_6406);
xnor U8876 (N_8876,N_7441,N_6898);
nor U8877 (N_8877,N_7845,N_7181);
nand U8878 (N_8878,N_6303,N_6815);
and U8879 (N_8879,N_6300,N_6876);
xnor U8880 (N_8880,N_7722,N_6353);
nand U8881 (N_8881,N_6116,N_7386);
or U8882 (N_8882,N_6850,N_6486);
nand U8883 (N_8883,N_7329,N_7094);
nand U8884 (N_8884,N_7451,N_6492);
xor U8885 (N_8885,N_6738,N_7690);
and U8886 (N_8886,N_6449,N_6381);
nand U8887 (N_8887,N_6199,N_7384);
xnor U8888 (N_8888,N_7717,N_6145);
nor U8889 (N_8889,N_7273,N_7478);
nor U8890 (N_8890,N_6685,N_7422);
nand U8891 (N_8891,N_7391,N_6071);
and U8892 (N_8892,N_7471,N_7158);
and U8893 (N_8893,N_6149,N_6841);
or U8894 (N_8894,N_6729,N_6497);
and U8895 (N_8895,N_6536,N_7797);
and U8896 (N_8896,N_6009,N_7794);
and U8897 (N_8897,N_6063,N_6024);
nand U8898 (N_8898,N_6385,N_7576);
and U8899 (N_8899,N_6646,N_7282);
xnor U8900 (N_8900,N_6342,N_7883);
nor U8901 (N_8901,N_7791,N_7628);
nand U8902 (N_8902,N_6584,N_6205);
or U8903 (N_8903,N_7980,N_7296);
xor U8904 (N_8904,N_6539,N_6425);
nor U8905 (N_8905,N_6683,N_6991);
xor U8906 (N_8906,N_6301,N_6855);
nand U8907 (N_8907,N_6789,N_7798);
nand U8908 (N_8908,N_7001,N_7634);
xnor U8909 (N_8909,N_7616,N_6142);
nand U8910 (N_8910,N_6891,N_7246);
or U8911 (N_8911,N_6735,N_6939);
or U8912 (N_8912,N_6292,N_6420);
or U8913 (N_8913,N_6788,N_7216);
and U8914 (N_8914,N_6908,N_6611);
or U8915 (N_8915,N_7449,N_7705);
or U8916 (N_8916,N_6612,N_7398);
and U8917 (N_8917,N_6115,N_7713);
or U8918 (N_8918,N_6059,N_7206);
nand U8919 (N_8919,N_6733,N_7808);
nor U8920 (N_8920,N_7090,N_6309);
and U8921 (N_8921,N_7243,N_7467);
nand U8922 (N_8922,N_6297,N_6538);
nor U8923 (N_8923,N_7895,N_7515);
or U8924 (N_8924,N_7166,N_6986);
xor U8925 (N_8925,N_6770,N_7749);
xnor U8926 (N_8926,N_7448,N_7318);
or U8927 (N_8927,N_7691,N_7123);
xnor U8928 (N_8928,N_6419,N_6971);
nand U8929 (N_8929,N_6944,N_7179);
and U8930 (N_8930,N_6544,N_6417);
nand U8931 (N_8931,N_6761,N_7198);
xor U8932 (N_8932,N_6472,N_7455);
and U8933 (N_8933,N_7078,N_6262);
nand U8934 (N_8934,N_7361,N_7126);
or U8935 (N_8935,N_7142,N_6873);
xnor U8936 (N_8936,N_7162,N_7862);
and U8937 (N_8937,N_7430,N_7251);
xor U8938 (N_8938,N_6267,N_6531);
nor U8939 (N_8939,N_6545,N_7473);
xnor U8940 (N_8940,N_7091,N_7501);
and U8941 (N_8941,N_6496,N_7667);
and U8942 (N_8942,N_6056,N_6007);
or U8943 (N_8943,N_6938,N_7741);
and U8944 (N_8944,N_6240,N_6132);
nand U8945 (N_8945,N_6552,N_7859);
nor U8946 (N_8946,N_7528,N_7402);
and U8947 (N_8947,N_6198,N_6095);
xor U8948 (N_8948,N_7831,N_7531);
or U8949 (N_8949,N_6023,N_7633);
or U8950 (N_8950,N_7129,N_6226);
and U8951 (N_8951,N_7901,N_7823);
nor U8952 (N_8952,N_7116,N_7943);
nand U8953 (N_8953,N_6824,N_6792);
or U8954 (N_8954,N_7210,N_7821);
xnor U8955 (N_8955,N_6829,N_7559);
nor U8956 (N_8956,N_6501,N_6312);
xnor U8957 (N_8957,N_7247,N_7945);
and U8958 (N_8958,N_7054,N_6459);
xnor U8959 (N_8959,N_7556,N_7351);
or U8960 (N_8960,N_7418,N_6328);
nand U8961 (N_8961,N_7714,N_7354);
or U8962 (N_8962,N_7711,N_7227);
xor U8963 (N_8963,N_7520,N_7017);
nor U8964 (N_8964,N_7919,N_6701);
or U8965 (N_8965,N_6111,N_6793);
or U8966 (N_8966,N_7737,N_7598);
xnor U8967 (N_8967,N_6203,N_7867);
or U8968 (N_8968,N_7041,N_6595);
or U8969 (N_8969,N_6817,N_6987);
nor U8970 (N_8970,N_6543,N_6166);
and U8971 (N_8971,N_7656,N_6371);
or U8972 (N_8972,N_6587,N_7013);
xnor U8973 (N_8973,N_6900,N_6676);
and U8974 (N_8974,N_6379,N_6212);
and U8975 (N_8975,N_7880,N_6962);
or U8976 (N_8976,N_7757,N_7270);
and U8977 (N_8977,N_7819,N_6298);
nand U8978 (N_8978,N_7679,N_6603);
and U8979 (N_8979,N_7852,N_6750);
nor U8980 (N_8980,N_7215,N_6641);
and U8981 (N_8981,N_7695,N_7437);
nand U8982 (N_8982,N_6386,N_6857);
nor U8983 (N_8983,N_7237,N_6772);
nor U8984 (N_8984,N_6645,N_6244);
or U8985 (N_8985,N_6369,N_7495);
xnor U8986 (N_8986,N_6714,N_7929);
nor U8987 (N_8987,N_6078,N_7432);
and U8988 (N_8988,N_7076,N_6275);
and U8989 (N_8989,N_7579,N_6443);
nand U8990 (N_8990,N_7196,N_7720);
nor U8991 (N_8991,N_6700,N_6696);
nand U8992 (N_8992,N_7267,N_6365);
xnor U8993 (N_8993,N_6602,N_7171);
and U8994 (N_8994,N_7278,N_6377);
xor U8995 (N_8995,N_7375,N_6008);
xnor U8996 (N_8996,N_6269,N_6747);
nand U8997 (N_8997,N_7582,N_6375);
or U8998 (N_8998,N_7489,N_7352);
and U8999 (N_8999,N_7055,N_6333);
xnor U9000 (N_9000,N_6068,N_6981);
and U9001 (N_9001,N_6653,N_7188);
and U9002 (N_9002,N_7734,N_7033);
or U9003 (N_9003,N_7169,N_6229);
and U9004 (N_9004,N_6349,N_7469);
nand U9005 (N_9005,N_7541,N_7152);
nand U9006 (N_9006,N_7871,N_6088);
or U9007 (N_9007,N_7932,N_6271);
xnor U9008 (N_9008,N_7219,N_6044);
and U9009 (N_9009,N_7977,N_6616);
xnor U9010 (N_9010,N_6887,N_6994);
xnor U9011 (N_9011,N_7315,N_7933);
nor U9012 (N_9012,N_7395,N_6554);
nand U9013 (N_9013,N_6216,N_7142);
xnor U9014 (N_9014,N_7254,N_6028);
xnor U9015 (N_9015,N_6367,N_6645);
and U9016 (N_9016,N_7228,N_6084);
and U9017 (N_9017,N_6035,N_7246);
xor U9018 (N_9018,N_6017,N_6790);
and U9019 (N_9019,N_6032,N_6959);
xnor U9020 (N_9020,N_6750,N_7277);
nand U9021 (N_9021,N_7140,N_6897);
nor U9022 (N_9022,N_6085,N_6190);
nor U9023 (N_9023,N_6299,N_7761);
nor U9024 (N_9024,N_7918,N_6885);
and U9025 (N_9025,N_7742,N_7071);
and U9026 (N_9026,N_7138,N_7487);
nor U9027 (N_9027,N_6830,N_6923);
and U9028 (N_9028,N_6067,N_7799);
nand U9029 (N_9029,N_7805,N_7945);
nand U9030 (N_9030,N_7935,N_7931);
nand U9031 (N_9031,N_7310,N_6659);
xor U9032 (N_9032,N_6609,N_7800);
xnor U9033 (N_9033,N_6507,N_6101);
nand U9034 (N_9034,N_7188,N_7245);
and U9035 (N_9035,N_6936,N_7401);
xnor U9036 (N_9036,N_7897,N_7177);
or U9037 (N_9037,N_7878,N_7940);
xnor U9038 (N_9038,N_6734,N_6266);
and U9039 (N_9039,N_6990,N_7806);
and U9040 (N_9040,N_6996,N_7503);
and U9041 (N_9041,N_6978,N_6527);
xnor U9042 (N_9042,N_6488,N_7194);
and U9043 (N_9043,N_6603,N_6936);
or U9044 (N_9044,N_7573,N_7804);
nor U9045 (N_9045,N_6858,N_6898);
nor U9046 (N_9046,N_6010,N_6163);
nand U9047 (N_9047,N_6984,N_6826);
and U9048 (N_9048,N_6552,N_7406);
nor U9049 (N_9049,N_7261,N_7473);
and U9050 (N_9050,N_7049,N_7372);
xor U9051 (N_9051,N_6082,N_7827);
nor U9052 (N_9052,N_6454,N_6749);
nand U9053 (N_9053,N_6084,N_7162);
or U9054 (N_9054,N_6284,N_6414);
xor U9055 (N_9055,N_6082,N_6469);
or U9056 (N_9056,N_6637,N_7763);
xnor U9057 (N_9057,N_6632,N_6981);
nor U9058 (N_9058,N_7863,N_7903);
nand U9059 (N_9059,N_6536,N_6879);
and U9060 (N_9060,N_7202,N_7143);
and U9061 (N_9061,N_6874,N_7809);
nand U9062 (N_9062,N_7071,N_7351);
nor U9063 (N_9063,N_7646,N_7146);
nor U9064 (N_9064,N_6473,N_7843);
nor U9065 (N_9065,N_6790,N_6415);
nor U9066 (N_9066,N_6896,N_6932);
or U9067 (N_9067,N_7408,N_7518);
or U9068 (N_9068,N_7504,N_7209);
or U9069 (N_9069,N_6378,N_7993);
nor U9070 (N_9070,N_7895,N_7114);
or U9071 (N_9071,N_6872,N_6368);
nor U9072 (N_9072,N_7542,N_7348);
and U9073 (N_9073,N_6195,N_7829);
nor U9074 (N_9074,N_6408,N_7504);
nand U9075 (N_9075,N_6654,N_7783);
nor U9076 (N_9076,N_6050,N_6888);
nor U9077 (N_9077,N_6528,N_6305);
nand U9078 (N_9078,N_7966,N_6570);
nand U9079 (N_9079,N_7949,N_6268);
nand U9080 (N_9080,N_7275,N_7672);
nor U9081 (N_9081,N_6539,N_7956);
xnor U9082 (N_9082,N_6055,N_6805);
nand U9083 (N_9083,N_6122,N_6898);
or U9084 (N_9084,N_7395,N_6460);
and U9085 (N_9085,N_6264,N_6181);
nand U9086 (N_9086,N_7818,N_6461);
or U9087 (N_9087,N_6463,N_6257);
or U9088 (N_9088,N_6899,N_7478);
and U9089 (N_9089,N_6878,N_6646);
and U9090 (N_9090,N_6229,N_6262);
xnor U9091 (N_9091,N_6048,N_7169);
or U9092 (N_9092,N_6738,N_6273);
nor U9093 (N_9093,N_7970,N_7045);
nor U9094 (N_9094,N_7223,N_7499);
nor U9095 (N_9095,N_6068,N_6771);
xnor U9096 (N_9096,N_6162,N_6646);
or U9097 (N_9097,N_6639,N_7181);
xor U9098 (N_9098,N_7108,N_7059);
and U9099 (N_9099,N_6310,N_6694);
nand U9100 (N_9100,N_6141,N_7808);
or U9101 (N_9101,N_6646,N_7677);
xor U9102 (N_9102,N_7615,N_6152);
or U9103 (N_9103,N_7412,N_7518);
and U9104 (N_9104,N_6085,N_6106);
xor U9105 (N_9105,N_7314,N_6083);
nor U9106 (N_9106,N_7821,N_7710);
or U9107 (N_9107,N_6118,N_6103);
and U9108 (N_9108,N_7637,N_6973);
nor U9109 (N_9109,N_6221,N_7545);
or U9110 (N_9110,N_7763,N_6725);
or U9111 (N_9111,N_6916,N_6244);
and U9112 (N_9112,N_6027,N_7100);
xor U9113 (N_9113,N_6542,N_6342);
nor U9114 (N_9114,N_6833,N_7796);
and U9115 (N_9115,N_7470,N_6132);
nand U9116 (N_9116,N_7583,N_6153);
and U9117 (N_9117,N_6992,N_6776);
nand U9118 (N_9118,N_7828,N_6118);
nand U9119 (N_9119,N_7273,N_6059);
nor U9120 (N_9120,N_6448,N_6640);
and U9121 (N_9121,N_7127,N_6027);
or U9122 (N_9122,N_6664,N_6249);
or U9123 (N_9123,N_6390,N_7787);
and U9124 (N_9124,N_7619,N_6555);
xor U9125 (N_9125,N_6700,N_7738);
xnor U9126 (N_9126,N_7527,N_7573);
or U9127 (N_9127,N_7457,N_6542);
and U9128 (N_9128,N_6568,N_7894);
and U9129 (N_9129,N_6650,N_7744);
xnor U9130 (N_9130,N_7794,N_7217);
xor U9131 (N_9131,N_6966,N_7936);
or U9132 (N_9132,N_6587,N_6229);
xor U9133 (N_9133,N_7956,N_7889);
nand U9134 (N_9134,N_7590,N_7530);
xor U9135 (N_9135,N_6235,N_7637);
nand U9136 (N_9136,N_6511,N_7192);
and U9137 (N_9137,N_7621,N_7254);
or U9138 (N_9138,N_6609,N_7819);
nor U9139 (N_9139,N_6011,N_7788);
or U9140 (N_9140,N_6360,N_6712);
nand U9141 (N_9141,N_6838,N_6656);
or U9142 (N_9142,N_7161,N_7934);
nor U9143 (N_9143,N_6949,N_6134);
nand U9144 (N_9144,N_6669,N_6617);
nor U9145 (N_9145,N_7981,N_6145);
or U9146 (N_9146,N_6650,N_6460);
and U9147 (N_9147,N_6267,N_6301);
or U9148 (N_9148,N_6622,N_7419);
nand U9149 (N_9149,N_6310,N_6089);
xnor U9150 (N_9150,N_6069,N_7493);
and U9151 (N_9151,N_7405,N_6092);
nor U9152 (N_9152,N_6346,N_6929);
and U9153 (N_9153,N_6015,N_7603);
or U9154 (N_9154,N_6031,N_6540);
or U9155 (N_9155,N_6431,N_6751);
nor U9156 (N_9156,N_6121,N_7035);
or U9157 (N_9157,N_6007,N_7551);
nand U9158 (N_9158,N_6649,N_7768);
nor U9159 (N_9159,N_7078,N_7431);
or U9160 (N_9160,N_7080,N_7559);
nor U9161 (N_9161,N_6951,N_6584);
xnor U9162 (N_9162,N_7916,N_6092);
nand U9163 (N_9163,N_7543,N_6851);
or U9164 (N_9164,N_6161,N_6456);
nor U9165 (N_9165,N_7767,N_6090);
xnor U9166 (N_9166,N_6671,N_7324);
or U9167 (N_9167,N_6829,N_6787);
xnor U9168 (N_9168,N_7864,N_6689);
nor U9169 (N_9169,N_7150,N_7883);
or U9170 (N_9170,N_6972,N_6261);
nor U9171 (N_9171,N_7740,N_7297);
xnor U9172 (N_9172,N_6673,N_7360);
nand U9173 (N_9173,N_6952,N_6850);
nand U9174 (N_9174,N_7766,N_6142);
nor U9175 (N_9175,N_7266,N_6089);
nand U9176 (N_9176,N_6334,N_6418);
and U9177 (N_9177,N_7663,N_7756);
nor U9178 (N_9178,N_7689,N_6448);
or U9179 (N_9179,N_6730,N_7853);
nand U9180 (N_9180,N_7868,N_7828);
nand U9181 (N_9181,N_7842,N_7023);
xnor U9182 (N_9182,N_6696,N_6505);
nor U9183 (N_9183,N_6283,N_6345);
nand U9184 (N_9184,N_6883,N_7312);
and U9185 (N_9185,N_6430,N_6925);
xnor U9186 (N_9186,N_7668,N_6919);
nor U9187 (N_9187,N_6073,N_6016);
nand U9188 (N_9188,N_7159,N_7913);
xnor U9189 (N_9189,N_7152,N_6558);
and U9190 (N_9190,N_7793,N_6852);
nand U9191 (N_9191,N_7134,N_7871);
nor U9192 (N_9192,N_6067,N_6977);
nor U9193 (N_9193,N_7782,N_6474);
nand U9194 (N_9194,N_7017,N_6121);
nand U9195 (N_9195,N_7957,N_6934);
or U9196 (N_9196,N_6588,N_6682);
or U9197 (N_9197,N_6172,N_6780);
nand U9198 (N_9198,N_7690,N_6091);
xnor U9199 (N_9199,N_7801,N_6559);
or U9200 (N_9200,N_6284,N_7687);
nand U9201 (N_9201,N_7702,N_6909);
nor U9202 (N_9202,N_7832,N_6035);
and U9203 (N_9203,N_6573,N_7882);
and U9204 (N_9204,N_6715,N_7925);
nor U9205 (N_9205,N_6473,N_6545);
xor U9206 (N_9206,N_6388,N_7069);
xor U9207 (N_9207,N_6992,N_6115);
or U9208 (N_9208,N_6965,N_6197);
nand U9209 (N_9209,N_7683,N_7249);
and U9210 (N_9210,N_6698,N_7054);
nor U9211 (N_9211,N_7122,N_6107);
xor U9212 (N_9212,N_6834,N_6238);
and U9213 (N_9213,N_6337,N_7162);
nor U9214 (N_9214,N_6321,N_6540);
or U9215 (N_9215,N_6848,N_7706);
nand U9216 (N_9216,N_6490,N_6942);
xor U9217 (N_9217,N_6857,N_7614);
and U9218 (N_9218,N_7366,N_6056);
nor U9219 (N_9219,N_6938,N_7510);
xnor U9220 (N_9220,N_6886,N_7495);
xnor U9221 (N_9221,N_6469,N_7686);
nor U9222 (N_9222,N_6938,N_7967);
nor U9223 (N_9223,N_6303,N_6756);
xnor U9224 (N_9224,N_7674,N_7592);
nor U9225 (N_9225,N_7863,N_6026);
xnor U9226 (N_9226,N_7409,N_7191);
nor U9227 (N_9227,N_7525,N_7065);
nor U9228 (N_9228,N_6975,N_7588);
nor U9229 (N_9229,N_7980,N_7470);
nand U9230 (N_9230,N_6609,N_6758);
xor U9231 (N_9231,N_6090,N_7947);
xor U9232 (N_9232,N_7490,N_6645);
nor U9233 (N_9233,N_6201,N_6541);
and U9234 (N_9234,N_7899,N_6650);
nor U9235 (N_9235,N_6129,N_7738);
nand U9236 (N_9236,N_7527,N_7983);
nand U9237 (N_9237,N_6856,N_7422);
nor U9238 (N_9238,N_7658,N_6097);
or U9239 (N_9239,N_6704,N_7472);
or U9240 (N_9240,N_6006,N_6104);
nand U9241 (N_9241,N_6086,N_6208);
xnor U9242 (N_9242,N_7062,N_6949);
nor U9243 (N_9243,N_6284,N_7123);
xnor U9244 (N_9244,N_7816,N_6028);
nand U9245 (N_9245,N_7228,N_7043);
xnor U9246 (N_9246,N_7066,N_6773);
nand U9247 (N_9247,N_6361,N_6371);
nor U9248 (N_9248,N_7076,N_7530);
nor U9249 (N_9249,N_6961,N_6862);
xnor U9250 (N_9250,N_7213,N_7194);
nor U9251 (N_9251,N_7438,N_6219);
nor U9252 (N_9252,N_7990,N_7860);
or U9253 (N_9253,N_6020,N_6304);
xnor U9254 (N_9254,N_6820,N_6706);
xnor U9255 (N_9255,N_6628,N_7381);
xor U9256 (N_9256,N_7613,N_7397);
xnor U9257 (N_9257,N_7065,N_7040);
or U9258 (N_9258,N_6466,N_7714);
or U9259 (N_9259,N_6508,N_6849);
nor U9260 (N_9260,N_7867,N_6526);
nor U9261 (N_9261,N_6907,N_6800);
and U9262 (N_9262,N_6271,N_7768);
or U9263 (N_9263,N_7777,N_7985);
or U9264 (N_9264,N_7112,N_6718);
nor U9265 (N_9265,N_6825,N_7801);
nand U9266 (N_9266,N_6757,N_6840);
nand U9267 (N_9267,N_6240,N_6241);
or U9268 (N_9268,N_7774,N_6598);
xor U9269 (N_9269,N_7148,N_7914);
or U9270 (N_9270,N_6470,N_6706);
nand U9271 (N_9271,N_6794,N_7110);
nand U9272 (N_9272,N_6987,N_6431);
xnor U9273 (N_9273,N_7669,N_6555);
xnor U9274 (N_9274,N_6778,N_6615);
or U9275 (N_9275,N_6260,N_6037);
nor U9276 (N_9276,N_6760,N_6492);
xnor U9277 (N_9277,N_6301,N_6787);
nor U9278 (N_9278,N_7133,N_7701);
nor U9279 (N_9279,N_7243,N_7198);
or U9280 (N_9280,N_7428,N_7936);
and U9281 (N_9281,N_7756,N_6164);
and U9282 (N_9282,N_7418,N_7393);
or U9283 (N_9283,N_6196,N_7737);
nor U9284 (N_9284,N_6135,N_6377);
and U9285 (N_9285,N_7296,N_7511);
nand U9286 (N_9286,N_6154,N_7590);
nand U9287 (N_9287,N_7490,N_6596);
nand U9288 (N_9288,N_7284,N_7818);
nand U9289 (N_9289,N_6774,N_6485);
nor U9290 (N_9290,N_6899,N_6473);
or U9291 (N_9291,N_7530,N_7419);
nand U9292 (N_9292,N_7967,N_6400);
and U9293 (N_9293,N_7939,N_7910);
and U9294 (N_9294,N_6411,N_6046);
xnor U9295 (N_9295,N_6784,N_6181);
and U9296 (N_9296,N_6469,N_7478);
xor U9297 (N_9297,N_7999,N_6151);
nand U9298 (N_9298,N_7470,N_6161);
xnor U9299 (N_9299,N_6145,N_7001);
and U9300 (N_9300,N_7441,N_7582);
xnor U9301 (N_9301,N_6641,N_6048);
xor U9302 (N_9302,N_7794,N_6659);
nor U9303 (N_9303,N_7416,N_6706);
nand U9304 (N_9304,N_6089,N_6081);
and U9305 (N_9305,N_6175,N_6773);
and U9306 (N_9306,N_6971,N_7272);
nand U9307 (N_9307,N_7529,N_7547);
nand U9308 (N_9308,N_7651,N_6989);
or U9309 (N_9309,N_6247,N_6653);
nor U9310 (N_9310,N_7447,N_6223);
and U9311 (N_9311,N_6401,N_7412);
xnor U9312 (N_9312,N_6427,N_7098);
and U9313 (N_9313,N_7136,N_6054);
nor U9314 (N_9314,N_7738,N_7353);
xnor U9315 (N_9315,N_6834,N_6929);
nand U9316 (N_9316,N_6191,N_7437);
and U9317 (N_9317,N_6682,N_7564);
xnor U9318 (N_9318,N_7972,N_6576);
nand U9319 (N_9319,N_6914,N_6014);
nand U9320 (N_9320,N_7267,N_6904);
xnor U9321 (N_9321,N_6871,N_7883);
or U9322 (N_9322,N_6583,N_7619);
and U9323 (N_9323,N_7086,N_6097);
and U9324 (N_9324,N_7323,N_6662);
nand U9325 (N_9325,N_7573,N_6173);
and U9326 (N_9326,N_6759,N_7120);
nand U9327 (N_9327,N_6605,N_7962);
or U9328 (N_9328,N_7354,N_6079);
or U9329 (N_9329,N_6965,N_6092);
xor U9330 (N_9330,N_7364,N_6528);
and U9331 (N_9331,N_6681,N_7921);
xor U9332 (N_9332,N_7752,N_6246);
nor U9333 (N_9333,N_7786,N_6199);
and U9334 (N_9334,N_6252,N_6373);
and U9335 (N_9335,N_6187,N_7980);
and U9336 (N_9336,N_7435,N_7889);
xnor U9337 (N_9337,N_6585,N_7654);
xor U9338 (N_9338,N_6084,N_7321);
and U9339 (N_9339,N_7366,N_6305);
xnor U9340 (N_9340,N_7757,N_6698);
or U9341 (N_9341,N_7110,N_7199);
nor U9342 (N_9342,N_6937,N_6932);
and U9343 (N_9343,N_7306,N_6016);
xor U9344 (N_9344,N_6401,N_6429);
or U9345 (N_9345,N_6328,N_7416);
nand U9346 (N_9346,N_6176,N_7974);
nor U9347 (N_9347,N_7118,N_7475);
nor U9348 (N_9348,N_7667,N_6981);
or U9349 (N_9349,N_6486,N_7038);
nand U9350 (N_9350,N_6127,N_6059);
nor U9351 (N_9351,N_7004,N_6452);
nand U9352 (N_9352,N_6430,N_6698);
nor U9353 (N_9353,N_7932,N_7429);
nor U9354 (N_9354,N_6514,N_7448);
nand U9355 (N_9355,N_7575,N_6627);
or U9356 (N_9356,N_7170,N_7212);
xor U9357 (N_9357,N_7462,N_6450);
and U9358 (N_9358,N_6125,N_6785);
nor U9359 (N_9359,N_6588,N_7592);
xor U9360 (N_9360,N_7522,N_6340);
and U9361 (N_9361,N_6766,N_7501);
xor U9362 (N_9362,N_7418,N_7645);
and U9363 (N_9363,N_7127,N_6884);
xnor U9364 (N_9364,N_7556,N_6669);
nor U9365 (N_9365,N_6829,N_6708);
and U9366 (N_9366,N_7284,N_7805);
nand U9367 (N_9367,N_6594,N_6983);
nand U9368 (N_9368,N_6307,N_7537);
nand U9369 (N_9369,N_7513,N_7281);
nor U9370 (N_9370,N_6326,N_7965);
xor U9371 (N_9371,N_6881,N_6439);
and U9372 (N_9372,N_6680,N_7057);
and U9373 (N_9373,N_7072,N_7581);
or U9374 (N_9374,N_6837,N_6164);
and U9375 (N_9375,N_7348,N_6323);
nand U9376 (N_9376,N_6775,N_6073);
and U9377 (N_9377,N_6245,N_7455);
nor U9378 (N_9378,N_7830,N_6560);
nand U9379 (N_9379,N_6601,N_7497);
or U9380 (N_9380,N_6370,N_6706);
nand U9381 (N_9381,N_6731,N_7280);
and U9382 (N_9382,N_7973,N_6289);
nand U9383 (N_9383,N_6622,N_7167);
nand U9384 (N_9384,N_6083,N_6135);
or U9385 (N_9385,N_6155,N_6757);
xor U9386 (N_9386,N_6293,N_6158);
nand U9387 (N_9387,N_7475,N_7398);
and U9388 (N_9388,N_7264,N_7683);
or U9389 (N_9389,N_6275,N_7780);
nand U9390 (N_9390,N_6823,N_7051);
nor U9391 (N_9391,N_7409,N_7550);
nand U9392 (N_9392,N_6548,N_6604);
nand U9393 (N_9393,N_7837,N_7097);
and U9394 (N_9394,N_6792,N_7471);
nor U9395 (N_9395,N_7800,N_6523);
xnor U9396 (N_9396,N_6548,N_6939);
nand U9397 (N_9397,N_7934,N_6090);
and U9398 (N_9398,N_6045,N_7120);
nand U9399 (N_9399,N_6372,N_7022);
and U9400 (N_9400,N_6088,N_7629);
xor U9401 (N_9401,N_7388,N_7097);
nor U9402 (N_9402,N_7855,N_7123);
and U9403 (N_9403,N_7308,N_6719);
or U9404 (N_9404,N_6866,N_7825);
nor U9405 (N_9405,N_6200,N_7587);
nor U9406 (N_9406,N_6268,N_7800);
nand U9407 (N_9407,N_7800,N_7140);
xor U9408 (N_9408,N_6069,N_6236);
nor U9409 (N_9409,N_7083,N_6154);
nor U9410 (N_9410,N_7224,N_7764);
nand U9411 (N_9411,N_6246,N_7091);
and U9412 (N_9412,N_6498,N_6394);
or U9413 (N_9413,N_7278,N_6247);
or U9414 (N_9414,N_7111,N_7449);
and U9415 (N_9415,N_6793,N_7283);
and U9416 (N_9416,N_7261,N_7881);
and U9417 (N_9417,N_6647,N_6367);
and U9418 (N_9418,N_6538,N_6579);
and U9419 (N_9419,N_7637,N_7727);
xnor U9420 (N_9420,N_6953,N_6271);
nand U9421 (N_9421,N_7997,N_6334);
xor U9422 (N_9422,N_6602,N_7136);
xor U9423 (N_9423,N_6270,N_7369);
xor U9424 (N_9424,N_7124,N_7382);
nand U9425 (N_9425,N_6900,N_7493);
or U9426 (N_9426,N_6792,N_7843);
nor U9427 (N_9427,N_6679,N_6705);
or U9428 (N_9428,N_7322,N_6169);
and U9429 (N_9429,N_6982,N_7283);
or U9430 (N_9430,N_7618,N_7904);
and U9431 (N_9431,N_7258,N_6975);
nor U9432 (N_9432,N_6614,N_7914);
and U9433 (N_9433,N_6087,N_6740);
xor U9434 (N_9434,N_6521,N_7554);
xor U9435 (N_9435,N_6442,N_7586);
nand U9436 (N_9436,N_6748,N_7067);
nand U9437 (N_9437,N_6479,N_7910);
xnor U9438 (N_9438,N_6461,N_6361);
nor U9439 (N_9439,N_6577,N_6845);
or U9440 (N_9440,N_7229,N_6787);
xor U9441 (N_9441,N_7845,N_7560);
and U9442 (N_9442,N_6236,N_6145);
xnor U9443 (N_9443,N_7550,N_7560);
or U9444 (N_9444,N_7076,N_6138);
xor U9445 (N_9445,N_6864,N_6374);
nand U9446 (N_9446,N_6140,N_7329);
or U9447 (N_9447,N_6518,N_7295);
xor U9448 (N_9448,N_7272,N_6076);
and U9449 (N_9449,N_6681,N_6153);
nor U9450 (N_9450,N_6123,N_6458);
nand U9451 (N_9451,N_7902,N_6604);
xor U9452 (N_9452,N_7068,N_6324);
nor U9453 (N_9453,N_6725,N_7146);
and U9454 (N_9454,N_6107,N_7787);
or U9455 (N_9455,N_7368,N_6591);
nor U9456 (N_9456,N_7469,N_7603);
xnor U9457 (N_9457,N_6929,N_7710);
xor U9458 (N_9458,N_6900,N_6417);
or U9459 (N_9459,N_7363,N_7708);
xor U9460 (N_9460,N_6250,N_7307);
xnor U9461 (N_9461,N_6283,N_7913);
nand U9462 (N_9462,N_6652,N_7445);
nand U9463 (N_9463,N_6238,N_7857);
xnor U9464 (N_9464,N_7348,N_7037);
or U9465 (N_9465,N_6002,N_6823);
or U9466 (N_9466,N_6795,N_7681);
or U9467 (N_9467,N_6010,N_6793);
nor U9468 (N_9468,N_7826,N_6788);
nor U9469 (N_9469,N_6163,N_7734);
nor U9470 (N_9470,N_7809,N_6008);
and U9471 (N_9471,N_6383,N_6777);
xnor U9472 (N_9472,N_6576,N_6324);
or U9473 (N_9473,N_6084,N_7082);
nand U9474 (N_9474,N_6373,N_7578);
and U9475 (N_9475,N_6396,N_6375);
or U9476 (N_9476,N_7522,N_6282);
and U9477 (N_9477,N_6367,N_6685);
and U9478 (N_9478,N_7401,N_7073);
nor U9479 (N_9479,N_6733,N_7494);
xor U9480 (N_9480,N_7222,N_7205);
nor U9481 (N_9481,N_6552,N_7902);
or U9482 (N_9482,N_6600,N_7082);
and U9483 (N_9483,N_6779,N_6562);
and U9484 (N_9484,N_7115,N_7913);
and U9485 (N_9485,N_7929,N_6003);
nand U9486 (N_9486,N_7317,N_7399);
or U9487 (N_9487,N_7982,N_6943);
nand U9488 (N_9488,N_6955,N_7746);
and U9489 (N_9489,N_6338,N_7606);
and U9490 (N_9490,N_6889,N_7224);
nand U9491 (N_9491,N_6785,N_7668);
nor U9492 (N_9492,N_7196,N_6885);
and U9493 (N_9493,N_7349,N_6289);
nand U9494 (N_9494,N_7981,N_6210);
or U9495 (N_9495,N_6157,N_7313);
xor U9496 (N_9496,N_7735,N_7469);
nor U9497 (N_9497,N_7937,N_6366);
xor U9498 (N_9498,N_6586,N_7968);
nand U9499 (N_9499,N_6050,N_6769);
or U9500 (N_9500,N_7164,N_6832);
nor U9501 (N_9501,N_6091,N_6720);
nand U9502 (N_9502,N_7108,N_7843);
nand U9503 (N_9503,N_7605,N_6435);
nor U9504 (N_9504,N_6647,N_6312);
or U9505 (N_9505,N_7756,N_6719);
or U9506 (N_9506,N_6826,N_7609);
or U9507 (N_9507,N_7569,N_7950);
nor U9508 (N_9508,N_6910,N_6839);
nand U9509 (N_9509,N_7265,N_7261);
nor U9510 (N_9510,N_7098,N_6600);
xor U9511 (N_9511,N_6822,N_7404);
and U9512 (N_9512,N_6658,N_7044);
nor U9513 (N_9513,N_7703,N_7457);
or U9514 (N_9514,N_6672,N_7791);
nand U9515 (N_9515,N_6265,N_7683);
nor U9516 (N_9516,N_7189,N_7882);
and U9517 (N_9517,N_6272,N_7479);
nor U9518 (N_9518,N_7172,N_7415);
xor U9519 (N_9519,N_6686,N_6400);
xor U9520 (N_9520,N_6685,N_6871);
or U9521 (N_9521,N_6174,N_6914);
and U9522 (N_9522,N_7488,N_7947);
nor U9523 (N_9523,N_7422,N_7993);
nor U9524 (N_9524,N_7291,N_7732);
nand U9525 (N_9525,N_7826,N_7726);
and U9526 (N_9526,N_6927,N_6049);
and U9527 (N_9527,N_7091,N_6433);
xnor U9528 (N_9528,N_7174,N_6367);
nor U9529 (N_9529,N_7683,N_6791);
xor U9530 (N_9530,N_6836,N_6899);
nor U9531 (N_9531,N_7729,N_6859);
and U9532 (N_9532,N_7692,N_7066);
xor U9533 (N_9533,N_7382,N_7101);
and U9534 (N_9534,N_7354,N_7327);
and U9535 (N_9535,N_7140,N_7952);
and U9536 (N_9536,N_7845,N_7741);
xor U9537 (N_9537,N_7672,N_6787);
nor U9538 (N_9538,N_6546,N_6143);
or U9539 (N_9539,N_6267,N_7562);
or U9540 (N_9540,N_6306,N_6638);
xnor U9541 (N_9541,N_6211,N_6434);
or U9542 (N_9542,N_6453,N_6459);
xor U9543 (N_9543,N_6261,N_7380);
xnor U9544 (N_9544,N_7927,N_6828);
nand U9545 (N_9545,N_6831,N_7993);
or U9546 (N_9546,N_7491,N_7854);
xor U9547 (N_9547,N_6299,N_6833);
nand U9548 (N_9548,N_7705,N_7060);
nand U9549 (N_9549,N_6571,N_7524);
and U9550 (N_9550,N_7642,N_6102);
and U9551 (N_9551,N_6821,N_6848);
xor U9552 (N_9552,N_7808,N_6796);
and U9553 (N_9553,N_6361,N_6078);
or U9554 (N_9554,N_7301,N_7657);
nor U9555 (N_9555,N_7613,N_7730);
nand U9556 (N_9556,N_7145,N_7122);
nand U9557 (N_9557,N_7767,N_7331);
nand U9558 (N_9558,N_7592,N_7591);
nor U9559 (N_9559,N_6896,N_7123);
xnor U9560 (N_9560,N_6155,N_7443);
nand U9561 (N_9561,N_6902,N_7544);
and U9562 (N_9562,N_6649,N_6850);
nand U9563 (N_9563,N_7439,N_6316);
or U9564 (N_9564,N_6720,N_7726);
nand U9565 (N_9565,N_7224,N_7115);
xnor U9566 (N_9566,N_7278,N_6484);
nor U9567 (N_9567,N_7232,N_7260);
nand U9568 (N_9568,N_6577,N_7171);
xnor U9569 (N_9569,N_6881,N_7014);
nand U9570 (N_9570,N_7101,N_7277);
xor U9571 (N_9571,N_7760,N_6005);
nand U9572 (N_9572,N_7987,N_7286);
nand U9573 (N_9573,N_7841,N_6112);
nor U9574 (N_9574,N_6269,N_6587);
or U9575 (N_9575,N_7050,N_7944);
nand U9576 (N_9576,N_6624,N_7843);
xnor U9577 (N_9577,N_7295,N_6169);
xnor U9578 (N_9578,N_7535,N_7213);
and U9579 (N_9579,N_7543,N_6933);
nand U9580 (N_9580,N_6824,N_7708);
and U9581 (N_9581,N_7490,N_6306);
nor U9582 (N_9582,N_7453,N_7279);
or U9583 (N_9583,N_6791,N_6161);
xnor U9584 (N_9584,N_7327,N_7274);
and U9585 (N_9585,N_7033,N_7312);
nor U9586 (N_9586,N_7725,N_7699);
xnor U9587 (N_9587,N_6456,N_6457);
and U9588 (N_9588,N_6457,N_6017);
xor U9589 (N_9589,N_6408,N_6604);
or U9590 (N_9590,N_7305,N_7494);
xor U9591 (N_9591,N_6736,N_7409);
nand U9592 (N_9592,N_7100,N_7572);
nor U9593 (N_9593,N_7336,N_6380);
xnor U9594 (N_9594,N_6915,N_7094);
and U9595 (N_9595,N_6656,N_6516);
nor U9596 (N_9596,N_7845,N_6463);
xnor U9597 (N_9597,N_6921,N_6897);
nand U9598 (N_9598,N_7237,N_6341);
and U9599 (N_9599,N_7178,N_7084);
xor U9600 (N_9600,N_7768,N_7196);
nand U9601 (N_9601,N_6832,N_6050);
or U9602 (N_9602,N_6394,N_6597);
nor U9603 (N_9603,N_6740,N_7420);
nand U9604 (N_9604,N_6725,N_7110);
and U9605 (N_9605,N_6892,N_7866);
xnor U9606 (N_9606,N_7713,N_7480);
nor U9607 (N_9607,N_6233,N_7738);
nor U9608 (N_9608,N_6080,N_6796);
and U9609 (N_9609,N_7934,N_6411);
nor U9610 (N_9610,N_7935,N_7821);
or U9611 (N_9611,N_6872,N_7124);
xor U9612 (N_9612,N_6039,N_7802);
or U9613 (N_9613,N_6745,N_6177);
xnor U9614 (N_9614,N_7658,N_7454);
nor U9615 (N_9615,N_6062,N_7226);
xnor U9616 (N_9616,N_7239,N_6662);
nand U9617 (N_9617,N_6460,N_7956);
nor U9618 (N_9618,N_7605,N_7773);
xor U9619 (N_9619,N_7529,N_6322);
xor U9620 (N_9620,N_7996,N_6555);
nand U9621 (N_9621,N_7551,N_7665);
xor U9622 (N_9622,N_6340,N_6406);
or U9623 (N_9623,N_7010,N_6664);
nor U9624 (N_9624,N_7258,N_6504);
xnor U9625 (N_9625,N_7592,N_6618);
and U9626 (N_9626,N_7420,N_6123);
and U9627 (N_9627,N_6713,N_6478);
or U9628 (N_9628,N_7858,N_6235);
xor U9629 (N_9629,N_7930,N_7276);
nand U9630 (N_9630,N_6494,N_7260);
nand U9631 (N_9631,N_7267,N_6440);
xor U9632 (N_9632,N_6713,N_6856);
nand U9633 (N_9633,N_7564,N_7406);
and U9634 (N_9634,N_6926,N_6985);
xor U9635 (N_9635,N_7271,N_6451);
and U9636 (N_9636,N_7581,N_6384);
xnor U9637 (N_9637,N_6281,N_7532);
or U9638 (N_9638,N_7799,N_6211);
nor U9639 (N_9639,N_7651,N_6359);
nand U9640 (N_9640,N_6164,N_6039);
nor U9641 (N_9641,N_6476,N_6493);
nand U9642 (N_9642,N_7043,N_6464);
xor U9643 (N_9643,N_6234,N_7658);
xor U9644 (N_9644,N_6710,N_6827);
or U9645 (N_9645,N_6072,N_6479);
and U9646 (N_9646,N_7255,N_6722);
and U9647 (N_9647,N_6374,N_7755);
nor U9648 (N_9648,N_7068,N_7661);
or U9649 (N_9649,N_7139,N_7377);
nor U9650 (N_9650,N_7193,N_6876);
xnor U9651 (N_9651,N_6105,N_7781);
and U9652 (N_9652,N_6406,N_7022);
or U9653 (N_9653,N_6399,N_6871);
or U9654 (N_9654,N_7550,N_6779);
xnor U9655 (N_9655,N_7858,N_7384);
or U9656 (N_9656,N_7473,N_7681);
or U9657 (N_9657,N_6211,N_7531);
nand U9658 (N_9658,N_7650,N_6969);
or U9659 (N_9659,N_6331,N_7397);
nor U9660 (N_9660,N_6390,N_7091);
and U9661 (N_9661,N_6268,N_6411);
nand U9662 (N_9662,N_7050,N_6364);
or U9663 (N_9663,N_6871,N_7514);
xnor U9664 (N_9664,N_6648,N_6245);
nand U9665 (N_9665,N_6650,N_7217);
nand U9666 (N_9666,N_7115,N_6068);
xor U9667 (N_9667,N_6378,N_7590);
and U9668 (N_9668,N_7751,N_6219);
or U9669 (N_9669,N_6007,N_7924);
and U9670 (N_9670,N_7396,N_6511);
and U9671 (N_9671,N_6512,N_6681);
nand U9672 (N_9672,N_6953,N_6632);
or U9673 (N_9673,N_7222,N_6049);
nor U9674 (N_9674,N_7798,N_7228);
or U9675 (N_9675,N_6747,N_6674);
xor U9676 (N_9676,N_7376,N_6573);
xnor U9677 (N_9677,N_7636,N_6259);
xor U9678 (N_9678,N_6021,N_6046);
nand U9679 (N_9679,N_7495,N_7653);
nor U9680 (N_9680,N_6053,N_6251);
or U9681 (N_9681,N_6622,N_6092);
xor U9682 (N_9682,N_7508,N_7235);
or U9683 (N_9683,N_7451,N_7295);
xor U9684 (N_9684,N_6459,N_6312);
nand U9685 (N_9685,N_6175,N_6239);
nor U9686 (N_9686,N_6797,N_7003);
nor U9687 (N_9687,N_7295,N_7971);
xnor U9688 (N_9688,N_7317,N_7105);
or U9689 (N_9689,N_7220,N_6188);
and U9690 (N_9690,N_6212,N_6317);
xor U9691 (N_9691,N_6647,N_7330);
xor U9692 (N_9692,N_6781,N_6123);
nand U9693 (N_9693,N_7391,N_7262);
and U9694 (N_9694,N_7343,N_6108);
nor U9695 (N_9695,N_6022,N_7227);
and U9696 (N_9696,N_7038,N_6367);
nor U9697 (N_9697,N_6181,N_6617);
nand U9698 (N_9698,N_6266,N_7860);
and U9699 (N_9699,N_7547,N_7394);
nand U9700 (N_9700,N_7488,N_6679);
and U9701 (N_9701,N_6685,N_6732);
and U9702 (N_9702,N_6497,N_7432);
xor U9703 (N_9703,N_7236,N_7738);
nand U9704 (N_9704,N_6003,N_6726);
and U9705 (N_9705,N_6119,N_7727);
nand U9706 (N_9706,N_6481,N_7924);
or U9707 (N_9707,N_6948,N_6604);
nand U9708 (N_9708,N_7819,N_7826);
or U9709 (N_9709,N_6523,N_7129);
nor U9710 (N_9710,N_7919,N_7619);
or U9711 (N_9711,N_6204,N_7839);
nand U9712 (N_9712,N_7840,N_7143);
nor U9713 (N_9713,N_7506,N_7046);
and U9714 (N_9714,N_6260,N_6522);
xnor U9715 (N_9715,N_7492,N_6841);
and U9716 (N_9716,N_7346,N_6007);
nor U9717 (N_9717,N_7660,N_7919);
xnor U9718 (N_9718,N_6762,N_7714);
nor U9719 (N_9719,N_6169,N_7187);
or U9720 (N_9720,N_6162,N_7111);
nor U9721 (N_9721,N_7515,N_6916);
and U9722 (N_9722,N_6104,N_7057);
or U9723 (N_9723,N_6726,N_7313);
nor U9724 (N_9724,N_7063,N_6089);
nand U9725 (N_9725,N_6172,N_6161);
xor U9726 (N_9726,N_7268,N_6495);
and U9727 (N_9727,N_6462,N_7418);
and U9728 (N_9728,N_7948,N_7822);
xnor U9729 (N_9729,N_6002,N_7457);
or U9730 (N_9730,N_6767,N_6151);
xnor U9731 (N_9731,N_7610,N_7319);
nor U9732 (N_9732,N_7870,N_7930);
xor U9733 (N_9733,N_6806,N_6220);
xnor U9734 (N_9734,N_6118,N_7511);
or U9735 (N_9735,N_6224,N_7176);
xnor U9736 (N_9736,N_6562,N_7612);
and U9737 (N_9737,N_7268,N_6056);
nor U9738 (N_9738,N_7786,N_6270);
and U9739 (N_9739,N_6436,N_7458);
nand U9740 (N_9740,N_6382,N_7185);
nand U9741 (N_9741,N_7026,N_6965);
and U9742 (N_9742,N_7887,N_7732);
nor U9743 (N_9743,N_7913,N_6837);
nor U9744 (N_9744,N_7188,N_6529);
xor U9745 (N_9745,N_6103,N_6212);
nor U9746 (N_9746,N_7804,N_6470);
xnor U9747 (N_9747,N_7979,N_7288);
xor U9748 (N_9748,N_7132,N_7847);
xnor U9749 (N_9749,N_6347,N_6116);
nor U9750 (N_9750,N_7905,N_7204);
nand U9751 (N_9751,N_6461,N_6333);
nand U9752 (N_9752,N_7342,N_7505);
xor U9753 (N_9753,N_6528,N_7345);
xnor U9754 (N_9754,N_6074,N_7476);
xnor U9755 (N_9755,N_7823,N_7185);
nor U9756 (N_9756,N_7329,N_6951);
nor U9757 (N_9757,N_7255,N_6729);
or U9758 (N_9758,N_7137,N_6793);
nor U9759 (N_9759,N_6973,N_7320);
and U9760 (N_9760,N_6491,N_7812);
nor U9761 (N_9761,N_7115,N_7571);
or U9762 (N_9762,N_6156,N_6097);
xnor U9763 (N_9763,N_6505,N_7190);
xnor U9764 (N_9764,N_7039,N_7577);
nor U9765 (N_9765,N_7742,N_7947);
xnor U9766 (N_9766,N_7698,N_7155);
or U9767 (N_9767,N_6077,N_6127);
or U9768 (N_9768,N_7046,N_7341);
and U9769 (N_9769,N_7445,N_7335);
or U9770 (N_9770,N_6187,N_7669);
xor U9771 (N_9771,N_6206,N_7437);
and U9772 (N_9772,N_6802,N_7093);
xor U9773 (N_9773,N_7593,N_7374);
nor U9774 (N_9774,N_6057,N_7881);
nor U9775 (N_9775,N_6668,N_7327);
nor U9776 (N_9776,N_7776,N_7766);
nand U9777 (N_9777,N_6760,N_6382);
or U9778 (N_9778,N_6939,N_7254);
xnor U9779 (N_9779,N_6135,N_7313);
nor U9780 (N_9780,N_6477,N_7347);
xor U9781 (N_9781,N_7774,N_7012);
nand U9782 (N_9782,N_6598,N_7308);
and U9783 (N_9783,N_7837,N_6108);
nand U9784 (N_9784,N_6531,N_7164);
nand U9785 (N_9785,N_7622,N_7603);
nand U9786 (N_9786,N_7942,N_6863);
or U9787 (N_9787,N_7615,N_6321);
or U9788 (N_9788,N_7767,N_6708);
nor U9789 (N_9789,N_6851,N_7501);
or U9790 (N_9790,N_6386,N_6419);
nor U9791 (N_9791,N_7034,N_6215);
or U9792 (N_9792,N_7670,N_7691);
xnor U9793 (N_9793,N_6848,N_7514);
and U9794 (N_9794,N_6874,N_7970);
and U9795 (N_9795,N_6983,N_6800);
nor U9796 (N_9796,N_6468,N_7091);
or U9797 (N_9797,N_6899,N_6864);
and U9798 (N_9798,N_6158,N_6375);
or U9799 (N_9799,N_7099,N_6996);
nor U9800 (N_9800,N_7351,N_6814);
nor U9801 (N_9801,N_6222,N_7310);
and U9802 (N_9802,N_7932,N_7494);
nor U9803 (N_9803,N_7855,N_7635);
or U9804 (N_9804,N_7501,N_6059);
and U9805 (N_9805,N_6949,N_6474);
and U9806 (N_9806,N_6830,N_6646);
nor U9807 (N_9807,N_6967,N_6162);
and U9808 (N_9808,N_7015,N_6720);
and U9809 (N_9809,N_7696,N_7571);
xor U9810 (N_9810,N_6247,N_6841);
and U9811 (N_9811,N_7010,N_6159);
xnor U9812 (N_9812,N_6730,N_7591);
xnor U9813 (N_9813,N_7354,N_6623);
nor U9814 (N_9814,N_6308,N_7735);
and U9815 (N_9815,N_7327,N_6196);
or U9816 (N_9816,N_6272,N_6443);
nor U9817 (N_9817,N_6777,N_6317);
or U9818 (N_9818,N_7585,N_7163);
nand U9819 (N_9819,N_6212,N_7576);
and U9820 (N_9820,N_6764,N_7991);
and U9821 (N_9821,N_7283,N_6172);
or U9822 (N_9822,N_7154,N_7885);
and U9823 (N_9823,N_6842,N_7067);
or U9824 (N_9824,N_6442,N_7604);
nor U9825 (N_9825,N_6904,N_7003);
and U9826 (N_9826,N_6575,N_6998);
nand U9827 (N_9827,N_6671,N_6170);
nand U9828 (N_9828,N_6777,N_7846);
nand U9829 (N_9829,N_6340,N_7640);
or U9830 (N_9830,N_7733,N_6998);
and U9831 (N_9831,N_7753,N_6656);
nand U9832 (N_9832,N_6012,N_7668);
and U9833 (N_9833,N_7702,N_7291);
nor U9834 (N_9834,N_6609,N_6904);
xor U9835 (N_9835,N_7975,N_7566);
nand U9836 (N_9836,N_7459,N_7754);
and U9837 (N_9837,N_6591,N_7823);
and U9838 (N_9838,N_7718,N_6340);
xnor U9839 (N_9839,N_7326,N_7399);
and U9840 (N_9840,N_7778,N_6510);
xor U9841 (N_9841,N_6285,N_6889);
and U9842 (N_9842,N_7138,N_6459);
and U9843 (N_9843,N_7982,N_6471);
xor U9844 (N_9844,N_7211,N_6786);
nand U9845 (N_9845,N_6461,N_6726);
nor U9846 (N_9846,N_7425,N_6019);
xnor U9847 (N_9847,N_7387,N_6146);
nor U9848 (N_9848,N_6661,N_6143);
nand U9849 (N_9849,N_7484,N_6999);
nand U9850 (N_9850,N_7103,N_7131);
or U9851 (N_9851,N_7610,N_6122);
nand U9852 (N_9852,N_6995,N_6030);
xnor U9853 (N_9853,N_6243,N_6189);
xnor U9854 (N_9854,N_7696,N_6784);
xor U9855 (N_9855,N_7569,N_7125);
nor U9856 (N_9856,N_7596,N_7944);
nand U9857 (N_9857,N_6337,N_7559);
xnor U9858 (N_9858,N_6472,N_6549);
or U9859 (N_9859,N_7210,N_6663);
xnor U9860 (N_9860,N_6359,N_6986);
xnor U9861 (N_9861,N_6223,N_7104);
xnor U9862 (N_9862,N_7163,N_6096);
nand U9863 (N_9863,N_7523,N_6728);
xnor U9864 (N_9864,N_6639,N_6110);
nor U9865 (N_9865,N_7607,N_6722);
or U9866 (N_9866,N_7160,N_6464);
xor U9867 (N_9867,N_7887,N_7104);
xor U9868 (N_9868,N_6779,N_6125);
or U9869 (N_9869,N_7405,N_6848);
nor U9870 (N_9870,N_7046,N_6734);
xor U9871 (N_9871,N_6974,N_7521);
or U9872 (N_9872,N_6718,N_6600);
or U9873 (N_9873,N_7245,N_7741);
nand U9874 (N_9874,N_7865,N_7997);
or U9875 (N_9875,N_7863,N_7535);
nor U9876 (N_9876,N_6571,N_7872);
nand U9877 (N_9877,N_7592,N_7748);
nand U9878 (N_9878,N_7643,N_7910);
nand U9879 (N_9879,N_7482,N_7772);
nand U9880 (N_9880,N_6838,N_7439);
xnor U9881 (N_9881,N_6150,N_6454);
xor U9882 (N_9882,N_7421,N_6499);
xor U9883 (N_9883,N_7414,N_6858);
nand U9884 (N_9884,N_6390,N_6910);
nor U9885 (N_9885,N_6456,N_7179);
and U9886 (N_9886,N_6498,N_6819);
nand U9887 (N_9887,N_6799,N_7999);
nand U9888 (N_9888,N_6580,N_7826);
and U9889 (N_9889,N_6917,N_7183);
nand U9890 (N_9890,N_6521,N_7237);
nand U9891 (N_9891,N_7012,N_6202);
xor U9892 (N_9892,N_6442,N_6897);
and U9893 (N_9893,N_7893,N_7719);
and U9894 (N_9894,N_7339,N_7210);
xor U9895 (N_9895,N_6978,N_7011);
and U9896 (N_9896,N_7603,N_7053);
nor U9897 (N_9897,N_6008,N_6835);
nand U9898 (N_9898,N_7762,N_6617);
or U9899 (N_9899,N_6588,N_7720);
or U9900 (N_9900,N_6495,N_7777);
nand U9901 (N_9901,N_7910,N_6830);
nand U9902 (N_9902,N_7431,N_6647);
or U9903 (N_9903,N_7782,N_7945);
or U9904 (N_9904,N_6831,N_7125);
nand U9905 (N_9905,N_6399,N_6575);
or U9906 (N_9906,N_7175,N_7030);
or U9907 (N_9907,N_6849,N_7718);
nor U9908 (N_9908,N_7494,N_6701);
xor U9909 (N_9909,N_7447,N_7542);
nor U9910 (N_9910,N_7640,N_6990);
nor U9911 (N_9911,N_6232,N_7587);
or U9912 (N_9912,N_6195,N_6196);
nor U9913 (N_9913,N_6074,N_7044);
nor U9914 (N_9914,N_7485,N_7478);
nand U9915 (N_9915,N_6256,N_7761);
and U9916 (N_9916,N_6668,N_6923);
nand U9917 (N_9917,N_6156,N_6003);
xor U9918 (N_9918,N_6532,N_6869);
nor U9919 (N_9919,N_7908,N_7909);
nand U9920 (N_9920,N_6182,N_6762);
and U9921 (N_9921,N_7406,N_6212);
nand U9922 (N_9922,N_7554,N_7641);
or U9923 (N_9923,N_6213,N_6721);
and U9924 (N_9924,N_7073,N_7674);
and U9925 (N_9925,N_7867,N_6787);
nand U9926 (N_9926,N_6975,N_6523);
or U9927 (N_9927,N_6188,N_7949);
or U9928 (N_9928,N_7887,N_6106);
nor U9929 (N_9929,N_7024,N_6444);
xor U9930 (N_9930,N_7293,N_6450);
nand U9931 (N_9931,N_6700,N_7576);
nor U9932 (N_9932,N_7908,N_6245);
or U9933 (N_9933,N_6083,N_6804);
and U9934 (N_9934,N_6807,N_7612);
and U9935 (N_9935,N_7983,N_6053);
and U9936 (N_9936,N_6953,N_6829);
nor U9937 (N_9937,N_6804,N_7212);
and U9938 (N_9938,N_7581,N_6091);
or U9939 (N_9939,N_6044,N_6264);
nand U9940 (N_9940,N_7294,N_7354);
or U9941 (N_9941,N_7535,N_7601);
or U9942 (N_9942,N_7759,N_7188);
xor U9943 (N_9943,N_7227,N_7672);
or U9944 (N_9944,N_7160,N_6755);
nand U9945 (N_9945,N_6676,N_6546);
or U9946 (N_9946,N_6235,N_7049);
xor U9947 (N_9947,N_7896,N_6248);
or U9948 (N_9948,N_6433,N_6168);
nand U9949 (N_9949,N_6799,N_6301);
and U9950 (N_9950,N_7423,N_6261);
nand U9951 (N_9951,N_6005,N_7888);
and U9952 (N_9952,N_6559,N_7309);
and U9953 (N_9953,N_6639,N_7613);
or U9954 (N_9954,N_7612,N_7097);
or U9955 (N_9955,N_6689,N_6079);
xnor U9956 (N_9956,N_7135,N_6879);
nand U9957 (N_9957,N_7323,N_6715);
nor U9958 (N_9958,N_7653,N_7703);
xnor U9959 (N_9959,N_6815,N_6986);
nor U9960 (N_9960,N_6668,N_6027);
and U9961 (N_9961,N_6422,N_7433);
nand U9962 (N_9962,N_7400,N_7593);
nand U9963 (N_9963,N_7143,N_6563);
nor U9964 (N_9964,N_6527,N_6935);
xor U9965 (N_9965,N_6622,N_6137);
and U9966 (N_9966,N_6012,N_6599);
xor U9967 (N_9967,N_6173,N_7477);
nand U9968 (N_9968,N_7165,N_7337);
or U9969 (N_9969,N_7922,N_6564);
nor U9970 (N_9970,N_6093,N_7315);
nand U9971 (N_9971,N_6245,N_6418);
and U9972 (N_9972,N_6648,N_6539);
nor U9973 (N_9973,N_6035,N_6238);
or U9974 (N_9974,N_6237,N_7836);
nand U9975 (N_9975,N_7903,N_7127);
xnor U9976 (N_9976,N_6349,N_7970);
nor U9977 (N_9977,N_6459,N_7738);
or U9978 (N_9978,N_7763,N_6573);
xnor U9979 (N_9979,N_6741,N_6037);
xnor U9980 (N_9980,N_6412,N_7351);
nor U9981 (N_9981,N_7914,N_6579);
nor U9982 (N_9982,N_6842,N_7608);
nor U9983 (N_9983,N_6837,N_7954);
xnor U9984 (N_9984,N_7356,N_6976);
nor U9985 (N_9985,N_7363,N_7217);
and U9986 (N_9986,N_7411,N_6937);
xor U9987 (N_9987,N_7970,N_6551);
or U9988 (N_9988,N_6918,N_6876);
and U9989 (N_9989,N_6809,N_6293);
or U9990 (N_9990,N_7206,N_7502);
xor U9991 (N_9991,N_6736,N_6393);
nor U9992 (N_9992,N_6138,N_6978);
nand U9993 (N_9993,N_7112,N_6393);
nand U9994 (N_9994,N_6417,N_7275);
or U9995 (N_9995,N_6904,N_7820);
nor U9996 (N_9996,N_7243,N_6443);
xor U9997 (N_9997,N_7019,N_6238);
xnor U9998 (N_9998,N_6253,N_6930);
and U9999 (N_9999,N_6188,N_6730);
and U10000 (N_10000,N_9847,N_8299);
or U10001 (N_10001,N_8040,N_9693);
xor U10002 (N_10002,N_8292,N_9743);
xor U10003 (N_10003,N_8029,N_8275);
or U10004 (N_10004,N_8910,N_8894);
nor U10005 (N_10005,N_9642,N_9118);
xnor U10006 (N_10006,N_9413,N_9604);
or U10007 (N_10007,N_8016,N_8764);
xnor U10008 (N_10008,N_9956,N_9150);
and U10009 (N_10009,N_8484,N_8893);
and U10010 (N_10010,N_8466,N_8491);
nand U10011 (N_10011,N_9835,N_9176);
or U10012 (N_10012,N_9982,N_8436);
and U10013 (N_10013,N_8038,N_8816);
and U10014 (N_10014,N_8168,N_9860);
or U10015 (N_10015,N_8662,N_8081);
and U10016 (N_10016,N_8659,N_9997);
or U10017 (N_10017,N_8983,N_9893);
nor U10018 (N_10018,N_9426,N_8594);
or U10019 (N_10019,N_8953,N_8210);
nor U10020 (N_10020,N_9208,N_9363);
nand U10021 (N_10021,N_9650,N_9216);
and U10022 (N_10022,N_8214,N_8088);
nor U10023 (N_10023,N_9553,N_9653);
xnor U10024 (N_10024,N_8061,N_9040);
xnor U10025 (N_10025,N_9338,N_9065);
or U10026 (N_10026,N_8515,N_9283);
and U10027 (N_10027,N_8938,N_8544);
and U10028 (N_10028,N_8514,N_8243);
and U10029 (N_10029,N_9605,N_9629);
and U10030 (N_10030,N_8531,N_8701);
nor U10031 (N_10031,N_8858,N_9213);
and U10032 (N_10032,N_8915,N_8969);
xor U10033 (N_10033,N_8402,N_8583);
and U10034 (N_10034,N_9550,N_8854);
and U10035 (N_10035,N_9498,N_8830);
nand U10036 (N_10036,N_8826,N_8564);
or U10037 (N_10037,N_9073,N_9184);
xor U10038 (N_10038,N_8799,N_9350);
xor U10039 (N_10039,N_9038,N_8288);
nand U10040 (N_10040,N_8434,N_8385);
xor U10041 (N_10041,N_9549,N_9139);
or U10042 (N_10042,N_8154,N_9875);
xor U10043 (N_10043,N_9173,N_8178);
nand U10044 (N_10044,N_9069,N_8062);
or U10045 (N_10045,N_9648,N_9232);
xnor U10046 (N_10046,N_9053,N_9255);
xor U10047 (N_10047,N_8902,N_9037);
or U10048 (N_10048,N_8929,N_8669);
and U10049 (N_10049,N_9921,N_9298);
nor U10050 (N_10050,N_9108,N_9744);
or U10051 (N_10051,N_8539,N_8496);
nor U10052 (N_10052,N_8820,N_9671);
nor U10053 (N_10053,N_8831,N_8507);
or U10054 (N_10054,N_9010,N_8919);
and U10055 (N_10055,N_9947,N_9966);
nor U10056 (N_10056,N_9555,N_8080);
nand U10057 (N_10057,N_8879,N_9247);
or U10058 (N_10058,N_8312,N_8031);
and U10059 (N_10059,N_9480,N_8206);
and U10060 (N_10060,N_8440,N_9584);
xor U10061 (N_10061,N_8205,N_8304);
xor U10062 (N_10062,N_8828,N_9827);
or U10063 (N_10063,N_9696,N_8571);
xnor U10064 (N_10064,N_8432,N_8883);
nand U10065 (N_10065,N_9660,N_8093);
xor U10066 (N_10066,N_9048,N_9406);
nor U10067 (N_10067,N_9026,N_8842);
and U10068 (N_10068,N_8630,N_8503);
and U10069 (N_10069,N_8791,N_8837);
xor U10070 (N_10070,N_9189,N_8013);
or U10071 (N_10071,N_9709,N_9470);
nand U10072 (N_10072,N_9249,N_9858);
xor U10073 (N_10073,N_9017,N_8247);
and U10074 (N_10074,N_9345,N_9270);
and U10075 (N_10075,N_9513,N_9209);
or U10076 (N_10076,N_9282,N_8160);
nor U10077 (N_10077,N_8596,N_9427);
nand U10078 (N_10078,N_8321,N_8931);
nor U10079 (N_10079,N_9746,N_8073);
nor U10080 (N_10080,N_9986,N_8241);
nand U10081 (N_10081,N_8096,N_9909);
nor U10082 (N_10082,N_8132,N_8296);
xor U10083 (N_10083,N_9144,N_8251);
nand U10084 (N_10084,N_9439,N_8227);
and U10085 (N_10085,N_8020,N_9598);
nor U10086 (N_10086,N_8542,N_9075);
and U10087 (N_10087,N_9367,N_8665);
and U10088 (N_10088,N_9294,N_8649);
and U10089 (N_10089,N_8778,N_9083);
or U10090 (N_10090,N_8884,N_8957);
nor U10091 (N_10091,N_9664,N_9318);
nand U10092 (N_10092,N_8933,N_9940);
and U10093 (N_10093,N_8386,N_9867);
xnor U10094 (N_10094,N_9691,N_8360);
or U10095 (N_10095,N_9499,N_8454);
nand U10096 (N_10096,N_9911,N_9398);
and U10097 (N_10097,N_8116,N_9797);
xor U10098 (N_10098,N_8164,N_8054);
and U10099 (N_10099,N_8456,N_9347);
xnor U10100 (N_10100,N_8927,N_8761);
and U10101 (N_10101,N_8622,N_9391);
xnor U10102 (N_10102,N_8954,N_8217);
or U10103 (N_10103,N_8125,N_8479);
nor U10104 (N_10104,N_9475,N_9715);
xnor U10105 (N_10105,N_8122,N_8334);
nor U10106 (N_10106,N_8129,N_9561);
nand U10107 (N_10107,N_8234,N_8283);
nor U10108 (N_10108,N_8417,N_8808);
nor U10109 (N_10109,N_9519,N_9640);
nand U10110 (N_10110,N_8203,N_9755);
xnor U10111 (N_10111,N_9431,N_9225);
nand U10112 (N_10112,N_9938,N_9064);
xnor U10113 (N_10113,N_8091,N_9292);
xor U10114 (N_10114,N_8173,N_9131);
nand U10115 (N_10115,N_8332,N_8645);
nor U10116 (N_10116,N_8448,N_8476);
xnor U10117 (N_10117,N_9996,N_9933);
and U10118 (N_10118,N_8414,N_9138);
or U10119 (N_10119,N_8975,N_8433);
nor U10120 (N_10120,N_9082,N_9865);
nor U10121 (N_10121,N_9424,N_8625);
and U10122 (N_10122,N_9264,N_9178);
xor U10123 (N_10123,N_9133,N_8782);
and U10124 (N_10124,N_9222,N_8555);
and U10125 (N_10125,N_8736,N_9528);
nand U10126 (N_10126,N_8924,N_8756);
and U10127 (N_10127,N_9975,N_8779);
nor U10128 (N_10128,N_8770,N_8917);
or U10129 (N_10129,N_9870,N_9397);
xor U10130 (N_10130,N_9685,N_9830);
xnor U10131 (N_10131,N_9182,N_9285);
and U10132 (N_10132,N_9957,N_9171);
xor U10133 (N_10133,N_8302,N_8875);
xor U10134 (N_10134,N_9316,N_9370);
or U10135 (N_10135,N_9541,N_9085);
or U10136 (N_10136,N_9136,N_9912);
and U10137 (N_10137,N_9942,N_8474);
nor U10138 (N_10138,N_8303,N_9885);
or U10139 (N_10139,N_8968,N_8568);
nand U10140 (N_10140,N_9240,N_8987);
nor U10141 (N_10141,N_8813,N_9889);
nand U10142 (N_10142,N_9970,N_8690);
nand U10143 (N_10143,N_8030,N_8404);
nor U10144 (N_10144,N_9362,N_9619);
or U10145 (N_10145,N_8477,N_9497);
xor U10146 (N_10146,N_8997,N_8546);
nor U10147 (N_10147,N_8469,N_8082);
and U10148 (N_10148,N_9055,N_9606);
and U10149 (N_10149,N_9522,N_8011);
nor U10150 (N_10150,N_9521,N_8783);
nor U10151 (N_10151,N_8156,N_9608);
nor U10152 (N_10152,N_9525,N_8365);
nor U10153 (N_10153,N_9977,N_8726);
xnor U10154 (N_10154,N_9575,N_8811);
xor U10155 (N_10155,N_9032,N_8223);
and U10156 (N_10156,N_8376,N_9121);
nor U10157 (N_10157,N_8950,N_9461);
nand U10158 (N_10158,N_8790,N_8904);
and U10159 (N_10159,N_8516,N_8856);
nand U10160 (N_10160,N_9379,N_9631);
or U10161 (N_10161,N_8518,N_9654);
xnor U10162 (N_10162,N_8259,N_8089);
or U10163 (N_10163,N_8485,N_9899);
and U10164 (N_10164,N_8486,N_9158);
xor U10165 (N_10165,N_8489,N_9481);
nand U10166 (N_10166,N_8406,N_8827);
or U10167 (N_10167,N_9905,N_9188);
and U10168 (N_10168,N_9116,N_8754);
nor U10169 (N_10169,N_9109,N_9446);
or U10170 (N_10170,N_8814,N_9983);
xnor U10171 (N_10171,N_8990,N_8520);
nand U10172 (N_10172,N_8780,N_8991);
and U10173 (N_10173,N_8429,N_9688);
nand U10174 (N_10174,N_8700,N_8834);
nor U10175 (N_10175,N_9348,N_9624);
and U10176 (N_10176,N_8866,N_9887);
and U10177 (N_10177,N_9679,N_9015);
nor U10178 (N_10178,N_8051,N_9339);
nand U10179 (N_10179,N_8566,N_8102);
nor U10180 (N_10180,N_8960,N_8114);
nor U10181 (N_10181,N_8728,N_8447);
and U10182 (N_10182,N_9502,N_8242);
nor U10183 (N_10183,N_8500,N_8166);
xnor U10184 (N_10184,N_9708,N_9290);
xor U10185 (N_10185,N_8674,N_9365);
or U10186 (N_10186,N_9340,N_8972);
xnor U10187 (N_10187,N_8262,N_8996);
xor U10188 (N_10188,N_8578,N_9813);
or U10189 (N_10189,N_9193,N_9652);
and U10190 (N_10190,N_8608,N_8235);
and U10191 (N_10191,N_9218,N_9934);
xnor U10192 (N_10192,N_9310,N_9273);
and U10193 (N_10193,N_9459,N_8776);
nand U10194 (N_10194,N_9465,N_9980);
xnor U10195 (N_10195,N_8180,N_8956);
or U10196 (N_10196,N_8993,N_9871);
nand U10197 (N_10197,N_8058,N_9241);
and U10198 (N_10198,N_9143,N_8718);
and U10199 (N_10199,N_9455,N_8068);
xor U10200 (N_10200,N_9449,N_9711);
xor U10201 (N_10201,N_8188,N_8677);
nor U10202 (N_10202,N_9198,N_9493);
nor U10203 (N_10203,N_8079,N_8633);
and U10204 (N_10204,N_9412,N_8716);
xnor U10205 (N_10205,N_9422,N_9333);
nand U10206 (N_10206,N_8959,N_8570);
xnor U10207 (N_10207,N_9358,N_8631);
or U10208 (N_10208,N_8139,N_8059);
xor U10209 (N_10209,N_9914,N_8257);
and U10210 (N_10210,N_9160,N_9945);
nand U10211 (N_10211,N_9731,N_9236);
nor U10212 (N_10212,N_8735,N_8090);
and U10213 (N_10213,N_8437,N_8268);
nor U10214 (N_10214,N_9562,N_9842);
xor U10215 (N_10215,N_8724,N_9312);
nand U10216 (N_10216,N_9395,N_9949);
nor U10217 (N_10217,N_9008,N_8336);
and U10218 (N_10218,N_8995,N_8287);
and U10219 (N_10219,N_9181,N_8258);
xor U10220 (N_10220,N_9783,N_9353);
or U10221 (N_10221,N_9665,N_8273);
xnor U10222 (N_10222,N_9487,N_8053);
nand U10223 (N_10223,N_8920,N_8260);
xnor U10224 (N_10224,N_8657,N_9132);
nand U10225 (N_10225,N_9741,N_8939);
and U10226 (N_10226,N_8575,N_8679);
xor U10227 (N_10227,N_8313,N_8238);
nand U10228 (N_10228,N_9873,N_9836);
xor U10229 (N_10229,N_8117,N_8098);
and U10230 (N_10230,N_9712,N_9751);
nor U10231 (N_10231,N_8732,N_8423);
nor U10232 (N_10232,N_8561,N_8601);
and U10233 (N_10233,N_9306,N_9718);
nor U10234 (N_10234,N_9451,N_8322);
nand U10235 (N_10235,N_8453,N_8052);
or U10236 (N_10236,N_8379,N_9594);
nand U10237 (N_10237,N_9080,N_9421);
nand U10238 (N_10238,N_9866,N_9265);
or U10239 (N_10239,N_9752,N_9898);
and U10240 (N_10240,N_9284,N_9355);
and U10241 (N_10241,N_8451,N_9666);
or U10242 (N_10242,N_9592,N_8552);
or U10243 (N_10243,N_8353,N_9662);
and U10244 (N_10244,N_8643,N_8747);
or U10245 (N_10245,N_8352,N_9915);
or U10246 (N_10246,N_8994,N_8399);
nand U10247 (N_10247,N_9260,N_8841);
nand U10248 (N_10248,N_9419,N_9523);
xnor U10249 (N_10249,N_8638,N_9786);
or U10250 (N_10250,N_9588,N_9503);
or U10251 (N_10251,N_9689,N_9296);
or U10252 (N_10252,N_9684,N_8855);
and U10253 (N_10253,N_9482,N_9354);
or U10254 (N_10254,N_9617,N_8743);
and U10255 (N_10255,N_9372,N_9563);
xor U10256 (N_10256,N_9926,N_9700);
or U10257 (N_10257,N_8762,N_8339);
and U10258 (N_10258,N_8100,N_9200);
xnor U10259 (N_10259,N_8343,N_8985);
nand U10260 (N_10260,N_9954,N_8192);
or U10261 (N_10261,N_8951,N_9878);
nand U10262 (N_10262,N_8301,N_9096);
and U10263 (N_10263,N_9201,N_9364);
nor U10264 (N_10264,N_8508,N_9719);
xor U10265 (N_10265,N_9995,N_9599);
nor U10266 (N_10266,N_9287,N_8420);
nor U10267 (N_10267,N_9389,N_8310);
or U10268 (N_10268,N_8396,N_9163);
and U10269 (N_10269,N_9066,N_8668);
nor U10270 (N_10270,N_9432,N_9990);
nor U10271 (N_10271,N_8163,N_9177);
xor U10272 (N_10272,N_9840,N_9018);
and U10273 (N_10273,N_9917,N_8525);
or U10274 (N_10274,N_9235,N_8263);
or U10275 (N_10275,N_9515,N_8306);
xnor U10276 (N_10276,N_9972,N_8133);
nor U10277 (N_10277,N_8557,N_8347);
and U10278 (N_10278,N_9441,N_9998);
xnor U10279 (N_10279,N_8593,N_8586);
nor U10280 (N_10280,N_9692,N_9377);
xor U10281 (N_10281,N_9979,N_9924);
xnor U10282 (N_10282,N_8300,N_9361);
nand U10283 (N_10283,N_9855,N_9180);
nor U10284 (N_10284,N_9237,N_9854);
and U10285 (N_10285,N_8430,N_8768);
or U10286 (N_10286,N_9103,N_8579);
nor U10287 (N_10287,N_8534,N_8597);
xnor U10288 (N_10288,N_8916,N_9518);
nor U10289 (N_10289,N_9047,N_8124);
and U10290 (N_10290,N_8978,N_8908);
xor U10291 (N_10291,N_9102,N_9552);
xnor U10292 (N_10292,N_8443,N_8545);
xnor U10293 (N_10293,N_9556,N_8295);
nand U10294 (N_10294,N_9376,N_8707);
nor U10295 (N_10295,N_9778,N_9477);
nor U10296 (N_10296,N_8528,N_9929);
nor U10297 (N_10297,N_8853,N_9618);
xor U10298 (N_10298,N_8237,N_8463);
xor U10299 (N_10299,N_9174,N_8078);
xor U10300 (N_10300,N_8829,N_8183);
nor U10301 (N_10301,N_9988,N_8219);
nor U10302 (N_10302,N_8532,N_8725);
nor U10303 (N_10303,N_8197,N_9936);
nor U10304 (N_10304,N_9764,N_9020);
nor U10305 (N_10305,N_8802,N_9438);
nand U10306 (N_10306,N_9039,N_8729);
nand U10307 (N_10307,N_8194,N_9420);
or U10308 (N_10308,N_9777,N_9454);
or U10309 (N_10309,N_8248,N_8146);
xnor U10310 (N_10310,N_8371,N_9027);
nor U10311 (N_10311,N_9076,N_8757);
and U10312 (N_10312,N_8846,N_9922);
nor U10313 (N_10313,N_8070,N_8758);
or U10314 (N_10314,N_9068,N_8825);
xnor U10315 (N_10315,N_9167,N_8943);
and U10316 (N_10316,N_9614,N_8097);
xor U10317 (N_10317,N_8870,N_8445);
or U10318 (N_10318,N_8652,N_8635);
nand U10319 (N_10319,N_8873,N_9051);
or U10320 (N_10320,N_8121,N_8592);
and U10321 (N_10321,N_9702,N_9742);
nand U10322 (N_10322,N_8558,N_8499);
nor U10323 (N_10323,N_9403,N_8517);
nor U10324 (N_10324,N_9033,N_8621);
nand U10325 (N_10325,N_8107,N_8961);
nand U10326 (N_10326,N_8005,N_9307);
xnor U10327 (N_10327,N_9001,N_8792);
nand U10328 (N_10328,N_8676,N_8424);
and U10329 (N_10329,N_9733,N_8291);
xnor U10330 (N_10330,N_9050,N_9124);
nand U10331 (N_10331,N_9821,N_8976);
or U10332 (N_10332,N_8822,N_9574);
or U10333 (N_10333,N_9590,N_9545);
or U10334 (N_10334,N_9485,N_9634);
xor U10335 (N_10335,N_8838,N_8656);
xor U10336 (N_10336,N_9378,N_9128);
or U10337 (N_10337,N_9399,N_8582);
nand U10338 (N_10338,N_9360,N_9576);
or U10339 (N_10339,N_8319,N_8108);
nor U10340 (N_10340,N_9321,N_8942);
xor U10341 (N_10341,N_8986,N_9879);
or U10342 (N_10342,N_9295,N_8144);
and U10343 (N_10343,N_9701,N_8141);
xnor U10344 (N_10344,N_8465,N_9831);
and U10345 (N_10345,N_9568,N_9002);
or U10346 (N_10346,N_8882,N_8602);
nand U10347 (N_10347,N_8106,N_8245);
nand U10348 (N_10348,N_8979,N_8523);
nor U10349 (N_10349,N_9463,N_9205);
nor U10350 (N_10350,N_9645,N_8413);
or U10351 (N_10351,N_9334,N_8207);
nand U10352 (N_10352,N_8265,N_9627);
xor U10353 (N_10353,N_8548,N_8905);
nor U10354 (N_10354,N_9309,N_9526);
xor U10355 (N_10355,N_8171,N_8087);
xnor U10356 (N_10356,N_8039,N_8022);
xnor U10357 (N_10357,N_9041,N_8229);
nor U10358 (N_10358,N_8177,N_9514);
and U10359 (N_10359,N_8026,N_8346);
and U10360 (N_10360,N_8766,N_8236);
nand U10361 (N_10361,N_9301,N_9190);
nor U10362 (N_10362,N_8760,N_9621);
and U10363 (N_10363,N_9596,N_8709);
or U10364 (N_10364,N_8755,N_9567);
nor U10365 (N_10365,N_9387,N_8786);
and U10366 (N_10366,N_9233,N_8230);
and U10367 (N_10367,N_9759,N_8581);
and U10368 (N_10368,N_9100,N_9279);
and U10369 (N_10369,N_8890,N_9531);
nor U10370 (N_10370,N_8023,N_9165);
and U10371 (N_10371,N_8042,N_8658);
nor U10372 (N_10372,N_8712,N_8045);
nor U10373 (N_10373,N_8462,N_8613);
nor U10374 (N_10374,N_8519,N_8439);
or U10375 (N_10375,N_9678,N_9919);
and U10376 (N_10376,N_9856,N_9636);
and U10377 (N_10377,N_9823,N_9952);
and U10378 (N_10378,N_8573,N_9229);
and U10379 (N_10379,N_9841,N_9770);
and U10380 (N_10380,N_9400,N_9587);
nand U10381 (N_10381,N_9371,N_8111);
xnor U10382 (N_10382,N_8971,N_9810);
or U10383 (N_10383,N_9386,N_9024);
xor U10384 (N_10384,N_9071,N_9196);
or U10385 (N_10385,N_8599,N_8785);
nand U10386 (N_10386,N_9509,N_8158);
nor U10387 (N_10387,N_9543,N_9450);
xor U10388 (N_10388,N_9090,N_9935);
nand U10389 (N_10389,N_8992,N_8127);
nor U10390 (N_10390,N_8267,N_9444);
nand U10391 (N_10391,N_9573,N_8472);
nor U10392 (N_10392,N_8427,N_9863);
xor U10393 (N_10393,N_8105,N_8749);
nand U10394 (N_10394,N_8232,N_9226);
nand U10395 (N_10395,N_9056,N_8033);
xnor U10396 (N_10396,N_9794,N_8113);
or U10397 (N_10397,N_8974,N_8615);
xnor U10398 (N_10398,N_9591,N_9862);
and U10399 (N_10399,N_8112,N_9837);
nand U10400 (N_10400,N_8043,N_8293);
nor U10401 (N_10401,N_8845,N_9610);
or U10402 (N_10402,N_8182,N_9437);
and U10403 (N_10403,N_9559,N_8024);
xnor U10404 (N_10404,N_9532,N_8307);
or U10405 (N_10405,N_9723,N_8748);
nand U10406 (N_10406,N_8684,N_9331);
nand U10407 (N_10407,N_8682,N_9675);
and U10408 (N_10408,N_9097,N_8641);
nor U10409 (N_10409,N_9884,N_8636);
nand U10410 (N_10410,N_9114,N_9130);
or U10411 (N_10411,N_9787,N_9806);
and U10412 (N_10412,N_8199,N_8903);
xor U10413 (N_10413,N_9941,N_9845);
nor U10414 (N_10414,N_9433,N_8378);
and U10415 (N_10415,N_8988,N_8442);
nand U10416 (N_10416,N_9336,N_8254);
nor U10417 (N_10417,N_8308,N_9713);
xnor U10418 (N_10418,N_8001,N_9829);
and U10419 (N_10419,N_8285,N_9390);
nor U10420 (N_10420,N_9874,N_9882);
and U10421 (N_10421,N_8314,N_9994);
nor U10422 (N_10422,N_9724,N_9299);
or U10423 (N_10423,N_9635,N_9478);
xnor U10424 (N_10424,N_9607,N_8450);
and U10425 (N_10425,N_9542,N_9800);
nor U10426 (N_10426,N_8934,N_9643);
nor U10427 (N_10427,N_9824,N_8727);
or U10428 (N_10428,N_9495,N_9655);
xor U10429 (N_10429,N_9892,N_9886);
xor U10430 (N_10430,N_9802,N_9440);
nor U10431 (N_10431,N_9939,N_8590);
xor U10432 (N_10432,N_9323,N_8891);
xor U10433 (N_10433,N_9900,N_9697);
and U10434 (N_10434,N_9093,N_9079);
or U10435 (N_10435,N_9099,N_9145);
nor U10436 (N_10436,N_9135,N_9245);
xnor U10437 (N_10437,N_9036,N_8935);
nor U10438 (N_10438,N_8867,N_8798);
xor U10439 (N_10439,N_8069,N_9782);
nand U10440 (N_10440,N_9021,N_9254);
or U10441 (N_10441,N_8553,N_8461);
or U10442 (N_10442,N_9560,N_8711);
nor U10443 (N_10443,N_9325,N_9221);
nor U10444 (N_10444,N_9302,N_8806);
or U10445 (N_10445,N_9828,N_8409);
and U10446 (N_10446,N_8289,N_8666);
xnor U10447 (N_10447,N_8812,N_9058);
xnor U10448 (N_10448,N_8769,N_8928);
or U10449 (N_10449,N_8136,N_9094);
or U10450 (N_10450,N_9680,N_9156);
nor U10451 (N_10451,N_8401,N_9435);
xnor U10452 (N_10452,N_8218,N_9819);
xnor U10453 (N_10453,N_9714,N_8865);
or U10454 (N_10454,N_8007,N_8901);
nor U10455 (N_10455,N_8713,N_8179);
nor U10456 (N_10456,N_9796,N_8877);
and U10457 (N_10457,N_8266,N_9848);
nor U10458 (N_10458,N_9937,N_8817);
nor U10459 (N_10459,N_9570,N_9330);
or U10460 (N_10460,N_8984,N_9566);
or U10461 (N_10461,N_9374,N_9207);
and U10462 (N_10462,N_8277,N_8370);
and U10463 (N_10463,N_8533,N_8655);
xnor U10464 (N_10464,N_9798,N_9763);
and U10465 (N_10465,N_8176,N_8400);
and U10466 (N_10466,N_9661,N_8646);
nor U10467 (N_10467,N_9641,N_9262);
nor U10468 (N_10468,N_8535,N_9571);
and U10469 (N_10469,N_9572,N_8055);
nor U10470 (N_10470,N_9637,N_9029);
or U10471 (N_10471,N_9375,N_8004);
nand U10472 (N_10472,N_8387,N_8467);
xnor U10473 (N_10473,N_9647,N_9547);
nor U10474 (N_10474,N_9231,N_8200);
and U10475 (N_10475,N_9872,N_8731);
and U10476 (N_10476,N_8793,N_8264);
nand U10477 (N_10477,N_8428,N_8603);
xor U10478 (N_10478,N_9407,N_9272);
nor U10479 (N_10479,N_9603,N_9005);
nor U10480 (N_10480,N_8464,N_8772);
nor U10481 (N_10481,N_8576,N_9185);
nand U10482 (N_10482,N_8216,N_8274);
or U10483 (N_10483,N_8473,N_8459);
nor U10484 (N_10484,N_8252,N_8233);
nand U10485 (N_10485,N_8940,N_9586);
and U10486 (N_10486,N_9757,N_9125);
and U10487 (N_10487,N_8692,N_9928);
nand U10488 (N_10488,N_9028,N_9293);
nor U10489 (N_10489,N_8074,N_9266);
and U10490 (N_10490,N_8949,N_9335);
nor U10491 (N_10491,N_9960,N_8495);
nor U10492 (N_10492,N_8704,N_8872);
and U10493 (N_10493,N_8746,N_9826);
nand U10494 (N_10494,N_8067,N_9142);
xnor U10495 (N_10495,N_8538,N_8560);
and U10496 (N_10496,N_9944,N_9057);
or U10497 (N_10497,N_9259,N_8703);
nor U10498 (N_10498,N_9535,N_9516);
xnor U10499 (N_10499,N_9238,N_8624);
and U10500 (N_10500,N_8955,N_9626);
or U10501 (N_10501,N_8368,N_9901);
or U10502 (N_10502,N_8839,N_9447);
nand U10503 (N_10503,N_9916,N_8092);
nand U10504 (N_10504,N_9554,N_8046);
nand U10505 (N_10505,N_8390,N_9955);
or U10506 (N_10506,N_8490,N_9043);
and U10507 (N_10507,N_9506,N_8367);
nand U10508 (N_10508,N_8419,N_8836);
and U10509 (N_10509,N_8738,N_9890);
xnor U10510 (N_10510,N_8311,N_8383);
nand U10511 (N_10511,N_9583,N_9127);
nand U10512 (N_10512,N_8228,N_8691);
or U10513 (N_10513,N_8941,N_9638);
nand U10514 (N_10514,N_9203,N_8497);
and U10515 (N_10515,N_8809,N_9352);
nand U10516 (N_10516,N_8374,N_8403);
xnor U10517 (N_10517,N_9989,N_8165);
xnor U10518 (N_10518,N_9342,N_8338);
nand U10519 (N_10519,N_8511,N_8708);
nand U10520 (N_10520,N_8222,N_9261);
xnor U10521 (N_10521,N_8962,N_9169);
nand U10522 (N_10522,N_9738,N_8025);
xor U10523 (N_10523,N_9206,N_9443);
nand U10524 (N_10524,N_8261,N_9170);
or U10525 (N_10525,N_9971,N_8759);
nor U10526 (N_10526,N_8686,N_9223);
nor U10527 (N_10527,N_9319,N_9773);
xnor U10528 (N_10528,N_9978,N_9857);
nand U10529 (N_10529,N_9529,N_9081);
and U10530 (N_10530,N_9468,N_9849);
or U10531 (N_10531,N_8175,N_8320);
and U10532 (N_10532,N_8480,N_9750);
nor U10533 (N_10533,N_8372,N_9834);
xnor U10534 (N_10534,N_9699,N_8355);
nor U10535 (N_10535,N_9197,N_9492);
xor U10536 (N_10536,N_8600,N_9278);
nand U10537 (N_10537,N_9600,N_8487);
nor U10538 (N_10538,N_8921,N_9242);
and U10539 (N_10539,N_9667,N_8781);
or U10540 (N_10540,N_9869,N_8118);
nand U10541 (N_10541,N_8504,N_8906);
nor U10542 (N_10542,N_9760,N_8642);
nand U10543 (N_10543,N_9149,N_9725);
nand U10544 (N_10544,N_9357,N_8000);
and U10545 (N_10545,N_9888,N_9324);
xor U10546 (N_10546,N_9172,N_9258);
xor U10547 (N_10547,N_9805,N_9280);
xor U10548 (N_10548,N_9537,N_8598);
xnor U10549 (N_10549,N_9344,N_9153);
nand U10550 (N_10550,N_9137,N_8130);
xnor U10551 (N_10551,N_9428,N_8914);
nor U10552 (N_10552,N_8681,N_9414);
nor U10553 (N_10553,N_8337,N_8823);
nand U10554 (N_10554,N_8694,N_9062);
nor U10555 (N_10555,N_9859,N_9186);
or U10556 (N_10556,N_8394,N_9098);
and U10557 (N_10557,N_8398,N_9019);
or U10558 (N_10558,N_8632,N_9467);
or U10559 (N_10559,N_8330,N_8012);
nand U10560 (N_10560,N_8076,N_9148);
nand U10561 (N_10561,N_9781,N_9488);
nor U10562 (N_10562,N_9313,N_9224);
xnor U10563 (N_10563,N_9676,N_9483);
xnor U10564 (N_10564,N_8881,N_9595);
xnor U10565 (N_10565,N_9981,N_8416);
nand U10566 (N_10566,N_8618,N_9925);
or U10567 (N_10567,N_8147,N_9252);
or U10568 (N_10568,N_9356,N_8815);
or U10569 (N_10569,N_9923,N_8084);
nor U10570 (N_10570,N_8973,N_8821);
or U10571 (N_10571,N_8326,N_8619);
nand U10572 (N_10572,N_9716,N_8966);
nor U10573 (N_10573,N_8455,N_9286);
or U10574 (N_10574,N_8889,N_8281);
xor U10575 (N_10575,N_9327,N_9609);
xor U10576 (N_10576,N_8869,N_9052);
or U10577 (N_10577,N_9095,N_9007);
and U10578 (N_10578,N_9740,N_9146);
and U10579 (N_10579,N_9993,N_9219);
or U10580 (N_10580,N_8543,N_8348);
or U10581 (N_10581,N_9948,N_9720);
or U10582 (N_10582,N_9507,N_9215);
nor U10583 (N_10583,N_8185,N_9694);
or U10584 (N_10584,N_8110,N_8871);
nand U10585 (N_10585,N_9393,N_8137);
nor U10586 (N_10586,N_9927,N_8134);
and U10587 (N_10587,N_8270,N_8696);
xor U10588 (N_10588,N_9876,N_8407);
xnor U10589 (N_10589,N_8697,N_9409);
or U10590 (N_10590,N_8588,N_9602);
nand U10591 (N_10591,N_8737,N_8109);
xnor U10592 (N_10592,N_9088,N_9394);
or U10593 (N_10593,N_9612,N_9120);
xor U10594 (N_10594,N_9154,N_8064);
nand U10595 (N_10595,N_8710,N_8685);
or U10596 (N_10596,N_9546,N_9877);
xor U10597 (N_10597,N_8614,N_9418);
nand U10598 (N_10598,N_9668,N_8661);
or U10599 (N_10599,N_9651,N_8626);
xor U10600 (N_10600,N_9411,N_9000);
xor U10601 (N_10601,N_8008,N_8526);
or U10602 (N_10602,N_8750,N_8449);
nor U10603 (N_10603,N_9087,N_9943);
and U10604 (N_10604,N_8506,N_8221);
or U10605 (N_10605,N_8309,N_8126);
and U10606 (N_10606,N_9268,N_8123);
nor U10607 (N_10607,N_9639,N_8693);
nand U10608 (N_10608,N_8739,N_9122);
and U10609 (N_10609,N_8611,N_9054);
nor U10610 (N_10610,N_9060,N_8019);
nor U10611 (N_10611,N_9107,N_9788);
or U10612 (N_10612,N_8835,N_8591);
or U10613 (N_10613,N_9155,N_9687);
or U10614 (N_10614,N_8341,N_8617);
or U10615 (N_10615,N_8181,N_8559);
nand U10616 (N_10616,N_8475,N_8840);
nand U10617 (N_10617,N_8876,N_8278);
nor U10618 (N_10618,N_8280,N_9034);
xor U10619 (N_10619,N_9536,N_9366);
nor U10620 (N_10620,N_8190,N_9698);
or U10621 (N_10621,N_8284,N_8138);
xnor U10622 (N_10622,N_8498,N_9745);
xnor U10623 (N_10623,N_9410,N_9179);
or U10624 (N_10624,N_9351,N_9722);
or U10625 (N_10625,N_9851,N_8115);
and U10626 (N_10626,N_8565,N_9368);
or U10627 (N_10627,N_8551,N_9382);
nand U10628 (N_10628,N_8148,N_9508);
nand U10629 (N_10629,N_8777,N_9540);
xnor U10630 (N_10630,N_9895,N_9346);
or U10631 (N_10631,N_8272,N_8819);
nand U10632 (N_10632,N_9288,N_9303);
and U10633 (N_10633,N_9765,N_9649);
and U10634 (N_10634,N_8721,N_8412);
nor U10635 (N_10635,N_8239,N_8077);
nand U10636 (N_10636,N_8244,N_9214);
and U10637 (N_10637,N_8664,N_9625);
xor U10638 (N_10638,N_9151,N_8153);
xor U10639 (N_10639,N_8009,N_8391);
nor U10640 (N_10640,N_9267,N_9695);
xnor U10641 (N_10641,N_9657,N_8805);
xor U10642 (N_10642,N_8833,N_8255);
or U10643 (N_10643,N_9402,N_8897);
or U10644 (N_10644,N_9274,N_8094);
xor U10645 (N_10645,N_9022,N_9721);
xor U10646 (N_10646,N_9117,N_8787);
and U10647 (N_10647,N_9767,N_8587);
or U10648 (N_10648,N_9953,N_8609);
nand U10649 (N_10649,N_9656,N_9091);
and U10650 (N_10650,N_9013,N_9234);
nor U10651 (N_10651,N_9946,N_8140);
or U10652 (N_10652,N_9464,N_9811);
nor U10653 (N_10653,N_8859,N_8715);
nor U10654 (N_10654,N_8329,N_8964);
nor U10655 (N_10655,N_8104,N_9795);
nor U10656 (N_10656,N_8521,N_9496);
nand U10657 (N_10657,N_8395,N_9808);
and U10658 (N_10658,N_9727,N_9119);
and U10659 (N_10659,N_9257,N_8673);
and U10660 (N_10660,N_8947,N_8422);
nand U10661 (N_10661,N_8324,N_9838);
and U10662 (N_10662,N_8471,N_8874);
or U10663 (N_10663,N_8730,N_8946);
or U10664 (N_10664,N_8536,N_8202);
or U10665 (N_10665,N_8807,N_8095);
nand U10666 (N_10666,N_9726,N_9785);
nand U10667 (N_10667,N_8733,N_8027);
and U10668 (N_10668,N_8784,N_9380);
xor U10669 (N_10669,N_8753,N_8193);
or U10670 (N_10670,N_9059,N_9703);
nor U10671 (N_10671,N_9896,N_9517);
nand U10672 (N_10672,N_9084,N_8028);
and U10673 (N_10673,N_8159,N_8279);
xor U10674 (N_10674,N_8810,N_8589);
and U10675 (N_10675,N_8907,N_8298);
and U10676 (N_10676,N_9166,N_8269);
or U10677 (N_10677,N_9633,N_9958);
nand U10678 (N_10678,N_9902,N_9505);
xnor U10679 (N_10679,N_8010,N_8253);
and U10680 (N_10680,N_9964,N_9404);
nor U10681 (N_10681,N_9305,N_8794);
and U10682 (N_10682,N_8678,N_8860);
nor U10683 (N_10683,N_8926,N_9530);
or U10684 (N_10684,N_8675,N_9453);
or U10685 (N_10685,N_9430,N_8358);
xor U10686 (N_10686,N_9864,N_9392);
nor U10687 (N_10687,N_8361,N_9458);
nand U10688 (N_10688,N_8066,N_9077);
and U10689 (N_10689,N_8204,N_9969);
nand U10690 (N_10690,N_9950,N_8509);
or U10691 (N_10691,N_9736,N_8103);
xnor U10692 (N_10692,N_8408,N_8550);
nand U10693 (N_10693,N_9670,N_9511);
nand U10694 (N_10694,N_9320,N_8572);
nor U10695 (N_10695,N_8212,N_8530);
or U10696 (N_10696,N_9775,N_8801);
or U10697 (N_10697,N_9771,N_9512);
nor U10698 (N_10698,N_9105,N_8388);
or U10699 (N_10699,N_9799,N_9192);
nand U10700 (N_10700,N_9558,N_8502);
nand U10701 (N_10701,N_9615,N_8282);
or U10702 (N_10702,N_9078,N_9484);
nand U10703 (N_10703,N_9728,N_8861);
and U10704 (N_10704,N_8667,N_9396);
nor U10705 (N_10705,N_9070,N_8909);
xnor U10706 (N_10706,N_9613,N_8512);
xor U10707 (N_10707,N_8898,N_9825);
or U10708 (N_10708,N_8057,N_8880);
or U10709 (N_10709,N_8637,N_8529);
and U10710 (N_10710,N_8441,N_9814);
or U10711 (N_10711,N_8612,N_9025);
nor U10712 (N_10712,N_8918,N_9551);
nand U10713 (N_10713,N_8982,N_8377);
nor U10714 (N_10714,N_8389,N_9967);
and U10715 (N_10715,N_9987,N_8363);
or U10716 (N_10716,N_8824,N_9479);
and U10717 (N_10717,N_9271,N_8318);
or U10718 (N_10718,N_8044,N_9682);
or U10719 (N_10719,N_9832,N_9623);
nor U10720 (N_10720,N_8470,N_8384);
nand U10721 (N_10721,N_8580,N_9489);
nand U10722 (N_10722,N_8071,N_8359);
and U10723 (N_10723,N_9779,N_8350);
nand U10724 (N_10724,N_8060,N_8958);
xor U10725 (N_10725,N_9754,N_8912);
or U10726 (N_10726,N_8340,N_8540);
nor U10727 (N_10727,N_9920,N_9747);
nor U10728 (N_10728,N_9417,N_9141);
or U10729 (N_10729,N_9349,N_8695);
and U10730 (N_10730,N_8751,N_8211);
nand U10731 (N_10731,N_9275,N_9159);
nor U10732 (N_10732,N_8457,N_8050);
nor U10733 (N_10733,N_8297,N_8847);
nand U10734 (N_10734,N_8198,N_8771);
or U10735 (N_10735,N_9959,N_8654);
xor U10736 (N_10736,N_8705,N_9436);
nor U10737 (N_10737,N_8294,N_9861);
xor U10738 (N_10738,N_9585,N_8209);
and U10739 (N_10739,N_8848,N_8980);
nor U10740 (N_10740,N_9168,N_8392);
nand U10741 (N_10741,N_8325,N_9500);
nor U10742 (N_10742,N_8017,N_8315);
and U10743 (N_10743,N_9239,N_9520);
xor U10744 (N_10744,N_8765,N_8483);
nand U10745 (N_10745,N_8843,N_9737);
nand U10746 (N_10746,N_9883,N_9717);
nand U10747 (N_10747,N_8513,N_9843);
and U10748 (N_10748,N_9129,N_8796);
xnor U10749 (N_10749,N_9730,N_8952);
nand U10750 (N_10750,N_9734,N_9308);
nand U10751 (N_10751,N_9044,N_8965);
nand U10752 (N_10752,N_9669,N_9973);
xnor U10753 (N_10753,N_9147,N_8014);
and U10754 (N_10754,N_8036,N_8648);
and U10755 (N_10755,N_9581,N_8788);
xor U10756 (N_10756,N_8345,N_9227);
xnor U10757 (N_10757,N_9780,N_8567);
nand U10758 (N_10758,N_9904,N_9729);
xnor U10759 (N_10759,N_8932,N_9792);
or U10760 (N_10760,N_8863,N_8689);
xnor U10761 (N_10761,N_9003,N_8150);
or U10762 (N_10762,N_8857,N_9210);
nor U10763 (N_10763,N_9672,N_9253);
and U10764 (N_10764,N_8634,N_9991);
nand U10765 (N_10765,N_8563,N_9030);
or U10766 (N_10766,N_9442,N_9202);
xnor U10767 (N_10767,N_9822,N_9220);
xnor U10768 (N_10768,N_8482,N_9183);
and U10769 (N_10769,N_8047,N_8623);
or U10770 (N_10770,N_9582,N_8547);
xnor U10771 (N_10771,N_8936,N_8415);
nand U10772 (N_10772,N_9817,N_8037);
or U10773 (N_10773,N_9868,N_9332);
nand U10774 (N_10774,N_9228,N_9557);
nor U10775 (N_10775,N_8650,N_9776);
xnor U10776 (N_10776,N_9565,N_8680);
and U10777 (N_10777,N_8196,N_9906);
and U10778 (N_10778,N_8944,N_9601);
and U10779 (N_10779,N_8989,N_9739);
and U10780 (N_10780,N_9191,N_9897);
or U10781 (N_10781,N_9791,N_9962);
nand U10782 (N_10782,N_9974,N_9126);
nand U10783 (N_10783,N_9012,N_9006);
nand U10784 (N_10784,N_8286,N_9630);
and U10785 (N_10785,N_9686,N_9908);
and U10786 (N_10786,N_9918,N_8034);
nor U10787 (N_10787,N_9839,N_9175);
or U10788 (N_10788,N_9462,N_8911);
nand U10789 (N_10789,N_9732,N_9425);
or U10790 (N_10790,N_8864,N_8653);
and U10791 (N_10791,N_8421,N_8688);
nor U10792 (N_10792,N_9683,N_8610);
nor U10793 (N_10793,N_8003,N_8142);
nor U10794 (N_10794,N_8446,N_9115);
and U10795 (N_10795,N_8305,N_9804);
nand U10796 (N_10796,N_9405,N_8999);
or U10797 (N_10797,N_8967,N_8723);
or U10798 (N_10798,N_8021,N_9758);
nand U10799 (N_10799,N_8015,N_9111);
nand U10800 (N_10800,N_8717,N_9538);
nor U10801 (N_10801,N_9891,N_9046);
or U10802 (N_10802,N_8458,N_8444);
nor U10803 (N_10803,N_8767,N_8167);
or U10804 (N_10804,N_8672,N_8945);
and U10805 (N_10805,N_9011,N_8522);
xnor U10806 (N_10806,N_9474,N_9456);
nor U10807 (N_10807,N_9317,N_9251);
xor U10808 (N_10808,N_8832,N_8128);
nand U10809 (N_10809,N_8930,N_9844);
xor U10810 (N_10810,N_9277,N_8162);
nand U10811 (N_10811,N_8892,N_9388);
xnor U10812 (N_10812,N_8549,N_8505);
xor U10813 (N_10813,N_8397,N_8702);
and U10814 (N_10814,N_9793,N_8849);
xnor U10815 (N_10815,N_9589,N_8981);
or U10816 (N_10816,N_9063,N_9045);
xnor U10817 (N_10817,N_8191,N_9256);
and U10818 (N_10818,N_8492,N_8032);
xnor U10819 (N_10819,N_8605,N_8606);
nor U10820 (N_10820,N_9315,N_9992);
nand U10821 (N_10821,N_8744,N_8256);
nor U10822 (N_10822,N_9373,N_8628);
nand U10823 (N_10823,N_9472,N_9999);
xnor U10824 (N_10824,N_8393,N_8373);
and U10825 (N_10825,N_9023,N_8225);
xnor U10826 (N_10826,N_8083,N_9833);
or U10827 (N_10827,N_9016,N_8640);
and U10828 (N_10828,N_8155,N_8431);
nand U10829 (N_10829,N_9112,N_9784);
nor U10830 (N_10830,N_8425,N_8170);
and U10831 (N_10831,N_8720,N_9494);
nor U10832 (N_10832,N_8041,N_8556);
nand U10833 (N_10833,N_9772,N_9297);
nor U10834 (N_10834,N_9846,N_9457);
xnor U10835 (N_10835,N_8970,N_8101);
nor U10836 (N_10836,N_8627,N_8670);
and U10837 (N_10837,N_9162,N_9510);
or U10838 (N_10838,N_9789,N_8290);
and U10839 (N_10839,N_9429,N_9263);
xor U10840 (N_10840,N_9646,N_8527);
and U10841 (N_10841,N_9524,N_9152);
or U10842 (N_10842,N_8271,N_8584);
and U10843 (N_10843,N_8763,N_9704);
and U10844 (N_10844,N_9101,N_9616);
and U10845 (N_10845,N_8493,N_9473);
nand U10846 (N_10846,N_8585,N_8629);
xnor U10847 (N_10847,N_9212,N_9749);
nand U10848 (N_10848,N_8616,N_8510);
xor U10849 (N_10849,N_8683,N_9269);
nor U10850 (N_10850,N_9194,N_8501);
nand U10851 (N_10851,N_9476,N_9161);
or U10852 (N_10852,N_8438,N_8888);
nand U10853 (N_10853,N_9548,N_9381);
and U10854 (N_10854,N_8356,N_8722);
or U10855 (N_10855,N_9504,N_8862);
and U10856 (N_10856,N_9818,N_9074);
or U10857 (N_10857,N_8844,N_9881);
or U10858 (N_10858,N_8213,N_9434);
or U10859 (N_10859,N_9620,N_9815);
xnor U10860 (N_10860,N_9762,N_9031);
nand U10861 (N_10861,N_9951,N_8478);
nor U10862 (N_10862,N_9801,N_8687);
and U10863 (N_10863,N_8231,N_9968);
and U10864 (N_10864,N_9768,N_8201);
or U10865 (N_10865,N_8035,N_8460);
nand U10866 (N_10866,N_8187,N_8006);
nand U10867 (N_10867,N_8804,N_9976);
nor U10868 (N_10868,N_8380,N_8488);
nand U10869 (N_10869,N_8569,N_9663);
and U10870 (N_10870,N_8998,N_8595);
nand U10871 (N_10871,N_9674,N_9564);
xor U10872 (N_10872,N_8351,N_9359);
xor U10873 (N_10873,N_9673,N_9187);
xor U10874 (N_10874,N_8925,N_8468);
nor U10875 (N_10875,N_9913,N_9491);
nand U10876 (N_10876,N_8886,N_9705);
and U10877 (N_10877,N_8742,N_8174);
nor U10878 (N_10878,N_8426,N_8328);
or U10879 (N_10879,N_8537,N_9853);
xnor U10880 (N_10880,N_9930,N_9774);
nand U10881 (N_10881,N_8323,N_9593);
nand U10882 (N_10882,N_8852,N_8620);
xor U10883 (N_10883,N_9539,N_9300);
nor U10884 (N_10884,N_8663,N_8172);
nand U10885 (N_10885,N_9123,N_8977);
nand U10886 (N_10886,N_9250,N_9690);
nor U10887 (N_10887,N_8186,N_8276);
nand U10888 (N_10888,N_8887,N_8850);
or U10889 (N_10889,N_8382,N_8331);
nand U10890 (N_10890,N_8316,N_9415);
or U10891 (N_10891,N_8145,N_9490);
xor U10892 (N_10892,N_9710,N_8405);
or U10893 (N_10893,N_9803,N_9756);
or U10894 (N_10894,N_8002,N_9460);
xnor U10895 (N_10895,N_9681,N_9246);
and U10896 (N_10896,N_9311,N_8362);
xor U10897 (N_10897,N_8344,N_8913);
nand U10898 (N_10898,N_9580,N_9471);
and U10899 (N_10899,N_9328,N_8937);
or U10900 (N_10900,N_8072,N_9622);
nand U10901 (N_10901,N_8086,N_9534);
nor U10902 (N_10902,N_8800,N_9416);
nor U10903 (N_10903,N_9243,N_9659);
nand U10904 (N_10904,N_8607,N_8418);
nor U10905 (N_10905,N_8773,N_8149);
nor U10906 (N_10906,N_8752,N_9314);
nor U10907 (N_10907,N_9211,N_8152);
and U10908 (N_10908,N_8899,N_9423);
or U10909 (N_10909,N_8246,N_9164);
nand U10910 (N_10910,N_9072,N_9466);
and U10911 (N_10911,N_9577,N_8878);
and U10912 (N_10912,N_8922,N_8775);
xnor U10913 (N_10913,N_9852,N_9812);
and U10914 (N_10914,N_8366,N_8335);
nand U10915 (N_10915,N_9963,N_8948);
nand U10916 (N_10916,N_8745,N_8699);
nand U10917 (N_10917,N_8161,N_9337);
or U10918 (N_10918,N_8797,N_9369);
nor U10919 (N_10919,N_8342,N_9134);
nor U10920 (N_10920,N_8494,N_8195);
and U10921 (N_10921,N_9304,N_8644);
and U10922 (N_10922,N_8357,N_8604);
xor U10923 (N_10923,N_9106,N_9469);
and U10924 (N_10924,N_9644,N_9527);
nand U10925 (N_10925,N_9281,N_9384);
nor U10926 (N_10926,N_8734,N_8524);
or U10927 (N_10927,N_9907,N_8818);
nand U10928 (N_10928,N_9533,N_8085);
nor U10929 (N_10929,N_9042,N_8220);
and U10930 (N_10930,N_9448,N_8048);
or U10931 (N_10931,N_8660,N_8706);
nor U10932 (N_10932,N_8647,N_9009);
and U10933 (N_10933,N_9932,N_9597);
nor U10934 (N_10934,N_9067,N_9113);
and U10935 (N_10935,N_9910,N_9501);
nand U10936 (N_10936,N_9677,N_8410);
nand U10937 (N_10937,N_9341,N_9486);
or U10938 (N_10938,N_9230,N_9049);
nand U10939 (N_10939,N_9984,N_8651);
nor U10940 (N_10940,N_9385,N_8226);
nand U10941 (N_10941,N_9014,N_8184);
xnor U10942 (N_10942,N_9766,N_8774);
or U10943 (N_10943,N_9110,N_8698);
nand U10944 (N_10944,N_9291,N_9816);
xor U10945 (N_10945,N_8714,N_8740);
or U10946 (N_10946,N_9244,N_8639);
nand U10947 (N_10947,N_9965,N_9329);
nand U10948 (N_10948,N_8719,N_8963);
or U10949 (N_10949,N_9383,N_8349);
or U10950 (N_10950,N_9035,N_9195);
and U10951 (N_10951,N_9769,N_8250);
or U10952 (N_10952,N_8868,N_9961);
and U10953 (N_10953,N_8143,N_8896);
or U10954 (N_10954,N_8900,N_8240);
xnor U10955 (N_10955,N_9104,N_9445);
and U10956 (N_10956,N_8063,N_9735);
or U10957 (N_10957,N_9140,N_9753);
nand U10958 (N_10958,N_8135,N_8369);
or U10959 (N_10959,N_9217,N_8452);
or U10960 (N_10960,N_8923,N_9579);
or U10961 (N_10961,N_8224,N_8375);
xnor U10962 (N_10962,N_8249,N_8169);
and U10963 (N_10963,N_8208,N_8364);
xor U10964 (N_10964,N_8157,N_9289);
and U10965 (N_10965,N_9061,N_9086);
nand U10966 (N_10966,N_8151,N_9343);
nor U10967 (N_10967,N_8803,N_9611);
xnor U10968 (N_10968,N_8741,N_8075);
nor U10969 (N_10969,N_8018,N_8795);
nand U10970 (N_10970,N_9276,N_8131);
or U10971 (N_10971,N_9931,N_9985);
and U10972 (N_10972,N_8895,N_9850);
nand U10973 (N_10973,N_9761,N_9903);
nand U10974 (N_10974,N_9157,N_8065);
nor U10975 (N_10975,N_9658,N_8671);
xnor U10976 (N_10976,N_9809,N_9748);
nor U10977 (N_10977,N_8049,N_9707);
and U10978 (N_10978,N_8215,N_8189);
and U10979 (N_10979,N_8574,N_9322);
nand U10980 (N_10980,N_8411,N_8327);
nor U10981 (N_10981,N_8481,N_9204);
nor U10982 (N_10982,N_8056,N_9632);
and U10983 (N_10983,N_9248,N_8562);
xnor U10984 (N_10984,N_9880,N_9544);
and U10985 (N_10985,N_9408,N_9199);
and U10986 (N_10986,N_8119,N_9401);
and U10987 (N_10987,N_8541,N_8554);
nor U10988 (N_10988,N_8885,N_9092);
or U10989 (N_10989,N_9569,N_8317);
and U10990 (N_10990,N_9089,N_8381);
and U10991 (N_10991,N_8333,N_9820);
nand U10992 (N_10992,N_9578,N_8099);
and U10993 (N_10993,N_8851,N_9807);
nand U10994 (N_10994,N_8435,N_9452);
nand U10995 (N_10995,N_9894,N_9326);
or U10996 (N_10996,N_9790,N_8354);
or U10997 (N_10997,N_8120,N_9004);
and U10998 (N_10998,N_8789,N_9706);
or U10999 (N_10999,N_8577,N_9628);
and U11000 (N_11000,N_8620,N_9787);
nand U11001 (N_11001,N_8256,N_8908);
nand U11002 (N_11002,N_8078,N_8443);
nor U11003 (N_11003,N_8510,N_9732);
xor U11004 (N_11004,N_9094,N_9622);
nor U11005 (N_11005,N_8795,N_8443);
xor U11006 (N_11006,N_8594,N_9207);
and U11007 (N_11007,N_9759,N_9243);
nor U11008 (N_11008,N_9184,N_9403);
xor U11009 (N_11009,N_9579,N_8181);
nand U11010 (N_11010,N_9262,N_9819);
xor U11011 (N_11011,N_8559,N_9036);
xnor U11012 (N_11012,N_8913,N_8923);
nand U11013 (N_11013,N_8820,N_9910);
or U11014 (N_11014,N_8073,N_8623);
or U11015 (N_11015,N_9542,N_9168);
or U11016 (N_11016,N_8764,N_9001);
xor U11017 (N_11017,N_8425,N_8526);
or U11018 (N_11018,N_8520,N_9753);
nand U11019 (N_11019,N_9126,N_8198);
nor U11020 (N_11020,N_9545,N_9396);
and U11021 (N_11021,N_8774,N_9771);
nor U11022 (N_11022,N_9801,N_8056);
nor U11023 (N_11023,N_9979,N_9293);
xnor U11024 (N_11024,N_9816,N_8238);
nand U11025 (N_11025,N_9597,N_8202);
and U11026 (N_11026,N_9483,N_9476);
and U11027 (N_11027,N_8163,N_9962);
or U11028 (N_11028,N_9835,N_8444);
nand U11029 (N_11029,N_8538,N_8626);
nand U11030 (N_11030,N_9821,N_8466);
and U11031 (N_11031,N_9847,N_8045);
nand U11032 (N_11032,N_9573,N_8770);
xnor U11033 (N_11033,N_8695,N_8797);
or U11034 (N_11034,N_8371,N_8176);
and U11035 (N_11035,N_8819,N_8716);
nor U11036 (N_11036,N_8745,N_8134);
or U11037 (N_11037,N_9130,N_9389);
or U11038 (N_11038,N_8358,N_8721);
or U11039 (N_11039,N_8324,N_8621);
xor U11040 (N_11040,N_8545,N_9214);
and U11041 (N_11041,N_8670,N_8459);
xor U11042 (N_11042,N_8843,N_9743);
nand U11043 (N_11043,N_9840,N_8248);
nand U11044 (N_11044,N_9878,N_9298);
xor U11045 (N_11045,N_9915,N_9369);
or U11046 (N_11046,N_8302,N_9146);
and U11047 (N_11047,N_8235,N_9292);
or U11048 (N_11048,N_8384,N_9072);
and U11049 (N_11049,N_8588,N_8059);
nor U11050 (N_11050,N_8981,N_9170);
nand U11051 (N_11051,N_8801,N_8305);
or U11052 (N_11052,N_9408,N_8263);
and U11053 (N_11053,N_8499,N_8935);
nand U11054 (N_11054,N_9196,N_8439);
nor U11055 (N_11055,N_9206,N_9931);
xor U11056 (N_11056,N_8234,N_9387);
and U11057 (N_11057,N_8109,N_9331);
nor U11058 (N_11058,N_9843,N_9004);
nand U11059 (N_11059,N_9893,N_9164);
nor U11060 (N_11060,N_8993,N_8458);
nand U11061 (N_11061,N_9939,N_8110);
nand U11062 (N_11062,N_8120,N_9561);
or U11063 (N_11063,N_8225,N_9710);
nor U11064 (N_11064,N_8447,N_8472);
nor U11065 (N_11065,N_9133,N_8655);
nand U11066 (N_11066,N_9822,N_9913);
or U11067 (N_11067,N_8583,N_9416);
xor U11068 (N_11068,N_8616,N_9129);
xnor U11069 (N_11069,N_9986,N_9681);
nand U11070 (N_11070,N_8310,N_8035);
or U11071 (N_11071,N_9922,N_9690);
xnor U11072 (N_11072,N_9867,N_9778);
xor U11073 (N_11073,N_8471,N_9735);
nor U11074 (N_11074,N_9568,N_9815);
nor U11075 (N_11075,N_9361,N_9196);
nand U11076 (N_11076,N_9185,N_9914);
and U11077 (N_11077,N_9210,N_9147);
and U11078 (N_11078,N_8294,N_9625);
or U11079 (N_11079,N_8597,N_8288);
nor U11080 (N_11080,N_8185,N_9511);
nand U11081 (N_11081,N_8149,N_8872);
xnor U11082 (N_11082,N_8232,N_8606);
xor U11083 (N_11083,N_9255,N_8917);
nand U11084 (N_11084,N_9761,N_9465);
xor U11085 (N_11085,N_8645,N_8765);
nor U11086 (N_11086,N_9545,N_8547);
nand U11087 (N_11087,N_8414,N_8375);
and U11088 (N_11088,N_8107,N_8135);
and U11089 (N_11089,N_8960,N_8785);
nor U11090 (N_11090,N_9295,N_9239);
nor U11091 (N_11091,N_9615,N_8280);
xor U11092 (N_11092,N_9234,N_9191);
nor U11093 (N_11093,N_8780,N_8998);
nand U11094 (N_11094,N_8392,N_8339);
nand U11095 (N_11095,N_9425,N_9610);
xor U11096 (N_11096,N_9119,N_8317);
nand U11097 (N_11097,N_8316,N_8422);
xor U11098 (N_11098,N_8181,N_8399);
xnor U11099 (N_11099,N_9804,N_9912);
nand U11100 (N_11100,N_8334,N_9418);
xnor U11101 (N_11101,N_9913,N_9902);
or U11102 (N_11102,N_9098,N_8614);
nor U11103 (N_11103,N_9299,N_8732);
xor U11104 (N_11104,N_9193,N_8691);
or U11105 (N_11105,N_9493,N_9078);
nand U11106 (N_11106,N_8550,N_9799);
nor U11107 (N_11107,N_9488,N_8753);
nand U11108 (N_11108,N_8570,N_8421);
and U11109 (N_11109,N_9537,N_8166);
xor U11110 (N_11110,N_9474,N_9579);
nor U11111 (N_11111,N_9897,N_9809);
xnor U11112 (N_11112,N_9388,N_9674);
nor U11113 (N_11113,N_9818,N_8949);
and U11114 (N_11114,N_9488,N_8595);
and U11115 (N_11115,N_8507,N_8430);
and U11116 (N_11116,N_9314,N_8126);
and U11117 (N_11117,N_8171,N_8644);
or U11118 (N_11118,N_9685,N_9925);
xnor U11119 (N_11119,N_9685,N_8296);
or U11120 (N_11120,N_8731,N_9327);
and U11121 (N_11121,N_8216,N_8658);
and U11122 (N_11122,N_8218,N_9393);
or U11123 (N_11123,N_8488,N_8565);
nand U11124 (N_11124,N_8066,N_9216);
nor U11125 (N_11125,N_9408,N_8285);
xor U11126 (N_11126,N_8311,N_9645);
xnor U11127 (N_11127,N_8541,N_9123);
nand U11128 (N_11128,N_9580,N_8178);
xnor U11129 (N_11129,N_8015,N_8385);
xnor U11130 (N_11130,N_8080,N_8413);
xor U11131 (N_11131,N_8497,N_8910);
xnor U11132 (N_11132,N_8792,N_9632);
or U11133 (N_11133,N_8557,N_9016);
nand U11134 (N_11134,N_9301,N_9770);
and U11135 (N_11135,N_9744,N_9043);
nand U11136 (N_11136,N_9088,N_8961);
nand U11137 (N_11137,N_8804,N_8213);
nor U11138 (N_11138,N_8305,N_8106);
xnor U11139 (N_11139,N_9432,N_9101);
or U11140 (N_11140,N_9332,N_9611);
xor U11141 (N_11141,N_9966,N_9207);
xor U11142 (N_11142,N_8381,N_8807);
nand U11143 (N_11143,N_9341,N_8284);
nand U11144 (N_11144,N_9271,N_8901);
and U11145 (N_11145,N_8800,N_9421);
nand U11146 (N_11146,N_9830,N_8015);
or U11147 (N_11147,N_8931,N_9826);
or U11148 (N_11148,N_8459,N_9353);
and U11149 (N_11149,N_9066,N_8715);
and U11150 (N_11150,N_8214,N_8821);
and U11151 (N_11151,N_9868,N_8537);
and U11152 (N_11152,N_8242,N_9007);
and U11153 (N_11153,N_9349,N_8147);
and U11154 (N_11154,N_8291,N_8511);
or U11155 (N_11155,N_9304,N_8788);
nand U11156 (N_11156,N_8189,N_9188);
and U11157 (N_11157,N_8237,N_9397);
or U11158 (N_11158,N_8709,N_8396);
nor U11159 (N_11159,N_9442,N_9440);
or U11160 (N_11160,N_8778,N_8717);
nand U11161 (N_11161,N_9573,N_8183);
xor U11162 (N_11162,N_9298,N_9970);
or U11163 (N_11163,N_9890,N_9904);
and U11164 (N_11164,N_8364,N_8181);
or U11165 (N_11165,N_8966,N_9741);
nor U11166 (N_11166,N_9582,N_9852);
or U11167 (N_11167,N_9482,N_8832);
nand U11168 (N_11168,N_8069,N_8918);
nand U11169 (N_11169,N_9290,N_9381);
xnor U11170 (N_11170,N_8732,N_9663);
and U11171 (N_11171,N_8494,N_8740);
or U11172 (N_11172,N_9075,N_9566);
xnor U11173 (N_11173,N_8565,N_9894);
nor U11174 (N_11174,N_8981,N_8939);
and U11175 (N_11175,N_8602,N_9051);
nor U11176 (N_11176,N_9936,N_9948);
and U11177 (N_11177,N_9884,N_9914);
and U11178 (N_11178,N_9526,N_9944);
or U11179 (N_11179,N_9459,N_9914);
nand U11180 (N_11180,N_9396,N_8045);
or U11181 (N_11181,N_9108,N_8980);
and U11182 (N_11182,N_9290,N_8283);
or U11183 (N_11183,N_9208,N_9430);
nor U11184 (N_11184,N_9813,N_8001);
or U11185 (N_11185,N_8093,N_9296);
or U11186 (N_11186,N_9926,N_8858);
or U11187 (N_11187,N_8584,N_9707);
or U11188 (N_11188,N_8150,N_8825);
nand U11189 (N_11189,N_8066,N_9116);
xnor U11190 (N_11190,N_9109,N_8319);
or U11191 (N_11191,N_9579,N_8653);
xnor U11192 (N_11192,N_9062,N_9777);
nor U11193 (N_11193,N_9778,N_8117);
nor U11194 (N_11194,N_9957,N_8679);
nand U11195 (N_11195,N_8608,N_9173);
nand U11196 (N_11196,N_8154,N_9301);
and U11197 (N_11197,N_8781,N_8200);
and U11198 (N_11198,N_9568,N_8658);
nand U11199 (N_11199,N_8593,N_8838);
nor U11200 (N_11200,N_8389,N_9529);
xor U11201 (N_11201,N_9321,N_9038);
xor U11202 (N_11202,N_8317,N_8659);
and U11203 (N_11203,N_9175,N_8185);
nand U11204 (N_11204,N_9438,N_9684);
nor U11205 (N_11205,N_8002,N_9977);
nand U11206 (N_11206,N_9376,N_8059);
nor U11207 (N_11207,N_9259,N_8148);
xor U11208 (N_11208,N_8763,N_9769);
nand U11209 (N_11209,N_8740,N_9243);
nand U11210 (N_11210,N_8804,N_9582);
nand U11211 (N_11211,N_8388,N_9446);
nor U11212 (N_11212,N_8528,N_9270);
and U11213 (N_11213,N_8000,N_8482);
or U11214 (N_11214,N_8883,N_8195);
or U11215 (N_11215,N_8548,N_8379);
nand U11216 (N_11216,N_9062,N_8239);
nor U11217 (N_11217,N_9476,N_8011);
nor U11218 (N_11218,N_8138,N_8149);
nand U11219 (N_11219,N_9086,N_8279);
nand U11220 (N_11220,N_9688,N_8515);
nor U11221 (N_11221,N_9378,N_8273);
or U11222 (N_11222,N_9701,N_9042);
and U11223 (N_11223,N_8939,N_9468);
nand U11224 (N_11224,N_9058,N_8381);
nor U11225 (N_11225,N_9750,N_9769);
or U11226 (N_11226,N_9912,N_9135);
nand U11227 (N_11227,N_9798,N_9483);
and U11228 (N_11228,N_9124,N_8269);
or U11229 (N_11229,N_9045,N_8971);
nor U11230 (N_11230,N_8592,N_8839);
nand U11231 (N_11231,N_8905,N_8181);
xor U11232 (N_11232,N_9425,N_9744);
xnor U11233 (N_11233,N_8189,N_9231);
or U11234 (N_11234,N_9767,N_9752);
nor U11235 (N_11235,N_8971,N_9128);
and U11236 (N_11236,N_8834,N_8219);
nor U11237 (N_11237,N_9705,N_9771);
and U11238 (N_11238,N_8226,N_9243);
xor U11239 (N_11239,N_8044,N_8038);
and U11240 (N_11240,N_8523,N_9447);
nand U11241 (N_11241,N_8442,N_9778);
nand U11242 (N_11242,N_9704,N_8527);
nor U11243 (N_11243,N_8180,N_9076);
xor U11244 (N_11244,N_9354,N_9777);
nand U11245 (N_11245,N_9572,N_8049);
and U11246 (N_11246,N_8106,N_8104);
xnor U11247 (N_11247,N_9460,N_8741);
xnor U11248 (N_11248,N_8583,N_9614);
xnor U11249 (N_11249,N_9565,N_8976);
nand U11250 (N_11250,N_9053,N_9425);
and U11251 (N_11251,N_9222,N_9781);
and U11252 (N_11252,N_9031,N_9131);
or U11253 (N_11253,N_8318,N_8462);
and U11254 (N_11254,N_8449,N_9246);
and U11255 (N_11255,N_9670,N_8210);
nor U11256 (N_11256,N_9897,N_9675);
and U11257 (N_11257,N_8501,N_9285);
nor U11258 (N_11258,N_9097,N_8976);
nand U11259 (N_11259,N_9760,N_8411);
xnor U11260 (N_11260,N_9596,N_8238);
nand U11261 (N_11261,N_9546,N_9489);
or U11262 (N_11262,N_8820,N_9948);
or U11263 (N_11263,N_8020,N_8154);
xnor U11264 (N_11264,N_8879,N_9112);
nand U11265 (N_11265,N_8016,N_9181);
xor U11266 (N_11266,N_9261,N_9582);
xnor U11267 (N_11267,N_8857,N_9695);
or U11268 (N_11268,N_9048,N_9398);
or U11269 (N_11269,N_9754,N_9719);
nor U11270 (N_11270,N_8423,N_9970);
and U11271 (N_11271,N_8156,N_9688);
and U11272 (N_11272,N_9535,N_9749);
and U11273 (N_11273,N_8532,N_9707);
xnor U11274 (N_11274,N_9547,N_9003);
xor U11275 (N_11275,N_8089,N_8023);
nor U11276 (N_11276,N_8231,N_8065);
nor U11277 (N_11277,N_8068,N_9272);
xor U11278 (N_11278,N_9778,N_9134);
and U11279 (N_11279,N_8878,N_9000);
or U11280 (N_11280,N_9622,N_8624);
xnor U11281 (N_11281,N_8180,N_8453);
nand U11282 (N_11282,N_8256,N_9951);
or U11283 (N_11283,N_8623,N_9485);
or U11284 (N_11284,N_8546,N_9420);
xor U11285 (N_11285,N_8971,N_8021);
nor U11286 (N_11286,N_9807,N_9830);
and U11287 (N_11287,N_9857,N_9880);
nand U11288 (N_11288,N_9869,N_9799);
xnor U11289 (N_11289,N_9213,N_9395);
xnor U11290 (N_11290,N_8970,N_8787);
xnor U11291 (N_11291,N_9987,N_9659);
nor U11292 (N_11292,N_9094,N_8276);
nand U11293 (N_11293,N_9877,N_8633);
nand U11294 (N_11294,N_8328,N_9504);
nor U11295 (N_11295,N_8851,N_9061);
and U11296 (N_11296,N_8070,N_8812);
or U11297 (N_11297,N_8222,N_9245);
nor U11298 (N_11298,N_9902,N_9492);
and U11299 (N_11299,N_9433,N_8870);
nand U11300 (N_11300,N_8813,N_9667);
nand U11301 (N_11301,N_8262,N_8381);
xnor U11302 (N_11302,N_9043,N_9732);
nor U11303 (N_11303,N_8425,N_8699);
or U11304 (N_11304,N_8514,N_9688);
or U11305 (N_11305,N_9944,N_8592);
nor U11306 (N_11306,N_8073,N_8562);
xor U11307 (N_11307,N_8145,N_9913);
xnor U11308 (N_11308,N_8958,N_8345);
nand U11309 (N_11309,N_8833,N_9899);
nor U11310 (N_11310,N_9582,N_8745);
nand U11311 (N_11311,N_8749,N_8670);
and U11312 (N_11312,N_9207,N_9433);
and U11313 (N_11313,N_8520,N_9155);
nand U11314 (N_11314,N_8189,N_9798);
and U11315 (N_11315,N_8266,N_8490);
nor U11316 (N_11316,N_9909,N_8902);
or U11317 (N_11317,N_9333,N_8331);
and U11318 (N_11318,N_9294,N_9916);
nand U11319 (N_11319,N_9682,N_8163);
nor U11320 (N_11320,N_8065,N_8920);
xor U11321 (N_11321,N_9858,N_8617);
xnor U11322 (N_11322,N_9575,N_9294);
xnor U11323 (N_11323,N_8078,N_8990);
nor U11324 (N_11324,N_8895,N_8522);
or U11325 (N_11325,N_9164,N_9463);
xnor U11326 (N_11326,N_9345,N_9899);
xnor U11327 (N_11327,N_9794,N_8562);
nor U11328 (N_11328,N_9555,N_8675);
nand U11329 (N_11329,N_8727,N_9494);
nor U11330 (N_11330,N_9934,N_9346);
or U11331 (N_11331,N_9760,N_9429);
nand U11332 (N_11332,N_8340,N_9606);
nand U11333 (N_11333,N_8026,N_8079);
nand U11334 (N_11334,N_8796,N_8893);
xor U11335 (N_11335,N_9544,N_9099);
xnor U11336 (N_11336,N_8374,N_9264);
xor U11337 (N_11337,N_9550,N_9551);
and U11338 (N_11338,N_9937,N_8992);
or U11339 (N_11339,N_9339,N_8449);
nor U11340 (N_11340,N_8700,N_8742);
or U11341 (N_11341,N_8739,N_9290);
xor U11342 (N_11342,N_9696,N_9150);
nor U11343 (N_11343,N_9129,N_8336);
nand U11344 (N_11344,N_9665,N_8497);
nor U11345 (N_11345,N_9791,N_8191);
nand U11346 (N_11346,N_9683,N_9228);
nand U11347 (N_11347,N_9252,N_8908);
nor U11348 (N_11348,N_8806,N_9243);
or U11349 (N_11349,N_9097,N_9716);
or U11350 (N_11350,N_8865,N_9691);
or U11351 (N_11351,N_9211,N_9560);
or U11352 (N_11352,N_9487,N_9802);
and U11353 (N_11353,N_9855,N_8224);
or U11354 (N_11354,N_9834,N_8635);
nand U11355 (N_11355,N_9254,N_9308);
or U11356 (N_11356,N_9754,N_8686);
and U11357 (N_11357,N_9865,N_9553);
xnor U11358 (N_11358,N_9345,N_9949);
xor U11359 (N_11359,N_8222,N_8117);
and U11360 (N_11360,N_9567,N_9627);
nand U11361 (N_11361,N_8313,N_8765);
and U11362 (N_11362,N_8678,N_8671);
or U11363 (N_11363,N_8884,N_8492);
nand U11364 (N_11364,N_8157,N_9346);
or U11365 (N_11365,N_9522,N_8010);
nand U11366 (N_11366,N_9657,N_8629);
xor U11367 (N_11367,N_8142,N_9536);
or U11368 (N_11368,N_9437,N_8530);
xnor U11369 (N_11369,N_8335,N_8713);
and U11370 (N_11370,N_8775,N_8310);
nand U11371 (N_11371,N_9433,N_9598);
and U11372 (N_11372,N_9414,N_9253);
nor U11373 (N_11373,N_8457,N_9425);
and U11374 (N_11374,N_9474,N_9954);
nand U11375 (N_11375,N_8671,N_8608);
xor U11376 (N_11376,N_8535,N_9220);
and U11377 (N_11377,N_8194,N_9489);
nor U11378 (N_11378,N_9584,N_9741);
or U11379 (N_11379,N_8396,N_8962);
nand U11380 (N_11380,N_8940,N_8939);
xnor U11381 (N_11381,N_9086,N_8055);
or U11382 (N_11382,N_8981,N_9009);
and U11383 (N_11383,N_8581,N_8671);
or U11384 (N_11384,N_9531,N_8273);
xor U11385 (N_11385,N_9034,N_9000);
nand U11386 (N_11386,N_8951,N_8815);
or U11387 (N_11387,N_9523,N_9516);
xnor U11388 (N_11388,N_9730,N_8730);
and U11389 (N_11389,N_8603,N_9405);
xnor U11390 (N_11390,N_9829,N_8245);
or U11391 (N_11391,N_9800,N_9497);
nor U11392 (N_11392,N_8324,N_8586);
and U11393 (N_11393,N_9682,N_9053);
nor U11394 (N_11394,N_9760,N_8694);
nor U11395 (N_11395,N_8952,N_8331);
xnor U11396 (N_11396,N_9334,N_9773);
or U11397 (N_11397,N_8378,N_8425);
and U11398 (N_11398,N_9060,N_8581);
and U11399 (N_11399,N_9493,N_9937);
and U11400 (N_11400,N_9995,N_8551);
nor U11401 (N_11401,N_8609,N_9491);
xor U11402 (N_11402,N_8892,N_9573);
nand U11403 (N_11403,N_8676,N_9747);
xnor U11404 (N_11404,N_9354,N_9937);
nand U11405 (N_11405,N_8402,N_8151);
xnor U11406 (N_11406,N_9349,N_9631);
and U11407 (N_11407,N_8107,N_8949);
nor U11408 (N_11408,N_9737,N_8967);
xor U11409 (N_11409,N_9367,N_8514);
nor U11410 (N_11410,N_8463,N_8772);
nand U11411 (N_11411,N_8664,N_9601);
xnor U11412 (N_11412,N_8398,N_8984);
or U11413 (N_11413,N_8988,N_8431);
nor U11414 (N_11414,N_8172,N_8658);
nand U11415 (N_11415,N_9974,N_8250);
xor U11416 (N_11416,N_8520,N_8200);
and U11417 (N_11417,N_9414,N_8976);
xor U11418 (N_11418,N_9709,N_9958);
xor U11419 (N_11419,N_8185,N_8016);
nand U11420 (N_11420,N_8467,N_9316);
and U11421 (N_11421,N_9097,N_9972);
or U11422 (N_11422,N_8629,N_8083);
or U11423 (N_11423,N_8909,N_8245);
or U11424 (N_11424,N_9720,N_8079);
nor U11425 (N_11425,N_9086,N_9610);
xnor U11426 (N_11426,N_8916,N_9913);
xnor U11427 (N_11427,N_8530,N_9452);
or U11428 (N_11428,N_9883,N_9160);
and U11429 (N_11429,N_9377,N_9786);
xor U11430 (N_11430,N_9639,N_8660);
or U11431 (N_11431,N_9933,N_9909);
nor U11432 (N_11432,N_9577,N_8406);
nand U11433 (N_11433,N_8500,N_8440);
or U11434 (N_11434,N_8222,N_9389);
nand U11435 (N_11435,N_8572,N_9233);
and U11436 (N_11436,N_8202,N_8273);
nand U11437 (N_11437,N_8453,N_9148);
and U11438 (N_11438,N_8851,N_8517);
and U11439 (N_11439,N_8203,N_8137);
or U11440 (N_11440,N_8158,N_9867);
or U11441 (N_11441,N_8674,N_8029);
xnor U11442 (N_11442,N_8676,N_8728);
or U11443 (N_11443,N_8692,N_9765);
xnor U11444 (N_11444,N_8016,N_9691);
xnor U11445 (N_11445,N_9635,N_9046);
nand U11446 (N_11446,N_8504,N_8766);
nand U11447 (N_11447,N_9385,N_8911);
or U11448 (N_11448,N_9673,N_9568);
and U11449 (N_11449,N_9474,N_8903);
xor U11450 (N_11450,N_9347,N_9409);
or U11451 (N_11451,N_8362,N_9519);
nor U11452 (N_11452,N_9873,N_9807);
and U11453 (N_11453,N_9379,N_8822);
and U11454 (N_11454,N_8410,N_9850);
and U11455 (N_11455,N_9481,N_9000);
nor U11456 (N_11456,N_8981,N_8108);
xnor U11457 (N_11457,N_9407,N_9993);
or U11458 (N_11458,N_9804,N_8653);
nor U11459 (N_11459,N_8181,N_8608);
nor U11460 (N_11460,N_8423,N_9786);
nand U11461 (N_11461,N_8374,N_9779);
nor U11462 (N_11462,N_8286,N_8824);
or U11463 (N_11463,N_9348,N_8358);
nor U11464 (N_11464,N_9688,N_8210);
nor U11465 (N_11465,N_8788,N_8175);
nand U11466 (N_11466,N_9973,N_8766);
nand U11467 (N_11467,N_8378,N_9456);
nand U11468 (N_11468,N_9625,N_8858);
nand U11469 (N_11469,N_9182,N_8728);
or U11470 (N_11470,N_9050,N_9802);
or U11471 (N_11471,N_8050,N_8468);
nor U11472 (N_11472,N_8353,N_8069);
or U11473 (N_11473,N_8817,N_9398);
nand U11474 (N_11474,N_8222,N_8376);
nand U11475 (N_11475,N_8716,N_8118);
xor U11476 (N_11476,N_8546,N_9606);
or U11477 (N_11477,N_9599,N_8953);
xnor U11478 (N_11478,N_8038,N_8837);
and U11479 (N_11479,N_9603,N_9963);
nor U11480 (N_11480,N_9552,N_9298);
xnor U11481 (N_11481,N_8812,N_8041);
xor U11482 (N_11482,N_9363,N_9654);
or U11483 (N_11483,N_9607,N_9032);
and U11484 (N_11484,N_8484,N_9802);
nor U11485 (N_11485,N_8306,N_9609);
and U11486 (N_11486,N_9144,N_9172);
or U11487 (N_11487,N_8880,N_9084);
xnor U11488 (N_11488,N_9324,N_9696);
or U11489 (N_11489,N_9463,N_9572);
xor U11490 (N_11490,N_8218,N_8455);
nor U11491 (N_11491,N_9626,N_8857);
or U11492 (N_11492,N_8897,N_8063);
nand U11493 (N_11493,N_8864,N_8876);
xnor U11494 (N_11494,N_8305,N_8431);
xnor U11495 (N_11495,N_9138,N_8572);
or U11496 (N_11496,N_8981,N_9420);
nor U11497 (N_11497,N_9641,N_9025);
nor U11498 (N_11498,N_8928,N_8407);
nand U11499 (N_11499,N_8274,N_9454);
nor U11500 (N_11500,N_8884,N_9026);
nand U11501 (N_11501,N_8373,N_9289);
or U11502 (N_11502,N_9500,N_9945);
and U11503 (N_11503,N_8347,N_8507);
nand U11504 (N_11504,N_9946,N_8649);
nor U11505 (N_11505,N_8588,N_9799);
xnor U11506 (N_11506,N_9647,N_8732);
nand U11507 (N_11507,N_9051,N_9717);
nor U11508 (N_11508,N_8285,N_9799);
xor U11509 (N_11509,N_9320,N_9020);
or U11510 (N_11510,N_9169,N_8296);
or U11511 (N_11511,N_8807,N_9444);
xor U11512 (N_11512,N_8108,N_9551);
or U11513 (N_11513,N_9223,N_8019);
nand U11514 (N_11514,N_8706,N_8351);
or U11515 (N_11515,N_8732,N_9650);
and U11516 (N_11516,N_9381,N_8586);
or U11517 (N_11517,N_9068,N_8583);
nor U11518 (N_11518,N_9454,N_9400);
nand U11519 (N_11519,N_8980,N_8323);
nor U11520 (N_11520,N_8226,N_9757);
nor U11521 (N_11521,N_9059,N_9062);
and U11522 (N_11522,N_9386,N_9265);
or U11523 (N_11523,N_9079,N_9601);
or U11524 (N_11524,N_8544,N_8780);
xnor U11525 (N_11525,N_9204,N_9584);
nand U11526 (N_11526,N_9598,N_9730);
xor U11527 (N_11527,N_8782,N_9525);
and U11528 (N_11528,N_8915,N_8258);
or U11529 (N_11529,N_9483,N_8527);
nor U11530 (N_11530,N_8727,N_8358);
or U11531 (N_11531,N_9423,N_9989);
and U11532 (N_11532,N_8898,N_9866);
or U11533 (N_11533,N_9268,N_8271);
and U11534 (N_11534,N_9414,N_8636);
nand U11535 (N_11535,N_8575,N_9891);
or U11536 (N_11536,N_9090,N_8892);
and U11537 (N_11537,N_8554,N_9570);
or U11538 (N_11538,N_8227,N_9809);
xnor U11539 (N_11539,N_9330,N_9181);
or U11540 (N_11540,N_9632,N_9335);
or U11541 (N_11541,N_8763,N_9703);
nand U11542 (N_11542,N_9519,N_8939);
nand U11543 (N_11543,N_8943,N_8373);
and U11544 (N_11544,N_8414,N_8396);
nand U11545 (N_11545,N_9659,N_9382);
nand U11546 (N_11546,N_9844,N_9886);
nand U11547 (N_11547,N_9776,N_8157);
nor U11548 (N_11548,N_8764,N_8398);
and U11549 (N_11549,N_8021,N_8611);
nor U11550 (N_11550,N_9405,N_9494);
nand U11551 (N_11551,N_8759,N_9417);
and U11552 (N_11552,N_8254,N_8392);
and U11553 (N_11553,N_9698,N_9010);
nor U11554 (N_11554,N_8360,N_9858);
or U11555 (N_11555,N_8782,N_9063);
or U11556 (N_11556,N_8377,N_9522);
nor U11557 (N_11557,N_9177,N_9132);
or U11558 (N_11558,N_9360,N_9201);
or U11559 (N_11559,N_8372,N_8353);
nor U11560 (N_11560,N_8421,N_9411);
xnor U11561 (N_11561,N_8859,N_8231);
nor U11562 (N_11562,N_8059,N_8359);
or U11563 (N_11563,N_8333,N_8210);
nand U11564 (N_11564,N_9159,N_8374);
nand U11565 (N_11565,N_9581,N_8042);
xnor U11566 (N_11566,N_8088,N_8411);
or U11567 (N_11567,N_8523,N_8079);
nand U11568 (N_11568,N_9958,N_9322);
and U11569 (N_11569,N_8770,N_8359);
and U11570 (N_11570,N_9875,N_9580);
and U11571 (N_11571,N_8459,N_9517);
nor U11572 (N_11572,N_8447,N_9712);
and U11573 (N_11573,N_9382,N_8051);
nand U11574 (N_11574,N_8986,N_9116);
xor U11575 (N_11575,N_9482,N_9526);
or U11576 (N_11576,N_9590,N_9936);
nor U11577 (N_11577,N_8501,N_9407);
xor U11578 (N_11578,N_9396,N_9264);
nand U11579 (N_11579,N_9099,N_8795);
or U11580 (N_11580,N_8962,N_9644);
and U11581 (N_11581,N_8699,N_9869);
xor U11582 (N_11582,N_8296,N_8801);
or U11583 (N_11583,N_9403,N_9949);
xnor U11584 (N_11584,N_9144,N_8608);
nor U11585 (N_11585,N_8514,N_9504);
or U11586 (N_11586,N_8888,N_8539);
xnor U11587 (N_11587,N_9370,N_8437);
xnor U11588 (N_11588,N_8541,N_8924);
xnor U11589 (N_11589,N_8292,N_9009);
xnor U11590 (N_11590,N_9135,N_8611);
nor U11591 (N_11591,N_9478,N_8195);
xnor U11592 (N_11592,N_8275,N_8506);
nand U11593 (N_11593,N_8644,N_9076);
or U11594 (N_11594,N_8361,N_9468);
xor U11595 (N_11595,N_8815,N_8862);
and U11596 (N_11596,N_9534,N_9809);
or U11597 (N_11597,N_9340,N_8783);
and U11598 (N_11598,N_8385,N_9557);
nor U11599 (N_11599,N_8690,N_8716);
nand U11600 (N_11600,N_9507,N_9367);
nor U11601 (N_11601,N_9676,N_9639);
or U11602 (N_11602,N_8419,N_9171);
xor U11603 (N_11603,N_9437,N_9236);
and U11604 (N_11604,N_9163,N_8952);
nand U11605 (N_11605,N_9760,N_9734);
nor U11606 (N_11606,N_8874,N_9584);
xor U11607 (N_11607,N_9308,N_8311);
xor U11608 (N_11608,N_8546,N_9265);
or U11609 (N_11609,N_9292,N_8723);
xor U11610 (N_11610,N_8619,N_9335);
nor U11611 (N_11611,N_8536,N_8663);
and U11612 (N_11612,N_8007,N_9990);
and U11613 (N_11613,N_8789,N_8278);
nor U11614 (N_11614,N_9003,N_9226);
xnor U11615 (N_11615,N_8328,N_9533);
nor U11616 (N_11616,N_9195,N_8144);
nand U11617 (N_11617,N_9754,N_8368);
or U11618 (N_11618,N_9747,N_8137);
nor U11619 (N_11619,N_8570,N_9134);
or U11620 (N_11620,N_8411,N_8542);
xnor U11621 (N_11621,N_8388,N_9445);
nand U11622 (N_11622,N_8240,N_9824);
nor U11623 (N_11623,N_8876,N_9886);
or U11624 (N_11624,N_9247,N_9783);
nor U11625 (N_11625,N_9974,N_8806);
or U11626 (N_11626,N_9748,N_8483);
and U11627 (N_11627,N_8858,N_8035);
xor U11628 (N_11628,N_9917,N_9468);
nor U11629 (N_11629,N_8279,N_8529);
xor U11630 (N_11630,N_9240,N_8028);
nand U11631 (N_11631,N_9530,N_8882);
nand U11632 (N_11632,N_8631,N_9440);
nand U11633 (N_11633,N_9786,N_8593);
and U11634 (N_11634,N_8884,N_9890);
nor U11635 (N_11635,N_9292,N_8422);
nor U11636 (N_11636,N_8253,N_8101);
nand U11637 (N_11637,N_8561,N_8769);
or U11638 (N_11638,N_9926,N_9108);
and U11639 (N_11639,N_9307,N_8439);
or U11640 (N_11640,N_8856,N_9995);
xnor U11641 (N_11641,N_8842,N_9048);
and U11642 (N_11642,N_9754,N_9523);
or U11643 (N_11643,N_8137,N_9993);
nand U11644 (N_11644,N_9645,N_8832);
nand U11645 (N_11645,N_8919,N_9665);
or U11646 (N_11646,N_9013,N_9127);
xnor U11647 (N_11647,N_8400,N_8325);
nor U11648 (N_11648,N_9831,N_8632);
nor U11649 (N_11649,N_9107,N_8663);
and U11650 (N_11650,N_8381,N_8823);
and U11651 (N_11651,N_9726,N_8666);
and U11652 (N_11652,N_8703,N_8766);
or U11653 (N_11653,N_8988,N_9604);
or U11654 (N_11654,N_8740,N_9164);
nor U11655 (N_11655,N_9542,N_9984);
or U11656 (N_11656,N_9994,N_8401);
nand U11657 (N_11657,N_8290,N_9104);
or U11658 (N_11658,N_8529,N_8632);
and U11659 (N_11659,N_9496,N_8076);
and U11660 (N_11660,N_8721,N_9527);
xor U11661 (N_11661,N_8143,N_8358);
xor U11662 (N_11662,N_9658,N_8537);
or U11663 (N_11663,N_9789,N_9512);
nand U11664 (N_11664,N_8431,N_9497);
nor U11665 (N_11665,N_8102,N_9312);
nor U11666 (N_11666,N_8192,N_9507);
or U11667 (N_11667,N_9537,N_8639);
and U11668 (N_11668,N_9098,N_9301);
and U11669 (N_11669,N_8856,N_9871);
nand U11670 (N_11670,N_8804,N_8660);
nand U11671 (N_11671,N_9635,N_8538);
or U11672 (N_11672,N_8942,N_9896);
xor U11673 (N_11673,N_8082,N_9803);
nand U11674 (N_11674,N_8390,N_9155);
nor U11675 (N_11675,N_9120,N_8675);
or U11676 (N_11676,N_9626,N_9509);
xor U11677 (N_11677,N_9995,N_9246);
nor U11678 (N_11678,N_8248,N_8296);
xor U11679 (N_11679,N_9431,N_8485);
or U11680 (N_11680,N_9577,N_8082);
nor U11681 (N_11681,N_9670,N_9603);
nand U11682 (N_11682,N_9784,N_8308);
or U11683 (N_11683,N_9288,N_8402);
xnor U11684 (N_11684,N_8139,N_8593);
xor U11685 (N_11685,N_9413,N_9713);
nand U11686 (N_11686,N_9560,N_9299);
nand U11687 (N_11687,N_8372,N_9452);
xor U11688 (N_11688,N_9630,N_9185);
nor U11689 (N_11689,N_8092,N_9318);
and U11690 (N_11690,N_8203,N_8967);
nand U11691 (N_11691,N_9139,N_9283);
or U11692 (N_11692,N_9828,N_8709);
xor U11693 (N_11693,N_9006,N_8950);
nand U11694 (N_11694,N_9873,N_9510);
nand U11695 (N_11695,N_8703,N_8839);
nand U11696 (N_11696,N_8468,N_9035);
nand U11697 (N_11697,N_9112,N_8587);
or U11698 (N_11698,N_9201,N_8519);
or U11699 (N_11699,N_8688,N_9303);
xnor U11700 (N_11700,N_9447,N_9082);
or U11701 (N_11701,N_8528,N_8800);
xnor U11702 (N_11702,N_8690,N_8321);
nor U11703 (N_11703,N_9894,N_9124);
xnor U11704 (N_11704,N_8786,N_9482);
xnor U11705 (N_11705,N_9581,N_8944);
xnor U11706 (N_11706,N_9428,N_8005);
xor U11707 (N_11707,N_9198,N_8180);
nand U11708 (N_11708,N_8147,N_9303);
or U11709 (N_11709,N_9294,N_8407);
nor U11710 (N_11710,N_8178,N_9514);
nor U11711 (N_11711,N_9134,N_9031);
nand U11712 (N_11712,N_9450,N_8950);
xor U11713 (N_11713,N_9401,N_9035);
xor U11714 (N_11714,N_8448,N_8649);
nor U11715 (N_11715,N_9757,N_8228);
and U11716 (N_11716,N_8561,N_8052);
xnor U11717 (N_11717,N_8955,N_9755);
and U11718 (N_11718,N_9191,N_9150);
nand U11719 (N_11719,N_8275,N_8867);
nor U11720 (N_11720,N_9117,N_9143);
nand U11721 (N_11721,N_9636,N_9815);
and U11722 (N_11722,N_8671,N_8509);
and U11723 (N_11723,N_9881,N_9394);
and U11724 (N_11724,N_8917,N_8407);
or U11725 (N_11725,N_9252,N_8853);
xnor U11726 (N_11726,N_9678,N_8120);
and U11727 (N_11727,N_9923,N_8073);
or U11728 (N_11728,N_9074,N_9058);
and U11729 (N_11729,N_9647,N_9486);
xor U11730 (N_11730,N_9159,N_8687);
and U11731 (N_11731,N_8561,N_9718);
nand U11732 (N_11732,N_9806,N_8710);
nor U11733 (N_11733,N_8476,N_8016);
and U11734 (N_11734,N_8269,N_9815);
nor U11735 (N_11735,N_8404,N_9521);
nor U11736 (N_11736,N_9133,N_8776);
nand U11737 (N_11737,N_9963,N_9036);
nor U11738 (N_11738,N_9823,N_8458);
and U11739 (N_11739,N_8972,N_8513);
nand U11740 (N_11740,N_9617,N_8325);
nand U11741 (N_11741,N_9332,N_8752);
and U11742 (N_11742,N_8831,N_9788);
or U11743 (N_11743,N_8474,N_9822);
nor U11744 (N_11744,N_8312,N_9363);
nand U11745 (N_11745,N_8760,N_8098);
nand U11746 (N_11746,N_8929,N_9148);
nor U11747 (N_11747,N_8629,N_8147);
or U11748 (N_11748,N_9394,N_9779);
nand U11749 (N_11749,N_8513,N_9169);
or U11750 (N_11750,N_8540,N_8744);
xnor U11751 (N_11751,N_8333,N_9713);
or U11752 (N_11752,N_9764,N_9751);
nor U11753 (N_11753,N_9125,N_9461);
and U11754 (N_11754,N_9379,N_9641);
or U11755 (N_11755,N_8754,N_8332);
nand U11756 (N_11756,N_9791,N_9171);
and U11757 (N_11757,N_8288,N_8745);
or U11758 (N_11758,N_8445,N_9944);
or U11759 (N_11759,N_9536,N_9066);
nand U11760 (N_11760,N_9149,N_8822);
xor U11761 (N_11761,N_8098,N_8418);
xnor U11762 (N_11762,N_9329,N_9534);
and U11763 (N_11763,N_8176,N_8402);
xor U11764 (N_11764,N_9739,N_9279);
or U11765 (N_11765,N_8937,N_8222);
and U11766 (N_11766,N_8055,N_9262);
xor U11767 (N_11767,N_9057,N_9942);
or U11768 (N_11768,N_9060,N_9664);
or U11769 (N_11769,N_9320,N_8910);
and U11770 (N_11770,N_8884,N_9768);
or U11771 (N_11771,N_8357,N_9329);
nor U11772 (N_11772,N_9167,N_9129);
or U11773 (N_11773,N_8965,N_9827);
nor U11774 (N_11774,N_9026,N_8722);
nor U11775 (N_11775,N_8813,N_8537);
xor U11776 (N_11776,N_9361,N_8759);
xor U11777 (N_11777,N_9770,N_9702);
and U11778 (N_11778,N_9355,N_8339);
xnor U11779 (N_11779,N_9266,N_8966);
nor U11780 (N_11780,N_8072,N_9165);
or U11781 (N_11781,N_8765,N_8288);
or U11782 (N_11782,N_9863,N_9727);
and U11783 (N_11783,N_8925,N_8613);
nor U11784 (N_11784,N_8137,N_8248);
xor U11785 (N_11785,N_8001,N_8018);
or U11786 (N_11786,N_8209,N_9171);
nor U11787 (N_11787,N_8716,N_9689);
xnor U11788 (N_11788,N_8688,N_8949);
nor U11789 (N_11789,N_9737,N_8715);
xnor U11790 (N_11790,N_8979,N_9518);
or U11791 (N_11791,N_9501,N_9623);
and U11792 (N_11792,N_9990,N_9077);
xor U11793 (N_11793,N_8318,N_9436);
and U11794 (N_11794,N_9644,N_9377);
or U11795 (N_11795,N_8951,N_9602);
xnor U11796 (N_11796,N_9701,N_9598);
and U11797 (N_11797,N_8376,N_9877);
xor U11798 (N_11798,N_9281,N_9101);
nor U11799 (N_11799,N_8397,N_9898);
and U11800 (N_11800,N_9966,N_9238);
nand U11801 (N_11801,N_9405,N_9037);
xnor U11802 (N_11802,N_8376,N_8118);
and U11803 (N_11803,N_9502,N_8180);
and U11804 (N_11804,N_9735,N_9100);
nor U11805 (N_11805,N_9951,N_8174);
and U11806 (N_11806,N_8197,N_9174);
xnor U11807 (N_11807,N_8065,N_9999);
and U11808 (N_11808,N_8371,N_8423);
nand U11809 (N_11809,N_8555,N_9027);
xnor U11810 (N_11810,N_9129,N_9783);
or U11811 (N_11811,N_9106,N_9096);
or U11812 (N_11812,N_9275,N_8367);
and U11813 (N_11813,N_9780,N_9428);
and U11814 (N_11814,N_8672,N_9335);
or U11815 (N_11815,N_8274,N_9093);
nor U11816 (N_11816,N_9957,N_8986);
and U11817 (N_11817,N_8993,N_8029);
or U11818 (N_11818,N_9342,N_8703);
nor U11819 (N_11819,N_8391,N_8103);
nor U11820 (N_11820,N_9490,N_8364);
or U11821 (N_11821,N_9386,N_8566);
nand U11822 (N_11822,N_8795,N_8178);
and U11823 (N_11823,N_9403,N_8574);
nor U11824 (N_11824,N_8750,N_8950);
or U11825 (N_11825,N_8352,N_8104);
nor U11826 (N_11826,N_9332,N_8391);
xnor U11827 (N_11827,N_8177,N_8973);
and U11828 (N_11828,N_9923,N_8971);
nand U11829 (N_11829,N_9883,N_9379);
nor U11830 (N_11830,N_9107,N_9998);
nand U11831 (N_11831,N_9685,N_9510);
and U11832 (N_11832,N_8349,N_9594);
xnor U11833 (N_11833,N_9031,N_8104);
and U11834 (N_11834,N_8598,N_8319);
xor U11835 (N_11835,N_8267,N_9864);
and U11836 (N_11836,N_8114,N_9389);
xnor U11837 (N_11837,N_9107,N_9710);
and U11838 (N_11838,N_8579,N_8071);
nand U11839 (N_11839,N_9318,N_9868);
and U11840 (N_11840,N_8386,N_9776);
xnor U11841 (N_11841,N_9862,N_9435);
and U11842 (N_11842,N_8988,N_8882);
nand U11843 (N_11843,N_8150,N_9704);
nor U11844 (N_11844,N_8666,N_8578);
or U11845 (N_11845,N_8031,N_8043);
nand U11846 (N_11846,N_9296,N_8568);
xor U11847 (N_11847,N_9589,N_9270);
and U11848 (N_11848,N_9180,N_9442);
xor U11849 (N_11849,N_8823,N_9948);
nor U11850 (N_11850,N_9254,N_9339);
nand U11851 (N_11851,N_8753,N_8627);
nand U11852 (N_11852,N_8831,N_8352);
nand U11853 (N_11853,N_8744,N_8240);
nor U11854 (N_11854,N_9741,N_8424);
xnor U11855 (N_11855,N_8630,N_9761);
nor U11856 (N_11856,N_9851,N_9893);
and U11857 (N_11857,N_9087,N_8870);
xor U11858 (N_11858,N_8048,N_8626);
nand U11859 (N_11859,N_8422,N_8778);
and U11860 (N_11860,N_9296,N_9726);
and U11861 (N_11861,N_8300,N_9007);
nand U11862 (N_11862,N_9599,N_9750);
nand U11863 (N_11863,N_8071,N_9057);
and U11864 (N_11864,N_9384,N_8045);
nor U11865 (N_11865,N_8495,N_8778);
and U11866 (N_11866,N_8135,N_8982);
nand U11867 (N_11867,N_8152,N_9857);
xor U11868 (N_11868,N_8939,N_9246);
xnor U11869 (N_11869,N_9862,N_9037);
xor U11870 (N_11870,N_9703,N_9876);
nor U11871 (N_11871,N_9249,N_9713);
or U11872 (N_11872,N_9276,N_9686);
and U11873 (N_11873,N_8763,N_8606);
and U11874 (N_11874,N_8616,N_8794);
nor U11875 (N_11875,N_8750,N_9582);
nand U11876 (N_11876,N_9323,N_9316);
nand U11877 (N_11877,N_8811,N_8517);
xor U11878 (N_11878,N_8814,N_9193);
or U11879 (N_11879,N_9443,N_9606);
nor U11880 (N_11880,N_8586,N_9480);
and U11881 (N_11881,N_9425,N_8759);
and U11882 (N_11882,N_9118,N_8992);
or U11883 (N_11883,N_8818,N_8315);
and U11884 (N_11884,N_9754,N_8298);
and U11885 (N_11885,N_9223,N_8107);
or U11886 (N_11886,N_9994,N_9709);
and U11887 (N_11887,N_8285,N_9774);
nand U11888 (N_11888,N_9978,N_8174);
xor U11889 (N_11889,N_9536,N_9512);
xor U11890 (N_11890,N_8392,N_9524);
nor U11891 (N_11891,N_8677,N_8018);
or U11892 (N_11892,N_8257,N_9531);
and U11893 (N_11893,N_9634,N_8915);
nand U11894 (N_11894,N_8094,N_9014);
nor U11895 (N_11895,N_9568,N_9244);
nor U11896 (N_11896,N_8230,N_9795);
and U11897 (N_11897,N_9907,N_9947);
nand U11898 (N_11898,N_8521,N_9370);
or U11899 (N_11899,N_9553,N_9418);
or U11900 (N_11900,N_9182,N_9425);
xor U11901 (N_11901,N_9541,N_8542);
xor U11902 (N_11902,N_8837,N_9901);
or U11903 (N_11903,N_8048,N_8023);
xor U11904 (N_11904,N_8602,N_8578);
nand U11905 (N_11905,N_9090,N_8393);
nand U11906 (N_11906,N_9601,N_8430);
xor U11907 (N_11907,N_9490,N_9453);
or U11908 (N_11908,N_8223,N_9459);
and U11909 (N_11909,N_8306,N_8031);
and U11910 (N_11910,N_9063,N_9523);
and U11911 (N_11911,N_8408,N_8913);
nor U11912 (N_11912,N_8788,N_8715);
xnor U11913 (N_11913,N_9103,N_9749);
or U11914 (N_11914,N_8248,N_9604);
nor U11915 (N_11915,N_9818,N_8708);
and U11916 (N_11916,N_8563,N_9512);
xor U11917 (N_11917,N_9908,N_9549);
and U11918 (N_11918,N_8978,N_8565);
nor U11919 (N_11919,N_9597,N_9348);
and U11920 (N_11920,N_8267,N_8542);
nor U11921 (N_11921,N_9591,N_9218);
xnor U11922 (N_11922,N_9917,N_9015);
nand U11923 (N_11923,N_9993,N_9753);
or U11924 (N_11924,N_8218,N_9151);
nand U11925 (N_11925,N_9507,N_9688);
nand U11926 (N_11926,N_8805,N_8889);
nor U11927 (N_11927,N_8760,N_8839);
and U11928 (N_11928,N_8420,N_8844);
nor U11929 (N_11929,N_9352,N_9609);
nor U11930 (N_11930,N_8818,N_9720);
xor U11931 (N_11931,N_9370,N_8368);
nand U11932 (N_11932,N_8177,N_8283);
xor U11933 (N_11933,N_8307,N_8912);
or U11934 (N_11934,N_8238,N_9817);
and U11935 (N_11935,N_9372,N_9989);
nor U11936 (N_11936,N_9362,N_8108);
or U11937 (N_11937,N_9420,N_8114);
nand U11938 (N_11938,N_8524,N_9315);
xor U11939 (N_11939,N_8367,N_9143);
and U11940 (N_11940,N_9430,N_9333);
and U11941 (N_11941,N_9008,N_9852);
nand U11942 (N_11942,N_9161,N_8004);
nor U11943 (N_11943,N_8331,N_8259);
or U11944 (N_11944,N_8634,N_9715);
or U11945 (N_11945,N_8247,N_9162);
nor U11946 (N_11946,N_8097,N_8077);
or U11947 (N_11947,N_9774,N_8266);
and U11948 (N_11948,N_8842,N_8424);
xnor U11949 (N_11949,N_8652,N_9588);
and U11950 (N_11950,N_8545,N_9796);
xor U11951 (N_11951,N_8353,N_8099);
and U11952 (N_11952,N_9140,N_8169);
nor U11953 (N_11953,N_9346,N_8076);
or U11954 (N_11954,N_9477,N_9687);
and U11955 (N_11955,N_8442,N_8284);
nor U11956 (N_11956,N_9598,N_8087);
and U11957 (N_11957,N_9287,N_8032);
nor U11958 (N_11958,N_9639,N_9451);
nor U11959 (N_11959,N_8477,N_8620);
and U11960 (N_11960,N_9479,N_9929);
nand U11961 (N_11961,N_9546,N_8757);
nand U11962 (N_11962,N_9841,N_8636);
and U11963 (N_11963,N_9630,N_8343);
and U11964 (N_11964,N_9425,N_8350);
nor U11965 (N_11965,N_8296,N_8109);
xor U11966 (N_11966,N_9072,N_9691);
nor U11967 (N_11967,N_8287,N_9870);
nand U11968 (N_11968,N_9932,N_9964);
and U11969 (N_11969,N_9795,N_8668);
xor U11970 (N_11970,N_8573,N_9321);
and U11971 (N_11971,N_8737,N_8849);
xor U11972 (N_11972,N_8735,N_8773);
xnor U11973 (N_11973,N_9018,N_9213);
nor U11974 (N_11974,N_9856,N_9423);
nor U11975 (N_11975,N_8829,N_9480);
nand U11976 (N_11976,N_9584,N_8155);
and U11977 (N_11977,N_8211,N_9547);
nand U11978 (N_11978,N_8373,N_8773);
or U11979 (N_11979,N_8219,N_9401);
nand U11980 (N_11980,N_9058,N_8577);
or U11981 (N_11981,N_8766,N_9475);
xor U11982 (N_11982,N_8608,N_8702);
nor U11983 (N_11983,N_8699,N_8211);
nor U11984 (N_11984,N_9738,N_9732);
nand U11985 (N_11985,N_9320,N_8059);
xnor U11986 (N_11986,N_8881,N_9146);
xnor U11987 (N_11987,N_8713,N_8846);
xor U11988 (N_11988,N_8707,N_9696);
nand U11989 (N_11989,N_9168,N_9751);
nor U11990 (N_11990,N_8370,N_8831);
and U11991 (N_11991,N_9859,N_8620);
or U11992 (N_11992,N_9293,N_9585);
xor U11993 (N_11993,N_8175,N_8899);
nand U11994 (N_11994,N_9711,N_8397);
nand U11995 (N_11995,N_8449,N_8054);
xor U11996 (N_11996,N_9140,N_9315);
nor U11997 (N_11997,N_9662,N_8757);
or U11998 (N_11998,N_8917,N_8688);
nand U11999 (N_11999,N_8297,N_8446);
nand U12000 (N_12000,N_11907,N_10335);
nand U12001 (N_12001,N_11514,N_10135);
and U12002 (N_12002,N_11697,N_11884);
nand U12003 (N_12003,N_10993,N_11572);
and U12004 (N_12004,N_10205,N_10535);
nor U12005 (N_12005,N_10833,N_10204);
xnor U12006 (N_12006,N_10911,N_10354);
nor U12007 (N_12007,N_10608,N_11401);
and U12008 (N_12008,N_11552,N_11836);
xor U12009 (N_12009,N_10018,N_10864);
or U12010 (N_12010,N_10572,N_11379);
nand U12011 (N_12011,N_11449,N_10991);
nand U12012 (N_12012,N_10656,N_11067);
xor U12013 (N_12013,N_11420,N_10471);
nand U12014 (N_12014,N_10464,N_10341);
nor U12015 (N_12015,N_10176,N_11002);
nor U12016 (N_12016,N_11911,N_11322);
and U12017 (N_12017,N_11868,N_11977);
nand U12018 (N_12018,N_11672,N_11016);
xnor U12019 (N_12019,N_11518,N_10006);
or U12020 (N_12020,N_10177,N_11240);
nand U12021 (N_12021,N_11460,N_10585);
and U12022 (N_12022,N_10104,N_11300);
or U12023 (N_12023,N_11490,N_11472);
xor U12024 (N_12024,N_10545,N_11849);
xor U12025 (N_12025,N_10754,N_11644);
xnor U12026 (N_12026,N_10769,N_11081);
and U12027 (N_12027,N_11660,N_11237);
nand U12028 (N_12028,N_11045,N_10131);
nor U12029 (N_12029,N_11835,N_11283);
nor U12030 (N_12030,N_11329,N_10939);
nor U12031 (N_12031,N_10450,N_11007);
xnor U12032 (N_12032,N_10706,N_11787);
nand U12033 (N_12033,N_10792,N_11422);
xor U12034 (N_12034,N_10718,N_10893);
nand U12035 (N_12035,N_11500,N_10343);
nand U12036 (N_12036,N_11064,N_10597);
and U12037 (N_12037,N_10404,N_11639);
or U12038 (N_12038,N_11469,N_11618);
and U12039 (N_12039,N_11436,N_11980);
or U12040 (N_12040,N_10857,N_10764);
nor U12041 (N_12041,N_11963,N_11171);
nand U12042 (N_12042,N_10897,N_11889);
and U12043 (N_12043,N_11194,N_11854);
xnor U12044 (N_12044,N_10870,N_10509);
nor U12045 (N_12045,N_10440,N_11990);
nor U12046 (N_12046,N_10869,N_10175);
nor U12047 (N_12047,N_10529,N_11954);
xor U12048 (N_12048,N_10125,N_11669);
or U12049 (N_12049,N_10133,N_11374);
nor U12050 (N_12050,N_10198,N_11904);
or U12051 (N_12051,N_10277,N_11798);
nor U12052 (N_12052,N_10802,N_10689);
nor U12053 (N_12053,N_11465,N_11871);
or U12054 (N_12054,N_11225,N_11192);
or U12055 (N_12055,N_11061,N_10673);
nor U12056 (N_12056,N_11381,N_11668);
xor U12057 (N_12057,N_10720,N_11955);
or U12058 (N_12058,N_10553,N_11933);
nor U12059 (N_12059,N_11456,N_10181);
xnor U12060 (N_12060,N_11321,N_10733);
or U12061 (N_12061,N_10919,N_10598);
xor U12062 (N_12062,N_11245,N_10069);
nor U12063 (N_12063,N_11914,N_11820);
xor U12064 (N_12064,N_11698,N_10022);
nand U12065 (N_12065,N_11020,N_11799);
xor U12066 (N_12066,N_11227,N_10308);
nand U12067 (N_12067,N_10820,N_10846);
nor U12068 (N_12068,N_11768,N_11367);
and U12069 (N_12069,N_11804,N_11785);
and U12070 (N_12070,N_11855,N_11615);
nor U12071 (N_12071,N_11119,N_11177);
and U12072 (N_12072,N_10452,N_11471);
and U12073 (N_12073,N_11372,N_11291);
nand U12074 (N_12074,N_11675,N_10514);
and U12075 (N_12075,N_10194,N_11583);
and U12076 (N_12076,N_10881,N_10155);
xor U12077 (N_12077,N_11896,N_10167);
nor U12078 (N_12078,N_11579,N_10504);
or U12079 (N_12079,N_11637,N_10490);
or U12080 (N_12080,N_10945,N_10542);
and U12081 (N_12081,N_10537,N_11663);
and U12082 (N_12082,N_10587,N_11488);
nor U12083 (N_12083,N_10770,N_11478);
xnor U12084 (N_12084,N_11450,N_10879);
nor U12085 (N_12085,N_10562,N_10650);
and U12086 (N_12086,N_10639,N_11997);
nor U12087 (N_12087,N_11247,N_11519);
nor U12088 (N_12088,N_11666,N_11203);
and U12089 (N_12089,N_11094,N_10146);
and U12090 (N_12090,N_11805,N_10474);
xnor U12091 (N_12091,N_10653,N_10121);
and U12092 (N_12092,N_10613,N_10189);
xnor U12093 (N_12093,N_11426,N_11215);
xor U12094 (N_12094,N_10842,N_11320);
or U12095 (N_12095,N_10551,N_11221);
nor U12096 (N_12096,N_11130,N_11921);
nand U12097 (N_12097,N_10749,N_11585);
xnor U12098 (N_12098,N_10352,N_10703);
xnor U12099 (N_12099,N_11342,N_11968);
or U12100 (N_12100,N_10560,N_10226);
nand U12101 (N_12101,N_10465,N_10491);
or U12102 (N_12102,N_11695,N_11416);
and U12103 (N_12103,N_10307,N_10238);
xnor U12104 (N_12104,N_10264,N_10375);
xor U12105 (N_12105,N_10372,N_10259);
or U12106 (N_12106,N_11197,N_10654);
or U12107 (N_12107,N_10616,N_11040);
or U12108 (N_12108,N_11485,N_11333);
or U12109 (N_12109,N_11984,N_11605);
nand U12110 (N_12110,N_11959,N_11070);
nand U12111 (N_12111,N_11285,N_10975);
nand U12112 (N_12112,N_11818,N_10547);
xor U12113 (N_12113,N_10351,N_11096);
or U12114 (N_12114,N_10959,N_10324);
nand U12115 (N_12115,N_10056,N_10643);
nor U12116 (N_12116,N_11512,N_10583);
nor U12117 (N_12117,N_10461,N_10215);
nor U12118 (N_12118,N_10773,N_11793);
xor U12119 (N_12119,N_10149,N_10822);
and U12120 (N_12120,N_11920,N_10012);
and U12121 (N_12121,N_10274,N_10139);
nand U12122 (N_12122,N_11011,N_11995);
and U12123 (N_12123,N_10419,N_10309);
and U12124 (N_12124,N_11009,N_10065);
nand U12125 (N_12125,N_10291,N_11112);
xor U12126 (N_12126,N_11147,N_11101);
nand U12127 (N_12127,N_10969,N_11674);
and U12128 (N_12128,N_10000,N_11159);
nand U12129 (N_12129,N_10541,N_10891);
nor U12130 (N_12130,N_10719,N_11358);
or U12131 (N_12131,N_10029,N_10449);
or U12132 (N_12132,N_10632,N_11025);
and U12133 (N_12133,N_10861,N_11445);
or U12134 (N_12134,N_11763,N_10921);
and U12135 (N_12135,N_11391,N_11457);
and U12136 (N_12136,N_11684,N_10809);
nand U12137 (N_12137,N_10457,N_11761);
nand U12138 (N_12138,N_10142,N_11719);
xor U12139 (N_12139,N_10928,N_11625);
xnor U12140 (N_12140,N_10637,N_11577);
and U12141 (N_12141,N_10326,N_11392);
xor U12142 (N_12142,N_11330,N_11410);
xor U12143 (N_12143,N_11287,N_10297);
or U12144 (N_12144,N_11417,N_10401);
or U12145 (N_12145,N_10625,N_11802);
and U12146 (N_12146,N_10768,N_10025);
xor U12147 (N_12147,N_10112,N_11468);
and U12148 (N_12148,N_10377,N_10912);
xnor U12149 (N_12149,N_10564,N_10480);
or U12150 (N_12150,N_10340,N_11250);
xor U12151 (N_12151,N_11738,N_11305);
xor U12152 (N_12152,N_11759,N_10827);
and U12153 (N_12153,N_11275,N_11754);
or U12154 (N_12154,N_10527,N_11459);
or U12155 (N_12155,N_10365,N_10859);
xor U12156 (N_12156,N_10217,N_10031);
or U12157 (N_12157,N_10954,N_11442);
nor U12158 (N_12158,N_11753,N_11875);
nand U12159 (N_12159,N_11090,N_10477);
nor U12160 (N_12160,N_10096,N_11125);
nand U12161 (N_12161,N_11857,N_10977);
and U12162 (N_12162,N_11053,N_11279);
and U12163 (N_12163,N_11630,N_10120);
or U12164 (N_12164,N_10400,N_10624);
nand U12165 (N_12165,N_10698,N_11217);
xor U12166 (N_12166,N_11923,N_10294);
nor U12167 (N_12167,N_10552,N_11302);
nand U12168 (N_12168,N_11492,N_10426);
or U12169 (N_12169,N_10323,N_11777);
and U12170 (N_12170,N_10874,N_10390);
and U12171 (N_12171,N_10479,N_11715);
xnor U12172 (N_12172,N_11794,N_11981);
nand U12173 (N_12173,N_10392,N_10575);
or U12174 (N_12174,N_11455,N_10038);
or U12175 (N_12175,N_10618,N_10011);
nand U12176 (N_12176,N_10684,N_11109);
or U12177 (N_12177,N_11035,N_10851);
or U12178 (N_12178,N_10866,N_10638);
nand U12179 (N_12179,N_11246,N_10856);
or U12180 (N_12180,N_11852,N_11945);
nand U12181 (N_12181,N_10787,N_11735);
nand U12182 (N_12182,N_10523,N_11386);
nand U12183 (N_12183,N_11729,N_11862);
xor U12184 (N_12184,N_10434,N_10243);
nor U12185 (N_12185,N_11876,N_10248);
nand U12186 (N_12186,N_11551,N_10708);
or U12187 (N_12187,N_10399,N_10116);
xnor U12188 (N_12188,N_11652,N_11328);
nor U12189 (N_12189,N_11208,N_11758);
or U12190 (N_12190,N_11614,N_10492);
or U12191 (N_12191,N_11253,N_10686);
and U12192 (N_12192,N_10994,N_10699);
or U12193 (N_12193,N_11567,N_11860);
or U12194 (N_12194,N_11676,N_11545);
nor U12195 (N_12195,N_10060,N_11654);
or U12196 (N_12196,N_11202,N_10130);
xnor U12197 (N_12197,N_11093,N_11178);
or U12198 (N_12198,N_11702,N_10843);
or U12199 (N_12199,N_11057,N_11557);
nor U12200 (N_12200,N_10990,N_11865);
nand U12201 (N_12201,N_11494,N_10301);
and U12202 (N_12202,N_10091,N_11710);
nand U12203 (N_12203,N_11778,N_11937);
nor U12204 (N_12204,N_11408,N_10070);
nor U12205 (N_12205,N_10900,N_10152);
xnor U12206 (N_12206,N_10321,N_11581);
xnor U12207 (N_12207,N_11462,N_10383);
nor U12208 (N_12208,N_11277,N_11947);
and U12209 (N_12209,N_11791,N_11482);
xnor U12210 (N_12210,N_11063,N_10315);
xor U12211 (N_12211,N_11601,N_11620);
or U12212 (N_12212,N_11789,N_10207);
nand U12213 (N_12213,N_11730,N_10772);
or U12214 (N_12214,N_11176,N_11306);
or U12215 (N_12215,N_10953,N_10935);
and U12216 (N_12216,N_10019,N_10561);
nor U12217 (N_12217,N_11080,N_11304);
xnor U12218 (N_12218,N_10493,N_10995);
nand U12219 (N_12219,N_11726,N_10791);
nor U12220 (N_12220,N_11993,N_11931);
or U12221 (N_12221,N_11878,N_10310);
and U12222 (N_12222,N_10111,N_11623);
xnor U12223 (N_12223,N_11788,N_10532);
nor U12224 (N_12224,N_10077,N_11260);
nand U12225 (N_12225,N_11099,N_10565);
and U12226 (N_12226,N_11095,N_11207);
nand U12227 (N_12227,N_11434,N_10105);
xnor U12228 (N_12228,N_10909,N_11111);
nor U12229 (N_12229,N_11925,N_10089);
xnor U12230 (N_12230,N_10412,N_11236);
nor U12231 (N_12231,N_11999,N_11262);
nand U12232 (N_12232,N_10807,N_10735);
nand U12233 (N_12233,N_10408,N_10320);
xnor U12234 (N_12234,N_11017,N_10166);
and U12235 (N_12235,N_10800,N_11167);
nor U12236 (N_12236,N_11256,N_10360);
xor U12237 (N_12237,N_10732,N_11932);
xor U12238 (N_12238,N_11983,N_11022);
or U12239 (N_12239,N_11812,N_11430);
nor U12240 (N_12240,N_11191,N_11604);
nor U12241 (N_12241,N_11748,N_10405);
nand U12242 (N_12242,N_11476,N_10244);
nor U12243 (N_12243,N_11319,N_11389);
or U12244 (N_12244,N_11106,N_11909);
nor U12245 (N_12245,N_10968,N_11866);
nor U12246 (N_12246,N_10629,N_11743);
xnor U12247 (N_12247,N_11830,N_10593);
nor U12248 (N_12248,N_11506,N_11324);
and U12249 (N_12249,N_11446,N_11104);
or U12250 (N_12250,N_10236,N_11251);
nor U12251 (N_12251,N_11559,N_11633);
and U12252 (N_12252,N_10495,N_11964);
and U12253 (N_12253,N_10611,N_11635);
nand U12254 (N_12254,N_10898,N_10314);
xor U12255 (N_12255,N_10222,N_10270);
nor U12256 (N_12256,N_11419,N_11882);
or U12257 (N_12257,N_10905,N_10439);
nor U12258 (N_12258,N_11249,N_11072);
nand U12259 (N_12259,N_10781,N_10087);
nand U12260 (N_12260,N_11824,N_10299);
or U12261 (N_12261,N_10382,N_10290);
nand U12262 (N_12262,N_11004,N_10160);
nor U12263 (N_12263,N_11609,N_10536);
nor U12264 (N_12264,N_10132,N_11313);
xor U12265 (N_12265,N_10498,N_10469);
and U12266 (N_12266,N_10986,N_10026);
or U12267 (N_12267,N_11670,N_10403);
and U12268 (N_12268,N_11910,N_11575);
or U12269 (N_12269,N_11032,N_11483);
or U12270 (N_12270,N_10020,N_10860);
and U12271 (N_12271,N_11825,N_10978);
and U12272 (N_12272,N_10933,N_11948);
xor U12273 (N_12273,N_11438,N_11443);
nand U12274 (N_12274,N_11913,N_11523);
xnor U12275 (N_12275,N_11049,N_10963);
nor U12276 (N_12276,N_10162,N_10228);
xnor U12277 (N_12277,N_11412,N_11133);
or U12278 (N_12278,N_11394,N_10245);
nand U12279 (N_12279,N_11359,N_11731);
nand U12280 (N_12280,N_10811,N_11747);
nand U12281 (N_12281,N_11856,N_10473);
nor U12282 (N_12282,N_10088,N_10558);
nor U12283 (N_12283,N_10885,N_10159);
or U12284 (N_12284,N_11773,N_11607);
or U12285 (N_12285,N_10338,N_10080);
xnor U12286 (N_12286,N_11685,N_10771);
and U12287 (N_12287,N_11894,N_11077);
xnor U12288 (N_12288,N_11965,N_10714);
xor U12289 (N_12289,N_11509,N_11209);
xnor U12290 (N_12290,N_11037,N_10958);
nor U12291 (N_12291,N_11272,N_10119);
nor U12292 (N_12292,N_11254,N_11205);
or U12293 (N_12293,N_10203,N_11843);
nand U12294 (N_12294,N_10083,N_10927);
nand U12295 (N_12295,N_10701,N_11929);
nand U12296 (N_12296,N_11562,N_10154);
or U12297 (N_12297,N_10641,N_10141);
or U12298 (N_12298,N_10705,N_11346);
nor U12299 (N_12299,N_10946,N_10790);
and U12300 (N_12300,N_10191,N_10554);
or U12301 (N_12301,N_10917,N_11850);
and U12302 (N_12302,N_10023,N_10265);
nand U12303 (N_12303,N_10361,N_10630);
and U12304 (N_12304,N_11853,N_10128);
and U12305 (N_12305,N_10894,N_11421);
nor U12306 (N_12306,N_11396,N_10303);
or U12307 (N_12307,N_10016,N_10187);
xor U12308 (N_12308,N_10432,N_11881);
nor U12309 (N_12309,N_10455,N_11621);
or U12310 (N_12310,N_10284,N_10915);
and U12311 (N_12311,N_10559,N_11586);
nand U12312 (N_12312,N_10370,N_10153);
xor U12313 (N_12313,N_11645,N_11549);
xnor U12314 (N_12314,N_10193,N_11477);
or U12315 (N_12315,N_10039,N_11362);
nor U12316 (N_12316,N_11339,N_11949);
or U12317 (N_12317,N_10380,N_11829);
nor U12318 (N_12318,N_10224,N_10621);
and U12319 (N_12319,N_10180,N_11661);
xor U12320 (N_12320,N_10293,N_10985);
nand U12321 (N_12321,N_11001,N_11377);
or U12322 (N_12322,N_11951,N_11985);
xnor U12323 (N_12323,N_10633,N_10941);
or U12324 (N_12324,N_10431,N_10117);
nand U12325 (N_12325,N_11926,N_11629);
nor U12326 (N_12326,N_11382,N_10256);
and U12327 (N_12327,N_10635,N_11224);
or U12328 (N_12328,N_11640,N_10648);
and U12329 (N_12329,N_11718,N_10500);
nor U12330 (N_12330,N_11898,N_11594);
nor U12331 (N_12331,N_11173,N_11274);
nor U12332 (N_12332,N_10005,N_11164);
xor U12333 (N_12333,N_10662,N_11228);
and U12334 (N_12334,N_10818,N_10728);
nand U12335 (N_12335,N_11966,N_11636);
or U12336 (N_12336,N_10330,N_11535);
xor U12337 (N_12337,N_10093,N_10024);
xnor U12338 (N_12338,N_11501,N_11309);
xor U12339 (N_12339,N_11268,N_11239);
nand U12340 (N_12340,N_10430,N_11065);
or U12341 (N_12341,N_10930,N_11199);
nor U12342 (N_12342,N_10373,N_10084);
nor U12343 (N_12343,N_10694,N_10964);
and U12344 (N_12344,N_10589,N_10533);
nor U12345 (N_12345,N_11632,N_11344);
and U12346 (N_12346,N_10695,N_10973);
xor U12347 (N_12347,N_10410,N_10674);
nor U12348 (N_12348,N_10762,N_11352);
xor U12349 (N_12349,N_10592,N_11248);
nand U12350 (N_12350,N_11560,N_11043);
nand U12351 (N_12351,N_10336,N_10260);
nor U12352 (N_12352,N_10036,N_10712);
and U12353 (N_12353,N_10066,N_10126);
and U12354 (N_12354,N_11429,N_11529);
and U12355 (N_12355,N_10122,N_10669);
or U12356 (N_12356,N_11570,N_10258);
or U12357 (N_12357,N_10538,N_10055);
nor U12358 (N_12358,N_10609,N_10312);
xnor U12359 (N_12359,N_10346,N_10707);
nor U12360 (N_12360,N_11899,N_10148);
nor U12361 (N_12361,N_10200,N_11704);
nand U12362 (N_12362,N_11073,N_11839);
nor U12363 (N_12363,N_11796,N_11068);
nand U12364 (N_12364,N_10750,N_11941);
nand U12365 (N_12365,N_11656,N_11369);
nand U12366 (N_12366,N_11390,N_10233);
or U12367 (N_12367,N_10344,N_10483);
nor U12368 (N_12368,N_11517,N_11034);
nand U12369 (N_12369,N_10003,N_11678);
or U12370 (N_12370,N_11893,N_10569);
and U12371 (N_12371,N_11296,N_10640);
or U12372 (N_12372,N_10094,N_10447);
or U12373 (N_12373,N_11184,N_10257);
nor U12374 (N_12374,N_10685,N_11115);
and U12375 (N_12375,N_10852,N_11264);
or U12376 (N_12376,N_10984,N_10368);
nor U12377 (N_12377,N_11714,N_11091);
and U12378 (N_12378,N_11822,N_10584);
and U12379 (N_12379,N_11353,N_11387);
or U12380 (N_12380,N_10765,N_10044);
or U12381 (N_12381,N_10657,N_10378);
or U12382 (N_12382,N_11087,N_10748);
nand U12383 (N_12383,N_11513,N_11634);
and U12384 (N_12384,N_11781,N_11481);
nor U12385 (N_12385,N_10745,N_11271);
and U12386 (N_12386,N_10614,N_10053);
nor U12387 (N_12387,N_10758,N_10220);
xor U12388 (N_12388,N_11525,N_10878);
and U12389 (N_12389,N_11448,N_11922);
or U12390 (N_12390,N_10666,N_11784);
or U12391 (N_12391,N_10890,N_11026);
xnor U12392 (N_12392,N_11869,N_10234);
nand U12393 (N_12393,N_10980,N_11003);
nand U12394 (N_12394,N_11005,N_11771);
and U12395 (N_12395,N_11085,N_10406);
nor U12396 (N_12396,N_10626,N_11145);
or U12397 (N_12397,N_11044,N_10511);
or U12398 (N_12398,N_10348,N_10379);
nor U12399 (N_12399,N_10485,N_11846);
and U12400 (N_12400,N_11598,N_11891);
xnor U12401 (N_12401,N_10098,N_10418);
nor U12402 (N_12402,N_11234,N_10704);
nand U12403 (N_12403,N_10420,N_11902);
nor U12404 (N_12404,N_11595,N_10502);
nand U12405 (N_12405,N_11953,N_10042);
xnor U12406 (N_12406,N_10667,N_11019);
and U12407 (N_12407,N_11593,N_10337);
or U12408 (N_12408,N_11606,N_10828);
or U12409 (N_12409,N_10428,N_10389);
or U12410 (N_12410,N_10178,N_11780);
xor U12411 (N_12411,N_10286,N_11756);
and U12412 (N_12412,N_10475,N_10903);
xnor U12413 (N_12413,N_11255,N_11371);
nor U12414 (N_12414,N_11282,N_10332);
nand U12415 (N_12415,N_11102,N_10302);
and U12416 (N_12416,N_10460,N_11126);
or U12417 (N_12417,N_10729,N_11028);
or U12418 (N_12418,N_11453,N_10118);
xor U12419 (N_12419,N_11388,N_11827);
and U12420 (N_12420,N_10237,N_11404);
and U12421 (N_12421,N_10199,N_11566);
nand U12422 (N_12422,N_10844,N_11023);
or U12423 (N_12423,N_11803,N_11219);
xnor U12424 (N_12424,N_11548,N_10169);
and U12425 (N_12425,N_10407,N_11779);
nand U12426 (N_12426,N_11265,N_10906);
xor U12427 (N_12427,N_11974,N_11664);
nor U12428 (N_12428,N_10947,N_10806);
xor U12429 (N_12429,N_11357,N_10853);
xnor U12430 (N_12430,N_11622,N_10279);
nor U12431 (N_12431,N_11276,N_11181);
nand U12432 (N_12432,N_10845,N_11495);
nand U12433 (N_12433,N_10767,N_11074);
xnor U12434 (N_12434,N_10059,N_11540);
nand U12435 (N_12435,N_11918,N_11764);
xnor U12436 (N_12436,N_11834,N_10061);
xor U12437 (N_12437,N_10943,N_11493);
and U12438 (N_12438,N_10398,N_10040);
or U12439 (N_12439,N_10540,N_10867);
or U12440 (N_12440,N_11503,N_10700);
xnor U12441 (N_12441,N_11858,N_10350);
nand U12442 (N_12442,N_11659,N_10688);
nor U12443 (N_12443,N_10563,N_10496);
and U12444 (N_12444,N_11361,N_11008);
xor U12445 (N_12445,N_10358,N_11708);
nor U12446 (N_12446,N_10776,N_11479);
xnor U12447 (N_12447,N_11195,N_10796);
or U12448 (N_12448,N_10161,N_10318);
or U12449 (N_12449,N_10507,N_11936);
xor U12450 (N_12450,N_10550,N_10746);
xnor U12451 (N_12451,N_11750,N_10607);
xor U12452 (N_12452,N_11364,N_11703);
and U12453 (N_12453,N_11737,N_11840);
xnor U12454 (N_12454,N_11767,N_10381);
and U12455 (N_12455,N_11677,N_11516);
or U12456 (N_12456,N_11683,N_10513);
nor U12457 (N_12457,N_10937,N_11558);
nor U12458 (N_12458,N_11332,N_10218);
or U12459 (N_12459,N_10603,N_11723);
and U12460 (N_12460,N_11877,N_10009);
and U12461 (N_12461,N_10759,N_11169);
nand U12462 (N_12462,N_11757,N_10840);
or U12463 (N_12463,N_11244,N_10225);
xor U12464 (N_12464,N_10803,N_11079);
nor U12465 (N_12465,N_10268,N_11116);
and U12466 (N_12466,N_10795,N_10214);
nor U12467 (N_12467,N_10158,N_11334);
xnor U12468 (N_12468,N_11539,N_11870);
and U12469 (N_12469,N_10331,N_10106);
nand U12470 (N_12470,N_10539,N_10872);
nor U12471 (N_12471,N_11528,N_10725);
and U12472 (N_12472,N_11337,N_11325);
xnor U12473 (N_12473,N_10230,N_11497);
nor U12474 (N_12474,N_11290,N_11986);
nand U12475 (N_12475,N_10129,N_11363);
nor U12476 (N_12476,N_11163,N_10356);
nor U12477 (N_12477,N_10278,N_10170);
nand U12478 (N_12478,N_11589,N_11782);
nand U12479 (N_12479,N_10697,N_11837);
nand U12480 (N_12480,N_10936,N_10041);
nand U12481 (N_12481,N_10273,N_10548);
nor U12482 (N_12482,N_10249,N_11619);
nor U12483 (N_12483,N_11188,N_10466);
nand U12484 (N_12484,N_10942,N_11083);
and U12485 (N_12485,N_11576,N_11395);
or U12486 (N_12486,N_10325,N_10835);
or U12487 (N_12487,N_11924,N_11867);
nand U12488 (N_12488,N_10742,N_10863);
xnor U12489 (N_12489,N_10021,N_11069);
or U12490 (N_12490,N_10831,N_11452);
nor U12491 (N_12491,N_11284,N_11258);
xnor U12492 (N_12492,N_10517,N_11086);
and U12493 (N_12493,N_10213,N_11120);
nor U12494 (N_12494,N_11439,N_11491);
and U12495 (N_12495,N_10967,N_10197);
xnor U12496 (N_12496,N_10738,N_10459);
and U12497 (N_12497,N_10322,N_10821);
nand U12498 (N_12498,N_11458,N_10645);
nand U12499 (N_12499,N_10441,N_10384);
nand U12500 (N_12500,N_11801,N_10730);
nand U12501 (N_12501,N_10899,N_11734);
nor U12502 (N_12502,N_10185,N_10668);
xnor U12503 (N_12503,N_10892,N_11129);
or U12504 (N_12504,N_10266,N_10467);
nor U12505 (N_12505,N_11774,N_11821);
or U12506 (N_12506,N_11293,N_10034);
xnor U12507 (N_12507,N_11722,N_11817);
xor U12508 (N_12508,N_11238,N_10747);
and U12509 (N_12509,N_10288,N_10068);
or U12510 (N_12510,N_11331,N_11406);
and U12511 (N_12511,N_11689,N_11650);
nor U12512 (N_12512,N_11934,N_11505);
or U12513 (N_12513,N_11915,N_11489);
and U12514 (N_12514,N_10210,N_10409);
nor U12515 (N_12515,N_10642,N_10731);
or U12516 (N_12516,N_10115,N_11651);
xor U12517 (N_12517,N_11118,N_10202);
and U12518 (N_12518,N_10812,N_11912);
or U12519 (N_12519,N_11289,N_10201);
or U12520 (N_12520,N_11498,N_11873);
and U12521 (N_12521,N_11411,N_11693);
nand U12522 (N_12522,N_11484,N_10622);
and U12523 (N_12523,N_11373,N_10777);
xor U12524 (N_12524,N_10424,N_10989);
and U12525 (N_12525,N_10393,N_11084);
nand U12526 (N_12526,N_10168,N_10195);
nand U12527 (N_12527,N_11679,N_11988);
or U12528 (N_12528,N_10808,N_10814);
nor U12529 (N_12529,N_10134,N_11054);
xnor U12530 (N_12530,N_10680,N_11648);
nand U12531 (N_12531,N_11366,N_11943);
xnor U12532 (N_12532,N_10871,N_10524);
and U12533 (N_12533,N_11041,N_10952);
or U12534 (N_12534,N_10100,N_11561);
xor U12535 (N_12535,N_10574,N_10570);
or U12536 (N_12536,N_11270,N_11156);
and U12537 (N_12537,N_11602,N_10081);
nor U12538 (N_12538,N_10054,N_11014);
xor U12539 (N_12539,N_11146,N_10085);
xor U12540 (N_12540,N_11970,N_11301);
and U12541 (N_12541,N_11667,N_11349);
nand U12542 (N_12542,N_10140,N_10516);
nor U12543 (N_12543,N_11161,N_10785);
or U12544 (N_12544,N_11613,N_11744);
or U12545 (N_12545,N_11160,N_11554);
nand U12546 (N_12546,N_11991,N_11832);
and U12547 (N_12547,N_11646,N_10276);
nand U12548 (N_12548,N_11550,N_11864);
or U12549 (N_12549,N_10992,N_10797);
or U12550 (N_12550,N_10670,N_10164);
nand U12551 (N_12551,N_11281,N_10950);
and U12552 (N_12552,N_10227,N_11338);
nand U12553 (N_12553,N_11013,N_10580);
or U12554 (N_12554,N_10549,N_10934);
nor U12555 (N_12555,N_10751,N_10636);
nor U12556 (N_12556,N_11165,N_10875);
nand U12557 (N_12557,N_11257,N_10347);
nand U12558 (N_12558,N_10727,N_10615);
and U12559 (N_12559,N_10047,N_10456);
xnor U12560 (N_12560,N_11556,N_10655);
and U12561 (N_12561,N_11879,N_11380);
nand U12562 (N_12562,N_10590,N_11536);
nor U12563 (N_12563,N_10766,N_11823);
nand U12564 (N_12564,N_10503,N_10283);
nand U12565 (N_12565,N_11027,N_10102);
nand U12566 (N_12566,N_11790,N_11927);
nor U12567 (N_12567,N_10349,N_10287);
and U12568 (N_12568,N_11712,N_11880);
nand U12569 (N_12569,N_11792,N_11946);
and U12570 (N_12570,N_10252,N_10246);
xnor U12571 (N_12571,N_11467,N_11887);
xnor U12572 (N_12572,N_11335,N_11826);
or U12573 (N_12573,N_11716,N_10425);
nor U12574 (N_12574,N_10819,N_10017);
nor U12575 (N_12575,N_10940,N_10868);
xnor U12576 (N_12576,N_10702,N_11403);
xnor U12577 (N_12577,N_10304,N_11166);
nand U12578 (N_12578,N_11851,N_10910);
nand U12579 (N_12579,N_11775,N_11724);
nand U12580 (N_12580,N_10757,N_11762);
xnor U12581 (N_12581,N_11720,N_11987);
xnor U12582 (N_12582,N_10778,N_10071);
or U12583 (N_12583,N_10974,N_11546);
xor U12584 (N_12584,N_11259,N_11755);
xnor U12585 (N_12585,N_11341,N_11214);
nand U12586 (N_12586,N_10711,N_11012);
or U12587 (N_12587,N_10353,N_11596);
and U12588 (N_12588,N_10755,N_11134);
or U12589 (N_12589,N_11531,N_11348);
and U12590 (N_12590,N_10723,N_11603);
nor U12591 (N_12591,N_11261,N_10999);
and U12592 (N_12592,N_11435,N_10627);
and U12593 (N_12593,N_10644,N_10555);
nor U12594 (N_12594,N_10255,N_10110);
xor U12595 (N_12595,N_10062,N_10097);
nand U12596 (N_12596,N_10269,N_10679);
nor U12597 (N_12597,N_10376,N_10961);
xor U12598 (N_12598,N_11105,N_10956);
and U12599 (N_12599,N_11092,N_10171);
and U12600 (N_12600,N_11728,N_11196);
nor U12601 (N_12601,N_11957,N_10032);
nor U12602 (N_12602,N_11627,N_11892);
or U12603 (N_12603,N_10072,N_11307);
nand U12604 (N_12604,N_11733,N_11113);
and U12605 (N_12605,N_10008,N_11128);
xnor U12606 (N_12606,N_11969,N_10578);
nor U12607 (N_12607,N_10955,N_11243);
nand U12608 (N_12608,N_10415,N_11649);
nand U12609 (N_12609,N_11647,N_11496);
nand U12610 (N_12610,N_10687,N_11350);
or U12611 (N_12611,N_10660,N_11127);
xor U12612 (N_12612,N_10064,N_10825);
nor U12613 (N_12613,N_10522,N_10681);
nor U12614 (N_12614,N_11398,N_11267);
nand U12615 (N_12615,N_11814,N_10505);
or U12616 (N_12616,N_11547,N_10604);
xor U12617 (N_12617,N_11736,N_10394);
nor U12618 (N_12618,N_10960,N_11021);
xnor U12619 (N_12619,N_11591,N_10849);
or U12620 (N_12620,N_10355,N_11222);
nor U12621 (N_12621,N_10497,N_11694);
and U12622 (N_12622,N_10079,N_10519);
nand U12623 (N_12623,N_11600,N_10908);
or U12624 (N_12624,N_10413,N_10998);
and U12625 (N_12625,N_10896,N_11810);
or U12626 (N_12626,N_10817,N_10794);
nor U12627 (N_12627,N_11979,N_10137);
nor U12628 (N_12628,N_11982,N_11806);
nor U12629 (N_12629,N_10916,N_11418);
or U12630 (N_12630,N_11474,N_11233);
or U12631 (N_12631,N_11393,N_11563);
nand U12632 (N_12632,N_11241,N_11172);
nand U12633 (N_12633,N_11958,N_10628);
and U12634 (N_12634,N_11776,N_11414);
xnor U12635 (N_12635,N_11706,N_10371);
xnor U12636 (N_12636,N_11149,N_11286);
or U12637 (N_12637,N_11174,N_11580);
xor U12638 (N_12638,N_10395,N_11451);
nor U12639 (N_12639,N_10359,N_11573);
and U12640 (N_12640,N_11972,N_10599);
nor U12641 (N_12641,N_11808,N_11711);
and U12642 (N_12642,N_11427,N_11399);
xor U12643 (N_12643,N_11141,N_11908);
or U12644 (N_12644,N_10402,N_10010);
nor U12645 (N_12645,N_11180,N_11504);
nand U12646 (N_12646,N_10391,N_10693);
and U12647 (N_12647,N_10423,N_10506);
and U12648 (N_12648,N_10661,N_11961);
xnor U12649 (N_12649,N_10209,N_10521);
nand U12650 (N_12650,N_11150,N_10316);
xnor U12651 (N_12651,N_11464,N_10101);
and U12652 (N_12652,N_10223,N_10272);
or U12653 (N_12653,N_11082,N_11510);
nor U12654 (N_12654,N_10775,N_10736);
nor U12655 (N_12655,N_11721,N_10165);
or U12656 (N_12656,N_11511,N_10188);
nor U12657 (N_12657,N_11310,N_11185);
or U12658 (N_12658,N_11144,N_10211);
xnor U12659 (N_12659,N_10957,N_11066);
xnor U12660 (N_12660,N_11709,N_11280);
and U12661 (N_12661,N_10976,N_10683);
nor U12662 (N_12662,N_11611,N_10103);
nand U12663 (N_12663,N_11612,N_10696);
or U12664 (N_12664,N_11168,N_10854);
nand U12665 (N_12665,N_10678,N_10734);
or U12666 (N_12666,N_11641,N_10235);
and U12667 (N_12667,N_11318,N_11308);
nor U12668 (N_12668,N_10753,N_10388);
nand U12669 (N_12669,N_11592,N_11299);
xor U12670 (N_12670,N_11186,N_10841);
nor U12671 (N_12671,N_10605,N_10877);
or U12672 (N_12672,N_11345,N_11783);
nor U12673 (N_12673,N_10873,N_11971);
or U12674 (N_12674,N_10046,N_11356);
nor U12675 (N_12675,N_11378,N_10913);
or U12676 (N_12676,N_10004,N_10862);
nor U12677 (N_12677,N_11078,N_10987);
and U12678 (N_12678,N_10573,N_11466);
nor U12679 (N_12679,N_10582,N_10445);
nand U12680 (N_12680,N_11655,N_11232);
nor U12681 (N_12681,N_11230,N_11522);
xor U12682 (N_12682,N_11216,N_10342);
nand U12683 (N_12683,N_10007,N_11314);
nor U12684 (N_12684,N_10254,N_10932);
or U12685 (N_12685,N_11151,N_10907);
xor U12686 (N_12686,N_10557,N_11795);
nand U12687 (N_12687,N_10836,N_11897);
nor U12688 (N_12688,N_10443,N_11811);
or U12689 (N_12689,N_11696,N_11553);
and U12690 (N_12690,N_11475,N_10510);
or U12691 (N_12691,N_11542,N_10610);
nor U12692 (N_12692,N_11447,N_11048);
nand U12693 (N_12693,N_11555,N_10895);
nor U12694 (N_12694,N_11541,N_11229);
nand U12695 (N_12695,N_11204,N_11190);
or U12696 (N_12696,N_10813,N_11919);
xor U12697 (N_12697,N_10476,N_11425);
nand U12698 (N_12698,N_10619,N_10690);
nand U12699 (N_12699,N_11772,N_10676);
or U12700 (N_12700,N_10837,N_10571);
or U12701 (N_12701,N_10612,N_11976);
nand U12702 (N_12702,N_10212,N_11833);
xor U12703 (N_12703,N_10659,N_11108);
and U12704 (N_12704,N_10724,N_11874);
xor U12705 (N_12705,N_10451,N_11564);
nand U12706 (N_12706,N_11059,N_11688);
nand U12707 (N_12707,N_10970,N_11742);
nor U12708 (N_12708,N_11890,N_10397);
nand U12709 (N_12709,N_11231,N_10902);
or U12710 (N_12710,N_10923,N_10526);
nand U12711 (N_12711,N_10076,N_10109);
and U12712 (N_12712,N_10241,N_10438);
nor U12713 (N_12713,N_11786,N_10280);
xnor U12714 (N_12714,N_10345,N_10839);
nor U12715 (N_12715,N_11631,N_10515);
nand U12716 (N_12716,N_11140,N_10784);
nand U12717 (N_12717,N_11571,N_11935);
xnor U12718 (N_12718,N_11658,N_11643);
or U12719 (N_12719,N_10411,N_11705);
nor U12720 (N_12720,N_10601,N_10444);
and U12721 (N_12721,N_10931,N_11978);
xnor U12722 (N_12722,N_10546,N_11841);
xnor U12723 (N_12723,N_10051,N_11665);
nand U12724 (N_12724,N_11624,N_10357);
and U12725 (N_12725,N_10664,N_10150);
or U12726 (N_12726,N_10317,N_10924);
nor U12727 (N_12727,N_10453,N_11201);
and U12728 (N_12728,N_11917,N_11327);
and U12729 (N_12729,N_10463,N_10013);
nand U12730 (N_12730,N_11323,N_10073);
or U12731 (N_12731,N_11432,N_10804);
nand U12732 (N_12732,N_10173,N_11292);
nand U12733 (N_12733,N_11423,N_11537);
nor U12734 (N_12734,N_10508,N_10481);
and U12735 (N_12735,N_10876,N_10422);
xor U12736 (N_12736,N_10887,N_11143);
nand U12737 (N_12737,N_10436,N_11527);
nor U12738 (N_12738,N_11610,N_10824);
nor U12739 (N_12739,N_11354,N_11098);
nand U12740 (N_12740,N_11749,N_11608);
or U12741 (N_12741,N_10793,N_10092);
xnor U12742 (N_12742,N_10030,N_11681);
nand U12743 (N_12743,N_10544,N_10339);
xor U12744 (N_12744,N_11888,N_10275);
nor U12745 (N_12745,N_11444,N_11463);
nor U12746 (N_12746,N_11375,N_10219);
and U12747 (N_12747,N_10501,N_10815);
and U12748 (N_12748,N_11956,N_11872);
nand U12749 (N_12749,N_10530,N_11903);
or U12750 (N_12750,N_11950,N_10884);
xnor U12751 (N_12751,N_10446,N_11686);
or U12752 (N_12752,N_10904,N_11424);
xnor U12753 (N_12753,N_11526,N_10367);
and U12754 (N_12754,N_10938,N_11901);
nor U12755 (N_12755,N_11252,N_11746);
or U12756 (N_12756,N_11062,N_10744);
xor U12757 (N_12757,N_10334,N_10595);
nor U12758 (N_12758,N_11124,N_11587);
nor U12759 (N_12759,N_10179,N_10594);
and U12760 (N_12760,N_10739,N_10567);
or U12761 (N_12761,N_10716,N_11152);
nand U12762 (N_12762,N_10829,N_11582);
xnor U12763 (N_12763,N_10027,N_10888);
and U12764 (N_12764,N_10665,N_10163);
nand U12765 (N_12765,N_11502,N_10606);
or U12766 (N_12766,N_10028,N_10292);
xor U12767 (N_12767,N_10996,N_11816);
xor U12768 (N_12768,N_10838,N_11189);
xor U12769 (N_12769,N_11193,N_11039);
or U12770 (N_12770,N_10306,N_10682);
and U12771 (N_12771,N_10886,N_10858);
xnor U12772 (N_12772,N_11294,N_10414);
nand U12773 (N_12773,N_10525,N_10184);
or U12774 (N_12774,N_11653,N_10328);
nand U12775 (N_12775,N_10090,N_10675);
nor U12776 (N_12776,N_10623,N_10740);
xor U12777 (N_12777,N_11198,N_10454);
nand U12778 (N_12778,N_11508,N_10327);
nand U12779 (N_12779,N_11402,N_11136);
xor U12780 (N_12780,N_10901,N_11701);
or U12781 (N_12781,N_11657,N_10289);
and U12782 (N_12782,N_10591,N_10127);
nand U12783 (N_12783,N_10568,N_10780);
xor U12784 (N_12784,N_10035,N_10602);
nand U12785 (N_12785,N_11538,N_10114);
xnor U12786 (N_12786,N_11569,N_10417);
nor U12787 (N_12787,N_11515,N_10634);
xor U12788 (N_12788,N_10847,N_10588);
or U12789 (N_12789,N_11110,N_11815);
nand U12790 (N_12790,N_11042,N_11691);
xnor U12791 (N_12791,N_10926,N_11507);
or U12792 (N_12792,N_11713,N_11155);
or U12793 (N_12793,N_10721,N_11928);
nand U12794 (N_12794,N_10880,N_11278);
and U12795 (N_12795,N_11295,N_10216);
and U12796 (N_12796,N_10651,N_10494);
and U12797 (N_12797,N_11967,N_10782);
or U12798 (N_12798,N_10285,N_10512);
nor U12799 (N_12799,N_10889,N_10671);
and U12800 (N_12800,N_11861,N_11312);
nand U12801 (N_12801,N_10948,N_11015);
or U12802 (N_12802,N_11942,N_10247);
nand U12803 (N_12803,N_10830,N_11883);
or U12804 (N_12804,N_11939,N_11905);
or U12805 (N_12805,N_11431,N_10600);
nand U12806 (N_12806,N_11142,N_11809);
nand U12807 (N_12807,N_11532,N_11533);
nand U12808 (N_12808,N_11962,N_11158);
or U12809 (N_12809,N_11437,N_10581);
nor U12810 (N_12810,N_10099,N_10798);
or U12811 (N_12811,N_10075,N_10617);
xnor U12812 (N_12812,N_11326,N_11838);
xor U12813 (N_12813,N_11692,N_11355);
nand U12814 (N_12814,N_10646,N_11031);
nand U12815 (N_12815,N_11480,N_11521);
and U12816 (N_12816,N_10988,N_11642);
or U12817 (N_12817,N_10472,N_10363);
or U12818 (N_12818,N_10192,N_10113);
nor U12819 (N_12819,N_11998,N_11385);
xor U12820 (N_12820,N_11298,N_10095);
or U12821 (N_12821,N_11409,N_10543);
nor U12822 (N_12822,N_10920,N_11973);
or U12823 (N_12823,N_11994,N_11470);
xnor U12824 (N_12824,N_11863,N_11121);
nor U12825 (N_12825,N_10966,N_11000);
or U12826 (N_12826,N_11828,N_10834);
and U12827 (N_12827,N_10437,N_10487);
and U12828 (N_12828,N_11616,N_11139);
or U12829 (N_12829,N_11590,N_11384);
or U12830 (N_12830,N_10577,N_11347);
nand U12831 (N_12831,N_11154,N_11046);
or U12832 (N_12832,N_11938,N_10364);
or U12833 (N_12833,N_10997,N_11218);
and U12834 (N_12834,N_11940,N_11071);
or U12835 (N_12835,N_10489,N_11340);
and U12836 (N_12836,N_11131,N_10737);
xor U12837 (N_12837,N_11413,N_11170);
nor U12838 (N_12838,N_10442,N_11739);
and U12839 (N_12839,N_11223,N_10647);
xor U12840 (N_12840,N_10722,N_10045);
and U12841 (N_12841,N_10458,N_11845);
nand U12842 (N_12842,N_10271,N_11842);
xor U12843 (N_12843,N_11376,N_11187);
or U12844 (N_12844,N_10231,N_11400);
xnor U12845 (N_12845,N_10715,N_11210);
or U12846 (N_12846,N_11138,N_10965);
or U12847 (N_12847,N_10741,N_10482);
nor U12848 (N_12848,N_10037,N_11461);
or U12849 (N_12849,N_10319,N_10805);
nor U12850 (N_12850,N_11343,N_11717);
and U12851 (N_12851,N_10239,N_10387);
nand U12852 (N_12852,N_11052,N_10366);
xnor U12853 (N_12853,N_11212,N_11960);
and U12854 (N_12854,N_10138,N_11578);
and U12855 (N_12855,N_10486,N_11235);
xor U12856 (N_12856,N_10783,N_11311);
nand U12857 (N_12857,N_10850,N_10296);
nor U12858 (N_12858,N_10182,N_11226);
nand U12859 (N_12859,N_10311,N_11687);
xnor U12860 (N_12860,N_11831,N_11114);
nand U12861 (N_12861,N_10250,N_11752);
nand U12862 (N_12862,N_10232,N_10049);
and U12863 (N_12863,N_11975,N_11848);
and U12864 (N_12864,N_11269,N_10556);
nor U12865 (N_12865,N_10786,N_10710);
and U12866 (N_12866,N_11175,N_11440);
xor U12867 (N_12867,N_10001,N_10014);
and U12868 (N_12868,N_10883,N_10206);
and U12869 (N_12869,N_11103,N_11499);
nand U12870 (N_12870,N_11740,N_11297);
and U12871 (N_12871,N_11047,N_11996);
xnor U12872 (N_12872,N_11303,N_10918);
and U12873 (N_12873,N_10251,N_10982);
and U12874 (N_12874,N_11770,N_11433);
nor U12875 (N_12875,N_11700,N_11117);
or U12876 (N_12876,N_11680,N_10760);
nor U12877 (N_12877,N_10979,N_11673);
or U12878 (N_12878,N_10253,N_11800);
and U12879 (N_12879,N_10048,N_11819);
nand U12880 (N_12880,N_11060,N_11807);
and U12881 (N_12881,N_11288,N_10823);
xor U12882 (N_12882,N_10261,N_11565);
nand U12883 (N_12883,N_11263,N_11760);
xor U12884 (N_12884,N_10448,N_10462);
or U12885 (N_12885,N_11682,N_11157);
and U12886 (N_12886,N_11766,N_11524);
and U12887 (N_12887,N_10374,N_10157);
xnor U12888 (N_12888,N_11638,N_11588);
or U12889 (N_12889,N_10124,N_10281);
nor U12890 (N_12890,N_10763,N_10386);
xnor U12891 (N_12891,N_10078,N_11123);
nand U12892 (N_12892,N_11405,N_11765);
nand U12893 (N_12893,N_11885,N_11051);
nor U12894 (N_12894,N_10520,N_10313);
nand U12895 (N_12895,N_10262,N_11574);
nand U12896 (N_12896,N_10972,N_10183);
nand U12897 (N_12897,N_11088,N_11132);
nor U12898 (N_12898,N_11543,N_10186);
nor U12899 (N_12899,N_10329,N_11916);
or U12900 (N_12900,N_11699,N_10649);
or U12901 (N_12901,N_10063,N_10435);
nor U12902 (N_12902,N_11952,N_10240);
and U12903 (N_12903,N_10658,N_10147);
and U12904 (N_12904,N_10576,N_10082);
and U12905 (N_12905,N_11847,N_11441);
and U12906 (N_12906,N_10156,N_10267);
or U12907 (N_12907,N_11122,N_11266);
and U12908 (N_12908,N_10531,N_10362);
and U12909 (N_12909,N_10043,N_10058);
xor U12910 (N_12910,N_10752,N_10385);
or U12911 (N_12911,N_10761,N_11368);
nand U12912 (N_12912,N_11690,N_11568);
nand U12913 (N_12913,N_10663,N_11153);
and U12914 (N_12914,N_10305,N_10929);
xnor U12915 (N_12915,N_11397,N_10882);
xnor U12916 (N_12916,N_11030,N_11707);
nor U12917 (N_12917,N_11617,N_11530);
xor U12918 (N_12918,N_11944,N_10652);
xnor U12919 (N_12919,N_10691,N_11137);
and U12920 (N_12920,N_11097,N_11895);
or U12921 (N_12921,N_11056,N_10855);
nand U12922 (N_12922,N_10015,N_10229);
or U12923 (N_12923,N_11336,N_11628);
and U12924 (N_12924,N_11725,N_11107);
and U12925 (N_12925,N_11732,N_10962);
nand U12926 (N_12926,N_10208,N_11989);
nand U12927 (N_12927,N_10488,N_11544);
and U12928 (N_12928,N_10172,N_11859);
nand U12929 (N_12929,N_11534,N_11407);
xnor U12930 (N_12930,N_10086,N_11360);
or U12931 (N_12931,N_10484,N_11018);
and U12932 (N_12932,N_11024,N_10145);
nor U12933 (N_12933,N_10057,N_11415);
xor U12934 (N_12934,N_11428,N_10108);
nand U12935 (N_12935,N_10002,N_10416);
and U12936 (N_12936,N_10925,N_11769);
or U12937 (N_12937,N_11100,N_11089);
nor U12938 (N_12938,N_10421,N_11473);
nor U12939 (N_12939,N_10726,N_11179);
or U12940 (N_12940,N_10333,N_11886);
nor U12941 (N_12941,N_10282,N_10949);
nor U12942 (N_12942,N_10586,N_10816);
and U12943 (N_12943,N_10174,N_11813);
xnor U12944 (N_12944,N_10369,N_11520);
xnor U12945 (N_12945,N_10151,N_10789);
nor U12946 (N_12946,N_11741,N_11662);
nand U12947 (N_12947,N_11597,N_11010);
nand U12948 (N_12948,N_10427,N_10713);
nor U12949 (N_12949,N_10528,N_11727);
xnor U12950 (N_12950,N_10136,N_10983);
nor U12951 (N_12951,N_10620,N_11316);
xor U12952 (N_12952,N_11487,N_10971);
and U12953 (N_12953,N_10826,N_10470);
and U12954 (N_12954,N_10300,N_10190);
xor U12955 (N_12955,N_10242,N_10756);
nand U12956 (N_12956,N_10221,N_10743);
or U12957 (N_12957,N_11200,N_10468);
nand U12958 (N_12958,N_10074,N_10810);
or U12959 (N_12959,N_10144,N_11273);
nor U12960 (N_12960,N_11900,N_11383);
and U12961 (N_12961,N_10692,N_11242);
and U12962 (N_12962,N_10677,N_10944);
nor U12963 (N_12963,N_10107,N_11148);
and U12964 (N_12964,N_10298,N_10396);
xnor U12965 (N_12965,N_11844,N_10052);
or U12966 (N_12966,N_10566,N_10518);
and U12967 (N_12967,N_10123,N_11351);
xnor U12968 (N_12968,N_11599,N_10779);
xnor U12969 (N_12969,N_10922,N_11050);
or U12970 (N_12970,N_11033,N_10433);
and U12971 (N_12971,N_11317,N_11076);
or U12972 (N_12972,N_10848,N_11182);
nand U12973 (N_12973,N_10951,N_11038);
xnor U12974 (N_12974,N_10631,N_11213);
xor U12975 (N_12975,N_10717,N_11183);
and U12976 (N_12976,N_11745,N_10799);
and U12977 (N_12977,N_10774,N_11135);
nor U12978 (N_12978,N_10709,N_10295);
or U12979 (N_12979,N_10832,N_10534);
and U12980 (N_12980,N_11992,N_11055);
or U12981 (N_12981,N_10914,N_11036);
nand U12982 (N_12982,N_11454,N_11930);
nor U12983 (N_12983,N_10050,N_10499);
and U12984 (N_12984,N_10067,N_10143);
or U12985 (N_12985,N_11220,N_10596);
xor U12986 (N_12986,N_11584,N_11797);
nand U12987 (N_12987,N_10033,N_10865);
and U12988 (N_12988,N_11058,N_11006);
xor U12989 (N_12989,N_11486,N_11626);
or U12990 (N_12990,N_10196,N_10478);
xnor U12991 (N_12991,N_11029,N_11075);
nand U12992 (N_12992,N_10263,N_11370);
nor U12993 (N_12993,N_11671,N_11906);
xor U12994 (N_12994,N_11751,N_11211);
or U12995 (N_12995,N_10672,N_10788);
or U12996 (N_12996,N_11365,N_10981);
nor U12997 (N_12997,N_11162,N_10801);
and U12998 (N_12998,N_10429,N_11206);
xnor U12999 (N_12999,N_11315,N_10579);
nand U13000 (N_13000,N_10824,N_10815);
nand U13001 (N_13001,N_11407,N_11158);
or U13002 (N_13002,N_10281,N_11237);
nand U13003 (N_13003,N_10861,N_11654);
or U13004 (N_13004,N_10081,N_11717);
xor U13005 (N_13005,N_11418,N_11450);
or U13006 (N_13006,N_10785,N_10992);
xnor U13007 (N_13007,N_11159,N_11349);
and U13008 (N_13008,N_11226,N_11954);
or U13009 (N_13009,N_11001,N_11611);
and U13010 (N_13010,N_11862,N_10481);
and U13011 (N_13011,N_11215,N_11898);
or U13012 (N_13012,N_10619,N_10265);
and U13013 (N_13013,N_10996,N_10253);
nor U13014 (N_13014,N_10696,N_10249);
nand U13015 (N_13015,N_11482,N_10130);
or U13016 (N_13016,N_11267,N_10269);
nand U13017 (N_13017,N_11058,N_10416);
nor U13018 (N_13018,N_11105,N_11047);
nand U13019 (N_13019,N_10872,N_10441);
nand U13020 (N_13020,N_10983,N_11258);
nand U13021 (N_13021,N_10427,N_11332);
nor U13022 (N_13022,N_11819,N_11670);
and U13023 (N_13023,N_10205,N_11634);
and U13024 (N_13024,N_11881,N_10283);
or U13025 (N_13025,N_10683,N_10365);
and U13026 (N_13026,N_10746,N_11964);
and U13027 (N_13027,N_11155,N_10233);
xor U13028 (N_13028,N_11996,N_10779);
and U13029 (N_13029,N_11205,N_10459);
or U13030 (N_13030,N_10271,N_10846);
or U13031 (N_13031,N_10603,N_10626);
xor U13032 (N_13032,N_10175,N_10153);
and U13033 (N_13033,N_11707,N_10566);
and U13034 (N_13034,N_10728,N_11621);
xnor U13035 (N_13035,N_11349,N_10353);
nand U13036 (N_13036,N_10879,N_10062);
nand U13037 (N_13037,N_11575,N_10561);
or U13038 (N_13038,N_10456,N_10760);
or U13039 (N_13039,N_10977,N_10090);
or U13040 (N_13040,N_10845,N_11409);
nand U13041 (N_13041,N_10595,N_10866);
xor U13042 (N_13042,N_11341,N_11200);
nand U13043 (N_13043,N_10458,N_11194);
or U13044 (N_13044,N_11165,N_10672);
nand U13045 (N_13045,N_11651,N_10062);
nand U13046 (N_13046,N_11470,N_11627);
nor U13047 (N_13047,N_11034,N_11873);
xnor U13048 (N_13048,N_11750,N_11321);
xor U13049 (N_13049,N_11278,N_10104);
and U13050 (N_13050,N_11417,N_11733);
xnor U13051 (N_13051,N_11064,N_10875);
xor U13052 (N_13052,N_11897,N_11654);
xnor U13053 (N_13053,N_10167,N_10678);
nor U13054 (N_13054,N_11258,N_11434);
xnor U13055 (N_13055,N_11065,N_10432);
nor U13056 (N_13056,N_10143,N_10791);
and U13057 (N_13057,N_10657,N_10189);
and U13058 (N_13058,N_10372,N_10893);
and U13059 (N_13059,N_10330,N_11033);
nand U13060 (N_13060,N_10784,N_11029);
xor U13061 (N_13061,N_10549,N_11903);
xor U13062 (N_13062,N_10616,N_11458);
xor U13063 (N_13063,N_10673,N_10550);
or U13064 (N_13064,N_10872,N_11574);
nand U13065 (N_13065,N_11654,N_10914);
nand U13066 (N_13066,N_10508,N_10977);
and U13067 (N_13067,N_11490,N_11108);
or U13068 (N_13068,N_10038,N_11899);
nor U13069 (N_13069,N_10066,N_11695);
nor U13070 (N_13070,N_10719,N_11184);
nor U13071 (N_13071,N_10661,N_10474);
xnor U13072 (N_13072,N_11320,N_11257);
nand U13073 (N_13073,N_10737,N_10209);
and U13074 (N_13074,N_11931,N_11193);
or U13075 (N_13075,N_10267,N_11132);
or U13076 (N_13076,N_11703,N_10773);
and U13077 (N_13077,N_10781,N_10671);
xor U13078 (N_13078,N_11378,N_11664);
nor U13079 (N_13079,N_10004,N_10826);
xnor U13080 (N_13080,N_10405,N_11071);
nand U13081 (N_13081,N_11854,N_11952);
nand U13082 (N_13082,N_10826,N_11342);
nor U13083 (N_13083,N_10103,N_10535);
or U13084 (N_13084,N_11256,N_11021);
or U13085 (N_13085,N_11407,N_11523);
nand U13086 (N_13086,N_10407,N_11084);
and U13087 (N_13087,N_10169,N_10130);
or U13088 (N_13088,N_11003,N_11478);
nor U13089 (N_13089,N_11410,N_11403);
and U13090 (N_13090,N_11595,N_11059);
nor U13091 (N_13091,N_11367,N_11700);
nand U13092 (N_13092,N_11035,N_10289);
nor U13093 (N_13093,N_11788,N_11215);
nor U13094 (N_13094,N_11709,N_10463);
or U13095 (N_13095,N_11281,N_11249);
and U13096 (N_13096,N_10610,N_11035);
nand U13097 (N_13097,N_11436,N_11625);
or U13098 (N_13098,N_10067,N_11319);
xor U13099 (N_13099,N_10330,N_10491);
nor U13100 (N_13100,N_10437,N_10043);
nor U13101 (N_13101,N_11071,N_10670);
xnor U13102 (N_13102,N_10794,N_10294);
nor U13103 (N_13103,N_11549,N_11727);
or U13104 (N_13104,N_10868,N_11957);
nand U13105 (N_13105,N_11057,N_11740);
nor U13106 (N_13106,N_10407,N_10846);
xnor U13107 (N_13107,N_10543,N_10202);
nor U13108 (N_13108,N_10863,N_10867);
xor U13109 (N_13109,N_10051,N_10458);
and U13110 (N_13110,N_10551,N_10623);
or U13111 (N_13111,N_11536,N_11592);
xor U13112 (N_13112,N_11231,N_10178);
and U13113 (N_13113,N_11026,N_10679);
and U13114 (N_13114,N_11466,N_11925);
or U13115 (N_13115,N_11779,N_11300);
and U13116 (N_13116,N_10725,N_10740);
nand U13117 (N_13117,N_11082,N_10042);
and U13118 (N_13118,N_10875,N_10750);
nand U13119 (N_13119,N_11598,N_10559);
nand U13120 (N_13120,N_11841,N_11645);
and U13121 (N_13121,N_11163,N_10345);
and U13122 (N_13122,N_11614,N_10085);
nand U13123 (N_13123,N_11952,N_10090);
xnor U13124 (N_13124,N_11512,N_11502);
nand U13125 (N_13125,N_10586,N_10954);
and U13126 (N_13126,N_11143,N_11182);
xnor U13127 (N_13127,N_10845,N_10037);
xor U13128 (N_13128,N_10824,N_10736);
and U13129 (N_13129,N_10908,N_11313);
nor U13130 (N_13130,N_10772,N_11507);
nand U13131 (N_13131,N_11315,N_11486);
nand U13132 (N_13132,N_11038,N_11100);
nor U13133 (N_13133,N_10260,N_10490);
and U13134 (N_13134,N_10636,N_11128);
and U13135 (N_13135,N_10600,N_11170);
nor U13136 (N_13136,N_10708,N_10665);
xnor U13137 (N_13137,N_10737,N_11176);
nor U13138 (N_13138,N_10328,N_11253);
xnor U13139 (N_13139,N_11922,N_11262);
nor U13140 (N_13140,N_11047,N_11125);
nand U13141 (N_13141,N_10743,N_11823);
or U13142 (N_13142,N_11072,N_10708);
nor U13143 (N_13143,N_10837,N_10084);
xor U13144 (N_13144,N_11624,N_10696);
xor U13145 (N_13145,N_11703,N_10990);
or U13146 (N_13146,N_11491,N_11160);
xnor U13147 (N_13147,N_10702,N_11013);
or U13148 (N_13148,N_11289,N_10761);
or U13149 (N_13149,N_11281,N_10625);
nor U13150 (N_13150,N_11879,N_11458);
nand U13151 (N_13151,N_10624,N_11952);
nand U13152 (N_13152,N_11394,N_11465);
nor U13153 (N_13153,N_10754,N_10702);
or U13154 (N_13154,N_11426,N_10861);
nand U13155 (N_13155,N_11785,N_10975);
xnor U13156 (N_13156,N_10719,N_11490);
and U13157 (N_13157,N_10280,N_11785);
xor U13158 (N_13158,N_10981,N_10852);
nand U13159 (N_13159,N_11628,N_10071);
nor U13160 (N_13160,N_11081,N_10195);
xor U13161 (N_13161,N_10589,N_10893);
and U13162 (N_13162,N_10917,N_10411);
nor U13163 (N_13163,N_11334,N_11670);
nand U13164 (N_13164,N_11666,N_11949);
xor U13165 (N_13165,N_11858,N_11871);
nor U13166 (N_13166,N_10245,N_11828);
nand U13167 (N_13167,N_10199,N_10097);
nor U13168 (N_13168,N_11436,N_11756);
nor U13169 (N_13169,N_10657,N_11909);
and U13170 (N_13170,N_11967,N_11671);
nand U13171 (N_13171,N_11912,N_10463);
xor U13172 (N_13172,N_10786,N_11071);
nand U13173 (N_13173,N_10423,N_11995);
nor U13174 (N_13174,N_11142,N_11865);
nor U13175 (N_13175,N_10144,N_11516);
xor U13176 (N_13176,N_10529,N_10245);
nor U13177 (N_13177,N_11750,N_11600);
xor U13178 (N_13178,N_11916,N_10457);
and U13179 (N_13179,N_11556,N_11248);
and U13180 (N_13180,N_10270,N_11751);
and U13181 (N_13181,N_11816,N_10394);
nor U13182 (N_13182,N_10689,N_11791);
and U13183 (N_13183,N_11705,N_11094);
and U13184 (N_13184,N_11192,N_10123);
nor U13185 (N_13185,N_11082,N_11854);
nor U13186 (N_13186,N_10510,N_11500);
xnor U13187 (N_13187,N_10088,N_10251);
nand U13188 (N_13188,N_10906,N_11449);
nand U13189 (N_13189,N_11608,N_10277);
xnor U13190 (N_13190,N_10457,N_11800);
xnor U13191 (N_13191,N_11333,N_11936);
and U13192 (N_13192,N_11992,N_10779);
nor U13193 (N_13193,N_10514,N_10123);
and U13194 (N_13194,N_11101,N_10992);
xor U13195 (N_13195,N_10375,N_10158);
or U13196 (N_13196,N_10472,N_11461);
nand U13197 (N_13197,N_11738,N_11031);
nand U13198 (N_13198,N_11812,N_10878);
nor U13199 (N_13199,N_11974,N_10950);
nand U13200 (N_13200,N_11400,N_11115);
nor U13201 (N_13201,N_10060,N_10269);
xor U13202 (N_13202,N_11060,N_11017);
nor U13203 (N_13203,N_11259,N_10566);
or U13204 (N_13204,N_11184,N_11464);
nor U13205 (N_13205,N_10209,N_10770);
nor U13206 (N_13206,N_11429,N_10694);
nand U13207 (N_13207,N_10025,N_11689);
nor U13208 (N_13208,N_11078,N_10134);
xor U13209 (N_13209,N_10087,N_11566);
nor U13210 (N_13210,N_10424,N_10716);
xnor U13211 (N_13211,N_11727,N_11525);
xor U13212 (N_13212,N_11031,N_10663);
nand U13213 (N_13213,N_11991,N_10706);
xor U13214 (N_13214,N_10841,N_10442);
or U13215 (N_13215,N_11818,N_11181);
xnor U13216 (N_13216,N_10267,N_11425);
nor U13217 (N_13217,N_10837,N_11050);
nor U13218 (N_13218,N_11964,N_10820);
nor U13219 (N_13219,N_10182,N_11251);
nand U13220 (N_13220,N_10778,N_10457);
nand U13221 (N_13221,N_10371,N_10261);
nor U13222 (N_13222,N_10600,N_11667);
or U13223 (N_13223,N_10813,N_11355);
nor U13224 (N_13224,N_11389,N_10147);
nor U13225 (N_13225,N_10494,N_10080);
nor U13226 (N_13226,N_10846,N_11728);
xor U13227 (N_13227,N_10214,N_11425);
nor U13228 (N_13228,N_10658,N_11238);
or U13229 (N_13229,N_11535,N_10038);
nor U13230 (N_13230,N_10977,N_11595);
or U13231 (N_13231,N_10367,N_11947);
xor U13232 (N_13232,N_10643,N_10956);
and U13233 (N_13233,N_10089,N_10212);
or U13234 (N_13234,N_10385,N_10310);
xor U13235 (N_13235,N_11577,N_11660);
xor U13236 (N_13236,N_10296,N_11257);
nand U13237 (N_13237,N_11921,N_11621);
and U13238 (N_13238,N_11848,N_11690);
nand U13239 (N_13239,N_10941,N_10606);
xor U13240 (N_13240,N_11873,N_10977);
and U13241 (N_13241,N_10462,N_11507);
and U13242 (N_13242,N_10131,N_10919);
or U13243 (N_13243,N_10965,N_10797);
nand U13244 (N_13244,N_10127,N_11723);
xnor U13245 (N_13245,N_11082,N_11554);
and U13246 (N_13246,N_10373,N_11917);
and U13247 (N_13247,N_10327,N_10876);
or U13248 (N_13248,N_10637,N_11937);
nand U13249 (N_13249,N_11972,N_11305);
or U13250 (N_13250,N_11078,N_10712);
nand U13251 (N_13251,N_11083,N_11583);
and U13252 (N_13252,N_11279,N_11304);
nand U13253 (N_13253,N_11026,N_10677);
nand U13254 (N_13254,N_10433,N_10041);
nand U13255 (N_13255,N_10277,N_10755);
or U13256 (N_13256,N_11183,N_10687);
nand U13257 (N_13257,N_10043,N_10523);
nor U13258 (N_13258,N_10439,N_10791);
xor U13259 (N_13259,N_10543,N_10159);
or U13260 (N_13260,N_10014,N_11124);
and U13261 (N_13261,N_11743,N_11364);
nand U13262 (N_13262,N_11818,N_10444);
or U13263 (N_13263,N_10911,N_11272);
or U13264 (N_13264,N_11820,N_11859);
nor U13265 (N_13265,N_11158,N_11493);
or U13266 (N_13266,N_10172,N_11012);
and U13267 (N_13267,N_10651,N_10291);
nor U13268 (N_13268,N_11955,N_11685);
nor U13269 (N_13269,N_10246,N_10110);
nor U13270 (N_13270,N_11099,N_11517);
or U13271 (N_13271,N_10602,N_11395);
and U13272 (N_13272,N_10295,N_10758);
nor U13273 (N_13273,N_11199,N_10890);
and U13274 (N_13274,N_11844,N_10600);
and U13275 (N_13275,N_10355,N_10428);
nand U13276 (N_13276,N_10004,N_11944);
or U13277 (N_13277,N_11926,N_10643);
and U13278 (N_13278,N_10503,N_11994);
nand U13279 (N_13279,N_11911,N_11791);
xnor U13280 (N_13280,N_11749,N_10270);
xor U13281 (N_13281,N_11127,N_11119);
nor U13282 (N_13282,N_10580,N_10000);
nor U13283 (N_13283,N_10380,N_10497);
nand U13284 (N_13284,N_10436,N_11278);
xnor U13285 (N_13285,N_10978,N_11865);
or U13286 (N_13286,N_10741,N_10267);
and U13287 (N_13287,N_10896,N_11940);
xnor U13288 (N_13288,N_11566,N_10031);
or U13289 (N_13289,N_11936,N_10315);
nand U13290 (N_13290,N_11975,N_11676);
xor U13291 (N_13291,N_10268,N_11010);
nor U13292 (N_13292,N_10700,N_10113);
and U13293 (N_13293,N_10966,N_10182);
and U13294 (N_13294,N_11880,N_11749);
nor U13295 (N_13295,N_10309,N_11144);
nor U13296 (N_13296,N_11522,N_10808);
nor U13297 (N_13297,N_11860,N_11924);
xor U13298 (N_13298,N_10395,N_10726);
and U13299 (N_13299,N_11864,N_10998);
nand U13300 (N_13300,N_10265,N_10538);
or U13301 (N_13301,N_10790,N_10748);
and U13302 (N_13302,N_10589,N_11471);
nor U13303 (N_13303,N_11925,N_10683);
and U13304 (N_13304,N_11090,N_10467);
and U13305 (N_13305,N_11485,N_10673);
xor U13306 (N_13306,N_11588,N_11410);
or U13307 (N_13307,N_10561,N_11740);
nor U13308 (N_13308,N_10489,N_11119);
xor U13309 (N_13309,N_10018,N_11952);
or U13310 (N_13310,N_10060,N_11198);
nor U13311 (N_13311,N_10777,N_10035);
or U13312 (N_13312,N_11682,N_11331);
xor U13313 (N_13313,N_10100,N_11566);
and U13314 (N_13314,N_11111,N_11420);
nor U13315 (N_13315,N_11189,N_11879);
xnor U13316 (N_13316,N_10070,N_10063);
xnor U13317 (N_13317,N_10195,N_11661);
xnor U13318 (N_13318,N_11926,N_10513);
or U13319 (N_13319,N_11418,N_10403);
or U13320 (N_13320,N_10740,N_10018);
and U13321 (N_13321,N_11316,N_11133);
nor U13322 (N_13322,N_11077,N_11757);
nand U13323 (N_13323,N_11113,N_11382);
nor U13324 (N_13324,N_11589,N_11209);
and U13325 (N_13325,N_10017,N_11124);
xnor U13326 (N_13326,N_10855,N_10994);
nor U13327 (N_13327,N_11229,N_11570);
and U13328 (N_13328,N_11267,N_11750);
xnor U13329 (N_13329,N_11049,N_11334);
and U13330 (N_13330,N_10111,N_11983);
or U13331 (N_13331,N_10519,N_11843);
or U13332 (N_13332,N_10799,N_11949);
and U13333 (N_13333,N_11721,N_11722);
nand U13334 (N_13334,N_10196,N_10042);
nand U13335 (N_13335,N_10151,N_11700);
and U13336 (N_13336,N_11592,N_10210);
and U13337 (N_13337,N_10571,N_10524);
xor U13338 (N_13338,N_11512,N_11554);
nand U13339 (N_13339,N_10509,N_10385);
or U13340 (N_13340,N_10396,N_11760);
or U13341 (N_13341,N_11174,N_11013);
nand U13342 (N_13342,N_11799,N_10463);
xor U13343 (N_13343,N_10292,N_10202);
xor U13344 (N_13344,N_10066,N_10386);
or U13345 (N_13345,N_11477,N_10716);
nand U13346 (N_13346,N_11695,N_10798);
xor U13347 (N_13347,N_10033,N_10165);
and U13348 (N_13348,N_11242,N_11035);
or U13349 (N_13349,N_11827,N_10820);
or U13350 (N_13350,N_11863,N_10084);
xor U13351 (N_13351,N_11326,N_11738);
nor U13352 (N_13352,N_11801,N_11395);
nor U13353 (N_13353,N_11312,N_11259);
and U13354 (N_13354,N_11074,N_11630);
xnor U13355 (N_13355,N_10876,N_10513);
or U13356 (N_13356,N_11321,N_10811);
nor U13357 (N_13357,N_11048,N_11520);
xnor U13358 (N_13358,N_11273,N_11130);
xnor U13359 (N_13359,N_10898,N_11789);
and U13360 (N_13360,N_11775,N_10120);
and U13361 (N_13361,N_11154,N_11885);
nor U13362 (N_13362,N_10144,N_10639);
and U13363 (N_13363,N_10499,N_10343);
nand U13364 (N_13364,N_10750,N_10650);
or U13365 (N_13365,N_11479,N_10395);
nand U13366 (N_13366,N_11965,N_10571);
and U13367 (N_13367,N_11632,N_10236);
or U13368 (N_13368,N_11882,N_10518);
nor U13369 (N_13369,N_11594,N_10368);
or U13370 (N_13370,N_10189,N_10377);
nor U13371 (N_13371,N_11092,N_10876);
or U13372 (N_13372,N_10923,N_11376);
nand U13373 (N_13373,N_11949,N_11338);
xnor U13374 (N_13374,N_10153,N_11961);
nor U13375 (N_13375,N_10881,N_10955);
and U13376 (N_13376,N_11431,N_10238);
nor U13377 (N_13377,N_10864,N_11713);
xnor U13378 (N_13378,N_11705,N_10635);
and U13379 (N_13379,N_10515,N_11580);
xor U13380 (N_13380,N_10205,N_10414);
xnor U13381 (N_13381,N_10344,N_10102);
and U13382 (N_13382,N_10115,N_10382);
nand U13383 (N_13383,N_10937,N_11804);
or U13384 (N_13384,N_11142,N_10539);
and U13385 (N_13385,N_10379,N_11398);
xor U13386 (N_13386,N_11980,N_10341);
nor U13387 (N_13387,N_10712,N_10898);
nand U13388 (N_13388,N_10263,N_11881);
and U13389 (N_13389,N_10003,N_11347);
and U13390 (N_13390,N_10555,N_10577);
nor U13391 (N_13391,N_11951,N_10830);
xnor U13392 (N_13392,N_10173,N_11110);
xor U13393 (N_13393,N_10861,N_11290);
nor U13394 (N_13394,N_10892,N_10215);
nor U13395 (N_13395,N_10421,N_10986);
or U13396 (N_13396,N_10232,N_10464);
nor U13397 (N_13397,N_11955,N_11050);
nor U13398 (N_13398,N_10653,N_11255);
or U13399 (N_13399,N_11591,N_11714);
or U13400 (N_13400,N_11801,N_11497);
xor U13401 (N_13401,N_11161,N_10403);
xnor U13402 (N_13402,N_11253,N_10856);
and U13403 (N_13403,N_11698,N_11300);
nor U13404 (N_13404,N_11605,N_11016);
nor U13405 (N_13405,N_11249,N_11925);
nor U13406 (N_13406,N_11674,N_11418);
and U13407 (N_13407,N_10690,N_10456);
nand U13408 (N_13408,N_10357,N_10583);
nand U13409 (N_13409,N_10219,N_10703);
xor U13410 (N_13410,N_10307,N_10544);
nor U13411 (N_13411,N_11909,N_11588);
and U13412 (N_13412,N_10236,N_11175);
or U13413 (N_13413,N_11213,N_10824);
or U13414 (N_13414,N_11486,N_10237);
and U13415 (N_13415,N_10045,N_10812);
nand U13416 (N_13416,N_11869,N_11671);
or U13417 (N_13417,N_10629,N_10948);
or U13418 (N_13418,N_10950,N_10525);
and U13419 (N_13419,N_11344,N_10838);
xnor U13420 (N_13420,N_10615,N_11061);
nand U13421 (N_13421,N_10182,N_10471);
nor U13422 (N_13422,N_11356,N_11504);
nand U13423 (N_13423,N_11323,N_10554);
nor U13424 (N_13424,N_10790,N_11539);
nand U13425 (N_13425,N_10011,N_11883);
nand U13426 (N_13426,N_11822,N_10918);
or U13427 (N_13427,N_10462,N_11892);
nor U13428 (N_13428,N_10042,N_11803);
xor U13429 (N_13429,N_10589,N_11415);
nand U13430 (N_13430,N_10333,N_11565);
xor U13431 (N_13431,N_11524,N_11554);
xor U13432 (N_13432,N_10202,N_10727);
or U13433 (N_13433,N_11027,N_11886);
or U13434 (N_13434,N_11269,N_10784);
and U13435 (N_13435,N_10825,N_10867);
and U13436 (N_13436,N_10279,N_10992);
and U13437 (N_13437,N_11858,N_10371);
and U13438 (N_13438,N_10308,N_10625);
or U13439 (N_13439,N_11341,N_10738);
and U13440 (N_13440,N_11847,N_11795);
and U13441 (N_13441,N_10938,N_10722);
and U13442 (N_13442,N_11014,N_11688);
xor U13443 (N_13443,N_11769,N_10057);
nor U13444 (N_13444,N_11258,N_11725);
and U13445 (N_13445,N_11236,N_10632);
nand U13446 (N_13446,N_11773,N_10624);
nor U13447 (N_13447,N_10125,N_10748);
and U13448 (N_13448,N_11456,N_10613);
xnor U13449 (N_13449,N_10981,N_11597);
xor U13450 (N_13450,N_10519,N_11155);
or U13451 (N_13451,N_10646,N_10141);
and U13452 (N_13452,N_11690,N_11224);
or U13453 (N_13453,N_10351,N_11711);
nand U13454 (N_13454,N_10389,N_10753);
nand U13455 (N_13455,N_11117,N_10245);
or U13456 (N_13456,N_11697,N_11721);
or U13457 (N_13457,N_10697,N_10401);
and U13458 (N_13458,N_10825,N_11982);
nand U13459 (N_13459,N_11878,N_11991);
xor U13460 (N_13460,N_10751,N_10705);
nand U13461 (N_13461,N_11160,N_10422);
nand U13462 (N_13462,N_10548,N_10238);
nand U13463 (N_13463,N_11818,N_10129);
nor U13464 (N_13464,N_10815,N_10884);
nor U13465 (N_13465,N_11141,N_11237);
xor U13466 (N_13466,N_11078,N_11971);
or U13467 (N_13467,N_11840,N_10209);
or U13468 (N_13468,N_11778,N_11409);
nor U13469 (N_13469,N_11029,N_11390);
and U13470 (N_13470,N_11574,N_11743);
xnor U13471 (N_13471,N_10303,N_11957);
and U13472 (N_13472,N_10534,N_11254);
or U13473 (N_13473,N_10741,N_10277);
nor U13474 (N_13474,N_10610,N_10431);
and U13475 (N_13475,N_11827,N_10818);
and U13476 (N_13476,N_10486,N_11969);
nor U13477 (N_13477,N_11307,N_10787);
and U13478 (N_13478,N_10503,N_11874);
and U13479 (N_13479,N_11766,N_11377);
or U13480 (N_13480,N_10082,N_11196);
and U13481 (N_13481,N_11549,N_11407);
xor U13482 (N_13482,N_11022,N_11649);
or U13483 (N_13483,N_10556,N_10399);
nor U13484 (N_13484,N_11320,N_11616);
and U13485 (N_13485,N_11090,N_11055);
xnor U13486 (N_13486,N_10216,N_11567);
nor U13487 (N_13487,N_11218,N_10484);
nor U13488 (N_13488,N_11437,N_10082);
nand U13489 (N_13489,N_11821,N_10973);
xor U13490 (N_13490,N_10288,N_10279);
xnor U13491 (N_13491,N_10102,N_11182);
xor U13492 (N_13492,N_11929,N_11907);
or U13493 (N_13493,N_11251,N_11398);
and U13494 (N_13494,N_10051,N_10241);
or U13495 (N_13495,N_11048,N_11849);
or U13496 (N_13496,N_11302,N_10493);
nor U13497 (N_13497,N_10346,N_10303);
and U13498 (N_13498,N_10539,N_10450);
and U13499 (N_13499,N_11034,N_10507);
or U13500 (N_13500,N_11335,N_10668);
or U13501 (N_13501,N_10993,N_10424);
nand U13502 (N_13502,N_11166,N_11984);
and U13503 (N_13503,N_11397,N_10098);
xnor U13504 (N_13504,N_10254,N_11286);
and U13505 (N_13505,N_10212,N_10201);
and U13506 (N_13506,N_11382,N_10275);
and U13507 (N_13507,N_10788,N_10630);
nor U13508 (N_13508,N_10583,N_11279);
and U13509 (N_13509,N_10299,N_10052);
xor U13510 (N_13510,N_11045,N_10751);
nor U13511 (N_13511,N_11631,N_11096);
nor U13512 (N_13512,N_11369,N_10155);
or U13513 (N_13513,N_11206,N_10587);
nand U13514 (N_13514,N_10661,N_11575);
and U13515 (N_13515,N_10398,N_11820);
or U13516 (N_13516,N_10510,N_10754);
nand U13517 (N_13517,N_10296,N_11993);
nand U13518 (N_13518,N_10040,N_11865);
and U13519 (N_13519,N_10100,N_11847);
and U13520 (N_13520,N_10886,N_10501);
nor U13521 (N_13521,N_10481,N_11422);
and U13522 (N_13522,N_11586,N_10438);
xnor U13523 (N_13523,N_10893,N_10359);
nand U13524 (N_13524,N_11049,N_10939);
or U13525 (N_13525,N_11563,N_10147);
nand U13526 (N_13526,N_10181,N_10136);
and U13527 (N_13527,N_11959,N_11793);
and U13528 (N_13528,N_11455,N_11669);
or U13529 (N_13529,N_10520,N_11427);
nand U13530 (N_13530,N_10939,N_10238);
or U13531 (N_13531,N_11449,N_11656);
nor U13532 (N_13532,N_11761,N_11424);
xor U13533 (N_13533,N_10812,N_10049);
xnor U13534 (N_13534,N_11284,N_10320);
nand U13535 (N_13535,N_10031,N_11246);
xnor U13536 (N_13536,N_11599,N_10531);
and U13537 (N_13537,N_11861,N_11044);
and U13538 (N_13538,N_11382,N_11598);
nor U13539 (N_13539,N_10179,N_10514);
and U13540 (N_13540,N_10383,N_11537);
nor U13541 (N_13541,N_10953,N_11603);
or U13542 (N_13542,N_11709,N_11471);
nor U13543 (N_13543,N_11793,N_10665);
nand U13544 (N_13544,N_11104,N_10724);
nand U13545 (N_13545,N_10327,N_10225);
nand U13546 (N_13546,N_11236,N_11210);
and U13547 (N_13547,N_10770,N_11310);
nand U13548 (N_13548,N_10472,N_11591);
nor U13549 (N_13549,N_10823,N_10504);
nand U13550 (N_13550,N_11601,N_10419);
nand U13551 (N_13551,N_11500,N_10048);
nor U13552 (N_13552,N_11957,N_11705);
nor U13553 (N_13553,N_10881,N_11948);
nand U13554 (N_13554,N_10471,N_10086);
or U13555 (N_13555,N_11731,N_10040);
or U13556 (N_13556,N_10847,N_10958);
xnor U13557 (N_13557,N_10182,N_11910);
nand U13558 (N_13558,N_10922,N_10389);
and U13559 (N_13559,N_10447,N_10448);
nand U13560 (N_13560,N_10049,N_10227);
xnor U13561 (N_13561,N_10147,N_11548);
nor U13562 (N_13562,N_10095,N_11385);
nor U13563 (N_13563,N_10487,N_10599);
nor U13564 (N_13564,N_10022,N_11600);
xnor U13565 (N_13565,N_11461,N_10026);
xor U13566 (N_13566,N_10583,N_10318);
and U13567 (N_13567,N_11537,N_11844);
nand U13568 (N_13568,N_11449,N_11847);
and U13569 (N_13569,N_10693,N_10329);
nand U13570 (N_13570,N_10591,N_10472);
nor U13571 (N_13571,N_10695,N_10858);
and U13572 (N_13572,N_11161,N_10863);
xnor U13573 (N_13573,N_11509,N_10916);
nor U13574 (N_13574,N_11249,N_10606);
nor U13575 (N_13575,N_10401,N_11509);
nor U13576 (N_13576,N_10531,N_11743);
nor U13577 (N_13577,N_11535,N_11903);
and U13578 (N_13578,N_11849,N_11349);
and U13579 (N_13579,N_10034,N_10702);
xnor U13580 (N_13580,N_10191,N_11952);
nor U13581 (N_13581,N_10818,N_11465);
nand U13582 (N_13582,N_11647,N_11928);
nor U13583 (N_13583,N_11469,N_11595);
xor U13584 (N_13584,N_11495,N_11332);
nor U13585 (N_13585,N_11783,N_10279);
and U13586 (N_13586,N_11235,N_10168);
nand U13587 (N_13587,N_11741,N_10976);
nor U13588 (N_13588,N_10791,N_10870);
nor U13589 (N_13589,N_10259,N_11204);
nand U13590 (N_13590,N_10554,N_11007);
nand U13591 (N_13591,N_10365,N_10986);
or U13592 (N_13592,N_10904,N_11669);
nand U13593 (N_13593,N_11242,N_10517);
nor U13594 (N_13594,N_10219,N_11675);
xor U13595 (N_13595,N_10053,N_11580);
xor U13596 (N_13596,N_11449,N_10409);
or U13597 (N_13597,N_11720,N_10928);
nand U13598 (N_13598,N_11727,N_11141);
and U13599 (N_13599,N_11758,N_10969);
nand U13600 (N_13600,N_11974,N_10661);
and U13601 (N_13601,N_11259,N_11941);
and U13602 (N_13602,N_10319,N_10663);
or U13603 (N_13603,N_10790,N_11348);
nand U13604 (N_13604,N_10902,N_10132);
xnor U13605 (N_13605,N_11000,N_10522);
nor U13606 (N_13606,N_11685,N_10042);
xor U13607 (N_13607,N_11265,N_10452);
nor U13608 (N_13608,N_10728,N_11532);
xnor U13609 (N_13609,N_11458,N_10812);
nand U13610 (N_13610,N_11503,N_11920);
nor U13611 (N_13611,N_11825,N_10044);
nor U13612 (N_13612,N_11241,N_10642);
nand U13613 (N_13613,N_11867,N_11336);
or U13614 (N_13614,N_10328,N_11085);
nand U13615 (N_13615,N_10871,N_11886);
xnor U13616 (N_13616,N_10877,N_10741);
nand U13617 (N_13617,N_10580,N_10109);
xor U13618 (N_13618,N_10355,N_11301);
xnor U13619 (N_13619,N_10437,N_10884);
nand U13620 (N_13620,N_10874,N_11225);
nor U13621 (N_13621,N_11899,N_10670);
nand U13622 (N_13622,N_10535,N_11012);
nor U13623 (N_13623,N_10664,N_11726);
nand U13624 (N_13624,N_10543,N_11448);
or U13625 (N_13625,N_11615,N_10091);
or U13626 (N_13626,N_11963,N_11463);
and U13627 (N_13627,N_11853,N_11711);
xor U13628 (N_13628,N_11126,N_11787);
or U13629 (N_13629,N_10551,N_11954);
nor U13630 (N_13630,N_10177,N_10371);
nand U13631 (N_13631,N_10118,N_10051);
nand U13632 (N_13632,N_10360,N_10666);
nand U13633 (N_13633,N_11918,N_11773);
and U13634 (N_13634,N_10387,N_11144);
xor U13635 (N_13635,N_11919,N_11838);
or U13636 (N_13636,N_11640,N_10148);
nand U13637 (N_13637,N_11467,N_11164);
xor U13638 (N_13638,N_10536,N_11371);
and U13639 (N_13639,N_11459,N_10819);
xnor U13640 (N_13640,N_10788,N_11974);
nor U13641 (N_13641,N_10586,N_11985);
nor U13642 (N_13642,N_11068,N_11280);
and U13643 (N_13643,N_10301,N_11386);
nor U13644 (N_13644,N_11787,N_11307);
or U13645 (N_13645,N_11064,N_11963);
or U13646 (N_13646,N_10480,N_10734);
and U13647 (N_13647,N_11115,N_10187);
nor U13648 (N_13648,N_11659,N_11792);
nor U13649 (N_13649,N_10235,N_11599);
nor U13650 (N_13650,N_11938,N_11207);
nor U13651 (N_13651,N_10564,N_10201);
or U13652 (N_13652,N_11833,N_11666);
nor U13653 (N_13653,N_10913,N_10399);
xor U13654 (N_13654,N_11004,N_11267);
or U13655 (N_13655,N_10671,N_11106);
and U13656 (N_13656,N_11948,N_11906);
nor U13657 (N_13657,N_10908,N_10847);
or U13658 (N_13658,N_11010,N_11547);
xnor U13659 (N_13659,N_11643,N_10086);
nand U13660 (N_13660,N_11877,N_10221);
or U13661 (N_13661,N_10496,N_11402);
and U13662 (N_13662,N_10224,N_10524);
and U13663 (N_13663,N_10048,N_11046);
xor U13664 (N_13664,N_10640,N_10324);
or U13665 (N_13665,N_10729,N_11699);
nor U13666 (N_13666,N_11956,N_10516);
or U13667 (N_13667,N_11631,N_10545);
and U13668 (N_13668,N_10129,N_11607);
xnor U13669 (N_13669,N_11874,N_11277);
nor U13670 (N_13670,N_11534,N_11953);
nor U13671 (N_13671,N_11858,N_11246);
or U13672 (N_13672,N_10610,N_10069);
nand U13673 (N_13673,N_11036,N_11330);
nand U13674 (N_13674,N_10860,N_11291);
xnor U13675 (N_13675,N_11804,N_11679);
or U13676 (N_13676,N_11114,N_11308);
xnor U13677 (N_13677,N_11301,N_10111);
xnor U13678 (N_13678,N_10196,N_10092);
nand U13679 (N_13679,N_10588,N_11512);
nor U13680 (N_13680,N_11425,N_10856);
and U13681 (N_13681,N_11828,N_11574);
nor U13682 (N_13682,N_10696,N_11934);
nor U13683 (N_13683,N_11636,N_11340);
nor U13684 (N_13684,N_10209,N_11650);
nor U13685 (N_13685,N_11274,N_10519);
nor U13686 (N_13686,N_10499,N_10555);
and U13687 (N_13687,N_11144,N_11631);
nand U13688 (N_13688,N_11701,N_10894);
nor U13689 (N_13689,N_11631,N_10110);
xnor U13690 (N_13690,N_11279,N_11704);
nand U13691 (N_13691,N_10896,N_11954);
nand U13692 (N_13692,N_10460,N_10434);
xnor U13693 (N_13693,N_10678,N_11198);
nand U13694 (N_13694,N_11668,N_10205);
and U13695 (N_13695,N_11296,N_10867);
or U13696 (N_13696,N_10241,N_11374);
nand U13697 (N_13697,N_11430,N_11259);
nand U13698 (N_13698,N_11513,N_11235);
and U13699 (N_13699,N_10601,N_11337);
xor U13700 (N_13700,N_10715,N_10784);
and U13701 (N_13701,N_11790,N_10930);
nor U13702 (N_13702,N_10730,N_10039);
and U13703 (N_13703,N_11898,N_11235);
and U13704 (N_13704,N_11887,N_11199);
nand U13705 (N_13705,N_10666,N_11812);
xor U13706 (N_13706,N_11612,N_10277);
nand U13707 (N_13707,N_10548,N_10440);
and U13708 (N_13708,N_11157,N_11744);
nor U13709 (N_13709,N_10262,N_10019);
or U13710 (N_13710,N_10514,N_10109);
or U13711 (N_13711,N_11247,N_10769);
and U13712 (N_13712,N_11757,N_10758);
xor U13713 (N_13713,N_10004,N_10144);
xor U13714 (N_13714,N_11959,N_10318);
xor U13715 (N_13715,N_10051,N_10820);
nand U13716 (N_13716,N_10011,N_11027);
xnor U13717 (N_13717,N_11306,N_10169);
nand U13718 (N_13718,N_10972,N_10840);
or U13719 (N_13719,N_10769,N_10212);
or U13720 (N_13720,N_11905,N_10025);
or U13721 (N_13721,N_11362,N_10413);
xnor U13722 (N_13722,N_10223,N_11859);
or U13723 (N_13723,N_11352,N_11068);
nand U13724 (N_13724,N_11624,N_11001);
xor U13725 (N_13725,N_10218,N_11516);
xor U13726 (N_13726,N_10631,N_11993);
and U13727 (N_13727,N_11625,N_11318);
nor U13728 (N_13728,N_11068,N_10415);
and U13729 (N_13729,N_11791,N_11688);
xor U13730 (N_13730,N_11080,N_10038);
xor U13731 (N_13731,N_11683,N_10198);
nand U13732 (N_13732,N_11850,N_11668);
nor U13733 (N_13733,N_11488,N_10850);
nand U13734 (N_13734,N_10863,N_11069);
or U13735 (N_13735,N_10779,N_10545);
or U13736 (N_13736,N_10383,N_11193);
nand U13737 (N_13737,N_11302,N_11348);
and U13738 (N_13738,N_10474,N_10153);
nand U13739 (N_13739,N_10086,N_10381);
xnor U13740 (N_13740,N_10419,N_10868);
and U13741 (N_13741,N_10328,N_11527);
or U13742 (N_13742,N_11645,N_11464);
nand U13743 (N_13743,N_10916,N_11996);
and U13744 (N_13744,N_10449,N_11664);
or U13745 (N_13745,N_10650,N_11428);
or U13746 (N_13746,N_10937,N_10894);
nand U13747 (N_13747,N_10576,N_11305);
xor U13748 (N_13748,N_10472,N_11146);
and U13749 (N_13749,N_10908,N_10786);
xor U13750 (N_13750,N_10869,N_11036);
xor U13751 (N_13751,N_10105,N_10000);
or U13752 (N_13752,N_10072,N_11150);
nand U13753 (N_13753,N_11924,N_10143);
or U13754 (N_13754,N_11649,N_11601);
or U13755 (N_13755,N_11413,N_10222);
nand U13756 (N_13756,N_10451,N_10844);
and U13757 (N_13757,N_10699,N_11862);
and U13758 (N_13758,N_11730,N_10137);
xor U13759 (N_13759,N_10770,N_10037);
nand U13760 (N_13760,N_10098,N_10282);
nand U13761 (N_13761,N_10534,N_11578);
or U13762 (N_13762,N_11842,N_10982);
and U13763 (N_13763,N_10250,N_10290);
or U13764 (N_13764,N_10665,N_10992);
or U13765 (N_13765,N_10310,N_11255);
xnor U13766 (N_13766,N_10212,N_10358);
nand U13767 (N_13767,N_10217,N_10027);
nand U13768 (N_13768,N_11153,N_10836);
and U13769 (N_13769,N_11688,N_11965);
nand U13770 (N_13770,N_10579,N_10329);
or U13771 (N_13771,N_10472,N_11778);
and U13772 (N_13772,N_10868,N_11017);
nand U13773 (N_13773,N_10452,N_11096);
nor U13774 (N_13774,N_10708,N_11712);
nor U13775 (N_13775,N_10761,N_11590);
or U13776 (N_13776,N_11531,N_11836);
nor U13777 (N_13777,N_11859,N_10198);
nor U13778 (N_13778,N_10546,N_11745);
nand U13779 (N_13779,N_11877,N_10950);
xnor U13780 (N_13780,N_11740,N_10245);
or U13781 (N_13781,N_10723,N_11762);
xor U13782 (N_13782,N_10936,N_10514);
xor U13783 (N_13783,N_10663,N_10527);
nor U13784 (N_13784,N_10868,N_11206);
xnor U13785 (N_13785,N_10553,N_11895);
nor U13786 (N_13786,N_11397,N_10575);
or U13787 (N_13787,N_10489,N_10956);
and U13788 (N_13788,N_11602,N_10395);
and U13789 (N_13789,N_10396,N_10366);
and U13790 (N_13790,N_11198,N_10810);
or U13791 (N_13791,N_11233,N_10737);
and U13792 (N_13792,N_10730,N_10164);
and U13793 (N_13793,N_10063,N_10269);
or U13794 (N_13794,N_11691,N_10583);
or U13795 (N_13795,N_10071,N_11886);
xor U13796 (N_13796,N_11578,N_10419);
nand U13797 (N_13797,N_11732,N_10697);
or U13798 (N_13798,N_10900,N_11835);
nand U13799 (N_13799,N_11118,N_10659);
nand U13800 (N_13800,N_11962,N_11786);
nor U13801 (N_13801,N_11043,N_11016);
nor U13802 (N_13802,N_11534,N_11814);
or U13803 (N_13803,N_11465,N_11791);
and U13804 (N_13804,N_11708,N_11440);
nor U13805 (N_13805,N_11141,N_11939);
nand U13806 (N_13806,N_10342,N_11912);
xnor U13807 (N_13807,N_10808,N_11519);
nand U13808 (N_13808,N_11235,N_11370);
nand U13809 (N_13809,N_10529,N_11794);
nand U13810 (N_13810,N_11193,N_11844);
nand U13811 (N_13811,N_10700,N_10727);
nor U13812 (N_13812,N_11651,N_11346);
and U13813 (N_13813,N_10222,N_11798);
and U13814 (N_13814,N_10939,N_11194);
or U13815 (N_13815,N_10723,N_10047);
nor U13816 (N_13816,N_10695,N_10071);
and U13817 (N_13817,N_10857,N_10688);
or U13818 (N_13818,N_11128,N_11394);
and U13819 (N_13819,N_11359,N_11065);
xnor U13820 (N_13820,N_11914,N_11559);
or U13821 (N_13821,N_10627,N_11324);
or U13822 (N_13822,N_11351,N_11266);
nor U13823 (N_13823,N_11352,N_11152);
nor U13824 (N_13824,N_11103,N_10376);
or U13825 (N_13825,N_10501,N_10167);
and U13826 (N_13826,N_11434,N_11572);
or U13827 (N_13827,N_10267,N_11168);
nor U13828 (N_13828,N_10744,N_10161);
and U13829 (N_13829,N_10504,N_11519);
nand U13830 (N_13830,N_11354,N_10280);
or U13831 (N_13831,N_10447,N_11379);
nand U13832 (N_13832,N_10734,N_10769);
nand U13833 (N_13833,N_10478,N_11835);
or U13834 (N_13834,N_11697,N_11061);
and U13835 (N_13835,N_10899,N_10694);
nor U13836 (N_13836,N_10060,N_10724);
nand U13837 (N_13837,N_11907,N_11115);
and U13838 (N_13838,N_11355,N_10997);
and U13839 (N_13839,N_11329,N_11917);
or U13840 (N_13840,N_10273,N_10082);
xnor U13841 (N_13841,N_10804,N_11357);
and U13842 (N_13842,N_11762,N_10555);
xnor U13843 (N_13843,N_11952,N_11099);
or U13844 (N_13844,N_10694,N_10596);
or U13845 (N_13845,N_11527,N_11283);
xnor U13846 (N_13846,N_11405,N_11491);
or U13847 (N_13847,N_11585,N_11414);
or U13848 (N_13848,N_11754,N_11016);
and U13849 (N_13849,N_11865,N_10279);
nand U13850 (N_13850,N_10012,N_11686);
or U13851 (N_13851,N_10046,N_11671);
xnor U13852 (N_13852,N_10485,N_10306);
and U13853 (N_13853,N_11774,N_11477);
xor U13854 (N_13854,N_11545,N_10548);
nand U13855 (N_13855,N_10341,N_10783);
nor U13856 (N_13856,N_11059,N_11019);
or U13857 (N_13857,N_11520,N_10789);
nor U13858 (N_13858,N_11555,N_10681);
nor U13859 (N_13859,N_10895,N_10817);
or U13860 (N_13860,N_10127,N_11568);
nor U13861 (N_13861,N_11123,N_11639);
nor U13862 (N_13862,N_10884,N_11373);
nand U13863 (N_13863,N_11955,N_10535);
xnor U13864 (N_13864,N_11795,N_11289);
nand U13865 (N_13865,N_10418,N_11330);
and U13866 (N_13866,N_11219,N_11380);
xnor U13867 (N_13867,N_10324,N_11312);
nor U13868 (N_13868,N_10979,N_11291);
and U13869 (N_13869,N_11315,N_10104);
or U13870 (N_13870,N_11649,N_11807);
nor U13871 (N_13871,N_10335,N_10406);
xnor U13872 (N_13872,N_11969,N_10270);
nor U13873 (N_13873,N_10493,N_10038);
or U13874 (N_13874,N_10428,N_10444);
nand U13875 (N_13875,N_11264,N_11604);
xnor U13876 (N_13876,N_10619,N_10833);
nand U13877 (N_13877,N_11748,N_10564);
and U13878 (N_13878,N_10080,N_10807);
nand U13879 (N_13879,N_10923,N_10776);
nor U13880 (N_13880,N_11732,N_11919);
xor U13881 (N_13881,N_11408,N_10449);
nor U13882 (N_13882,N_10894,N_11451);
nand U13883 (N_13883,N_10351,N_11648);
nor U13884 (N_13884,N_11580,N_10934);
nor U13885 (N_13885,N_11807,N_11925);
or U13886 (N_13886,N_11288,N_10879);
nor U13887 (N_13887,N_11923,N_10421);
or U13888 (N_13888,N_11952,N_10178);
xnor U13889 (N_13889,N_11619,N_10645);
xor U13890 (N_13890,N_10509,N_11936);
nor U13891 (N_13891,N_11261,N_10163);
nor U13892 (N_13892,N_11207,N_10774);
nand U13893 (N_13893,N_11241,N_10590);
and U13894 (N_13894,N_11876,N_11226);
xor U13895 (N_13895,N_10600,N_11430);
and U13896 (N_13896,N_11737,N_11232);
nor U13897 (N_13897,N_10140,N_11606);
xnor U13898 (N_13898,N_11283,N_10205);
and U13899 (N_13899,N_10665,N_10986);
nand U13900 (N_13900,N_10963,N_11834);
nor U13901 (N_13901,N_10026,N_10217);
or U13902 (N_13902,N_10727,N_10184);
or U13903 (N_13903,N_10560,N_11530);
nor U13904 (N_13904,N_10115,N_11892);
xor U13905 (N_13905,N_11040,N_10176);
or U13906 (N_13906,N_11405,N_10264);
nand U13907 (N_13907,N_10862,N_11069);
nor U13908 (N_13908,N_10934,N_10536);
nor U13909 (N_13909,N_11261,N_11735);
or U13910 (N_13910,N_11385,N_11902);
xor U13911 (N_13911,N_11928,N_11115);
and U13912 (N_13912,N_11012,N_10351);
or U13913 (N_13913,N_10627,N_10334);
nand U13914 (N_13914,N_11629,N_10098);
and U13915 (N_13915,N_10974,N_10633);
nor U13916 (N_13916,N_10432,N_11573);
or U13917 (N_13917,N_10206,N_10247);
nand U13918 (N_13918,N_10003,N_11136);
nand U13919 (N_13919,N_11947,N_10951);
and U13920 (N_13920,N_10256,N_10200);
and U13921 (N_13921,N_11610,N_11145);
or U13922 (N_13922,N_10174,N_11367);
xor U13923 (N_13923,N_11819,N_10660);
xnor U13924 (N_13924,N_11884,N_11317);
nand U13925 (N_13925,N_10559,N_10264);
nand U13926 (N_13926,N_11118,N_10622);
nand U13927 (N_13927,N_11201,N_11798);
nor U13928 (N_13928,N_10794,N_11504);
nor U13929 (N_13929,N_10895,N_10378);
and U13930 (N_13930,N_10848,N_11889);
xor U13931 (N_13931,N_10429,N_11969);
or U13932 (N_13932,N_10652,N_10824);
nand U13933 (N_13933,N_11631,N_11802);
nand U13934 (N_13934,N_10886,N_11369);
and U13935 (N_13935,N_10197,N_10156);
and U13936 (N_13936,N_10612,N_11116);
or U13937 (N_13937,N_10749,N_11859);
nand U13938 (N_13938,N_11948,N_10828);
xor U13939 (N_13939,N_10892,N_10019);
or U13940 (N_13940,N_10761,N_11095);
nor U13941 (N_13941,N_10329,N_10684);
xnor U13942 (N_13942,N_11980,N_11987);
and U13943 (N_13943,N_11556,N_11598);
xnor U13944 (N_13944,N_11586,N_11548);
or U13945 (N_13945,N_11624,N_10334);
and U13946 (N_13946,N_11382,N_11714);
nand U13947 (N_13947,N_11914,N_11745);
nand U13948 (N_13948,N_10317,N_10815);
or U13949 (N_13949,N_11744,N_10997);
and U13950 (N_13950,N_11371,N_11329);
nor U13951 (N_13951,N_10923,N_10915);
nand U13952 (N_13952,N_10918,N_10734);
nand U13953 (N_13953,N_10081,N_11502);
nand U13954 (N_13954,N_11049,N_11039);
or U13955 (N_13955,N_11634,N_11561);
or U13956 (N_13956,N_10116,N_10121);
or U13957 (N_13957,N_10745,N_10367);
and U13958 (N_13958,N_11086,N_11552);
or U13959 (N_13959,N_10415,N_11704);
nand U13960 (N_13960,N_11254,N_10753);
or U13961 (N_13961,N_11779,N_11001);
and U13962 (N_13962,N_11677,N_11411);
nand U13963 (N_13963,N_11452,N_10694);
nor U13964 (N_13964,N_10382,N_11504);
and U13965 (N_13965,N_11489,N_10023);
nor U13966 (N_13966,N_10132,N_11688);
xnor U13967 (N_13967,N_10417,N_11972);
nand U13968 (N_13968,N_10591,N_11684);
nand U13969 (N_13969,N_10709,N_10638);
and U13970 (N_13970,N_10719,N_10305);
and U13971 (N_13971,N_10794,N_11519);
nor U13972 (N_13972,N_11184,N_11305);
and U13973 (N_13973,N_10408,N_10198);
nor U13974 (N_13974,N_11889,N_10661);
nor U13975 (N_13975,N_10753,N_11590);
xnor U13976 (N_13976,N_11038,N_11743);
nor U13977 (N_13977,N_10604,N_11555);
xnor U13978 (N_13978,N_10840,N_11681);
or U13979 (N_13979,N_10520,N_11341);
or U13980 (N_13980,N_10403,N_11232);
nor U13981 (N_13981,N_11205,N_10389);
nand U13982 (N_13982,N_11970,N_11312);
xor U13983 (N_13983,N_11289,N_10348);
xor U13984 (N_13984,N_10965,N_11577);
xnor U13985 (N_13985,N_10100,N_10758);
xor U13986 (N_13986,N_10314,N_10661);
nand U13987 (N_13987,N_11738,N_10868);
or U13988 (N_13988,N_11848,N_11073);
nor U13989 (N_13989,N_11586,N_11445);
and U13990 (N_13990,N_11633,N_11883);
nor U13991 (N_13991,N_10886,N_10685);
nor U13992 (N_13992,N_11681,N_11527);
nor U13993 (N_13993,N_11825,N_10429);
nand U13994 (N_13994,N_10109,N_11477);
nand U13995 (N_13995,N_10736,N_10700);
nand U13996 (N_13996,N_10172,N_10899);
xnor U13997 (N_13997,N_10675,N_10153);
nand U13998 (N_13998,N_10158,N_11186);
and U13999 (N_13999,N_11079,N_10883);
and U14000 (N_14000,N_13447,N_12276);
nor U14001 (N_14001,N_12277,N_12397);
nand U14002 (N_14002,N_12543,N_12335);
nand U14003 (N_14003,N_12329,N_13179);
and U14004 (N_14004,N_12432,N_13481);
nor U14005 (N_14005,N_13333,N_12730);
nor U14006 (N_14006,N_12457,N_13293);
nor U14007 (N_14007,N_12932,N_12939);
and U14008 (N_14008,N_12944,N_12478);
xor U14009 (N_14009,N_13156,N_12090);
nand U14010 (N_14010,N_13160,N_13519);
nand U14011 (N_14011,N_12370,N_13269);
nand U14012 (N_14012,N_13327,N_12921);
nand U14013 (N_14013,N_13426,N_12127);
and U14014 (N_14014,N_12321,N_13994);
or U14015 (N_14015,N_12759,N_12157);
nand U14016 (N_14016,N_12264,N_12266);
and U14017 (N_14017,N_12624,N_13795);
nand U14018 (N_14018,N_13559,N_13243);
nand U14019 (N_14019,N_13092,N_12709);
and U14020 (N_14020,N_13338,N_13088);
and U14021 (N_14021,N_12684,N_13822);
and U14022 (N_14022,N_13261,N_13446);
xor U14023 (N_14023,N_12867,N_13251);
nand U14024 (N_14024,N_12604,N_13130);
nor U14025 (N_14025,N_12065,N_13820);
nor U14026 (N_14026,N_13964,N_12360);
and U14027 (N_14027,N_12030,N_13864);
and U14028 (N_14028,N_12561,N_12044);
nor U14029 (N_14029,N_13560,N_12871);
or U14030 (N_14030,N_12070,N_12627);
and U14031 (N_14031,N_12484,N_12280);
xor U14032 (N_14032,N_13692,N_13440);
nand U14033 (N_14033,N_13721,N_12510);
nor U14034 (N_14034,N_13104,N_13020);
nor U14035 (N_14035,N_12503,N_13655);
nor U14036 (N_14036,N_13277,N_12803);
or U14037 (N_14037,N_12783,N_13146);
xnor U14038 (N_14038,N_12073,N_13137);
xor U14039 (N_14039,N_13279,N_12592);
nor U14040 (N_14040,N_13922,N_12888);
nand U14041 (N_14041,N_12825,N_13352);
or U14042 (N_14042,N_13969,N_13726);
xnor U14043 (N_14043,N_12762,N_13660);
xor U14044 (N_14044,N_12590,N_13520);
nand U14045 (N_14045,N_13521,N_13834);
or U14046 (N_14046,N_13491,N_13400);
and U14047 (N_14047,N_12751,N_13363);
or U14048 (N_14048,N_13693,N_13851);
xor U14049 (N_14049,N_13295,N_13013);
and U14050 (N_14050,N_12663,N_12564);
or U14051 (N_14051,N_13948,N_12567);
and U14052 (N_14052,N_12823,N_13229);
and U14053 (N_14053,N_13696,N_12364);
or U14054 (N_14054,N_13956,N_13708);
and U14055 (N_14055,N_12128,N_13915);
nand U14056 (N_14056,N_12495,N_13935);
and U14057 (N_14057,N_13195,N_12801);
and U14058 (N_14058,N_13078,N_12525);
nor U14059 (N_14059,N_13443,N_13133);
xor U14060 (N_14060,N_13984,N_13030);
nor U14061 (N_14061,N_12753,N_12327);
and U14062 (N_14062,N_12454,N_12973);
or U14063 (N_14063,N_13397,N_13444);
nand U14064 (N_14064,N_12750,N_13373);
nand U14065 (N_14065,N_12602,N_13186);
nand U14066 (N_14066,N_13159,N_13100);
nand U14067 (N_14067,N_13334,N_12548);
and U14068 (N_14068,N_12497,N_12647);
nor U14069 (N_14069,N_12076,N_12284);
xor U14070 (N_14070,N_12047,N_13348);
nand U14071 (N_14071,N_13573,N_13758);
xnor U14072 (N_14072,N_12104,N_13052);
and U14073 (N_14073,N_12470,N_12930);
and U14074 (N_14074,N_12092,N_12231);
or U14075 (N_14075,N_12328,N_13585);
nor U14076 (N_14076,N_12173,N_13870);
nand U14077 (N_14077,N_12574,N_12075);
and U14078 (N_14078,N_12737,N_13194);
nand U14079 (N_14079,N_13533,N_12512);
nand U14080 (N_14080,N_12140,N_12797);
and U14081 (N_14081,N_12638,N_13061);
and U14082 (N_14082,N_13597,N_12630);
or U14083 (N_14083,N_13668,N_12441);
xor U14084 (N_14084,N_13752,N_13429);
or U14085 (N_14085,N_12527,N_13084);
and U14086 (N_14086,N_12203,N_12336);
xor U14087 (N_14087,N_12171,N_12131);
nand U14088 (N_14088,N_12225,N_13673);
or U14089 (N_14089,N_12198,N_13177);
nor U14090 (N_14090,N_13930,N_12752);
and U14091 (N_14091,N_13578,N_13152);
nor U14092 (N_14092,N_13147,N_12515);
or U14093 (N_14093,N_13980,N_13210);
nand U14094 (N_14094,N_13918,N_12694);
nor U14095 (N_14095,N_12887,N_13213);
nor U14096 (N_14096,N_13958,N_13891);
xor U14097 (N_14097,N_12387,N_12286);
or U14098 (N_14098,N_13477,N_12685);
nand U14099 (N_14099,N_13060,N_12051);
nand U14100 (N_14100,N_13472,N_13940);
nand U14101 (N_14101,N_12931,N_13292);
xnor U14102 (N_14102,N_12163,N_13244);
and U14103 (N_14103,N_12242,N_13503);
nand U14104 (N_14104,N_12582,N_12216);
or U14105 (N_14105,N_12540,N_13193);
nor U14106 (N_14106,N_13614,N_12062);
xnor U14107 (N_14107,N_12488,N_13392);
or U14108 (N_14108,N_12366,N_12431);
nand U14109 (N_14109,N_13385,N_13118);
and U14110 (N_14110,N_12905,N_13240);
and U14111 (N_14111,N_12642,N_13768);
and U14112 (N_14112,N_13157,N_13127);
and U14113 (N_14113,N_12236,N_12233);
nor U14114 (N_14114,N_13263,N_13996);
nor U14115 (N_14115,N_13063,N_12294);
nand U14116 (N_14116,N_12940,N_13110);
and U14117 (N_14117,N_13215,N_12367);
nor U14118 (N_14118,N_13467,N_13789);
or U14119 (N_14119,N_13530,N_13059);
nor U14120 (N_14120,N_13700,N_12608);
nor U14121 (N_14121,N_13753,N_13546);
nor U14122 (N_14122,N_13463,N_13608);
nor U14123 (N_14123,N_12086,N_13335);
nor U14124 (N_14124,N_13671,N_13459);
nor U14125 (N_14125,N_13670,N_12223);
nand U14126 (N_14126,N_13901,N_12342);
and U14127 (N_14127,N_13723,N_12584);
or U14128 (N_14128,N_12167,N_12283);
and U14129 (N_14129,N_13579,N_13469);
nor U14130 (N_14130,N_12977,N_13818);
nand U14131 (N_14131,N_13071,N_12320);
nor U14132 (N_14132,N_12831,N_13730);
or U14133 (N_14133,N_12442,N_13305);
and U14134 (N_14134,N_12889,N_13649);
xnor U14135 (N_14135,N_12997,N_13681);
xor U14136 (N_14136,N_12724,N_13647);
or U14137 (N_14137,N_13659,N_13878);
xor U14138 (N_14138,N_13867,N_13534);
xor U14139 (N_14139,N_13823,N_13912);
nor U14140 (N_14140,N_12813,N_12880);
nand U14141 (N_14141,N_13902,N_12956);
nand U14142 (N_14142,N_13086,N_12020);
and U14143 (N_14143,N_13316,N_13308);
nor U14144 (N_14144,N_12422,N_12145);
xnor U14145 (N_14145,N_12384,N_13114);
nor U14146 (N_14146,N_13771,N_13381);
nor U14147 (N_14147,N_13808,N_13238);
nand U14148 (N_14148,N_12463,N_13635);
or U14149 (N_14149,N_12066,N_12735);
nor U14150 (N_14150,N_13259,N_13920);
xor U14151 (N_14151,N_13065,N_13763);
nand U14152 (N_14152,N_12251,N_13553);
and U14153 (N_14153,N_12841,N_13970);
xor U14154 (N_14154,N_12617,N_12807);
or U14155 (N_14155,N_12784,N_13606);
nand U14156 (N_14156,N_12743,N_12015);
and U14157 (N_14157,N_13799,N_12810);
nand U14158 (N_14158,N_13264,N_13032);
nor U14159 (N_14159,N_12554,N_12411);
nand U14160 (N_14160,N_13642,N_13036);
xnor U14161 (N_14161,N_13347,N_12419);
nand U14162 (N_14162,N_13531,N_12502);
xnor U14163 (N_14163,N_12436,N_12227);
nand U14164 (N_14164,N_12183,N_12676);
and U14165 (N_14165,N_13070,N_12866);
nor U14166 (N_14166,N_12273,N_13372);
nand U14167 (N_14167,N_13946,N_13561);
and U14168 (N_14168,N_12244,N_12222);
or U14169 (N_14169,N_12691,N_13739);
nand U14170 (N_14170,N_12400,N_12974);
nand U14171 (N_14171,N_12846,N_12652);
and U14172 (N_14172,N_13034,N_12306);
xor U14173 (N_14173,N_12108,N_13234);
and U14174 (N_14174,N_13557,N_12493);
or U14175 (N_14175,N_12809,N_12501);
or U14176 (N_14176,N_12769,N_13171);
nor U14177 (N_14177,N_13005,N_13471);
xnor U14178 (N_14178,N_13786,N_13627);
nand U14179 (N_14179,N_13566,N_13054);
xnor U14180 (N_14180,N_12526,N_12395);
or U14181 (N_14181,N_13859,N_13377);
xor U14182 (N_14182,N_13022,N_12260);
xor U14183 (N_14183,N_12573,N_13968);
nor U14184 (N_14184,N_13665,N_13607);
and U14185 (N_14185,N_12068,N_13011);
nor U14186 (N_14186,N_12262,N_12137);
nor U14187 (N_14187,N_12847,N_12311);
xnor U14188 (N_14188,N_12088,N_13188);
nor U14189 (N_14189,N_12596,N_13260);
nor U14190 (N_14190,N_12146,N_13709);
nor U14191 (N_14191,N_13492,N_12105);
xor U14192 (N_14192,N_12742,N_12901);
xor U14193 (N_14193,N_12523,N_12178);
nand U14194 (N_14194,N_12172,N_12253);
xnor U14195 (N_14195,N_13149,N_13748);
nor U14196 (N_14196,N_13311,N_13417);
xnor U14197 (N_14197,N_13831,N_12927);
nand U14198 (N_14198,N_12275,N_13336);
nor U14199 (N_14199,N_12853,N_13214);
and U14200 (N_14200,N_13929,N_13778);
nor U14201 (N_14201,N_13782,N_13710);
nor U14202 (N_14202,N_12064,N_13053);
xor U14203 (N_14203,N_13488,N_13314);
nand U14204 (N_14204,N_12332,N_12291);
nand U14205 (N_14205,N_12918,N_13076);
or U14206 (N_14206,N_13258,N_13584);
and U14207 (N_14207,N_12597,N_12999);
nor U14208 (N_14208,N_13724,N_12412);
or U14209 (N_14209,N_13871,N_12628);
nor U14210 (N_14210,N_12374,N_12355);
nand U14211 (N_14211,N_13580,N_13605);
or U14212 (N_14212,N_13677,N_13618);
nor U14213 (N_14213,N_13565,N_12160);
xor U14214 (N_14214,N_13024,N_12469);
xnor U14215 (N_14215,N_12957,N_13325);
and U14216 (N_14216,N_12558,N_12996);
nor U14217 (N_14217,N_13398,N_13067);
nand U14218 (N_14218,N_13384,N_13082);
and U14219 (N_14219,N_13934,N_12498);
nor U14220 (N_14220,N_13266,N_13950);
nand U14221 (N_14221,N_12353,N_13880);
nand U14222 (N_14222,N_12705,N_13983);
nor U14223 (N_14223,N_12339,N_12000);
xor U14224 (N_14224,N_13543,N_13736);
and U14225 (N_14225,N_13456,N_13888);
xor U14226 (N_14226,N_12117,N_13493);
nor U14227 (N_14227,N_13802,N_13567);
nand U14228 (N_14228,N_13942,N_12755);
nor U14229 (N_14229,N_13840,N_13638);
nand U14230 (N_14230,N_12290,N_12677);
and U14231 (N_14231,N_13800,N_13887);
xnor U14232 (N_14232,N_12824,N_13705);
nor U14233 (N_14233,N_12465,N_13895);
xnor U14234 (N_14234,N_12696,N_13353);
and U14235 (N_14235,N_13897,N_12184);
nor U14236 (N_14236,N_13661,N_13976);
and U14237 (N_14237,N_13183,N_12878);
nor U14238 (N_14238,N_13781,N_12381);
nor U14239 (N_14239,N_12701,N_13174);
nand U14240 (N_14240,N_13466,N_13301);
or U14241 (N_14241,N_13866,N_13993);
nand U14242 (N_14242,N_13249,N_13847);
and U14243 (N_14243,N_13749,N_13702);
and U14244 (N_14244,N_12423,N_13675);
xnor U14245 (N_14245,N_13735,N_12961);
or U14246 (N_14246,N_13154,N_13703);
or U14247 (N_14247,N_13656,N_12153);
xnor U14248 (N_14248,N_13365,N_12891);
xor U14249 (N_14249,N_12008,N_13911);
nand U14250 (N_14250,N_12443,N_13882);
nor U14251 (N_14251,N_12710,N_13590);
nand U14252 (N_14252,N_13868,N_13109);
or U14253 (N_14253,N_13837,N_12844);
and U14254 (N_14254,N_13869,N_12874);
nor U14255 (N_14255,N_12588,N_12850);
xor U14256 (N_14256,N_12254,N_13073);
xor U14257 (N_14257,N_12832,N_12033);
or U14258 (N_14258,N_12272,N_12836);
xnor U14259 (N_14259,N_12544,N_12298);
nand U14260 (N_14260,N_12158,N_12027);
nor U14261 (N_14261,N_12224,N_12513);
and U14262 (N_14262,N_12461,N_13923);
nand U14263 (N_14263,N_12814,N_12933);
xnor U14264 (N_14264,N_13877,N_12792);
or U14265 (N_14265,N_12126,N_12886);
nor U14266 (N_14266,N_13512,N_13087);
nand U14267 (N_14267,N_13962,N_13204);
xor U14268 (N_14268,N_13207,N_13445);
or U14269 (N_14269,N_12586,N_12239);
or U14270 (N_14270,N_12645,N_12399);
and U14271 (N_14271,N_12972,N_13894);
nor U14272 (N_14272,N_12520,N_13187);
xnor U14273 (N_14273,N_12221,N_13502);
or U14274 (N_14274,N_13245,N_13226);
nand U14275 (N_14275,N_12271,N_13181);
xnor U14276 (N_14276,N_12130,N_13936);
xor U14277 (N_14277,N_13233,N_12220);
nor U14278 (N_14278,N_12169,N_12059);
and U14279 (N_14279,N_12585,N_13532);
nor U14280 (N_14280,N_13857,N_13354);
or U14281 (N_14281,N_12898,N_12672);
nor U14282 (N_14282,N_12711,N_12937);
or U14283 (N_14283,N_13439,N_13167);
xor U14284 (N_14284,N_12204,N_13641);
nand U14285 (N_14285,N_13138,N_12196);
nor U14286 (N_14286,N_12936,N_12613);
nand U14287 (N_14287,N_13835,N_13861);
or U14288 (N_14288,N_12714,N_12576);
and U14289 (N_14289,N_12806,N_13526);
nand U14290 (N_14290,N_13482,N_13284);
or U14291 (N_14291,N_12736,N_13914);
or U14292 (N_14292,N_13255,N_13538);
nor U14293 (N_14293,N_12919,N_12522);
and U14294 (N_14294,N_13192,N_12942);
nor U14295 (N_14295,N_13394,N_13939);
or U14296 (N_14296,N_13040,N_13003);
nand U14297 (N_14297,N_12912,N_13648);
and U14298 (N_14298,N_12528,N_12648);
xnor U14299 (N_14299,N_12777,N_12315);
nand U14300 (N_14300,N_13728,N_13657);
and U14301 (N_14301,N_13963,N_13960);
xnor U14302 (N_14302,N_12309,N_12869);
or U14303 (N_14303,N_12107,N_13809);
nor U14304 (N_14304,N_12418,N_13319);
nand U14305 (N_14305,N_13516,N_13402);
nor U14306 (N_14306,N_12098,N_13340);
nand U14307 (N_14307,N_13974,N_12349);
xor U14308 (N_14308,N_12719,N_12726);
or U14309 (N_14309,N_13345,N_13128);
nor U14310 (N_14310,N_12982,N_13297);
nand U14311 (N_14311,N_12096,N_13662);
and U14312 (N_14312,N_12829,N_12868);
xor U14313 (N_14313,N_12259,N_13568);
nand U14314 (N_14314,N_12804,N_13576);
and U14315 (N_14315,N_13805,N_12416);
nor U14316 (N_14316,N_12637,N_13632);
nor U14317 (N_14317,N_12965,N_12788);
and U14318 (N_14318,N_13272,N_12069);
nand U14319 (N_14319,N_12746,N_12848);
nand U14320 (N_14320,N_12211,N_12514);
xor U14321 (N_14321,N_13441,N_12634);
or U14322 (N_14322,N_12855,N_12344);
and U14323 (N_14323,N_12002,N_13825);
nor U14324 (N_14324,N_12174,N_13667);
nor U14325 (N_14325,N_12121,N_13037);
xnor U14326 (N_14326,N_12805,N_13883);
and U14327 (N_14327,N_13620,N_12671);
nand U14328 (N_14328,N_12885,N_13383);
nand U14329 (N_14329,N_12392,N_13628);
xor U14330 (N_14330,N_13932,N_12994);
nor U14331 (N_14331,N_13764,N_13380);
nand U14332 (N_14332,N_13720,N_12343);
and U14333 (N_14333,N_13913,N_12818);
nand U14334 (N_14334,N_13539,N_13158);
nand U14335 (N_14335,N_13884,N_13679);
or U14336 (N_14336,N_13995,N_12213);
nand U14337 (N_14337,N_12557,N_13563);
and U14338 (N_14338,N_12895,N_12626);
and U14339 (N_14339,N_12800,N_13746);
nor U14340 (N_14340,N_13241,N_13624);
and U14341 (N_14341,N_12383,N_12529);
xor U14342 (N_14342,N_12241,N_12718);
or U14343 (N_14343,N_13601,N_12960);
nor U14344 (N_14344,N_13672,N_13458);
nand U14345 (N_14345,N_13804,N_12669);
or U14346 (N_14346,N_13162,N_13613);
and U14347 (N_14347,N_12285,N_13682);
xnor U14348 (N_14348,N_13285,N_13905);
or U14349 (N_14349,N_12808,N_12427);
or U14350 (N_14350,N_12641,N_12281);
xor U14351 (N_14351,N_12689,N_12097);
or U14352 (N_14352,N_13023,N_13761);
nand U14353 (N_14353,N_12629,N_12838);
or U14354 (N_14354,N_13270,N_12012);
nand U14355 (N_14355,N_12976,N_13012);
nand U14356 (N_14356,N_13421,N_13784);
and U14357 (N_14357,N_13190,N_12908);
and U14358 (N_14358,N_13455,N_13433);
nand U14359 (N_14359,N_13548,N_12053);
nand U14360 (N_14360,N_12226,N_13414);
xor U14361 (N_14361,N_13688,N_13367);
and U14362 (N_14362,N_13569,N_12058);
nor U14363 (N_14363,N_12575,N_13437);
xnor U14364 (N_14364,N_12135,N_12894);
nand U14365 (N_14365,N_13115,N_13134);
nand U14366 (N_14366,N_12872,N_13166);
nor U14367 (N_14367,N_13701,N_12754);
nand U14368 (N_14368,N_12845,N_12700);
nor U14369 (N_14369,N_13296,N_13824);
and U14370 (N_14370,N_13302,N_13765);
or U14371 (N_14371,N_12560,N_13592);
or U14372 (N_14372,N_12029,N_13168);
nand U14373 (N_14373,N_13161,N_12858);
xor U14374 (N_14374,N_13273,N_12923);
xor U14375 (N_14375,N_12904,N_13219);
nor U14376 (N_14376,N_12005,N_13051);
xor U14377 (N_14377,N_13393,N_13132);
or U14378 (N_14378,N_13973,N_13315);
nor U14379 (N_14379,N_13714,N_13039);
xor U14380 (N_14380,N_12111,N_12625);
nor U14381 (N_14381,N_13949,N_12080);
and U14382 (N_14382,N_12425,N_13699);
and U14383 (N_14383,N_12545,N_13961);
and U14384 (N_14384,N_12317,N_13860);
or U14385 (N_14385,N_13630,N_13743);
nor U14386 (N_14386,N_12310,N_12028);
nand U14387 (N_14387,N_12490,N_12466);
or U14388 (N_14388,N_12313,N_13574);
or U14389 (N_14389,N_12352,N_12635);
nand U14390 (N_14390,N_13422,N_13103);
nand U14391 (N_14391,N_13798,N_12304);
nor U14392 (N_14392,N_13428,N_13170);
nand U14393 (N_14393,N_13031,N_13283);
xor U14394 (N_14394,N_13403,N_13035);
nand U14395 (N_14395,N_12506,N_13599);
nand U14396 (N_14396,N_13577,N_13379);
nor U14397 (N_14397,N_12969,N_13814);
xor U14398 (N_14398,N_13843,N_12319);
or U14399 (N_14399,N_13838,N_13797);
or U14400 (N_14400,N_12363,N_13136);
nand U14401 (N_14401,N_13986,N_12483);
nand U14402 (N_14402,N_12879,N_12667);
and U14403 (N_14403,N_12562,N_12083);
nand U14404 (N_14404,N_12843,N_13387);
and U14405 (N_14405,N_13903,N_13304);
nor U14406 (N_14406,N_13678,N_12067);
or U14407 (N_14407,N_13523,N_12893);
xor U14408 (N_14408,N_13411,N_12766);
xor U14409 (N_14409,N_12569,N_13077);
xnor U14410 (N_14410,N_12668,N_12039);
nand U14411 (N_14411,N_12738,N_13645);
nand U14412 (N_14412,N_13890,N_13680);
nor U14413 (N_14413,N_13788,N_13858);
xor U14414 (N_14414,N_12165,N_12600);
nor U14415 (N_14415,N_13211,N_13388);
xnor U14416 (N_14416,N_12968,N_13081);
xor U14417 (N_14417,N_13435,N_13529);
or U14418 (N_14418,N_13937,N_13364);
xnor U14419 (N_14419,N_12308,N_13487);
or U14420 (N_14420,N_13328,N_12408);
nor U14421 (N_14421,N_13998,N_13176);
nor U14422 (N_14422,N_12662,N_12900);
nor U14423 (N_14423,N_12857,N_13470);
nand U14424 (N_14424,N_12661,N_12394);
or U14425 (N_14425,N_12692,N_12162);
nor U14426 (N_14426,N_13683,N_13652);
and U14427 (N_14427,N_13898,N_12179);
and U14428 (N_14428,N_12152,N_12303);
nor U14429 (N_14429,N_12521,N_13107);
nand U14430 (N_14430,N_12606,N_12257);
and U14431 (N_14431,N_12048,N_13164);
nand U14432 (N_14432,N_13098,N_13275);
or U14433 (N_14433,N_12471,N_12420);
and U14434 (N_14434,N_12124,N_12690);
xnor U14435 (N_14435,N_13371,N_12118);
xnor U14436 (N_14436,N_12987,N_13536);
nand U14437 (N_14437,N_12365,N_12728);
or U14438 (N_14438,N_13346,N_13750);
and U14439 (N_14439,N_12820,N_12896);
nand U14440 (N_14440,N_13555,N_12757);
xnor U14441 (N_14441,N_12433,N_13817);
nor U14442 (N_14442,N_13148,N_12438);
nand U14443 (N_14443,N_13389,N_13990);
xnor U14444 (N_14444,N_12407,N_12357);
xor U14445 (N_14445,N_12147,N_12435);
xor U14446 (N_14446,N_12234,N_12269);
nand U14447 (N_14447,N_13633,N_12607);
nand U14448 (N_14448,N_12712,N_12734);
or U14449 (N_14449,N_13737,N_13423);
and U14450 (N_14450,N_12003,N_12300);
xor U14451 (N_14451,N_12486,N_13698);
nand U14452 (N_14452,N_12535,N_12538);
nor U14453 (N_14453,N_12713,N_13832);
nor U14454 (N_14454,N_12006,N_13408);
or U14455 (N_14455,N_12413,N_13089);
or U14456 (N_14456,N_13074,N_12534);
xor U14457 (N_14457,N_13007,N_12270);
nor U14458 (N_14458,N_12358,N_13664);
xor U14459 (N_14459,N_12980,N_13794);
xor U14460 (N_14460,N_13046,N_13331);
nor U14461 (N_14461,N_12881,N_12150);
nor U14462 (N_14462,N_12913,N_13291);
xnor U14463 (N_14463,N_13406,N_12761);
or U14464 (N_14464,N_12496,N_12289);
or U14465 (N_14465,N_13609,N_12322);
and U14466 (N_14466,N_13362,N_13775);
xnor U14467 (N_14467,N_13879,N_13615);
xnor U14468 (N_14468,N_13376,N_13265);
nand U14469 (N_14469,N_13904,N_13208);
xnor U14470 (N_14470,N_12106,N_12049);
nand U14471 (N_14471,N_12740,N_12346);
xor U14472 (N_14472,N_13791,N_12509);
nand U14473 (N_14473,N_13113,N_13839);
and U14474 (N_14474,N_13729,N_13189);
nand U14475 (N_14475,N_13959,N_12409);
nand U14476 (N_14476,N_12594,N_12375);
or U14477 (N_14477,N_13842,N_12212);
xor U14478 (N_14478,N_13055,N_13713);
or U14479 (N_14479,N_13228,N_13747);
nor U14480 (N_14480,N_13111,N_12731);
or U14481 (N_14481,N_12041,N_12018);
and U14482 (N_14482,N_12593,N_12084);
or U14483 (N_14483,N_13257,N_12890);
or U14484 (N_14484,N_12636,N_12477);
and U14485 (N_14485,N_12524,N_13390);
nor U14486 (N_14486,N_12149,N_13009);
nand U14487 (N_14487,N_13593,N_12359);
nand U14488 (N_14488,N_12612,N_13145);
and U14489 (N_14489,N_12386,N_12099);
xor U14490 (N_14490,N_12870,N_13066);
and U14491 (N_14491,N_13150,N_13821);
or U14492 (N_14492,N_12786,N_12430);
or U14493 (N_14493,N_13738,N_13725);
xor U14494 (N_14494,N_12610,N_12100);
and U14495 (N_14495,N_13436,N_13438);
or U14496 (N_14496,N_12016,N_12899);
xor U14497 (N_14497,N_13008,N_13570);
nor U14498 (N_14498,N_13827,N_13220);
nor U14499 (N_14499,N_12935,N_12389);
nand U14500 (N_14500,N_12708,N_13126);
nand U14501 (N_14501,N_13591,N_12771);
and U14502 (N_14502,N_13057,N_12492);
or U14503 (N_14503,N_12243,N_13992);
xor U14504 (N_14504,N_12052,N_12739);
nand U14505 (N_14505,N_12914,N_13987);
nand U14506 (N_14506,N_12715,N_12287);
and U14507 (N_14507,N_13357,N_12760);
nand U14508 (N_14508,N_12811,N_12385);
and U14509 (N_14509,N_12268,N_13595);
or U14510 (N_14510,N_12191,N_12673);
xnor U14511 (N_14511,N_13303,N_13716);
nand U14512 (N_14512,N_13787,N_13924);
nand U14513 (N_14513,N_13830,N_13489);
nor U14514 (N_14514,N_12219,N_13416);
xnor U14515 (N_14515,N_12653,N_13359);
xnor U14516 (N_14516,N_13217,N_13199);
nor U14517 (N_14517,N_13142,N_12391);
nand U14518 (N_14518,N_13102,N_12331);
and U14519 (N_14519,N_13571,N_13852);
nor U14520 (N_14520,N_12414,N_12729);
nand U14521 (N_14521,N_12744,N_12063);
nand U14522 (N_14522,N_13015,N_12799);
or U14523 (N_14523,N_12417,N_13919);
nand U14524 (N_14524,N_12134,N_13465);
or U14525 (N_14525,N_13513,N_12282);
or U14526 (N_14526,N_13218,N_13694);
nand U14527 (N_14527,N_13718,N_12440);
nand U14528 (N_14528,N_13342,N_13140);
or U14529 (N_14529,N_13200,N_13967);
nand U14530 (N_14530,N_12093,N_13461);
or U14531 (N_14531,N_12074,N_12902);
nor U14532 (N_14532,N_12482,N_12132);
nand U14533 (N_14533,N_13091,N_13953);
and U14534 (N_14534,N_12410,N_12201);
or U14535 (N_14535,N_12450,N_13815);
xnor U14536 (N_14536,N_13072,N_13121);
and U14537 (N_14537,N_12616,N_13318);
xnor U14538 (N_14538,N_12817,N_13783);
xnor U14539 (N_14539,N_13813,N_12656);
or U14540 (N_14540,N_12852,N_13223);
and U14541 (N_14541,N_13322,N_12568);
or U14542 (N_14542,N_13770,N_13262);
nor U14543 (N_14543,N_13779,N_12340);
nand U14544 (N_14544,N_13155,N_13732);
and U14545 (N_14545,N_12603,N_12565);
xnor U14546 (N_14546,N_12487,N_13224);
xnor U14547 (N_14547,N_13252,N_13287);
nor U14548 (N_14548,N_12581,N_12518);
or U14549 (N_14549,N_12209,N_12702);
xor U14550 (N_14550,N_12406,N_13727);
nand U14551 (N_14551,N_13988,N_12541);
nand U14552 (N_14552,N_12840,N_12833);
nand U14553 (N_14553,N_12341,N_13178);
nand U14554 (N_14554,N_12156,N_13623);
and U14555 (N_14555,N_13124,N_13125);
nand U14556 (N_14556,N_12741,N_13634);
or U14557 (N_14557,N_12706,N_13350);
and U14558 (N_14558,N_12622,N_13062);
and U14559 (N_14559,N_12141,N_12834);
nor U14560 (N_14560,N_12403,N_12054);
nor U14561 (N_14561,N_13129,N_13760);
or U14562 (N_14562,N_12816,N_13399);
and U14563 (N_14563,N_13027,N_12659);
nor U14564 (N_14564,N_12505,N_13462);
nor U14565 (N_14565,N_12032,N_13310);
nor U14566 (N_14566,N_12305,N_13651);
and U14567 (N_14567,N_13222,N_13478);
nor U14568 (N_14568,N_13141,N_12372);
nand U14569 (N_14569,N_13330,N_12330);
or U14570 (N_14570,N_12085,N_12265);
and U14571 (N_14571,N_12579,N_13910);
nor U14572 (N_14572,N_12632,N_13216);
and U14573 (N_14573,N_13957,N_13049);
or U14574 (N_14574,N_13772,N_13741);
nand U14575 (N_14575,N_13344,N_12113);
nor U14576 (N_14576,N_12369,N_13527);
or U14577 (N_14577,N_12217,N_12021);
nor U14578 (N_14578,N_13999,N_13480);
nor U14579 (N_14579,N_12324,N_12770);
nor U14580 (N_14580,N_13420,N_12765);
nand U14581 (N_14581,N_13836,N_12922);
and U14582 (N_14582,N_13021,N_13689);
and U14583 (N_14583,N_12601,N_13191);
nand U14584 (N_14584,N_13498,N_12046);
nor U14585 (N_14585,N_12546,N_13185);
or U14586 (N_14586,N_13985,N_12947);
nand U14587 (N_14587,N_13510,N_13617);
or U14588 (N_14588,N_12278,N_12464);
xor U14589 (N_14589,N_12380,N_13045);
xnor U14590 (N_14590,N_13368,N_12614);
nand U14591 (N_14591,N_12362,N_12963);
xor U14592 (N_14592,N_12314,N_13604);
and U14593 (N_14593,N_13629,N_13550);
nand U14594 (N_14594,N_13893,N_12424);
or U14595 (N_14595,N_13153,N_12447);
or U14596 (N_14596,N_13542,N_13766);
xor U14597 (N_14597,N_13375,N_13490);
xnor U14598 (N_14598,N_12687,N_13117);
nor U14599 (N_14599,N_13947,N_12795);
or U14600 (N_14600,N_13581,N_13221);
nor U14601 (N_14601,N_13558,N_12467);
and U14602 (N_14602,N_12964,N_12680);
nor U14603 (N_14603,N_12655,N_12650);
nor U14604 (N_14604,N_12082,N_13378);
xor U14605 (N_14605,N_12897,N_13281);
nand U14606 (N_14606,N_13889,N_13885);
and U14607 (N_14607,N_13686,N_13785);
xor U14608 (N_14608,N_12884,N_12697);
or U14609 (N_14609,N_12664,N_13979);
and U14610 (N_14610,N_12698,N_12725);
xnor U14611 (N_14611,N_13762,N_13180);
xnor U14612 (N_14612,N_13453,N_12168);
nor U14613 (N_14613,N_13139,N_12883);
nor U14614 (N_14614,N_12875,N_12876);
or U14615 (N_14615,N_12004,N_12536);
or U14616 (N_14616,N_12081,N_12301);
nand U14617 (N_14617,N_13324,N_12042);
and U14618 (N_14618,N_13742,N_13246);
xnor U14619 (N_14619,N_12188,N_12941);
and U14620 (N_14620,N_13906,N_12945);
nand U14621 (N_14621,N_13018,N_12077);
xor U14622 (N_14622,N_13300,N_13415);
nor U14623 (N_14623,N_13653,N_12489);
and U14624 (N_14624,N_13807,N_13409);
nand U14625 (N_14625,N_13712,N_13425);
or U14626 (N_14626,N_12851,N_13454);
xor U14627 (N_14627,N_13780,N_12499);
nor U14628 (N_14628,N_13276,N_12388);
nor U14629 (N_14629,N_13294,N_13099);
and U14630 (N_14630,N_12480,N_12703);
xor U14631 (N_14631,N_13019,N_12133);
and U14632 (N_14632,N_12102,N_12232);
nor U14633 (N_14633,N_13485,N_13684);
xor U14634 (N_14634,N_12356,N_12390);
and U14635 (N_14635,N_13704,N_13873);
or U14636 (N_14636,N_12325,N_13143);
xor U14637 (N_14637,N_13267,N_12998);
and U14638 (N_14638,N_12583,N_12556);
nor U14639 (N_14639,N_13135,N_12258);
and U14640 (N_14640,N_13594,N_13907);
nand U14641 (N_14641,N_12873,N_12155);
and U14642 (N_14642,N_13944,N_13419);
or U14643 (N_14643,N_12917,N_12542);
nand U14644 (N_14644,N_13846,N_12139);
and U14645 (N_14645,N_13144,N_13323);
nor U14646 (N_14646,N_12460,N_12979);
or U14647 (N_14647,N_13120,N_13080);
nor U14648 (N_14648,N_13881,N_12136);
and U14649 (N_14649,N_12240,N_13505);
nor U14650 (N_14650,N_13978,N_12519);
nand U14651 (N_14651,N_12686,N_12646);
xor U14652 (N_14652,N_12307,N_12318);
xnor U14653 (N_14653,N_13733,N_13744);
and U14654 (N_14654,N_12589,N_12449);
xor U14655 (N_14655,N_12681,N_13501);
and U14656 (N_14656,N_13551,N_12247);
or U14657 (N_14657,N_12621,N_13247);
xor U14658 (N_14658,N_12504,N_13603);
xnor U14659 (N_14659,N_13552,N_12620);
nor U14660 (N_14660,N_12245,N_12928);
xnor U14661 (N_14661,N_12148,N_12071);
nand U14662 (N_14662,N_12670,N_13464);
nand U14663 (N_14663,N_12733,N_12772);
or U14664 (N_14664,N_13583,N_13196);
or U14665 (N_14665,N_13639,N_13268);
or U14666 (N_14666,N_13351,N_12570);
or U14667 (N_14667,N_13774,N_13119);
or U14668 (N_14668,N_13596,N_13663);
xor U14669 (N_14669,N_13006,N_13042);
nor U14670 (N_14670,N_12827,N_12992);
xor U14671 (N_14671,N_13075,N_13016);
or U14672 (N_14672,N_12571,N_12142);
nor U14673 (N_14673,N_12337,N_12758);
and U14674 (N_14674,N_13202,N_12293);
xnor U14675 (N_14675,N_12302,N_12474);
nand U14676 (N_14676,N_13468,N_12929);
nor U14677 (N_14677,N_13290,N_12654);
xnor U14678 (N_14678,N_12040,N_13396);
and U14679 (N_14679,N_13955,N_12782);
or U14680 (N_14680,N_12368,N_12727);
nor U14681 (N_14681,N_12351,N_13239);
nand U14682 (N_14682,N_12911,N_13777);
and U14683 (N_14683,N_13360,N_12122);
and U14684 (N_14684,N_12345,N_13231);
nor U14685 (N_14685,N_12674,N_12180);
and U14686 (N_14686,N_13544,N_12651);
xor U14687 (N_14687,N_12297,N_13112);
nor U14688 (N_14688,N_13000,N_13850);
and U14689 (N_14689,N_13235,N_12246);
nor U14690 (N_14690,N_13405,N_13452);
nand U14691 (N_14691,N_12815,N_13511);
nor U14692 (N_14692,N_13844,N_12475);
and U14693 (N_14693,N_13954,N_12658);
nand U14694 (N_14694,N_12615,N_13674);
and U14695 (N_14695,N_12854,N_12468);
or U14696 (N_14696,N_13636,N_13524);
and U14697 (N_14697,N_12903,N_13321);
nand U14698 (N_14698,N_12214,N_12288);
or U14699 (N_14699,N_12682,N_13093);
nand U14700 (N_14700,N_12373,N_12025);
nand U14701 (N_14701,N_12494,N_13500);
or U14702 (N_14702,N_13209,N_12822);
nor U14703 (N_14703,N_12456,N_13010);
or U14704 (N_14704,N_12946,N_12458);
or U14705 (N_14705,N_12208,N_13163);
or U14706 (N_14706,N_12675,N_13965);
nand U14707 (N_14707,N_12078,N_13095);
xnor U14708 (N_14708,N_12906,N_12428);
or U14709 (N_14709,N_12190,N_12377);
and U14710 (N_14710,N_13026,N_12683);
xor U14711 (N_14711,N_12014,N_13449);
xor U14712 (N_14712,N_12237,N_13792);
nand U14713 (N_14713,N_13366,N_12533);
or U14714 (N_14714,N_13448,N_13598);
nand U14715 (N_14715,N_13058,N_13845);
nor U14716 (N_14716,N_13755,N_12228);
and U14717 (N_14717,N_12116,N_12550);
nor U14718 (N_14718,N_13926,N_12038);
xor U14719 (N_14719,N_13151,N_13280);
nor U14720 (N_14720,N_13927,N_12405);
or U14721 (N_14721,N_13622,N_13876);
nor U14722 (N_14722,N_12531,N_12206);
xor U14723 (N_14723,N_13205,N_13773);
nor U14724 (N_14724,N_13497,N_13044);
xor U14725 (N_14725,N_12170,N_13326);
or U14726 (N_14726,N_12001,N_12115);
xnor U14727 (N_14727,N_12455,N_12261);
xor U14728 (N_14728,N_13427,N_12695);
or U14729 (N_14729,N_12164,N_12763);
and U14730 (N_14730,N_13697,N_12479);
or U14731 (N_14731,N_13690,N_13943);
nor U14732 (N_14732,N_13374,N_12055);
nor U14733 (N_14733,N_12250,N_13654);
nand U14734 (N_14734,N_12207,N_12835);
nand U14735 (N_14735,N_12448,N_12907);
and U14736 (N_14736,N_12087,N_12549);
xnor U14737 (N_14737,N_13486,N_13855);
nor U14738 (N_14738,N_12704,N_13754);
xnor U14739 (N_14739,N_12796,N_13631);
xor U14740 (N_14740,N_13952,N_12707);
nor U14741 (N_14741,N_12379,N_13043);
nor U14742 (N_14742,N_13289,N_12453);
xnor U14743 (N_14743,N_13640,N_12256);
nand U14744 (N_14744,N_12348,N_13309);
and U14745 (N_14745,N_13556,N_12605);
or U14746 (N_14746,N_13506,N_13474);
and U14747 (N_14747,N_12948,N_12747);
and U14748 (N_14748,N_12773,N_13122);
nand U14749 (N_14749,N_13041,N_13863);
or U14750 (N_14750,N_13722,N_12267);
nand U14751 (N_14751,N_13225,N_13313);
and U14752 (N_14752,N_13806,N_12491);
and U14753 (N_14753,N_13793,N_12732);
or U14754 (N_14754,N_12017,N_13105);
and U14755 (N_14755,N_13951,N_12023);
or U14756 (N_14756,N_12166,N_13562);
nor U14757 (N_14757,N_13900,N_13286);
and U14758 (N_14758,N_13495,N_12326);
and U14759 (N_14759,N_13801,N_12181);
and U14760 (N_14760,N_12970,N_12112);
nand U14761 (N_14761,N_12347,N_12452);
nor U14762 (N_14762,N_13430,N_12507);
and U14763 (N_14763,N_13404,N_12192);
xor U14764 (N_14764,N_12229,N_13182);
or U14765 (N_14765,N_12316,N_13097);
nand U14766 (N_14766,N_12175,N_12129);
and U14767 (N_14767,N_12749,N_13068);
nor U14768 (N_14768,N_12312,N_13711);
or U14769 (N_14769,N_12079,N_12151);
nand U14770 (N_14770,N_12218,N_12473);
and U14771 (N_14771,N_13916,N_13612);
xor U14772 (N_14772,N_12756,N_12354);
nor U14773 (N_14773,N_13745,N_13756);
and U14774 (N_14774,N_12920,N_13997);
nor U14775 (N_14775,N_13769,N_13094);
or U14776 (N_14776,N_12120,N_12114);
or U14777 (N_14777,N_12720,N_12839);
xnor U14778 (N_14778,N_12790,N_12860);
nand U14779 (N_14779,N_12591,N_13757);
nand U14780 (N_14780,N_12193,N_13586);
xor U14781 (N_14781,N_12333,N_13734);
nor U14782 (N_14782,N_13412,N_13841);
or U14783 (N_14783,N_12338,N_12991);
xnor U14784 (N_14784,N_13029,N_12500);
xnor U14785 (N_14785,N_12031,N_13600);
nor U14786 (N_14786,N_13509,N_12775);
or U14787 (N_14787,N_13810,N_12396);
or U14788 (N_14788,N_12572,N_13611);
nor U14789 (N_14789,N_12609,N_13337);
or U14790 (N_14790,N_12864,N_12978);
or U14791 (N_14791,N_13349,N_13540);
or U14792 (N_14792,N_12187,N_13812);
or U14793 (N_14793,N_12983,N_13050);
xnor U14794 (N_14794,N_13206,N_13001);
nand U14795 (N_14795,N_13875,N_12802);
nor U14796 (N_14796,N_13460,N_12202);
xnor U14797 (N_14797,N_12197,N_12026);
nor U14798 (N_14798,N_13507,N_12437);
nand U14799 (N_14799,N_12971,N_13650);
nand U14800 (N_14800,N_12451,N_13541);
xor U14801 (N_14801,N_12439,N_12587);
nor U14802 (N_14802,N_12862,N_13274);
xor U14803 (N_14803,N_12279,N_12953);
and U14804 (N_14804,N_13717,N_13090);
or U14805 (N_14805,N_12402,N_12274);
nand U14806 (N_14806,N_12959,N_12826);
xor U14807 (N_14807,N_13587,N_12819);
or U14808 (N_14808,N_12909,N_13184);
nor U14809 (N_14809,N_13407,N_13014);
or U14810 (N_14810,N_13707,N_13828);
and U14811 (N_14811,N_13515,N_12962);
or U14812 (N_14812,N_12401,N_13833);
nor U14813 (N_14813,N_12791,N_13494);
and U14814 (N_14814,N_12619,N_12631);
xor U14815 (N_14815,N_13589,N_12037);
and U14816 (N_14816,N_12644,N_13826);
nor U14817 (N_14817,N_12200,N_13928);
nand U14818 (N_14818,N_13776,N_13339);
nor U14819 (N_14819,N_12793,N_12958);
nor U14820 (N_14820,N_13849,N_12195);
nor U14821 (N_14821,N_12013,N_12618);
xnor U14822 (N_14822,N_13496,N_12350);
and U14823 (N_14823,N_13343,N_13575);
nand U14824 (N_14824,N_13250,N_12462);
nor U14825 (N_14825,N_12842,N_12552);
and U14826 (N_14826,N_12555,N_12144);
and U14827 (N_14827,N_12415,N_13854);
or U14828 (N_14828,N_13938,N_13796);
xor U14829 (N_14829,N_12566,N_12019);
or U14830 (N_14830,N_13242,N_13108);
nand U14831 (N_14831,N_13253,N_12530);
nand U14832 (N_14832,N_13248,N_12299);
nand U14833 (N_14833,N_13856,N_13002);
nand U14834 (N_14834,N_12717,N_13038);
nand U14835 (N_14835,N_12943,N_13358);
or U14836 (N_14836,N_13504,N_12966);
and U14837 (N_14837,N_13271,N_12559);
nand U14838 (N_14838,N_13767,N_12837);
or U14839 (N_14839,N_12789,N_13982);
and U14840 (N_14840,N_12426,N_12665);
xnor U14841 (N_14841,N_13232,N_12990);
and U14842 (N_14842,N_12459,N_13312);
or U14843 (N_14843,N_13545,N_12981);
nand U14844 (N_14844,N_13395,N_12863);
nand U14845 (N_14845,N_12774,N_13169);
nand U14846 (N_14846,N_13450,N_13064);
and U14847 (N_14847,N_13522,N_13621);
xor U14848 (N_14848,N_12444,N_12511);
or U14849 (N_14849,N_12445,N_13227);
nor U14850 (N_14850,N_13256,N_12238);
or U14851 (N_14851,N_12926,N_12578);
xnor U14852 (N_14852,N_13341,N_13278);
and U14853 (N_14853,N_13872,N_12295);
or U14854 (N_14854,N_12119,N_12361);
nor U14855 (N_14855,N_13886,N_12421);
nand U14856 (N_14856,N_13691,N_12688);
and U14857 (N_14857,N_13028,N_13332);
or U14858 (N_14858,N_12050,N_13483);
nand U14859 (N_14859,N_13282,N_13564);
nor U14860 (N_14860,N_12882,N_13975);
or U14861 (N_14861,N_13085,N_13816);
and U14862 (N_14862,N_12623,N_13829);
or U14863 (N_14863,N_12666,N_12532);
and U14864 (N_14864,N_13434,N_13921);
and U14865 (N_14865,N_12089,N_12639);
and U14866 (N_14866,N_12094,N_12292);
xnor U14867 (N_14867,N_12161,N_13457);
or U14868 (N_14868,N_12539,N_13695);
or U14869 (N_14869,N_12798,N_12230);
and U14870 (N_14870,N_13473,N_13865);
xor U14871 (N_14871,N_13931,N_12185);
xnor U14872 (N_14872,N_12781,N_12949);
or U14873 (N_14873,N_13626,N_12434);
and U14874 (N_14874,N_13537,N_12095);
xor U14875 (N_14875,N_12159,N_12924);
nor U14876 (N_14876,N_12189,N_13514);
nor U14877 (N_14877,N_13048,N_13201);
and U14878 (N_14878,N_12334,N_12252);
xnor U14879 (N_14879,N_13549,N_13989);
or U14880 (N_14880,N_13751,N_12785);
and U14881 (N_14881,N_12143,N_13451);
and U14882 (N_14882,N_13172,N_13198);
or U14883 (N_14883,N_12235,N_12481);
nor U14884 (N_14884,N_13382,N_13386);
nand U14885 (N_14885,N_13853,N_12986);
nand U14886 (N_14886,N_12010,N_12024);
nor U14887 (N_14887,N_12176,N_12723);
or U14888 (N_14888,N_12123,N_12787);
or U14889 (N_14889,N_12060,N_13017);
nor U14890 (N_14890,N_13588,N_13669);
xor U14891 (N_14891,N_12022,N_12611);
nand U14892 (N_14892,N_12091,N_12780);
or U14893 (N_14893,N_12633,N_12101);
nand U14894 (N_14894,N_13554,N_13899);
and U14895 (N_14895,N_12011,N_13306);
or U14896 (N_14896,N_13069,N_12182);
or U14897 (N_14897,N_12194,N_13644);
xor U14898 (N_14898,N_12393,N_12856);
xor U14899 (N_14899,N_12072,N_13848);
or U14900 (N_14900,N_13361,N_13945);
and U14901 (N_14901,N_13528,N_12794);
xnor U14902 (N_14902,N_12915,N_13355);
and U14903 (N_14903,N_12849,N_13892);
or U14904 (N_14904,N_13476,N_12215);
and U14905 (N_14905,N_12925,N_13874);
nand U14906 (N_14906,N_12404,N_13484);
and U14907 (N_14907,N_12988,N_13547);
nand U14908 (N_14908,N_13811,N_13508);
or U14909 (N_14909,N_13991,N_12516);
nand U14910 (N_14910,N_12993,N_12580);
or U14911 (N_14911,N_12745,N_12249);
or U14912 (N_14912,N_13401,N_12954);
nor U14913 (N_14913,N_12828,N_13525);
and U14914 (N_14914,N_12382,N_12598);
xor U14915 (N_14915,N_13083,N_13203);
or U14916 (N_14916,N_12138,N_12984);
and U14917 (N_14917,N_13715,N_12778);
nand U14918 (N_14918,N_13933,N_13413);
xor U14919 (N_14919,N_12679,N_12035);
xnor U14920 (N_14920,N_13941,N_12547);
nand U14921 (N_14921,N_12934,N_12034);
nand U14922 (N_14922,N_12779,N_13925);
nor U14923 (N_14923,N_13972,N_13676);
and U14924 (N_14924,N_13687,N_13731);
xor U14925 (N_14925,N_12985,N_12721);
nor U14926 (N_14926,N_13499,N_12748);
and U14927 (N_14927,N_12371,N_12722);
and U14928 (N_14928,N_13410,N_13254);
or U14929 (N_14929,N_13004,N_12378);
xnor U14930 (N_14930,N_12967,N_13079);
and U14931 (N_14931,N_12508,N_12199);
xnor U14932 (N_14932,N_13298,N_13740);
nor U14933 (N_14933,N_12951,N_12446);
nand U14934 (N_14934,N_12045,N_13706);
nor U14935 (N_14935,N_13909,N_12296);
and U14936 (N_14936,N_12577,N_13173);
nand U14937 (N_14937,N_12429,N_12861);
nor U14938 (N_14938,N_12859,N_13123);
xnor U14939 (N_14939,N_13056,N_13047);
nor U14940 (N_14940,N_12767,N_12660);
xor U14941 (N_14941,N_12205,N_13106);
nor U14942 (N_14942,N_12177,N_13971);
nand U14943 (N_14943,N_12678,N_12865);
nand U14944 (N_14944,N_13862,N_13317);
or U14945 (N_14945,N_13165,N_13646);
nor U14946 (N_14946,N_13908,N_12812);
and U14947 (N_14947,N_13896,N_12649);
or U14948 (N_14948,N_13685,N_13759);
and U14949 (N_14949,N_13418,N_12955);
nor U14950 (N_14950,N_13917,N_12716);
and U14951 (N_14951,N_13610,N_13025);
xor U14952 (N_14952,N_13033,N_12398);
or U14953 (N_14953,N_12693,N_12551);
or U14954 (N_14954,N_13719,N_12950);
nor U14955 (N_14955,N_12517,N_12764);
nand U14956 (N_14956,N_12553,N_13236);
or U14957 (N_14957,N_12485,N_12995);
nand U14958 (N_14958,N_13432,N_13966);
nor U14959 (N_14959,N_13625,N_12830);
and U14960 (N_14960,N_12476,N_12376);
and U14961 (N_14961,N_12768,N_12563);
nand U14962 (N_14962,N_13369,N_12989);
nor U14963 (N_14963,N_13237,N_13116);
nand U14964 (N_14964,N_12776,N_12110);
nand U14965 (N_14965,N_12952,N_13602);
xor U14966 (N_14966,N_12154,N_13230);
or U14967 (N_14967,N_13299,N_13370);
and U14968 (N_14968,N_13175,N_12248);
nor U14969 (N_14969,N_13479,N_12255);
or U14970 (N_14970,N_12009,N_13518);
or U14971 (N_14971,N_13790,N_13582);
or U14972 (N_14972,N_12595,N_13212);
or U14973 (N_14973,N_13637,N_13096);
xor U14974 (N_14974,N_12892,N_13442);
nor U14975 (N_14975,N_13356,N_12643);
and U14976 (N_14976,N_12472,N_12657);
xor U14977 (N_14977,N_12699,N_12036);
and U14978 (N_14978,N_12263,N_12007);
nand U14979 (N_14979,N_13977,N_13424);
xor U14980 (N_14980,N_12056,N_12821);
nor U14981 (N_14981,N_13101,N_12210);
xor U14982 (N_14982,N_12877,N_12599);
nand U14983 (N_14983,N_12537,N_12975);
xnor U14984 (N_14984,N_13666,N_12109);
and U14985 (N_14985,N_13619,N_12916);
nor U14986 (N_14986,N_13307,N_12125);
or U14987 (N_14987,N_13643,N_13475);
and U14988 (N_14988,N_12061,N_12323);
xnor U14989 (N_14989,N_12103,N_13431);
nand U14990 (N_14990,N_13819,N_13658);
nand U14991 (N_14991,N_13131,N_13616);
and U14992 (N_14992,N_13197,N_13803);
and U14993 (N_14993,N_12057,N_13981);
nor U14994 (N_14994,N_13391,N_12938);
or U14995 (N_14995,N_13329,N_12043);
nand U14996 (N_14996,N_13320,N_13517);
nand U14997 (N_14997,N_13535,N_12640);
and U14998 (N_14998,N_13572,N_12910);
nor U14999 (N_14999,N_13288,N_12186);
and U15000 (N_15000,N_12646,N_13217);
xor U15001 (N_15001,N_13635,N_12900);
nand U15002 (N_15002,N_12786,N_13692);
or U15003 (N_15003,N_13286,N_13526);
nand U15004 (N_15004,N_13457,N_12398);
nor U15005 (N_15005,N_12546,N_13651);
nor U15006 (N_15006,N_12201,N_12268);
and U15007 (N_15007,N_12574,N_12585);
nand U15008 (N_15008,N_12165,N_12702);
or U15009 (N_15009,N_13816,N_12766);
nor U15010 (N_15010,N_13806,N_13895);
and U15011 (N_15011,N_12251,N_13809);
xor U15012 (N_15012,N_13966,N_12191);
or U15013 (N_15013,N_13263,N_12851);
xor U15014 (N_15014,N_12041,N_12577);
xor U15015 (N_15015,N_12404,N_12041);
nor U15016 (N_15016,N_13106,N_12124);
or U15017 (N_15017,N_12597,N_12483);
xor U15018 (N_15018,N_12545,N_13377);
or U15019 (N_15019,N_13057,N_12398);
xor U15020 (N_15020,N_13979,N_13500);
xnor U15021 (N_15021,N_12004,N_13827);
nand U15022 (N_15022,N_13104,N_13056);
and U15023 (N_15023,N_13871,N_13650);
nand U15024 (N_15024,N_12232,N_12639);
xor U15025 (N_15025,N_12782,N_12736);
nor U15026 (N_15026,N_12554,N_13774);
and U15027 (N_15027,N_12620,N_12822);
nor U15028 (N_15028,N_13414,N_12694);
or U15029 (N_15029,N_13078,N_12567);
nand U15030 (N_15030,N_13774,N_12037);
xor U15031 (N_15031,N_13616,N_12189);
nor U15032 (N_15032,N_12652,N_12570);
or U15033 (N_15033,N_13570,N_13793);
nor U15034 (N_15034,N_13917,N_13246);
nor U15035 (N_15035,N_13773,N_13286);
nand U15036 (N_15036,N_13154,N_13883);
nand U15037 (N_15037,N_12905,N_12337);
nand U15038 (N_15038,N_13401,N_12877);
nor U15039 (N_15039,N_12159,N_12652);
and U15040 (N_15040,N_12839,N_12330);
and U15041 (N_15041,N_13266,N_13943);
xnor U15042 (N_15042,N_12023,N_13185);
and U15043 (N_15043,N_12916,N_13540);
nor U15044 (N_15044,N_12973,N_12341);
nand U15045 (N_15045,N_12258,N_12710);
nor U15046 (N_15046,N_12707,N_12515);
and U15047 (N_15047,N_13125,N_13899);
or U15048 (N_15048,N_12901,N_13171);
and U15049 (N_15049,N_12790,N_12582);
xor U15050 (N_15050,N_12391,N_12332);
nand U15051 (N_15051,N_12691,N_12283);
or U15052 (N_15052,N_12369,N_12976);
nand U15053 (N_15053,N_12821,N_13829);
and U15054 (N_15054,N_13855,N_12613);
or U15055 (N_15055,N_12718,N_13489);
xor U15056 (N_15056,N_12860,N_13285);
nor U15057 (N_15057,N_13778,N_12167);
or U15058 (N_15058,N_13584,N_13686);
or U15059 (N_15059,N_13187,N_13489);
or U15060 (N_15060,N_13604,N_13498);
nand U15061 (N_15061,N_13138,N_13503);
nor U15062 (N_15062,N_13074,N_13568);
and U15063 (N_15063,N_13258,N_13924);
xnor U15064 (N_15064,N_12649,N_12983);
and U15065 (N_15065,N_12421,N_12839);
nand U15066 (N_15066,N_12451,N_12432);
and U15067 (N_15067,N_12179,N_13084);
and U15068 (N_15068,N_12235,N_13921);
nor U15069 (N_15069,N_12294,N_12289);
xnor U15070 (N_15070,N_13900,N_12421);
xnor U15071 (N_15071,N_12324,N_13755);
or U15072 (N_15072,N_13914,N_13165);
xor U15073 (N_15073,N_13196,N_13761);
nor U15074 (N_15074,N_12041,N_12637);
and U15075 (N_15075,N_12150,N_12262);
nand U15076 (N_15076,N_13964,N_13008);
nand U15077 (N_15077,N_13668,N_13860);
nand U15078 (N_15078,N_12146,N_12051);
xor U15079 (N_15079,N_12523,N_13661);
or U15080 (N_15080,N_13675,N_12157);
xor U15081 (N_15081,N_13834,N_12944);
and U15082 (N_15082,N_12791,N_13429);
nor U15083 (N_15083,N_13287,N_13982);
xor U15084 (N_15084,N_13439,N_12123);
nor U15085 (N_15085,N_13921,N_12820);
or U15086 (N_15086,N_13885,N_13456);
xnor U15087 (N_15087,N_12550,N_13793);
and U15088 (N_15088,N_13975,N_12721);
nor U15089 (N_15089,N_13286,N_13702);
or U15090 (N_15090,N_13474,N_13351);
xnor U15091 (N_15091,N_13833,N_13122);
or U15092 (N_15092,N_13771,N_12367);
nand U15093 (N_15093,N_13658,N_12040);
nand U15094 (N_15094,N_12479,N_13441);
xnor U15095 (N_15095,N_12360,N_13783);
xor U15096 (N_15096,N_12237,N_12601);
xnor U15097 (N_15097,N_12901,N_12878);
nor U15098 (N_15098,N_12987,N_12377);
nand U15099 (N_15099,N_13757,N_13869);
or U15100 (N_15100,N_13543,N_13303);
and U15101 (N_15101,N_13747,N_13052);
xor U15102 (N_15102,N_12650,N_13174);
and U15103 (N_15103,N_12594,N_13062);
and U15104 (N_15104,N_12289,N_13829);
and U15105 (N_15105,N_12485,N_12121);
nor U15106 (N_15106,N_13440,N_12154);
and U15107 (N_15107,N_13439,N_13690);
nand U15108 (N_15108,N_12933,N_12098);
nor U15109 (N_15109,N_12967,N_12270);
xor U15110 (N_15110,N_13728,N_12640);
or U15111 (N_15111,N_12574,N_12993);
nand U15112 (N_15112,N_12010,N_13319);
nor U15113 (N_15113,N_13422,N_12160);
and U15114 (N_15114,N_12097,N_12176);
xor U15115 (N_15115,N_12257,N_13779);
nor U15116 (N_15116,N_12932,N_12670);
nand U15117 (N_15117,N_13222,N_12786);
nor U15118 (N_15118,N_13711,N_12575);
nor U15119 (N_15119,N_12443,N_12531);
nand U15120 (N_15120,N_13682,N_12738);
xor U15121 (N_15121,N_12161,N_12407);
xnor U15122 (N_15122,N_12229,N_12290);
or U15123 (N_15123,N_13135,N_13678);
and U15124 (N_15124,N_13253,N_13219);
nand U15125 (N_15125,N_13933,N_12286);
or U15126 (N_15126,N_12735,N_13896);
xnor U15127 (N_15127,N_12776,N_13941);
or U15128 (N_15128,N_13005,N_12348);
xnor U15129 (N_15129,N_12958,N_12778);
nor U15130 (N_15130,N_13337,N_13773);
and U15131 (N_15131,N_13252,N_13963);
nand U15132 (N_15132,N_13400,N_12146);
nor U15133 (N_15133,N_12780,N_13291);
xor U15134 (N_15134,N_12605,N_12427);
xnor U15135 (N_15135,N_13113,N_12898);
xnor U15136 (N_15136,N_12839,N_13262);
nand U15137 (N_15137,N_12774,N_13151);
xor U15138 (N_15138,N_12848,N_12965);
nor U15139 (N_15139,N_13863,N_12707);
or U15140 (N_15140,N_13492,N_12396);
nand U15141 (N_15141,N_12844,N_13084);
xnor U15142 (N_15142,N_12025,N_13375);
nand U15143 (N_15143,N_12968,N_12127);
nand U15144 (N_15144,N_13703,N_12962);
nand U15145 (N_15145,N_12583,N_13962);
nand U15146 (N_15146,N_12585,N_12413);
and U15147 (N_15147,N_12529,N_13638);
nor U15148 (N_15148,N_12954,N_13314);
and U15149 (N_15149,N_12331,N_12179);
and U15150 (N_15150,N_13918,N_13414);
nand U15151 (N_15151,N_12376,N_13179);
xor U15152 (N_15152,N_13241,N_12829);
nand U15153 (N_15153,N_13493,N_12575);
nand U15154 (N_15154,N_12515,N_12563);
or U15155 (N_15155,N_12142,N_12482);
nor U15156 (N_15156,N_12869,N_13107);
and U15157 (N_15157,N_13900,N_13390);
and U15158 (N_15158,N_13634,N_12599);
nand U15159 (N_15159,N_13853,N_12641);
nor U15160 (N_15160,N_12097,N_13900);
xor U15161 (N_15161,N_13209,N_13293);
nor U15162 (N_15162,N_12976,N_13187);
nor U15163 (N_15163,N_13224,N_12362);
nand U15164 (N_15164,N_13750,N_12564);
and U15165 (N_15165,N_13629,N_12331);
xor U15166 (N_15166,N_13978,N_12993);
and U15167 (N_15167,N_12097,N_13558);
xor U15168 (N_15168,N_12997,N_13050);
and U15169 (N_15169,N_12810,N_12222);
nor U15170 (N_15170,N_12202,N_13483);
xnor U15171 (N_15171,N_12317,N_13981);
and U15172 (N_15172,N_13232,N_13770);
or U15173 (N_15173,N_12314,N_12467);
or U15174 (N_15174,N_12114,N_13967);
or U15175 (N_15175,N_13772,N_13613);
nand U15176 (N_15176,N_12718,N_13775);
nor U15177 (N_15177,N_12705,N_12500);
and U15178 (N_15178,N_12312,N_12169);
or U15179 (N_15179,N_12104,N_12882);
xor U15180 (N_15180,N_13302,N_12056);
or U15181 (N_15181,N_12887,N_13194);
or U15182 (N_15182,N_13538,N_12175);
or U15183 (N_15183,N_12137,N_12453);
or U15184 (N_15184,N_12039,N_12785);
and U15185 (N_15185,N_12469,N_12449);
nor U15186 (N_15186,N_13400,N_13554);
or U15187 (N_15187,N_12511,N_13214);
nand U15188 (N_15188,N_12854,N_12406);
nor U15189 (N_15189,N_13511,N_12228);
xor U15190 (N_15190,N_12089,N_12711);
nand U15191 (N_15191,N_13241,N_12010);
or U15192 (N_15192,N_12654,N_13954);
or U15193 (N_15193,N_12923,N_13533);
or U15194 (N_15194,N_12335,N_12444);
nand U15195 (N_15195,N_13326,N_13536);
nor U15196 (N_15196,N_13180,N_13131);
or U15197 (N_15197,N_13001,N_13472);
xnor U15198 (N_15198,N_12503,N_13426);
xor U15199 (N_15199,N_12089,N_12293);
or U15200 (N_15200,N_13726,N_13739);
or U15201 (N_15201,N_12652,N_12322);
or U15202 (N_15202,N_12369,N_13752);
or U15203 (N_15203,N_13647,N_12938);
nand U15204 (N_15204,N_12365,N_13947);
or U15205 (N_15205,N_13612,N_13732);
nand U15206 (N_15206,N_12041,N_13743);
nor U15207 (N_15207,N_13099,N_13633);
xnor U15208 (N_15208,N_12991,N_13058);
xnor U15209 (N_15209,N_13885,N_12202);
xor U15210 (N_15210,N_13311,N_13583);
nand U15211 (N_15211,N_12480,N_13215);
xor U15212 (N_15212,N_13364,N_12529);
or U15213 (N_15213,N_12585,N_13332);
or U15214 (N_15214,N_12966,N_12997);
nand U15215 (N_15215,N_13492,N_12824);
xnor U15216 (N_15216,N_13620,N_13514);
nand U15217 (N_15217,N_13253,N_13981);
nand U15218 (N_15218,N_12879,N_12693);
nand U15219 (N_15219,N_12519,N_12421);
xor U15220 (N_15220,N_12707,N_13878);
or U15221 (N_15221,N_12766,N_13412);
and U15222 (N_15222,N_13022,N_12934);
nand U15223 (N_15223,N_12207,N_13815);
nor U15224 (N_15224,N_12467,N_13442);
and U15225 (N_15225,N_13233,N_12320);
xor U15226 (N_15226,N_13550,N_13781);
nand U15227 (N_15227,N_13266,N_12921);
nor U15228 (N_15228,N_13379,N_12255);
and U15229 (N_15229,N_12726,N_13020);
nand U15230 (N_15230,N_12102,N_12025);
nand U15231 (N_15231,N_13480,N_13535);
or U15232 (N_15232,N_13888,N_12650);
nor U15233 (N_15233,N_13026,N_12818);
xor U15234 (N_15234,N_12461,N_13419);
xor U15235 (N_15235,N_13906,N_13987);
xnor U15236 (N_15236,N_13933,N_12928);
xnor U15237 (N_15237,N_12619,N_12134);
and U15238 (N_15238,N_13497,N_13056);
or U15239 (N_15239,N_13761,N_13197);
xor U15240 (N_15240,N_12786,N_13420);
nor U15241 (N_15241,N_13781,N_12193);
xor U15242 (N_15242,N_12055,N_12828);
xnor U15243 (N_15243,N_12381,N_12047);
xor U15244 (N_15244,N_12595,N_12610);
nor U15245 (N_15245,N_12452,N_13331);
nor U15246 (N_15246,N_12812,N_13363);
nor U15247 (N_15247,N_13302,N_12832);
xnor U15248 (N_15248,N_13890,N_12291);
nor U15249 (N_15249,N_13001,N_13559);
or U15250 (N_15250,N_13590,N_12386);
nor U15251 (N_15251,N_12516,N_12691);
xnor U15252 (N_15252,N_12013,N_12440);
and U15253 (N_15253,N_13582,N_12250);
nor U15254 (N_15254,N_13047,N_13326);
or U15255 (N_15255,N_12327,N_12216);
or U15256 (N_15256,N_13868,N_12159);
xor U15257 (N_15257,N_12370,N_12479);
nor U15258 (N_15258,N_12145,N_12066);
nor U15259 (N_15259,N_12321,N_12394);
and U15260 (N_15260,N_12473,N_12536);
nor U15261 (N_15261,N_13146,N_12319);
nor U15262 (N_15262,N_12036,N_13201);
nor U15263 (N_15263,N_12602,N_13606);
and U15264 (N_15264,N_12336,N_12098);
and U15265 (N_15265,N_12876,N_12805);
or U15266 (N_15266,N_12585,N_12394);
xnor U15267 (N_15267,N_13484,N_13648);
xnor U15268 (N_15268,N_13145,N_13361);
or U15269 (N_15269,N_13673,N_13993);
nor U15270 (N_15270,N_13211,N_12276);
and U15271 (N_15271,N_12757,N_13409);
xor U15272 (N_15272,N_12671,N_12378);
xor U15273 (N_15273,N_12926,N_12529);
and U15274 (N_15274,N_13552,N_12634);
xnor U15275 (N_15275,N_13357,N_12283);
xnor U15276 (N_15276,N_13923,N_13109);
nor U15277 (N_15277,N_13383,N_13855);
or U15278 (N_15278,N_13307,N_13268);
nor U15279 (N_15279,N_12384,N_13328);
or U15280 (N_15280,N_13076,N_13276);
nor U15281 (N_15281,N_13904,N_13826);
and U15282 (N_15282,N_12771,N_12642);
nor U15283 (N_15283,N_13998,N_13791);
nor U15284 (N_15284,N_13759,N_12336);
nand U15285 (N_15285,N_13552,N_12391);
and U15286 (N_15286,N_12489,N_13618);
xor U15287 (N_15287,N_13726,N_12847);
nor U15288 (N_15288,N_12277,N_13926);
and U15289 (N_15289,N_13141,N_12219);
and U15290 (N_15290,N_13602,N_12595);
nand U15291 (N_15291,N_13921,N_13950);
and U15292 (N_15292,N_13516,N_12603);
nor U15293 (N_15293,N_13240,N_13592);
nor U15294 (N_15294,N_13408,N_13036);
nor U15295 (N_15295,N_13869,N_12718);
nand U15296 (N_15296,N_12180,N_13262);
nor U15297 (N_15297,N_12124,N_12470);
nand U15298 (N_15298,N_13078,N_13689);
and U15299 (N_15299,N_13124,N_12166);
nand U15300 (N_15300,N_12414,N_13810);
nand U15301 (N_15301,N_13189,N_12168);
nor U15302 (N_15302,N_13600,N_13227);
and U15303 (N_15303,N_13865,N_13296);
nor U15304 (N_15304,N_13683,N_13639);
and U15305 (N_15305,N_12946,N_13145);
or U15306 (N_15306,N_12264,N_12082);
or U15307 (N_15307,N_13738,N_13166);
xnor U15308 (N_15308,N_13085,N_13789);
nand U15309 (N_15309,N_12624,N_12174);
nor U15310 (N_15310,N_13544,N_13087);
or U15311 (N_15311,N_13922,N_13619);
and U15312 (N_15312,N_13788,N_13320);
xnor U15313 (N_15313,N_13926,N_13869);
or U15314 (N_15314,N_13387,N_13770);
and U15315 (N_15315,N_13130,N_12990);
nand U15316 (N_15316,N_12739,N_13430);
nand U15317 (N_15317,N_12149,N_12262);
xnor U15318 (N_15318,N_13165,N_12783);
and U15319 (N_15319,N_13570,N_12354);
and U15320 (N_15320,N_12461,N_12062);
and U15321 (N_15321,N_13821,N_12266);
nor U15322 (N_15322,N_12534,N_13777);
nand U15323 (N_15323,N_12986,N_12012);
xor U15324 (N_15324,N_12908,N_13353);
or U15325 (N_15325,N_12431,N_13446);
and U15326 (N_15326,N_12235,N_13878);
and U15327 (N_15327,N_13052,N_13329);
nand U15328 (N_15328,N_12893,N_12913);
xnor U15329 (N_15329,N_13228,N_13214);
or U15330 (N_15330,N_13864,N_12796);
or U15331 (N_15331,N_13636,N_12172);
and U15332 (N_15332,N_12532,N_13339);
or U15333 (N_15333,N_12287,N_12448);
xnor U15334 (N_15334,N_13055,N_13035);
xor U15335 (N_15335,N_12181,N_12369);
or U15336 (N_15336,N_13862,N_13559);
xor U15337 (N_15337,N_12104,N_13888);
xnor U15338 (N_15338,N_12862,N_13037);
and U15339 (N_15339,N_13674,N_12849);
nand U15340 (N_15340,N_13044,N_13613);
xor U15341 (N_15341,N_12576,N_12933);
nand U15342 (N_15342,N_13503,N_12728);
and U15343 (N_15343,N_13131,N_12873);
xnor U15344 (N_15344,N_12503,N_12309);
or U15345 (N_15345,N_13625,N_12584);
xor U15346 (N_15346,N_12041,N_13455);
nor U15347 (N_15347,N_12554,N_13300);
xnor U15348 (N_15348,N_12924,N_12904);
nor U15349 (N_15349,N_12618,N_12328);
xor U15350 (N_15350,N_12427,N_12182);
nand U15351 (N_15351,N_13632,N_13604);
nor U15352 (N_15352,N_13978,N_12218);
or U15353 (N_15353,N_13568,N_12646);
nand U15354 (N_15354,N_13634,N_13971);
nor U15355 (N_15355,N_13555,N_13851);
xnor U15356 (N_15356,N_13236,N_12058);
nand U15357 (N_15357,N_13886,N_12783);
nand U15358 (N_15358,N_12269,N_13305);
or U15359 (N_15359,N_12795,N_13691);
xor U15360 (N_15360,N_12923,N_13194);
nor U15361 (N_15361,N_13820,N_12296);
or U15362 (N_15362,N_13245,N_12849);
nand U15363 (N_15363,N_13280,N_12494);
nor U15364 (N_15364,N_12616,N_12339);
or U15365 (N_15365,N_12624,N_12993);
nand U15366 (N_15366,N_12280,N_12664);
nor U15367 (N_15367,N_12885,N_13093);
and U15368 (N_15368,N_13410,N_13784);
nand U15369 (N_15369,N_13352,N_12949);
nand U15370 (N_15370,N_12741,N_12098);
and U15371 (N_15371,N_13497,N_13070);
xnor U15372 (N_15372,N_13165,N_12399);
and U15373 (N_15373,N_13834,N_13525);
and U15374 (N_15374,N_13804,N_13676);
nand U15375 (N_15375,N_13679,N_12209);
xor U15376 (N_15376,N_13400,N_13038);
nor U15377 (N_15377,N_12398,N_13463);
or U15378 (N_15378,N_13991,N_13173);
xor U15379 (N_15379,N_12184,N_12291);
and U15380 (N_15380,N_13916,N_12765);
nor U15381 (N_15381,N_13167,N_12467);
nor U15382 (N_15382,N_13377,N_12026);
and U15383 (N_15383,N_12146,N_13168);
nand U15384 (N_15384,N_12609,N_13540);
or U15385 (N_15385,N_12680,N_13511);
nand U15386 (N_15386,N_12908,N_12801);
xor U15387 (N_15387,N_13647,N_12123);
nand U15388 (N_15388,N_13747,N_13801);
nor U15389 (N_15389,N_12868,N_13378);
nand U15390 (N_15390,N_12259,N_12968);
nor U15391 (N_15391,N_12184,N_13527);
xor U15392 (N_15392,N_12010,N_12077);
xnor U15393 (N_15393,N_12997,N_12274);
nand U15394 (N_15394,N_13841,N_13665);
xnor U15395 (N_15395,N_12134,N_12352);
nor U15396 (N_15396,N_13562,N_13135);
nor U15397 (N_15397,N_12680,N_13353);
and U15398 (N_15398,N_12772,N_13278);
and U15399 (N_15399,N_12919,N_13453);
and U15400 (N_15400,N_13800,N_13592);
xor U15401 (N_15401,N_12158,N_12370);
xnor U15402 (N_15402,N_13262,N_12136);
or U15403 (N_15403,N_12212,N_12603);
and U15404 (N_15404,N_12295,N_13127);
xor U15405 (N_15405,N_12833,N_12595);
and U15406 (N_15406,N_12715,N_12008);
nor U15407 (N_15407,N_12439,N_13823);
nand U15408 (N_15408,N_13948,N_12841);
nor U15409 (N_15409,N_12214,N_12859);
and U15410 (N_15410,N_13687,N_13306);
nand U15411 (N_15411,N_13626,N_12932);
or U15412 (N_15412,N_12415,N_12837);
and U15413 (N_15413,N_13815,N_12525);
and U15414 (N_15414,N_13484,N_13876);
or U15415 (N_15415,N_13330,N_13075);
xor U15416 (N_15416,N_12492,N_13348);
or U15417 (N_15417,N_13398,N_12956);
xnor U15418 (N_15418,N_12073,N_12609);
nor U15419 (N_15419,N_13706,N_12468);
or U15420 (N_15420,N_13912,N_12101);
or U15421 (N_15421,N_13983,N_13514);
xor U15422 (N_15422,N_13007,N_12141);
nor U15423 (N_15423,N_12359,N_13834);
nand U15424 (N_15424,N_13332,N_12969);
nand U15425 (N_15425,N_12991,N_13505);
nor U15426 (N_15426,N_13875,N_12519);
or U15427 (N_15427,N_13056,N_12663);
nand U15428 (N_15428,N_13238,N_12036);
nand U15429 (N_15429,N_13696,N_12796);
xor U15430 (N_15430,N_12875,N_12326);
xnor U15431 (N_15431,N_12249,N_12079);
nand U15432 (N_15432,N_13812,N_13124);
nor U15433 (N_15433,N_12294,N_12828);
nor U15434 (N_15434,N_12195,N_12501);
xnor U15435 (N_15435,N_12561,N_12171);
nor U15436 (N_15436,N_12739,N_13115);
nand U15437 (N_15437,N_12822,N_13697);
nor U15438 (N_15438,N_13339,N_12644);
xnor U15439 (N_15439,N_12013,N_13395);
nand U15440 (N_15440,N_12185,N_13942);
or U15441 (N_15441,N_13583,N_12761);
nor U15442 (N_15442,N_13557,N_13341);
nor U15443 (N_15443,N_13848,N_13715);
nor U15444 (N_15444,N_13553,N_13048);
xor U15445 (N_15445,N_13813,N_13665);
nor U15446 (N_15446,N_12526,N_12207);
nor U15447 (N_15447,N_12487,N_12792);
nand U15448 (N_15448,N_12071,N_12916);
or U15449 (N_15449,N_12840,N_12937);
nor U15450 (N_15450,N_13428,N_12533);
xnor U15451 (N_15451,N_13774,N_13686);
or U15452 (N_15452,N_12864,N_12610);
nor U15453 (N_15453,N_13777,N_13449);
or U15454 (N_15454,N_13531,N_13919);
xnor U15455 (N_15455,N_12273,N_13250);
nand U15456 (N_15456,N_12737,N_13179);
nand U15457 (N_15457,N_13797,N_13902);
and U15458 (N_15458,N_12014,N_12889);
nor U15459 (N_15459,N_12900,N_12034);
and U15460 (N_15460,N_12268,N_12104);
or U15461 (N_15461,N_13315,N_13761);
or U15462 (N_15462,N_12502,N_13358);
nor U15463 (N_15463,N_13307,N_12900);
nor U15464 (N_15464,N_12831,N_13404);
or U15465 (N_15465,N_13771,N_12627);
or U15466 (N_15466,N_13366,N_13150);
nand U15467 (N_15467,N_13809,N_13643);
or U15468 (N_15468,N_13463,N_13276);
xor U15469 (N_15469,N_13528,N_12052);
and U15470 (N_15470,N_12151,N_12954);
or U15471 (N_15471,N_13982,N_13354);
and U15472 (N_15472,N_13669,N_12179);
nand U15473 (N_15473,N_13896,N_12650);
nand U15474 (N_15474,N_12480,N_13059);
and U15475 (N_15475,N_12840,N_12900);
xnor U15476 (N_15476,N_12949,N_12114);
and U15477 (N_15477,N_12118,N_12335);
and U15478 (N_15478,N_12989,N_12617);
xor U15479 (N_15479,N_12861,N_12754);
xor U15480 (N_15480,N_13513,N_13948);
and U15481 (N_15481,N_13477,N_13941);
or U15482 (N_15482,N_12192,N_12599);
and U15483 (N_15483,N_13905,N_13552);
nand U15484 (N_15484,N_12674,N_12348);
and U15485 (N_15485,N_13516,N_12991);
xor U15486 (N_15486,N_12943,N_12886);
or U15487 (N_15487,N_13965,N_13174);
and U15488 (N_15488,N_13461,N_13771);
and U15489 (N_15489,N_13859,N_12565);
xnor U15490 (N_15490,N_13470,N_12427);
xor U15491 (N_15491,N_13522,N_12089);
or U15492 (N_15492,N_12515,N_13735);
nand U15493 (N_15493,N_13313,N_12002);
nor U15494 (N_15494,N_13022,N_12807);
or U15495 (N_15495,N_12491,N_13041);
nor U15496 (N_15496,N_13110,N_13238);
or U15497 (N_15497,N_12257,N_13089);
nor U15498 (N_15498,N_13165,N_13900);
nand U15499 (N_15499,N_12124,N_13630);
or U15500 (N_15500,N_13931,N_12450);
nand U15501 (N_15501,N_13383,N_13295);
xor U15502 (N_15502,N_13875,N_13739);
nand U15503 (N_15503,N_12084,N_12433);
or U15504 (N_15504,N_13994,N_13541);
nand U15505 (N_15505,N_12057,N_12291);
nand U15506 (N_15506,N_12392,N_13707);
nor U15507 (N_15507,N_12314,N_13283);
and U15508 (N_15508,N_12824,N_12974);
nor U15509 (N_15509,N_12914,N_12894);
nand U15510 (N_15510,N_12759,N_13229);
and U15511 (N_15511,N_12308,N_13021);
or U15512 (N_15512,N_12187,N_13033);
or U15513 (N_15513,N_13085,N_12378);
xnor U15514 (N_15514,N_12523,N_13180);
xnor U15515 (N_15515,N_12483,N_13195);
and U15516 (N_15516,N_13221,N_13248);
and U15517 (N_15517,N_12374,N_12762);
or U15518 (N_15518,N_13892,N_12215);
and U15519 (N_15519,N_12723,N_12237);
nor U15520 (N_15520,N_12977,N_13269);
nand U15521 (N_15521,N_12395,N_12343);
nor U15522 (N_15522,N_13913,N_12364);
and U15523 (N_15523,N_12130,N_13090);
and U15524 (N_15524,N_12006,N_13303);
nand U15525 (N_15525,N_13177,N_13294);
or U15526 (N_15526,N_13912,N_13138);
and U15527 (N_15527,N_13592,N_12682);
nor U15528 (N_15528,N_12301,N_13385);
nand U15529 (N_15529,N_12887,N_13316);
and U15530 (N_15530,N_12471,N_12806);
nand U15531 (N_15531,N_12551,N_13714);
xnor U15532 (N_15532,N_12345,N_12439);
nor U15533 (N_15533,N_12388,N_12624);
nor U15534 (N_15534,N_13500,N_13684);
and U15535 (N_15535,N_12372,N_12581);
and U15536 (N_15536,N_13801,N_12748);
and U15537 (N_15537,N_13046,N_12808);
or U15538 (N_15538,N_12578,N_12408);
or U15539 (N_15539,N_12090,N_13553);
or U15540 (N_15540,N_12082,N_13963);
xnor U15541 (N_15541,N_13212,N_13527);
or U15542 (N_15542,N_13780,N_13765);
nor U15543 (N_15543,N_13328,N_12141);
nor U15544 (N_15544,N_13933,N_12835);
nand U15545 (N_15545,N_12902,N_13811);
nand U15546 (N_15546,N_12335,N_12430);
nor U15547 (N_15547,N_12266,N_13975);
nand U15548 (N_15548,N_12677,N_13387);
and U15549 (N_15549,N_13433,N_12196);
nand U15550 (N_15550,N_13883,N_12415);
xnor U15551 (N_15551,N_12410,N_13025);
nor U15552 (N_15552,N_13589,N_13800);
and U15553 (N_15553,N_13614,N_13790);
or U15554 (N_15554,N_13915,N_12336);
nor U15555 (N_15555,N_13078,N_12915);
or U15556 (N_15556,N_12477,N_13179);
xnor U15557 (N_15557,N_13745,N_12423);
xor U15558 (N_15558,N_13719,N_13506);
nand U15559 (N_15559,N_13291,N_13009);
xnor U15560 (N_15560,N_13117,N_13282);
xor U15561 (N_15561,N_13894,N_12474);
nand U15562 (N_15562,N_13728,N_13133);
or U15563 (N_15563,N_13671,N_12551);
xnor U15564 (N_15564,N_12843,N_12944);
nand U15565 (N_15565,N_12926,N_12361);
xor U15566 (N_15566,N_13551,N_12284);
or U15567 (N_15567,N_12180,N_12651);
and U15568 (N_15568,N_12253,N_12847);
and U15569 (N_15569,N_13290,N_13321);
and U15570 (N_15570,N_13249,N_13766);
nor U15571 (N_15571,N_13713,N_12791);
nor U15572 (N_15572,N_12223,N_12671);
nor U15573 (N_15573,N_13190,N_12820);
nand U15574 (N_15574,N_13896,N_12206);
nor U15575 (N_15575,N_12069,N_12832);
and U15576 (N_15576,N_12442,N_13408);
xor U15577 (N_15577,N_12480,N_12496);
xnor U15578 (N_15578,N_12144,N_13185);
xor U15579 (N_15579,N_13052,N_12326);
xor U15580 (N_15580,N_12809,N_13423);
xor U15581 (N_15581,N_13632,N_12904);
or U15582 (N_15582,N_13338,N_12499);
nor U15583 (N_15583,N_12184,N_12423);
and U15584 (N_15584,N_12095,N_12638);
or U15585 (N_15585,N_13647,N_12941);
nand U15586 (N_15586,N_13859,N_13246);
nor U15587 (N_15587,N_12084,N_12128);
xor U15588 (N_15588,N_13454,N_13996);
nand U15589 (N_15589,N_13273,N_13277);
xnor U15590 (N_15590,N_13110,N_13576);
nor U15591 (N_15591,N_13707,N_13838);
xnor U15592 (N_15592,N_12040,N_13987);
nor U15593 (N_15593,N_12386,N_13664);
xnor U15594 (N_15594,N_12320,N_13694);
nor U15595 (N_15595,N_12337,N_12507);
nand U15596 (N_15596,N_12571,N_13446);
nand U15597 (N_15597,N_13687,N_12823);
nor U15598 (N_15598,N_13555,N_12981);
nand U15599 (N_15599,N_13694,N_13997);
nor U15600 (N_15600,N_13759,N_13655);
or U15601 (N_15601,N_13968,N_12911);
xnor U15602 (N_15602,N_13241,N_13413);
xnor U15603 (N_15603,N_12455,N_13285);
xnor U15604 (N_15604,N_13783,N_12081);
or U15605 (N_15605,N_12880,N_12166);
and U15606 (N_15606,N_13678,N_12787);
nand U15607 (N_15607,N_13341,N_12364);
nor U15608 (N_15608,N_12794,N_12675);
nor U15609 (N_15609,N_13421,N_13536);
and U15610 (N_15610,N_13703,N_13501);
xor U15611 (N_15611,N_12674,N_13064);
nor U15612 (N_15612,N_13017,N_13952);
xnor U15613 (N_15613,N_12178,N_12984);
nand U15614 (N_15614,N_12232,N_12894);
or U15615 (N_15615,N_13051,N_12364);
xnor U15616 (N_15616,N_13889,N_13656);
nor U15617 (N_15617,N_12224,N_12834);
or U15618 (N_15618,N_13045,N_13595);
nand U15619 (N_15619,N_12449,N_13375);
or U15620 (N_15620,N_12439,N_12594);
and U15621 (N_15621,N_12072,N_13020);
or U15622 (N_15622,N_12531,N_13188);
and U15623 (N_15623,N_13343,N_12704);
and U15624 (N_15624,N_12105,N_13472);
and U15625 (N_15625,N_12354,N_12256);
nand U15626 (N_15626,N_12276,N_12899);
xor U15627 (N_15627,N_12224,N_13027);
or U15628 (N_15628,N_13055,N_13393);
nand U15629 (N_15629,N_12956,N_13411);
or U15630 (N_15630,N_13393,N_13488);
and U15631 (N_15631,N_12729,N_12919);
nand U15632 (N_15632,N_12367,N_13517);
nand U15633 (N_15633,N_12352,N_13983);
or U15634 (N_15634,N_12548,N_12442);
or U15635 (N_15635,N_12620,N_12933);
nand U15636 (N_15636,N_13882,N_12880);
nor U15637 (N_15637,N_12263,N_12427);
nand U15638 (N_15638,N_13554,N_12212);
nor U15639 (N_15639,N_13421,N_13499);
xor U15640 (N_15640,N_12106,N_12648);
or U15641 (N_15641,N_13878,N_13379);
or U15642 (N_15642,N_12209,N_13831);
xor U15643 (N_15643,N_12028,N_12523);
nor U15644 (N_15644,N_12333,N_13813);
xnor U15645 (N_15645,N_13909,N_13435);
nor U15646 (N_15646,N_13893,N_13372);
and U15647 (N_15647,N_13091,N_13261);
xor U15648 (N_15648,N_13615,N_13412);
or U15649 (N_15649,N_12612,N_12986);
nor U15650 (N_15650,N_12148,N_12723);
nor U15651 (N_15651,N_12961,N_12362);
and U15652 (N_15652,N_12864,N_12916);
and U15653 (N_15653,N_13122,N_13572);
nor U15654 (N_15654,N_13543,N_12114);
xnor U15655 (N_15655,N_13647,N_13677);
and U15656 (N_15656,N_13897,N_12000);
nand U15657 (N_15657,N_13378,N_12431);
nand U15658 (N_15658,N_12134,N_13204);
nor U15659 (N_15659,N_13292,N_13743);
nor U15660 (N_15660,N_13113,N_12724);
nand U15661 (N_15661,N_13716,N_13056);
and U15662 (N_15662,N_12353,N_13772);
nand U15663 (N_15663,N_13500,N_12651);
nand U15664 (N_15664,N_12811,N_13320);
and U15665 (N_15665,N_13594,N_13748);
nor U15666 (N_15666,N_12596,N_13140);
nor U15667 (N_15667,N_12851,N_13326);
xor U15668 (N_15668,N_13089,N_13627);
or U15669 (N_15669,N_12540,N_12777);
nand U15670 (N_15670,N_13382,N_13449);
and U15671 (N_15671,N_12402,N_12078);
nand U15672 (N_15672,N_12534,N_12085);
and U15673 (N_15673,N_12439,N_13405);
or U15674 (N_15674,N_12179,N_13963);
nand U15675 (N_15675,N_12326,N_12662);
and U15676 (N_15676,N_12186,N_12594);
or U15677 (N_15677,N_13619,N_12322);
xnor U15678 (N_15678,N_12290,N_12312);
nand U15679 (N_15679,N_13869,N_13751);
nor U15680 (N_15680,N_13506,N_13854);
and U15681 (N_15681,N_13252,N_12532);
xor U15682 (N_15682,N_12480,N_12360);
xnor U15683 (N_15683,N_13511,N_12699);
nor U15684 (N_15684,N_12838,N_13349);
and U15685 (N_15685,N_13879,N_12668);
and U15686 (N_15686,N_13964,N_12624);
xnor U15687 (N_15687,N_12345,N_13162);
or U15688 (N_15688,N_13714,N_13225);
or U15689 (N_15689,N_13628,N_13291);
and U15690 (N_15690,N_13206,N_12311);
nor U15691 (N_15691,N_12689,N_12422);
xor U15692 (N_15692,N_13614,N_13967);
xnor U15693 (N_15693,N_13487,N_12624);
or U15694 (N_15694,N_12522,N_13055);
xnor U15695 (N_15695,N_13383,N_12117);
xor U15696 (N_15696,N_12885,N_13252);
and U15697 (N_15697,N_13864,N_12384);
and U15698 (N_15698,N_13776,N_13027);
nor U15699 (N_15699,N_13402,N_13350);
and U15700 (N_15700,N_13614,N_12668);
and U15701 (N_15701,N_13155,N_12243);
and U15702 (N_15702,N_13349,N_13513);
and U15703 (N_15703,N_12513,N_13628);
xnor U15704 (N_15704,N_13699,N_12756);
xor U15705 (N_15705,N_13089,N_12245);
and U15706 (N_15706,N_12260,N_13639);
or U15707 (N_15707,N_13065,N_13174);
nor U15708 (N_15708,N_12564,N_12711);
nand U15709 (N_15709,N_12734,N_13405);
xnor U15710 (N_15710,N_12581,N_13486);
nor U15711 (N_15711,N_12983,N_13910);
or U15712 (N_15712,N_13912,N_12612);
nor U15713 (N_15713,N_12122,N_12235);
and U15714 (N_15714,N_13359,N_12163);
nand U15715 (N_15715,N_13831,N_12950);
nor U15716 (N_15716,N_12486,N_12914);
or U15717 (N_15717,N_13901,N_13758);
or U15718 (N_15718,N_12211,N_13789);
and U15719 (N_15719,N_13242,N_13927);
or U15720 (N_15720,N_12395,N_12380);
nand U15721 (N_15721,N_13558,N_12685);
and U15722 (N_15722,N_13705,N_12097);
nor U15723 (N_15723,N_12140,N_13898);
or U15724 (N_15724,N_13115,N_12278);
or U15725 (N_15725,N_13150,N_13074);
and U15726 (N_15726,N_12216,N_13041);
or U15727 (N_15727,N_12767,N_13503);
or U15728 (N_15728,N_13765,N_12126);
nor U15729 (N_15729,N_12355,N_12787);
nand U15730 (N_15730,N_12254,N_12690);
or U15731 (N_15731,N_12563,N_13547);
and U15732 (N_15732,N_12907,N_12175);
xor U15733 (N_15733,N_12927,N_13904);
nand U15734 (N_15734,N_12065,N_12614);
and U15735 (N_15735,N_13273,N_13519);
xnor U15736 (N_15736,N_13652,N_12614);
and U15737 (N_15737,N_12212,N_13702);
xnor U15738 (N_15738,N_12608,N_13851);
nand U15739 (N_15739,N_12896,N_13374);
or U15740 (N_15740,N_13084,N_13501);
and U15741 (N_15741,N_13710,N_13420);
or U15742 (N_15742,N_13187,N_13601);
and U15743 (N_15743,N_12977,N_13555);
or U15744 (N_15744,N_13288,N_13700);
nor U15745 (N_15745,N_13195,N_12866);
and U15746 (N_15746,N_13145,N_12289);
nor U15747 (N_15747,N_13248,N_13059);
nand U15748 (N_15748,N_12939,N_13053);
or U15749 (N_15749,N_13559,N_12511);
and U15750 (N_15750,N_13161,N_12683);
nor U15751 (N_15751,N_12889,N_13166);
nor U15752 (N_15752,N_13904,N_13903);
nand U15753 (N_15753,N_13318,N_13019);
nor U15754 (N_15754,N_13532,N_12194);
xnor U15755 (N_15755,N_12315,N_13256);
nor U15756 (N_15756,N_13303,N_12050);
xor U15757 (N_15757,N_12058,N_13662);
nand U15758 (N_15758,N_12992,N_13937);
and U15759 (N_15759,N_12467,N_13396);
nand U15760 (N_15760,N_12699,N_12275);
and U15761 (N_15761,N_13070,N_13164);
and U15762 (N_15762,N_12366,N_13943);
xor U15763 (N_15763,N_12923,N_12761);
xor U15764 (N_15764,N_12672,N_12805);
and U15765 (N_15765,N_13594,N_12908);
or U15766 (N_15766,N_12057,N_13519);
xor U15767 (N_15767,N_13429,N_12890);
nand U15768 (N_15768,N_13601,N_12617);
or U15769 (N_15769,N_13980,N_12272);
or U15770 (N_15770,N_12045,N_12426);
xnor U15771 (N_15771,N_13268,N_12813);
xnor U15772 (N_15772,N_12409,N_13564);
xnor U15773 (N_15773,N_13561,N_13047);
xor U15774 (N_15774,N_13223,N_12266);
nand U15775 (N_15775,N_12784,N_12982);
nand U15776 (N_15776,N_12758,N_12172);
and U15777 (N_15777,N_12122,N_13293);
or U15778 (N_15778,N_13990,N_12112);
nand U15779 (N_15779,N_13959,N_12578);
and U15780 (N_15780,N_13469,N_13549);
nor U15781 (N_15781,N_13557,N_13589);
nand U15782 (N_15782,N_12220,N_12231);
nand U15783 (N_15783,N_13090,N_13168);
or U15784 (N_15784,N_13300,N_12620);
or U15785 (N_15785,N_12167,N_12077);
and U15786 (N_15786,N_12177,N_13091);
and U15787 (N_15787,N_12144,N_12007);
xor U15788 (N_15788,N_13433,N_13910);
nor U15789 (N_15789,N_13309,N_12250);
xor U15790 (N_15790,N_12094,N_12549);
nand U15791 (N_15791,N_13556,N_13272);
nand U15792 (N_15792,N_12931,N_13220);
or U15793 (N_15793,N_12214,N_12469);
xor U15794 (N_15794,N_12140,N_13086);
nand U15795 (N_15795,N_12878,N_12535);
nand U15796 (N_15796,N_13189,N_12407);
or U15797 (N_15797,N_13858,N_13295);
xor U15798 (N_15798,N_13325,N_12738);
nand U15799 (N_15799,N_13205,N_12308);
or U15800 (N_15800,N_13314,N_13414);
nand U15801 (N_15801,N_12951,N_13973);
and U15802 (N_15802,N_13623,N_12228);
or U15803 (N_15803,N_12531,N_12367);
xnor U15804 (N_15804,N_12432,N_12371);
xor U15805 (N_15805,N_13356,N_13542);
nor U15806 (N_15806,N_12176,N_13723);
and U15807 (N_15807,N_13113,N_12747);
or U15808 (N_15808,N_12685,N_13863);
nand U15809 (N_15809,N_13272,N_12013);
xor U15810 (N_15810,N_13611,N_12671);
nand U15811 (N_15811,N_12559,N_12501);
nand U15812 (N_15812,N_12755,N_12620);
and U15813 (N_15813,N_12386,N_13485);
or U15814 (N_15814,N_12141,N_12954);
nand U15815 (N_15815,N_13916,N_12749);
or U15816 (N_15816,N_13337,N_12588);
nand U15817 (N_15817,N_12314,N_12277);
nor U15818 (N_15818,N_12676,N_12272);
nor U15819 (N_15819,N_12783,N_12772);
nor U15820 (N_15820,N_12605,N_13532);
nand U15821 (N_15821,N_13508,N_13157);
nand U15822 (N_15822,N_13189,N_12357);
xor U15823 (N_15823,N_12783,N_12813);
nand U15824 (N_15824,N_12742,N_13354);
nand U15825 (N_15825,N_12374,N_13112);
xnor U15826 (N_15826,N_12034,N_12616);
xor U15827 (N_15827,N_13181,N_13197);
nor U15828 (N_15828,N_13093,N_13654);
nand U15829 (N_15829,N_12005,N_13600);
or U15830 (N_15830,N_13563,N_13753);
or U15831 (N_15831,N_12531,N_12518);
nor U15832 (N_15832,N_13957,N_13367);
and U15833 (N_15833,N_12536,N_12461);
nand U15834 (N_15834,N_12341,N_12247);
or U15835 (N_15835,N_12556,N_12489);
and U15836 (N_15836,N_13738,N_13943);
or U15837 (N_15837,N_13970,N_13187);
nor U15838 (N_15838,N_13845,N_12350);
xnor U15839 (N_15839,N_13554,N_12772);
and U15840 (N_15840,N_12409,N_13881);
and U15841 (N_15841,N_12081,N_13979);
and U15842 (N_15842,N_13733,N_13472);
or U15843 (N_15843,N_13506,N_12763);
nor U15844 (N_15844,N_12726,N_12393);
or U15845 (N_15845,N_13724,N_12505);
nor U15846 (N_15846,N_12937,N_12236);
xor U15847 (N_15847,N_12550,N_12241);
xor U15848 (N_15848,N_12159,N_13566);
xnor U15849 (N_15849,N_13544,N_12815);
and U15850 (N_15850,N_13750,N_12233);
and U15851 (N_15851,N_12416,N_12002);
nor U15852 (N_15852,N_12533,N_13537);
xnor U15853 (N_15853,N_12488,N_13514);
nor U15854 (N_15854,N_13321,N_12174);
and U15855 (N_15855,N_13689,N_13975);
xor U15856 (N_15856,N_12024,N_12283);
nor U15857 (N_15857,N_12980,N_13952);
nand U15858 (N_15858,N_12838,N_12382);
or U15859 (N_15859,N_12164,N_13900);
or U15860 (N_15860,N_13741,N_13500);
or U15861 (N_15861,N_12151,N_12125);
nand U15862 (N_15862,N_13220,N_13117);
or U15863 (N_15863,N_12719,N_13674);
nand U15864 (N_15864,N_13388,N_12469);
xnor U15865 (N_15865,N_12254,N_13937);
and U15866 (N_15866,N_12458,N_13266);
nor U15867 (N_15867,N_13757,N_12543);
xnor U15868 (N_15868,N_12181,N_12923);
nand U15869 (N_15869,N_12014,N_12492);
and U15870 (N_15870,N_12180,N_13677);
nand U15871 (N_15871,N_13036,N_13001);
xnor U15872 (N_15872,N_12078,N_13413);
nand U15873 (N_15873,N_12565,N_12640);
nand U15874 (N_15874,N_12851,N_12885);
or U15875 (N_15875,N_12522,N_12358);
nand U15876 (N_15876,N_12158,N_12236);
or U15877 (N_15877,N_12792,N_12462);
nor U15878 (N_15878,N_12913,N_12088);
nand U15879 (N_15879,N_13585,N_13467);
nor U15880 (N_15880,N_13132,N_13515);
or U15881 (N_15881,N_13993,N_13513);
nor U15882 (N_15882,N_12321,N_12690);
or U15883 (N_15883,N_13672,N_13631);
nor U15884 (N_15884,N_12943,N_13014);
nor U15885 (N_15885,N_12216,N_13931);
or U15886 (N_15886,N_13883,N_12320);
nand U15887 (N_15887,N_13079,N_13908);
nand U15888 (N_15888,N_13963,N_12097);
nor U15889 (N_15889,N_12961,N_12054);
or U15890 (N_15890,N_13047,N_12552);
and U15891 (N_15891,N_13886,N_13958);
xor U15892 (N_15892,N_12928,N_13532);
nor U15893 (N_15893,N_12609,N_12454);
nand U15894 (N_15894,N_12187,N_12551);
and U15895 (N_15895,N_12596,N_13618);
or U15896 (N_15896,N_12004,N_12522);
or U15897 (N_15897,N_12864,N_13366);
nor U15898 (N_15898,N_13829,N_13503);
nand U15899 (N_15899,N_13547,N_12574);
nand U15900 (N_15900,N_12559,N_13869);
or U15901 (N_15901,N_12884,N_13293);
or U15902 (N_15902,N_12481,N_13402);
and U15903 (N_15903,N_12242,N_12717);
nor U15904 (N_15904,N_12781,N_13777);
nor U15905 (N_15905,N_13546,N_12450);
nor U15906 (N_15906,N_13943,N_13285);
xnor U15907 (N_15907,N_13399,N_12532);
or U15908 (N_15908,N_12893,N_13203);
and U15909 (N_15909,N_12328,N_12312);
or U15910 (N_15910,N_12603,N_12391);
or U15911 (N_15911,N_13247,N_12835);
xnor U15912 (N_15912,N_13019,N_12191);
or U15913 (N_15913,N_13836,N_13331);
nand U15914 (N_15914,N_13869,N_13206);
and U15915 (N_15915,N_13698,N_13325);
xor U15916 (N_15916,N_12454,N_13180);
or U15917 (N_15917,N_12677,N_12045);
xnor U15918 (N_15918,N_13265,N_13948);
and U15919 (N_15919,N_12235,N_12294);
or U15920 (N_15920,N_13424,N_12010);
nand U15921 (N_15921,N_12760,N_12997);
nor U15922 (N_15922,N_12376,N_12919);
xor U15923 (N_15923,N_12196,N_13556);
xnor U15924 (N_15924,N_13721,N_12250);
nor U15925 (N_15925,N_13792,N_13908);
and U15926 (N_15926,N_12090,N_13396);
or U15927 (N_15927,N_13714,N_13391);
xor U15928 (N_15928,N_12148,N_12620);
nor U15929 (N_15929,N_12178,N_12857);
xnor U15930 (N_15930,N_13135,N_12184);
xor U15931 (N_15931,N_12504,N_13660);
nand U15932 (N_15932,N_12731,N_13304);
and U15933 (N_15933,N_12520,N_12130);
and U15934 (N_15934,N_13102,N_13190);
or U15935 (N_15935,N_12141,N_12590);
or U15936 (N_15936,N_12274,N_13864);
nand U15937 (N_15937,N_13927,N_13258);
nor U15938 (N_15938,N_12875,N_12461);
or U15939 (N_15939,N_13712,N_13900);
nor U15940 (N_15940,N_13857,N_13629);
or U15941 (N_15941,N_13173,N_12314);
or U15942 (N_15942,N_12908,N_12886);
or U15943 (N_15943,N_12234,N_12554);
xor U15944 (N_15944,N_12983,N_12340);
nand U15945 (N_15945,N_13783,N_12197);
xnor U15946 (N_15946,N_13759,N_12919);
nand U15947 (N_15947,N_13287,N_12763);
and U15948 (N_15948,N_12099,N_12791);
nand U15949 (N_15949,N_13506,N_13787);
nor U15950 (N_15950,N_13465,N_13578);
nand U15951 (N_15951,N_12850,N_13008);
and U15952 (N_15952,N_12565,N_13365);
and U15953 (N_15953,N_12017,N_12253);
xnor U15954 (N_15954,N_12351,N_13480);
nand U15955 (N_15955,N_13715,N_13986);
xnor U15956 (N_15956,N_12077,N_13106);
nand U15957 (N_15957,N_12024,N_13831);
nand U15958 (N_15958,N_13201,N_12803);
or U15959 (N_15959,N_12793,N_12291);
or U15960 (N_15960,N_12624,N_13436);
xnor U15961 (N_15961,N_13590,N_13886);
or U15962 (N_15962,N_13891,N_13993);
xor U15963 (N_15963,N_12183,N_13892);
xnor U15964 (N_15964,N_12278,N_12026);
nor U15965 (N_15965,N_13508,N_12220);
or U15966 (N_15966,N_13915,N_13355);
nor U15967 (N_15967,N_12040,N_13970);
xor U15968 (N_15968,N_13531,N_12074);
and U15969 (N_15969,N_12562,N_12875);
and U15970 (N_15970,N_12391,N_13216);
nor U15971 (N_15971,N_12323,N_12461);
nor U15972 (N_15972,N_13506,N_13452);
and U15973 (N_15973,N_12008,N_13075);
xor U15974 (N_15974,N_13567,N_13133);
nand U15975 (N_15975,N_12408,N_13690);
and U15976 (N_15976,N_13574,N_13826);
nand U15977 (N_15977,N_13368,N_12266);
nand U15978 (N_15978,N_13263,N_13217);
xor U15979 (N_15979,N_13967,N_13291);
and U15980 (N_15980,N_12222,N_12776);
nand U15981 (N_15981,N_12361,N_13739);
xnor U15982 (N_15982,N_13866,N_12772);
nand U15983 (N_15983,N_13119,N_12413);
or U15984 (N_15984,N_13474,N_12452);
nor U15985 (N_15985,N_12218,N_13311);
and U15986 (N_15986,N_13267,N_13894);
nor U15987 (N_15987,N_12567,N_13179);
or U15988 (N_15988,N_12284,N_12475);
or U15989 (N_15989,N_13735,N_13110);
nor U15990 (N_15990,N_12436,N_12641);
nand U15991 (N_15991,N_13076,N_13097);
nor U15992 (N_15992,N_12493,N_13140);
nand U15993 (N_15993,N_12079,N_13698);
nand U15994 (N_15994,N_13320,N_12606);
xor U15995 (N_15995,N_12014,N_13151);
or U15996 (N_15996,N_12635,N_12178);
xnor U15997 (N_15997,N_13777,N_13523);
nand U15998 (N_15998,N_13266,N_12996);
and U15999 (N_15999,N_12060,N_12842);
xnor U16000 (N_16000,N_15956,N_14582);
and U16001 (N_16001,N_14735,N_14307);
nor U16002 (N_16002,N_15892,N_15242);
and U16003 (N_16003,N_14223,N_15780);
or U16004 (N_16004,N_15737,N_15464);
nand U16005 (N_16005,N_14451,N_15981);
nor U16006 (N_16006,N_15158,N_14071);
xnor U16007 (N_16007,N_15214,N_15059);
nand U16008 (N_16008,N_15677,N_15785);
xor U16009 (N_16009,N_15665,N_14885);
or U16010 (N_16010,N_15924,N_15832);
nor U16011 (N_16011,N_15592,N_14007);
xnor U16012 (N_16012,N_15836,N_15084);
or U16013 (N_16013,N_15881,N_15575);
and U16014 (N_16014,N_15484,N_15843);
and U16015 (N_16015,N_15585,N_14369);
nand U16016 (N_16016,N_15952,N_15531);
nand U16017 (N_16017,N_14993,N_15926);
xor U16018 (N_16018,N_14667,N_14992);
nor U16019 (N_16019,N_15745,N_15339);
and U16020 (N_16020,N_14415,N_14458);
or U16021 (N_16021,N_14937,N_15958);
or U16022 (N_16022,N_14665,N_15624);
or U16023 (N_16023,N_14359,N_15359);
nand U16024 (N_16024,N_14777,N_15269);
nand U16025 (N_16025,N_14465,N_14845);
xor U16026 (N_16026,N_15812,N_15847);
xnor U16027 (N_16027,N_14535,N_14767);
nor U16028 (N_16028,N_15860,N_15810);
xor U16029 (N_16029,N_14524,N_14076);
and U16030 (N_16030,N_14644,N_15577);
xnor U16031 (N_16031,N_15323,N_14306);
nand U16032 (N_16032,N_14343,N_14783);
nand U16033 (N_16033,N_15408,N_15070);
xor U16034 (N_16034,N_14599,N_15641);
nand U16035 (N_16035,N_14959,N_14372);
xor U16036 (N_16036,N_15985,N_14760);
nand U16037 (N_16037,N_14827,N_15186);
nand U16038 (N_16038,N_15420,N_15177);
nor U16039 (N_16039,N_14388,N_14921);
and U16040 (N_16040,N_14883,N_14002);
xor U16041 (N_16041,N_14635,N_14298);
and U16042 (N_16042,N_15324,N_15148);
nor U16043 (N_16043,N_14354,N_14390);
or U16044 (N_16044,N_14098,N_14420);
and U16045 (N_16045,N_14014,N_14593);
nand U16046 (N_16046,N_15435,N_14126);
or U16047 (N_16047,N_14199,N_14539);
or U16048 (N_16048,N_15698,N_14269);
and U16049 (N_16049,N_14419,N_15544);
nor U16050 (N_16050,N_15290,N_14036);
xnor U16051 (N_16051,N_15130,N_15009);
nand U16052 (N_16052,N_15377,N_14632);
nand U16053 (N_16053,N_15944,N_14443);
and U16054 (N_16054,N_14505,N_14228);
or U16055 (N_16055,N_14615,N_15425);
nor U16056 (N_16056,N_15440,N_14649);
and U16057 (N_16057,N_14942,N_15394);
or U16058 (N_16058,N_14965,N_15568);
nor U16059 (N_16059,N_15266,N_15416);
nand U16060 (N_16060,N_15548,N_15505);
nand U16061 (N_16061,N_14679,N_15406);
xor U16062 (N_16062,N_14797,N_15470);
xor U16063 (N_16063,N_15675,N_14472);
xnor U16064 (N_16064,N_14195,N_15795);
nor U16065 (N_16065,N_14448,N_14185);
or U16066 (N_16066,N_14802,N_15368);
or U16067 (N_16067,N_14115,N_15274);
and U16068 (N_16068,N_15788,N_15991);
nor U16069 (N_16069,N_14363,N_15529);
xnor U16070 (N_16070,N_15462,N_14313);
xor U16071 (N_16071,N_15216,N_15864);
xnor U16072 (N_16072,N_14880,N_14281);
or U16073 (N_16073,N_14967,N_15465);
xor U16074 (N_16074,N_15543,N_15581);
xnor U16075 (N_16075,N_15199,N_15128);
nand U16076 (N_16076,N_14863,N_14603);
nand U16077 (N_16077,N_14670,N_15508);
and U16078 (N_16078,N_15198,N_15649);
and U16079 (N_16079,N_14280,N_15532);
or U16080 (N_16080,N_15931,N_14994);
or U16081 (N_16081,N_14692,N_15626);
xnor U16082 (N_16082,N_14353,N_15671);
nor U16083 (N_16083,N_15871,N_15014);
or U16084 (N_16084,N_14858,N_14540);
and U16085 (N_16085,N_14497,N_15438);
nor U16086 (N_16086,N_15619,N_15397);
xor U16087 (N_16087,N_15280,N_15687);
or U16088 (N_16088,N_15841,N_14924);
nor U16089 (N_16089,N_15948,N_15605);
nand U16090 (N_16090,N_15026,N_14733);
nand U16091 (N_16091,N_15943,N_15413);
and U16092 (N_16092,N_15000,N_15825);
nand U16093 (N_16093,N_14500,N_14439);
and U16094 (N_16094,N_14013,N_14413);
nand U16095 (N_16095,N_15478,N_15371);
xor U16096 (N_16096,N_15419,N_15335);
nor U16097 (N_16097,N_15858,N_15630);
nand U16098 (N_16098,N_14889,N_14722);
nand U16099 (N_16099,N_15110,N_15923);
xnor U16100 (N_16100,N_15775,N_14042);
nor U16101 (N_16101,N_15264,N_15571);
xor U16102 (N_16102,N_14516,N_15092);
or U16103 (N_16103,N_14957,N_14550);
xnor U16104 (N_16104,N_14197,N_14918);
or U16105 (N_16105,N_15814,N_14303);
and U16106 (N_16106,N_14143,N_15082);
or U16107 (N_16107,N_14652,N_15513);
and U16108 (N_16108,N_15160,N_15447);
nand U16109 (N_16109,N_15297,N_15977);
xor U16110 (N_16110,N_15720,N_14188);
or U16111 (N_16111,N_15551,N_15352);
xnor U16112 (N_16112,N_14835,N_14431);
nand U16113 (N_16113,N_14435,N_14494);
and U16114 (N_16114,N_15786,N_14395);
or U16115 (N_16115,N_14606,N_14888);
nor U16116 (N_16116,N_15819,N_14460);
or U16117 (N_16117,N_15631,N_15247);
xnor U16118 (N_16118,N_14948,N_15121);
or U16119 (N_16119,N_15678,N_14341);
xor U16120 (N_16120,N_15370,N_15763);
or U16121 (N_16121,N_15719,N_15197);
or U16122 (N_16122,N_15741,N_14092);
xnor U16123 (N_16123,N_14962,N_15879);
and U16124 (N_16124,N_15751,N_14794);
and U16125 (N_16125,N_14689,N_14160);
or U16126 (N_16126,N_14850,N_14062);
xnor U16127 (N_16127,N_14044,N_15710);
xnor U16128 (N_16128,N_14252,N_15354);
xor U16129 (N_16129,N_14159,N_14742);
nor U16130 (N_16130,N_14112,N_15845);
xnor U16131 (N_16131,N_14805,N_14567);
nand U16132 (N_16132,N_14474,N_15385);
nor U16133 (N_16133,N_14440,N_14611);
nand U16134 (N_16134,N_14244,N_14816);
or U16135 (N_16135,N_14004,N_15765);
xnor U16136 (N_16136,N_15855,N_15898);
and U16137 (N_16137,N_15972,N_15866);
xor U16138 (N_16138,N_14301,N_14351);
nor U16139 (N_16139,N_15342,N_14236);
and U16140 (N_16140,N_15590,N_15584);
and U16141 (N_16141,N_15970,N_15444);
xor U16142 (N_16142,N_14642,N_15591);
or U16143 (N_16143,N_14607,N_15932);
xnor U16144 (N_16144,N_14952,N_14018);
nand U16145 (N_16145,N_15344,N_14400);
xor U16146 (N_16146,N_14067,N_14776);
nand U16147 (N_16147,N_15195,N_14931);
nand U16148 (N_16148,N_15143,N_15100);
and U16149 (N_16149,N_15697,N_15033);
or U16150 (N_16150,N_15383,N_14358);
nor U16151 (N_16151,N_15973,N_14614);
or U16152 (N_16152,N_15439,N_15379);
nor U16153 (N_16153,N_14789,N_14108);
and U16154 (N_16154,N_15363,N_14170);
nand U16155 (N_16155,N_15455,N_15979);
nor U16156 (N_16156,N_14140,N_14902);
nor U16157 (N_16157,N_14545,N_14374);
or U16158 (N_16158,N_14150,N_15011);
and U16159 (N_16159,N_15486,N_14547);
xnor U16160 (N_16160,N_14283,N_15052);
or U16161 (N_16161,N_14740,N_14501);
and U16162 (N_16162,N_15034,N_15154);
and U16163 (N_16163,N_15402,N_14565);
xor U16164 (N_16164,N_14158,N_14947);
and U16165 (N_16165,N_14037,N_14484);
nor U16166 (N_16166,N_15119,N_15752);
nor U16167 (N_16167,N_14254,N_15579);
or U16168 (N_16168,N_14741,N_15854);
and U16169 (N_16169,N_15239,N_14394);
or U16170 (N_16170,N_15491,N_15172);
or U16171 (N_16171,N_14914,N_14034);
nor U16172 (N_16172,N_14426,N_15246);
or U16173 (N_16173,N_15968,N_14174);
and U16174 (N_16174,N_14437,N_14398);
or U16175 (N_16175,N_14385,N_14754);
and U16176 (N_16176,N_14258,N_14983);
nor U16177 (N_16177,N_14862,N_14446);
nor U16178 (N_16178,N_15314,N_14790);
or U16179 (N_16179,N_15209,N_14799);
and U16180 (N_16180,N_14595,N_14731);
xor U16181 (N_16181,N_14519,N_14941);
nand U16182 (N_16182,N_15735,N_14526);
xnor U16183 (N_16183,N_14218,N_15840);
nand U16184 (N_16184,N_15602,N_14859);
and U16185 (N_16185,N_14318,N_15999);
nor U16186 (N_16186,N_14093,N_14536);
nor U16187 (N_16187,N_14459,N_15021);
or U16188 (N_16188,N_15906,N_15429);
or U16189 (N_16189,N_14659,N_15600);
nand U16190 (N_16190,N_14230,N_15389);
nand U16191 (N_16191,N_14422,N_14651);
nand U16192 (N_16192,N_14989,N_14806);
xnor U16193 (N_16193,N_15986,N_15567);
or U16194 (N_16194,N_14687,N_14700);
nand U16195 (N_16195,N_15882,N_14738);
nand U16196 (N_16196,N_14495,N_15768);
and U16197 (N_16197,N_15019,N_14339);
and U16198 (N_16198,N_14290,N_14909);
or U16199 (N_16199,N_14620,N_14214);
nor U16200 (N_16200,N_14096,N_15120);
or U16201 (N_16201,N_14421,N_14559);
nand U16202 (N_16202,N_15623,N_15450);
or U16203 (N_16203,N_14911,N_14424);
and U16204 (N_16204,N_14558,N_14148);
xnor U16205 (N_16205,N_14409,N_15949);
xor U16206 (N_16206,N_14499,N_15899);
nand U16207 (N_16207,N_15791,N_15813);
nor U16208 (N_16208,N_15807,N_14721);
or U16209 (N_16209,N_15181,N_15163);
and U16210 (N_16210,N_15200,N_14139);
xnor U16211 (N_16211,N_14674,N_14407);
nand U16212 (N_16212,N_14999,N_15682);
nor U16213 (N_16213,N_15422,N_14015);
nand U16214 (N_16214,N_15330,N_14685);
nand U16215 (N_16215,N_15707,N_15217);
xnor U16216 (N_16216,N_15736,N_14908);
nor U16217 (N_16217,N_15524,N_15661);
xor U16218 (N_16218,N_14376,N_14200);
nand U16219 (N_16219,N_14624,N_14661);
xnor U16220 (N_16220,N_14276,N_14346);
or U16221 (N_16221,N_14513,N_15477);
xnor U16222 (N_16222,N_15040,N_15012);
or U16223 (N_16223,N_14177,N_15129);
or U16224 (N_16224,N_15222,N_14479);
nand U16225 (N_16225,N_15310,N_15690);
or U16226 (N_16226,N_15495,N_14430);
xor U16227 (N_16227,N_15912,N_15069);
nand U16228 (N_16228,N_15224,N_15145);
xnor U16229 (N_16229,N_14896,N_15925);
or U16230 (N_16230,N_14824,N_15504);
nor U16231 (N_16231,N_14563,N_14489);
or U16232 (N_16232,N_15347,N_14775);
nor U16233 (N_16233,N_15565,N_14091);
xor U16234 (N_16234,N_14423,N_14755);
nand U16235 (N_16235,N_15828,N_15817);
nor U16236 (N_16236,N_15111,N_14347);
nor U16237 (N_16237,N_15555,N_15771);
xor U16238 (N_16238,N_15207,N_14444);
or U16239 (N_16239,N_15588,N_15095);
xor U16240 (N_16240,N_15421,N_14899);
and U16241 (N_16241,N_15920,N_14502);
nand U16242 (N_16242,N_15715,N_14566);
nor U16243 (N_16243,N_15051,N_15769);
or U16244 (N_16244,N_15941,N_14630);
xor U16245 (N_16245,N_15928,N_14712);
nor U16246 (N_16246,N_14569,N_14521);
nor U16247 (N_16247,N_15430,N_15183);
nor U16248 (N_16248,N_14345,N_15103);
and U16249 (N_16249,N_15168,N_15867);
and U16250 (N_16250,N_14552,N_15311);
nor U16251 (N_16251,N_15696,N_15512);
nand U16252 (N_16252,N_14976,N_14848);
or U16253 (N_16253,N_14627,N_15260);
or U16254 (N_16254,N_15960,N_14001);
and U16255 (N_16255,N_14382,N_14579);
and U16256 (N_16256,N_14145,N_14934);
xnor U16257 (N_16257,N_15896,N_15329);
nand U16258 (N_16258,N_14450,N_15996);
xnor U16259 (N_16259,N_15929,N_15407);
or U16260 (N_16260,N_14955,N_15079);
and U16261 (N_16261,N_14231,N_15176);
nand U16262 (N_16262,N_15445,N_15270);
or U16263 (N_16263,N_15456,N_15815);
xor U16264 (N_16264,N_15127,N_15793);
or U16265 (N_16265,N_15695,N_15672);
xor U16266 (N_16266,N_14168,N_14012);
nand U16267 (N_16267,N_15085,N_15481);
and U16268 (N_16268,N_15441,N_15794);
nor U16269 (N_16269,N_14930,N_15559);
xnor U16270 (N_16270,N_15490,N_15284);
xnor U16271 (N_16271,N_15865,N_14299);
nor U16272 (N_16272,N_15656,N_14541);
xor U16273 (N_16273,N_15534,N_14720);
nand U16274 (N_16274,N_14207,N_14074);
nand U16275 (N_16275,N_14672,N_14662);
nand U16276 (N_16276,N_15395,N_15541);
and U16277 (N_16277,N_14528,N_14602);
and U16278 (N_16278,N_15487,N_14527);
nand U16279 (N_16279,N_15617,N_14986);
nand U16280 (N_16280,N_14923,N_15171);
nand U16281 (N_16281,N_14633,N_15862);
nand U16282 (N_16282,N_14006,N_15992);
and U16283 (N_16283,N_14260,N_14716);
nor U16284 (N_16284,N_15073,N_14912);
xnor U16285 (N_16285,N_14548,N_15004);
or U16286 (N_16286,N_15404,N_15243);
and U16287 (N_16287,N_14564,N_14193);
xnor U16288 (N_16288,N_14153,N_15063);
xnor U16289 (N_16289,N_15538,N_14393);
or U16290 (N_16290,N_14945,N_15337);
nor U16291 (N_16291,N_15333,N_15888);
nor U16292 (N_16292,N_14568,N_15560);
nand U16293 (N_16293,N_14879,N_14471);
or U16294 (N_16294,N_14371,N_14123);
nand U16295 (N_16295,N_14154,N_14988);
xnor U16296 (N_16296,N_15753,N_14752);
nor U16297 (N_16297,N_15663,N_15834);
nand U16298 (N_16298,N_15152,N_14765);
nand U16299 (N_16299,N_15253,N_15552);
nor U16300 (N_16300,N_14588,N_15703);
nor U16301 (N_16301,N_15692,N_15578);
xnor U16302 (N_16302,N_15473,N_15277);
or U16303 (N_16303,N_15666,N_14637);
nand U16304 (N_16304,N_15178,N_14759);
nand U16305 (N_16305,N_14585,N_14979);
nor U16306 (N_16306,N_15468,N_14643);
xor U16307 (N_16307,N_14537,N_15414);
and U16308 (N_16308,N_14312,N_14613);
or U16309 (N_16309,N_14028,N_14723);
xor U16310 (N_16310,N_15963,N_15151);
nand U16311 (N_16311,N_14617,N_14938);
xnor U16312 (N_16312,N_14256,N_14830);
or U16313 (N_16313,N_15112,N_14708);
or U16314 (N_16314,N_14881,N_15637);
nand U16315 (N_16315,N_15709,N_15674);
nand U16316 (N_16316,N_14825,N_15002);
nor U16317 (N_16317,N_15366,N_15203);
nand U16318 (N_16318,N_15165,N_14717);
or U16319 (N_16319,N_15718,N_15915);
nand U16320 (N_16320,N_15770,N_15107);
and U16321 (N_16321,N_15787,N_14221);
nand U16322 (N_16322,N_14427,N_14151);
or U16323 (N_16323,N_15806,N_15460);
and U16324 (N_16324,N_15288,N_14784);
xnor U16325 (N_16325,N_14629,N_15679);
nor U16326 (N_16326,N_15459,N_15772);
xor U16327 (N_16327,N_14699,N_14447);
nor U16328 (N_16328,N_14077,N_15472);
nor U16329 (N_16329,N_14946,N_15937);
nor U16330 (N_16330,N_15933,N_15268);
nor U16331 (N_16331,N_15102,N_15667);
nor U16332 (N_16332,N_14250,N_14257);
nand U16333 (N_16333,N_15957,N_15580);
or U16334 (N_16334,N_14625,N_15146);
or U16335 (N_16335,N_15137,N_15756);
nand U16336 (N_16336,N_14102,N_14267);
nand U16337 (N_16337,N_15349,N_14972);
or U16338 (N_16338,N_15657,N_15283);
and U16339 (N_16339,N_14416,N_15766);
nand U16340 (N_16340,N_14043,N_15080);
or U16341 (N_16341,N_14073,N_15650);
xor U16342 (N_16342,N_15648,N_15976);
xnor U16343 (N_16343,N_14810,N_15939);
xnor U16344 (N_16344,N_14654,N_15028);
xor U16345 (N_16345,N_15616,N_14308);
xor U16346 (N_16346,N_14297,N_15849);
nand U16347 (N_16347,N_15811,N_15727);
and U16348 (N_16348,N_14414,N_15159);
nand U16349 (N_16349,N_14335,N_15747);
nor U16350 (N_16350,N_15842,N_15607);
nor U16351 (N_16351,N_15655,N_14890);
nand U16352 (N_16352,N_15259,N_14865);
or U16353 (N_16353,N_14828,N_14478);
nand U16354 (N_16354,N_14461,N_15360);
and U16355 (N_16355,N_15192,N_14523);
and U16356 (N_16356,N_14204,N_14184);
xor U16357 (N_16357,N_14833,N_15045);
nor U16358 (N_16358,N_15826,N_15320);
or U16359 (N_16359,N_14482,N_15184);
or U16360 (N_16360,N_15016,N_14418);
nand U16361 (N_16361,N_15803,N_14601);
nor U16362 (N_16362,N_15762,N_14476);
or U16363 (N_16363,N_15759,N_15820);
nor U16364 (N_16364,N_14048,N_15113);
and U16365 (N_16365,N_15036,N_15653);
or U16366 (N_16366,N_15098,N_15488);
nand U16367 (N_16367,N_15615,N_14453);
xor U16368 (N_16368,N_14905,N_15302);
and U16369 (N_16369,N_15308,N_15466);
nor U16370 (N_16370,N_15015,N_15701);
xor U16371 (N_16371,N_15437,N_14610);
nor U16372 (N_16372,N_14769,N_14876);
nor U16373 (N_16373,N_14097,N_15914);
xnor U16374 (N_16374,N_14340,N_15562);
or U16375 (N_16375,N_15273,N_14586);
nand U16376 (N_16376,N_14336,N_15554);
nand U16377 (N_16377,N_15646,N_14329);
and U16378 (N_16378,N_14406,N_14853);
nand U16379 (N_16379,N_14838,N_14025);
nand U16380 (N_16380,N_15878,N_15797);
nand U16381 (N_16381,N_15285,N_15729);
nor U16382 (N_16382,N_15528,N_15569);
or U16383 (N_16383,N_14818,N_15367);
nand U16384 (N_16384,N_15060,N_14491);
and U16385 (N_16385,N_15426,N_14518);
nand U16386 (N_16386,N_14141,N_15927);
xor U16387 (N_16387,N_14556,N_15993);
xnor U16388 (N_16388,N_14750,N_15068);
and U16389 (N_16389,N_14974,N_15921);
nor U16390 (N_16390,N_14366,N_14793);
xor U16391 (N_16391,N_14919,N_14688);
nor U16392 (N_16392,N_15506,N_15890);
nand U16393 (N_16393,N_15779,N_15256);
nand U16394 (N_16394,N_14984,N_14240);
and U16395 (N_16395,N_14739,N_15221);
nor U16396 (N_16396,N_14925,N_14234);
or U16397 (N_16397,N_14259,N_14105);
nor U16398 (N_16398,N_15700,N_14101);
and U16399 (N_16399,N_14412,N_15942);
and U16400 (N_16400,N_14323,N_15353);
or U16401 (N_16401,N_14287,N_15918);
or U16402 (N_16402,N_15078,N_15405);
nand U16403 (N_16403,N_15749,N_14330);
and U16404 (N_16404,N_14530,N_14991);
or U16405 (N_16405,N_15684,N_14000);
xor U16406 (N_16406,N_15180,N_15411);
nor U16407 (N_16407,N_14773,N_15652);
and U16408 (N_16408,N_14996,N_14581);
and U16409 (N_16409,N_15566,N_15583);
and U16410 (N_16410,N_15475,N_15587);
or U16411 (N_16411,N_14264,N_14864);
and U16412 (N_16412,N_14873,N_14008);
or U16413 (N_16413,N_15453,N_15075);
or U16414 (N_16414,N_15190,N_14094);
nand U16415 (N_16415,N_15851,N_14970);
or U16416 (N_16416,N_15248,N_15744);
or U16417 (N_16417,N_14171,N_15668);
nor U16418 (N_16418,N_15895,N_15317);
xnor U16419 (N_16419,N_15790,N_15123);
nand U16420 (N_16420,N_15090,N_15232);
or U16421 (N_16421,N_15714,N_15844);
or U16422 (N_16422,N_15193,N_14247);
and U16423 (N_16423,N_15573,N_15289);
xor U16424 (N_16424,N_14238,N_14576);
nand U16425 (N_16425,N_15194,N_15234);
nor U16426 (N_16426,N_14529,N_15332);
or U16427 (N_16427,N_15013,N_14026);
and U16428 (N_16428,N_15091,N_15106);
and U16429 (N_16429,N_14109,N_14035);
and U16430 (N_16430,N_14682,N_14227);
nor U16431 (N_16431,N_14737,N_14695);
or U16432 (N_16432,N_14626,N_15556);
or U16433 (N_16433,N_15046,N_15877);
nor U16434 (N_16434,N_15778,N_15596);
and U16435 (N_16435,N_14083,N_14373);
xor U16436 (N_16436,N_14401,N_15257);
and U16437 (N_16437,N_15427,N_15162);
or U16438 (N_16438,N_14127,N_14697);
xor U16439 (N_16439,N_15988,N_14445);
nand U16440 (N_16440,N_15699,N_15231);
nand U16441 (N_16441,N_15271,N_15237);
nor U16442 (N_16442,N_15537,N_14823);
xor U16443 (N_16443,N_15139,N_14022);
xor U16444 (N_16444,N_15919,N_14063);
nand U16445 (N_16445,N_14877,N_15117);
and U16446 (N_16446,N_14971,N_14634);
nand U16447 (N_16447,N_15185,N_15276);
nor U16448 (N_16448,N_14320,N_15831);
xnor U16449 (N_16449,N_14683,N_14844);
nand U16450 (N_16450,N_14121,N_14255);
xor U16451 (N_16451,N_15206,N_15022);
or U16452 (N_16452,N_14161,N_15801);
and U16453 (N_16453,N_15392,N_14872);
or U16454 (N_16454,N_15293,N_15328);
xor U16455 (N_16455,N_15156,N_15010);
xnor U16456 (N_16456,N_14842,N_14288);
xnor U16457 (N_16457,N_14144,N_15035);
nand U16458 (N_16458,N_15294,N_15066);
and U16459 (N_16459,N_15558,N_15030);
nand U16460 (N_16460,N_15664,N_14130);
nand U16461 (N_16461,N_15526,N_14981);
nor U16462 (N_16462,N_15415,N_14506);
and U16463 (N_16463,N_15296,N_14191);
nand U16464 (N_16464,N_14978,N_15983);
nand U16465 (N_16465,N_14829,N_15255);
nand U16466 (N_16466,N_14120,N_14949);
or U16467 (N_16467,N_14243,N_14295);
nand U16468 (N_16468,N_15767,N_14428);
or U16469 (N_16469,N_14782,N_15691);
nor U16470 (N_16470,N_15856,N_15547);
or U16471 (N_16471,N_14619,N_15125);
nand U16472 (N_16472,N_15595,N_14210);
or U16473 (N_16473,N_14657,N_14169);
xnor U16474 (N_16474,N_14932,N_14337);
and U16475 (N_16475,N_14886,N_15686);
xor U16476 (N_16476,N_15822,N_15612);
xnor U16477 (N_16477,N_14411,N_14532);
nor U16478 (N_16478,N_15443,N_14768);
nor U16479 (N_16479,N_15093,N_14892);
and U16480 (N_16480,N_15238,N_14761);
or U16481 (N_16481,N_15018,N_15776);
xor U16482 (N_16482,N_14819,N_15673);
and U16483 (N_16483,N_14709,N_15461);
xor U16484 (N_16484,N_15997,N_15292);
or U16485 (N_16485,N_15542,N_15062);
nand U16486 (N_16486,N_14294,N_15334);
or U16487 (N_16487,N_14289,N_15469);
and U16488 (N_16488,N_14003,N_14272);
nand U16489 (N_16489,N_14087,N_15638);
and U16490 (N_16490,N_15142,N_14577);
xnor U16491 (N_16491,N_14047,N_15399);
or U16492 (N_16492,N_15904,N_15809);
or U16493 (N_16493,N_14660,N_15319);
or U16494 (N_16494,N_14462,N_14747);
or U16495 (N_16495,N_14457,N_14557);
nor U16496 (N_16496,N_15628,N_14808);
nand U16497 (N_16497,N_14714,N_15312);
and U16498 (N_16498,N_15706,N_14349);
nor U16499 (N_16499,N_15321,N_15048);
or U16500 (N_16500,N_15676,N_14786);
nor U16501 (N_16501,N_14904,N_15507);
or U16502 (N_16502,N_15974,N_14669);
xor U16503 (N_16503,N_14417,N_15604);
nand U16504 (N_16504,N_14039,N_14935);
nand U16505 (N_16505,N_14095,N_14080);
nand U16506 (N_16506,N_14246,N_14870);
or U16507 (N_16507,N_14592,N_14609);
xor U16508 (N_16508,N_14762,N_15743);
or U16509 (N_16509,N_15777,N_15951);
xor U16510 (N_16510,N_14522,N_14425);
nor U16511 (N_16511,N_14404,N_14726);
or U16512 (N_16512,N_14915,N_14032);
nand U16513 (N_16513,N_14966,N_14673);
nand U16514 (N_16514,N_15728,N_14379);
or U16515 (N_16515,N_14392,N_15510);
xnor U16516 (N_16516,N_14176,N_14384);
or U16517 (N_16517,N_14334,N_15545);
nand U16518 (N_16518,N_14391,N_15410);
xor U16519 (N_16519,N_15227,N_14846);
nor U16520 (N_16520,N_14175,N_14009);
xnor U16521 (N_16521,N_15557,N_15886);
nor U16522 (N_16522,N_15982,N_14046);
and U16523 (N_16523,N_15829,N_14758);
xor U16524 (N_16524,N_15846,N_14855);
nand U16525 (N_16525,N_15436,N_15509);
nor U16526 (N_16526,N_14725,N_14106);
nor U16527 (N_16527,N_14263,N_15900);
and U16528 (N_16528,N_14572,N_15848);
and U16529 (N_16529,N_15739,N_14940);
xor U16530 (N_16530,N_15007,N_15109);
nor U16531 (N_16531,N_14597,N_15136);
nor U16532 (N_16532,N_14675,N_14854);
or U16533 (N_16533,N_15659,N_14676);
xnor U16534 (N_16534,N_15563,N_15304);
nor U16535 (N_16535,N_15356,N_14245);
xor U16536 (N_16536,N_15907,N_14326);
nor U16537 (N_16537,N_15250,N_14389);
or U16538 (N_16538,N_14894,N_15147);
xnor U16539 (N_16539,N_14114,N_14157);
nor U16540 (N_16540,N_15140,N_15116);
nor U16541 (N_16541,N_14798,N_15230);
nor U16542 (N_16542,N_15633,N_15527);
nor U16543 (N_16543,N_14555,N_15351);
nand U16544 (N_16544,N_15229,N_15476);
nor U16545 (N_16545,N_15621,N_15808);
xnor U16546 (N_16546,N_14405,N_15705);
nand U16547 (N_16547,N_14190,N_14059);
xnor U16548 (N_16548,N_15313,N_15967);
nand U16549 (N_16549,N_14005,N_15025);
or U16550 (N_16550,N_14533,N_14045);
xor U16551 (N_16551,N_15235,N_14311);
nor U16552 (N_16552,N_14578,N_15432);
nor U16553 (N_16553,N_14977,N_14958);
or U16554 (N_16554,N_15029,N_15634);
xnor U16555 (N_16555,N_15083,N_15774);
nor U16556 (N_16556,N_15713,N_15622);
or U16557 (N_16557,N_15969,N_14847);
xor U16558 (N_16558,N_15261,N_14694);
nor U16559 (N_16559,N_14814,N_15837);
nor U16560 (N_16560,N_14647,N_14100);
and U16561 (N_16561,N_14352,N_14348);
and U16562 (N_16562,N_15375,N_14746);
nor U16563 (N_16563,N_15821,N_15446);
or U16564 (N_16564,N_14693,N_14253);
nand U16565 (N_16565,N_14950,N_14317);
xnor U16566 (N_16566,N_15252,N_15994);
nor U16567 (N_16567,N_15835,N_15975);
nand U16568 (N_16568,N_15761,N_14205);
xor U16569 (N_16569,N_14402,N_15218);
or U16570 (N_16570,N_15220,N_14628);
nand U16571 (N_16571,N_14510,N_15511);
nand U16572 (N_16572,N_15384,N_14498);
xor U16573 (N_16573,N_14162,N_14328);
and U16574 (N_16574,N_14270,N_14142);
nor U16575 (N_16575,N_14213,N_15482);
and U16576 (N_16576,N_15228,N_15594);
nor U16577 (N_16577,N_14639,N_14490);
nand U16578 (N_16578,N_15149,N_14279);
and U16579 (N_16579,N_14757,N_14189);
xor U16580 (N_16580,N_14975,N_15731);
or U16581 (N_16581,N_15042,N_15564);
nor U16582 (N_16582,N_15708,N_14727);
nand U16583 (N_16583,N_15516,N_15364);
nor U16584 (N_16584,N_14364,N_14408);
nor U16585 (N_16585,N_14953,N_15361);
or U16586 (N_16586,N_14878,N_14365);
and U16587 (N_16587,N_15205,N_14748);
and U16588 (N_16588,N_14743,N_14655);
nor U16589 (N_16589,N_14903,N_15175);
xor U16590 (N_16590,N_14963,N_14487);
and U16591 (N_16591,N_15730,N_15804);
and U16592 (N_16592,N_15689,N_14186);
and U16593 (N_16593,N_15393,N_14900);
xnor U16594 (N_16594,N_14871,N_14812);
or U16595 (N_16595,N_15077,N_14362);
and U16596 (N_16596,N_15345,N_14271);
xnor U16597 (N_16597,N_14520,N_14172);
nor U16598 (N_16598,N_14248,N_14442);
nor U16599 (N_16599,N_15883,N_15182);
nand U16600 (N_16600,N_14485,N_14954);
nor U16601 (N_16601,N_14232,N_15114);
or U16602 (N_16602,N_15325,N_15945);
xor U16603 (N_16603,N_15704,N_15057);
and U16604 (N_16604,N_15189,N_15346);
xnor U16605 (N_16605,N_15824,N_14690);
nor U16606 (N_16606,N_15964,N_14982);
xor U16607 (N_16607,N_14274,N_14113);
xnor U16608 (N_16608,N_14286,N_14466);
xnor U16609 (N_16609,N_15398,N_15880);
and U16610 (N_16610,N_14261,N_14060);
and U16611 (N_16611,N_15173,N_15857);
nand U16612 (N_16612,N_15187,N_14711);
nor U16613 (N_16613,N_14898,N_14082);
nand U16614 (N_16614,N_14821,N_15887);
xnor U16615 (N_16615,N_14861,N_14017);
and U16616 (N_16616,N_15212,N_14893);
and U16617 (N_16617,N_14473,N_15910);
or U16618 (N_16618,N_14265,N_14696);
or U16619 (N_16619,N_15732,N_14396);
and U16620 (N_16620,N_15076,N_15097);
nor U16621 (N_16621,N_15764,N_14511);
or U16622 (N_16622,N_14192,N_15533);
nand U16623 (N_16623,N_14701,N_14496);
and U16624 (N_16624,N_14107,N_15167);
or U16625 (N_16625,N_15053,N_14691);
nand U16626 (N_16626,N_15299,N_15307);
nand U16627 (N_16627,N_14211,N_15303);
nand U16628 (N_16628,N_15380,N_15463);
nand U16629 (N_16629,N_14324,N_14070);
nor U16630 (N_16630,N_14222,N_15433);
xor U16631 (N_16631,N_14780,N_14021);
and U16632 (N_16632,N_15724,N_15990);
xnor U16633 (N_16633,N_14843,N_14636);
and U16634 (N_16634,N_14481,N_14718);
xor U16635 (N_16635,N_15315,N_15434);
or U16636 (N_16636,N_15418,N_14111);
xnor U16637 (N_16637,N_15947,N_15869);
nand U16638 (N_16638,N_15830,N_14350);
and U16639 (N_16639,N_15965,N_14117);
nor U16640 (N_16640,N_15244,N_15169);
and U16641 (N_16641,N_14387,N_14285);
or U16642 (N_16642,N_14668,N_14284);
or U16643 (N_16643,N_14710,N_14985);
nand U16644 (N_16644,N_15301,N_15525);
nor U16645 (N_16645,N_14594,N_14029);
xnor U16646 (N_16646,N_15959,N_15570);
nor U16647 (N_16647,N_14834,N_15316);
nand U16648 (N_16648,N_14867,N_14764);
xnor U16649 (N_16649,N_15483,N_15827);
xnor U16650 (N_16650,N_15449,N_15645);
or U16651 (N_16651,N_14016,N_15275);
nor U16652 (N_16652,N_15263,N_15327);
nand U16653 (N_16653,N_14041,N_14403);
and U16654 (N_16654,N_14826,N_14887);
and U16655 (N_16655,N_15940,N_14220);
xor U16656 (N_16656,N_15553,N_15267);
and U16657 (N_16657,N_15365,N_15839);
nor U16658 (N_16658,N_14973,N_14173);
xor U16659 (N_16659,N_15717,N_14208);
and U16660 (N_16660,N_14136,N_15474);
or U16661 (N_16661,N_15144,N_14551);
xnor U16662 (N_16662,N_14302,N_15174);
or U16663 (N_16663,N_14452,N_15272);
nand U16664 (N_16664,N_14468,N_14901);
or U16665 (N_16665,N_14706,N_14477);
and U16666 (N_16666,N_14866,N_14939);
nand U16667 (N_16667,N_14916,N_14310);
xor U16668 (N_16668,N_14956,N_15322);
and U16669 (N_16669,N_15196,N_15660);
or U16670 (N_16670,N_15213,N_15497);
xor U16671 (N_16671,N_15032,N_15278);
nor U16672 (N_16672,N_14131,N_14058);
nand U16673 (N_16673,N_15722,N_14732);
nor U16674 (N_16674,N_15501,N_14869);
and U16675 (N_16675,N_15598,N_14598);
xor U16676 (N_16676,N_15597,N_15502);
nor U16677 (N_16677,N_15071,N_14795);
nor U16678 (N_16678,N_15191,N_14381);
and U16679 (N_16679,N_15872,N_14553);
and U16680 (N_16680,N_15833,N_15295);
and U16681 (N_16681,N_15233,N_14605);
or U16682 (N_16682,N_15874,N_14249);
nor U16683 (N_16683,N_14583,N_14226);
and U16684 (N_16684,N_15823,N_14010);
nor U16685 (N_16685,N_14961,N_15350);
and U16686 (N_16686,N_15536,N_15008);
and U16687 (N_16687,N_14268,N_14011);
nand U16688 (N_16688,N_15606,N_15889);
xnor U16689 (N_16689,N_14832,N_14146);
and U16690 (N_16690,N_15105,N_15023);
or U16691 (N_16691,N_15721,N_14596);
xnor U16692 (N_16692,N_15041,N_15135);
nand U16693 (N_16693,N_15876,N_15391);
nand U16694 (N_16694,N_15680,N_15372);
xor U16695 (N_16695,N_14968,N_14215);
nor U16696 (N_16696,N_14124,N_15989);
and U16697 (N_16697,N_15514,N_14997);
xnor U16698 (N_16698,N_15796,N_14512);
nor U16699 (N_16699,N_15734,N_15431);
and U16700 (N_16700,N_14375,N_14183);
nand U16701 (N_16701,N_15043,N_14050);
xor U16702 (N_16702,N_15403,N_15118);
or U16703 (N_16703,N_15249,N_15027);
xor U16704 (N_16704,N_15336,N_15409);
or U16705 (N_16705,N_14203,N_14305);
nor U16706 (N_16706,N_15520,N_15067);
or U16707 (N_16707,N_15716,N_15357);
nand U16708 (N_16708,N_14698,N_15412);
and U16709 (N_16709,N_14503,N_15381);
and U16710 (N_16710,N_15451,N_15891);
xor U16711 (N_16711,N_14449,N_14587);
and U16712 (N_16712,N_14756,N_14282);
and U16713 (N_16713,N_14201,N_14891);
nand U16714 (N_16714,N_14397,N_15024);
xnor U16715 (N_16715,N_14383,N_15494);
and U16716 (N_16716,N_15618,N_14027);
and U16717 (N_16717,N_15223,N_14856);
nor U16718 (N_16718,N_15850,N_14641);
nand U16719 (N_16719,N_14180,N_14165);
xnor U16720 (N_16720,N_14075,N_14800);
and U16721 (N_16721,N_15614,N_14936);
or U16722 (N_16722,N_14574,N_14779);
and U16723 (N_16723,N_14357,N_14517);
and U16724 (N_16724,N_15800,N_14049);
xor U16725 (N_16725,N_15065,N_15240);
or U16726 (N_16726,N_15535,N_15913);
nand U16727 (N_16727,N_15150,N_14057);
and U16728 (N_16728,N_14291,N_15742);
nor U16729 (N_16729,N_15500,N_15417);
nor U16730 (N_16730,N_14119,N_15620);
nor U16731 (N_16731,N_14875,N_14315);
xor U16732 (N_16732,N_15632,N_15056);
or U16733 (N_16733,N_14703,N_15784);
or U16734 (N_16734,N_15115,N_15373);
nor U16735 (N_16735,N_14713,N_14913);
nand U16736 (N_16736,N_15020,N_14504);
or U16737 (N_16737,N_15400,N_15681);
nor U16738 (N_16738,N_14525,N_14129);
or U16739 (N_16739,N_15155,N_14906);
nor U16740 (N_16740,N_14155,N_15712);
nand U16741 (N_16741,N_15047,N_15961);
xnor U16742 (N_16742,N_14772,N_14122);
xnor U16743 (N_16743,N_15188,N_14163);
nor U16744 (N_16744,N_14841,N_14239);
xor U16745 (N_16745,N_15326,N_14410);
nor U16746 (N_16746,N_15903,N_15258);
or U16747 (N_16747,N_15530,N_15905);
xor U16748 (N_16748,N_15685,N_14069);
or U16749 (N_16749,N_14360,N_14702);
or U16750 (N_16750,N_14515,N_14817);
and U16751 (N_16751,N_14212,N_15601);
nand U16752 (N_16752,N_15953,N_15995);
and U16753 (N_16753,N_15251,N_15875);
nor U16754 (N_16754,N_14622,N_15442);
nor U16755 (N_16755,N_14030,N_15208);
or U16756 (N_16756,N_14377,N_15341);
or U16757 (N_16757,N_14874,N_14751);
xnor U16758 (N_16758,N_14796,N_14134);
and U16759 (N_16759,N_15693,N_15467);
nand U16760 (N_16760,N_15971,N_15873);
nand U16761 (N_16761,N_15911,N_15471);
and U16762 (N_16762,N_14194,N_14719);
or U16763 (N_16763,N_15286,N_14040);
xnor U16764 (N_16764,N_14433,N_15654);
nand U16765 (N_16765,N_14774,N_14327);
xnor U16766 (N_16766,N_14618,N_15503);
nand U16767 (N_16767,N_14744,N_15522);
and U16768 (N_16768,N_14133,N_14681);
xor U16769 (N_16769,N_14546,N_14235);
nor U16770 (N_16770,N_15396,N_15930);
and U16771 (N_16771,N_15966,N_14857);
nor U16772 (N_16772,N_15134,N_14809);
nor U16773 (N_16773,N_15424,N_14086);
and U16774 (N_16774,N_14590,N_15758);
nor U16775 (N_16775,N_14787,N_14182);
nand U16776 (N_16776,N_15593,N_15694);
xnor U16777 (N_16777,N_15760,N_14785);
nand U16778 (N_16778,N_14202,N_15518);
nand U16779 (N_16779,N_14771,N_14837);
nor U16780 (N_16780,N_14561,N_15044);
or U16781 (N_16781,N_14804,N_15058);
nor U16782 (N_16782,N_15521,N_14103);
and U16783 (N_16783,N_14454,N_14929);
xnor U16784 (N_16784,N_14486,N_15423);
xnor U16785 (N_16785,N_14852,N_14998);
and U16786 (N_16786,N_14770,N_15343);
nor U16787 (N_16787,N_14907,N_15838);
and U16788 (N_16788,N_14640,N_15853);
nand U16789 (N_16789,N_14766,N_15750);
and U16790 (N_16790,N_15740,N_15081);
xnor U16791 (N_16791,N_15783,N_15452);
nand U16792 (N_16792,N_14531,N_14580);
nor U16793 (N_16793,N_15017,N_15099);
nor U16794 (N_16794,N_14054,N_15984);
nand U16795 (N_16795,N_15226,N_14729);
xor U16796 (N_16796,N_14944,N_14509);
and U16797 (N_16797,N_14922,N_14233);
or U16798 (N_16798,N_14749,N_15515);
nand U16799 (N_16799,N_14024,N_14815);
xor U16800 (N_16800,N_14589,N_15279);
nand U16801 (N_16801,N_15202,N_14181);
and U16802 (N_16802,N_14704,N_14570);
or U16803 (N_16803,N_15298,N_15094);
xor U16804 (N_16804,N_15789,N_14897);
or U16805 (N_16805,N_15755,N_15669);
and U16806 (N_16806,N_14560,N_14584);
nor U16807 (N_16807,N_15683,N_14178);
or U16808 (N_16808,N_14332,N_15382);
nor U16809 (N_16809,N_15635,N_14677);
nand U16810 (N_16810,N_15519,N_14277);
nor U16811 (N_16811,N_15006,N_15309);
or U16812 (N_16812,N_15211,N_14068);
xnor U16813 (N_16813,N_15108,N_15582);
and U16814 (N_16814,N_15141,N_14072);
nand U16815 (N_16815,N_14217,N_14455);
xor U16816 (N_16816,N_15723,N_14820);
nor U16817 (N_16817,N_14138,N_15950);
nor U16818 (N_16818,N_15805,N_14325);
xnor U16819 (N_16819,N_14356,N_14831);
xnor U16820 (N_16820,N_15885,N_15388);
nor U16821 (N_16821,N_15348,N_15122);
nor U16822 (N_16822,N_15603,N_14380);
xor U16823 (N_16823,N_14084,N_15164);
nand U16824 (N_16824,N_14653,N_15893);
nand U16825 (N_16825,N_15153,N_15561);
nand U16826 (N_16826,N_14656,N_14621);
or U16827 (N_16827,N_15897,N_14266);
and U16828 (N_16828,N_15611,N_14137);
xnor U16829 (N_16829,N_14849,N_15651);
nor U16830 (N_16830,N_14573,N_15003);
and U16831 (N_16831,N_14399,N_15358);
xor U16832 (N_16832,N_14811,N_14469);
nor U16833 (N_16833,N_14378,N_14645);
nor U16834 (N_16834,N_15868,N_14367);
or U16835 (N_16835,N_15201,N_14179);
nand U16836 (N_16836,N_14128,N_14273);
and U16837 (N_16837,N_14839,N_14135);
nand U16838 (N_16838,N_15215,N_15523);
and U16839 (N_16839,N_15725,N_14623);
and U16840 (N_16840,N_15401,N_15087);
or U16841 (N_16841,N_14038,N_15818);
nand U16842 (N_16842,N_14344,N_14164);
nor U16843 (N_16843,N_15610,N_15005);
nand U16844 (N_16844,N_15726,N_15987);
or U16845 (N_16845,N_14508,N_14730);
nand U16846 (N_16846,N_15061,N_14686);
xor U16847 (N_16847,N_15088,N_15390);
xnor U16848 (N_16848,N_14355,N_14031);
nand U16849 (N_16849,N_14813,N_15086);
and U16850 (N_16850,N_14822,N_15387);
and U16851 (N_16851,N_15757,N_14917);
xnor U16852 (N_16852,N_14099,N_15241);
xor U16853 (N_16853,N_15870,N_15640);
or U16854 (N_16854,N_14314,N_14251);
and U16855 (N_16855,N_15935,N_15480);
nand U16856 (N_16856,N_15799,N_14055);
xor U16857 (N_16857,N_14275,N_15161);
nor U16858 (N_16858,N_14166,N_14156);
nor U16859 (N_16859,N_14053,N_14316);
and U16860 (N_16860,N_14331,N_14090);
or U16861 (N_16861,N_14736,N_14386);
and U16862 (N_16862,N_15448,N_15792);
or U16863 (N_16863,N_15901,N_14152);
or U16864 (N_16864,N_15236,N_15038);
or U16865 (N_16865,N_15550,N_14033);
xor U16866 (N_16866,N_14943,N_14884);
xor U16867 (N_16867,N_15738,N_15338);
nand U16868 (N_16868,N_14638,N_15031);
nand U16869 (N_16869,N_15639,N_14538);
and U16870 (N_16870,N_14616,N_14980);
xor U16871 (N_16871,N_15428,N_14753);
and U16872 (N_16872,N_15179,N_14229);
or U16873 (N_16873,N_14225,N_15608);
and U16874 (N_16874,N_14778,N_14434);
nor U16875 (N_16875,N_14209,N_14631);
and U16876 (N_16876,N_15539,N_15636);
and U16877 (N_16877,N_15493,N_15613);
and U16878 (N_16878,N_15496,N_15291);
xor U16879 (N_16879,N_14990,N_14544);
nand U16880 (N_16880,N_15265,N_14089);
or U16881 (N_16881,N_15748,N_15781);
nand U16882 (N_16882,N_15479,N_15754);
nand U16883 (N_16883,N_15138,N_14663);
xor U16884 (N_16884,N_15549,N_14300);
and U16885 (N_16885,N_14224,N_14608);
xor U16886 (N_16886,N_15936,N_14088);
nand U16887 (N_16887,N_15074,N_15998);
or U16888 (N_16888,N_15492,N_15574);
and U16889 (N_16889,N_15642,N_15572);
nand U16890 (N_16890,N_14470,N_15225);
or U16891 (N_16891,N_14110,N_14680);
and U16892 (N_16892,N_14926,N_15746);
nor U16893 (N_16893,N_14370,N_14507);
nand U16894 (N_16894,N_14910,N_14293);
xnor U16895 (N_16895,N_15170,N_14065);
nor U16896 (N_16896,N_14807,N_14514);
and U16897 (N_16897,N_14493,N_14019);
nand U16898 (N_16898,N_15386,N_15863);
or U16899 (N_16899,N_14803,N_14763);
and U16900 (N_16900,N_15376,N_14198);
nand U16901 (N_16901,N_15281,N_15254);
nor U16902 (N_16902,N_15733,N_15629);
and U16903 (N_16903,N_14020,N_15852);
nor U16904 (N_16904,N_14085,N_14840);
or U16905 (N_16905,N_14571,N_15625);
nor U16906 (N_16906,N_14147,N_14788);
nand U16907 (N_16907,N_14475,N_15884);
nand U16908 (N_16908,N_14081,N_14056);
nand U16909 (N_16909,N_15054,N_14438);
xor U16910 (N_16910,N_15861,N_14023);
nor U16911 (N_16911,N_15157,N_14237);
or U16912 (N_16912,N_14920,N_15050);
or U16913 (N_16913,N_15369,N_14436);
nand U16914 (N_16914,N_14951,N_15101);
or U16915 (N_16915,N_15210,N_14554);
nor U16916 (N_16916,N_14464,N_14149);
nand U16917 (N_16917,N_15282,N_15072);
nand U16918 (N_16918,N_14933,N_15978);
nand U16919 (N_16919,N_14219,N_15540);
nor U16920 (N_16920,N_15001,N_14534);
xor U16921 (N_16921,N_15374,N_15037);
or U16922 (N_16922,N_14467,N_14432);
or U16923 (N_16923,N_15499,N_14728);
or U16924 (N_16924,N_14969,N_14801);
or U16925 (N_16925,N_14646,N_15306);
and U16926 (N_16926,N_14995,N_15262);
nand U16927 (N_16927,N_15955,N_15305);
nand U16928 (N_16928,N_14061,N_14612);
nor U16929 (N_16929,N_15902,N_15287);
or U16930 (N_16930,N_15922,N_15457);
xor U16931 (N_16931,N_15131,N_14104);
and U16932 (N_16932,N_15458,N_14664);
nand U16933 (N_16933,N_14441,N_15816);
nor U16934 (N_16934,N_14591,N_15627);
nand U16935 (N_16935,N_15219,N_14333);
xor U16936 (N_16936,N_14116,N_15204);
xor U16937 (N_16937,N_14278,N_14296);
nor U16938 (N_16938,N_14648,N_15300);
or U16939 (N_16939,N_14542,N_14051);
and U16940 (N_16940,N_14549,N_15362);
nor U16941 (N_16941,N_14206,N_15124);
xnor U16942 (N_16942,N_14066,N_15489);
or U16943 (N_16943,N_15599,N_15782);
xnor U16944 (N_16944,N_14927,N_14715);
or U16945 (N_16945,N_15662,N_15245);
xor U16946 (N_16946,N_15355,N_15702);
or U16947 (N_16947,N_14987,N_14707);
nand U16948 (N_16948,N_15909,N_15644);
nand U16949 (N_16949,N_14118,N_15711);
xor U16950 (N_16950,N_15133,N_15064);
and U16951 (N_16951,N_15916,N_15589);
xnor U16952 (N_16952,N_15340,N_14851);
nor U16953 (N_16953,N_14342,N_14671);
xnor U16954 (N_16954,N_14492,N_15917);
and U16955 (N_16955,N_14562,N_14196);
xor U16956 (N_16956,N_14132,N_15908);
or U16957 (N_16957,N_15934,N_14483);
nand U16958 (N_16958,N_15643,N_14319);
nor U16959 (N_16959,N_14600,N_14079);
or U16960 (N_16960,N_15954,N_15498);
xnor U16961 (N_16961,N_15802,N_15586);
and U16962 (N_16962,N_14868,N_14724);
and U16963 (N_16963,N_14658,N_15773);
and U16964 (N_16964,N_15166,N_14322);
xnor U16965 (N_16965,N_15055,N_15132);
nand U16966 (N_16966,N_14052,N_14321);
or U16967 (N_16967,N_15647,N_14242);
nor U16968 (N_16968,N_15096,N_14650);
xnor U16969 (N_16969,N_14463,N_14304);
and U16970 (N_16970,N_15938,N_14309);
nand U16971 (N_16971,N_14262,N_15049);
or U16972 (N_16972,N_14791,N_15331);
xor U16973 (N_16973,N_14167,N_15859);
and U16974 (N_16974,N_14781,N_14964);
xnor U16975 (N_16975,N_14575,N_14960);
nand U16976 (N_16976,N_14488,N_15980);
nand U16977 (N_16977,N_14216,N_15039);
nand U16978 (N_16978,N_14456,N_15670);
xor U16979 (N_16979,N_15454,N_14836);
nand U16980 (N_16980,N_15485,N_15798);
xor U16981 (N_16981,N_14928,N_15658);
or U16982 (N_16982,N_14745,N_14368);
or U16983 (N_16983,N_14064,N_14860);
xor U16984 (N_16984,N_14078,N_15546);
and U16985 (N_16985,N_15104,N_14543);
nor U16986 (N_16986,N_15089,N_14792);
or U16987 (N_16987,N_14241,N_15609);
nor U16988 (N_16988,N_14895,N_14666);
xnor U16989 (N_16989,N_15946,N_15517);
or U16990 (N_16990,N_14361,N_15576);
or U16991 (N_16991,N_15126,N_15894);
nand U16992 (N_16992,N_14604,N_14480);
nor U16993 (N_16993,N_15378,N_14292);
or U16994 (N_16994,N_14678,N_14705);
xor U16995 (N_16995,N_14734,N_15688);
or U16996 (N_16996,N_14187,N_15962);
nand U16997 (N_16997,N_14338,N_14125);
nand U16998 (N_16998,N_14684,N_14882);
nand U16999 (N_16999,N_14429,N_15318);
and U17000 (N_17000,N_15003,N_15099);
nor U17001 (N_17001,N_14698,N_15889);
or U17002 (N_17002,N_15765,N_15604);
and U17003 (N_17003,N_15304,N_15270);
or U17004 (N_17004,N_15852,N_15425);
and U17005 (N_17005,N_15053,N_14217);
and U17006 (N_17006,N_14055,N_15972);
xor U17007 (N_17007,N_14325,N_15583);
and U17008 (N_17008,N_15101,N_14370);
and U17009 (N_17009,N_14403,N_14759);
or U17010 (N_17010,N_15657,N_14386);
xnor U17011 (N_17011,N_14234,N_15169);
nand U17012 (N_17012,N_14909,N_14272);
nand U17013 (N_17013,N_14250,N_14577);
or U17014 (N_17014,N_14362,N_15047);
nor U17015 (N_17015,N_15838,N_14458);
and U17016 (N_17016,N_15852,N_15153);
or U17017 (N_17017,N_14787,N_14530);
nor U17018 (N_17018,N_14722,N_15762);
or U17019 (N_17019,N_14429,N_15267);
or U17020 (N_17020,N_15389,N_15468);
and U17021 (N_17021,N_15427,N_15564);
or U17022 (N_17022,N_15111,N_14571);
or U17023 (N_17023,N_14484,N_14400);
nand U17024 (N_17024,N_14831,N_14168);
nand U17025 (N_17025,N_14087,N_15981);
and U17026 (N_17026,N_14330,N_14325);
and U17027 (N_17027,N_15643,N_14642);
or U17028 (N_17028,N_15527,N_14247);
nand U17029 (N_17029,N_14018,N_14666);
nand U17030 (N_17030,N_15751,N_15647);
xnor U17031 (N_17031,N_14967,N_14973);
nor U17032 (N_17032,N_15385,N_15605);
and U17033 (N_17033,N_14307,N_14093);
or U17034 (N_17034,N_15204,N_15085);
nor U17035 (N_17035,N_15098,N_15587);
nand U17036 (N_17036,N_15095,N_14497);
nor U17037 (N_17037,N_15686,N_15866);
nand U17038 (N_17038,N_15645,N_15097);
or U17039 (N_17039,N_15541,N_15110);
and U17040 (N_17040,N_15368,N_14524);
and U17041 (N_17041,N_14212,N_15430);
or U17042 (N_17042,N_15572,N_15637);
or U17043 (N_17043,N_14337,N_14623);
and U17044 (N_17044,N_15366,N_15334);
or U17045 (N_17045,N_15488,N_14274);
nand U17046 (N_17046,N_14944,N_15500);
and U17047 (N_17047,N_14433,N_15326);
nand U17048 (N_17048,N_15657,N_14498);
nand U17049 (N_17049,N_14457,N_15762);
nor U17050 (N_17050,N_14754,N_14047);
nor U17051 (N_17051,N_15784,N_15098);
xnor U17052 (N_17052,N_15322,N_14216);
or U17053 (N_17053,N_14276,N_15131);
nand U17054 (N_17054,N_14268,N_14877);
xor U17055 (N_17055,N_14608,N_15500);
xor U17056 (N_17056,N_15237,N_14648);
nor U17057 (N_17057,N_14996,N_14378);
or U17058 (N_17058,N_14606,N_15057);
nand U17059 (N_17059,N_15721,N_15185);
and U17060 (N_17060,N_15795,N_15399);
nand U17061 (N_17061,N_15332,N_14505);
xnor U17062 (N_17062,N_14430,N_14749);
or U17063 (N_17063,N_14393,N_14699);
and U17064 (N_17064,N_14278,N_14770);
or U17065 (N_17065,N_15167,N_14024);
or U17066 (N_17066,N_15229,N_14589);
nor U17067 (N_17067,N_15226,N_15898);
or U17068 (N_17068,N_15171,N_14690);
xnor U17069 (N_17069,N_15503,N_14194);
xnor U17070 (N_17070,N_15037,N_15382);
or U17071 (N_17071,N_15825,N_15305);
and U17072 (N_17072,N_15689,N_14939);
and U17073 (N_17073,N_15830,N_14727);
or U17074 (N_17074,N_15106,N_14221);
nor U17075 (N_17075,N_15871,N_15095);
xnor U17076 (N_17076,N_14270,N_14146);
nor U17077 (N_17077,N_14645,N_15934);
xnor U17078 (N_17078,N_14206,N_14021);
nand U17079 (N_17079,N_14376,N_15763);
nor U17080 (N_17080,N_15051,N_14824);
nand U17081 (N_17081,N_15526,N_14235);
nand U17082 (N_17082,N_14287,N_15472);
or U17083 (N_17083,N_14298,N_15877);
nand U17084 (N_17084,N_15403,N_15436);
nand U17085 (N_17085,N_14847,N_15415);
or U17086 (N_17086,N_15895,N_14483);
xnor U17087 (N_17087,N_14173,N_14214);
or U17088 (N_17088,N_14610,N_14564);
and U17089 (N_17089,N_15900,N_15064);
or U17090 (N_17090,N_14631,N_15149);
nand U17091 (N_17091,N_14691,N_14472);
nand U17092 (N_17092,N_14762,N_14005);
and U17093 (N_17093,N_14722,N_14111);
and U17094 (N_17094,N_14283,N_15251);
nor U17095 (N_17095,N_15846,N_15094);
nor U17096 (N_17096,N_14043,N_15992);
or U17097 (N_17097,N_14493,N_15360);
nor U17098 (N_17098,N_15277,N_15660);
or U17099 (N_17099,N_14899,N_15547);
xor U17100 (N_17100,N_14272,N_14154);
nand U17101 (N_17101,N_15492,N_15237);
xnor U17102 (N_17102,N_15745,N_14215);
and U17103 (N_17103,N_15931,N_14482);
nor U17104 (N_17104,N_14862,N_15783);
xnor U17105 (N_17105,N_14987,N_14750);
nor U17106 (N_17106,N_14081,N_15916);
xor U17107 (N_17107,N_14304,N_14538);
nor U17108 (N_17108,N_14660,N_14561);
nor U17109 (N_17109,N_14890,N_14620);
nand U17110 (N_17110,N_15674,N_15520);
nand U17111 (N_17111,N_15574,N_15021);
nor U17112 (N_17112,N_15175,N_15574);
or U17113 (N_17113,N_15732,N_14819);
or U17114 (N_17114,N_15075,N_15845);
xnor U17115 (N_17115,N_14269,N_14801);
nor U17116 (N_17116,N_14066,N_15416);
and U17117 (N_17117,N_14755,N_15075);
nor U17118 (N_17118,N_15805,N_14203);
or U17119 (N_17119,N_15431,N_15815);
and U17120 (N_17120,N_15481,N_14149);
or U17121 (N_17121,N_15319,N_15352);
nand U17122 (N_17122,N_14130,N_14951);
and U17123 (N_17123,N_14362,N_14056);
xnor U17124 (N_17124,N_14494,N_14556);
nand U17125 (N_17125,N_15658,N_15241);
xor U17126 (N_17126,N_14087,N_15740);
and U17127 (N_17127,N_15386,N_14978);
or U17128 (N_17128,N_15316,N_15759);
nor U17129 (N_17129,N_14881,N_15910);
nand U17130 (N_17130,N_15291,N_14496);
and U17131 (N_17131,N_14214,N_14830);
xor U17132 (N_17132,N_15408,N_15615);
xor U17133 (N_17133,N_14271,N_14226);
or U17134 (N_17134,N_15029,N_15133);
or U17135 (N_17135,N_14205,N_15333);
or U17136 (N_17136,N_14457,N_15087);
or U17137 (N_17137,N_14015,N_14957);
or U17138 (N_17138,N_15078,N_14188);
xor U17139 (N_17139,N_15393,N_15074);
nor U17140 (N_17140,N_15649,N_14234);
xor U17141 (N_17141,N_15484,N_14420);
or U17142 (N_17142,N_14817,N_15817);
nor U17143 (N_17143,N_14277,N_14340);
or U17144 (N_17144,N_14355,N_14772);
nor U17145 (N_17145,N_14957,N_15357);
or U17146 (N_17146,N_15751,N_15888);
and U17147 (N_17147,N_14011,N_15202);
nand U17148 (N_17148,N_15491,N_15798);
nand U17149 (N_17149,N_15151,N_14300);
nor U17150 (N_17150,N_15070,N_14110);
and U17151 (N_17151,N_15407,N_15453);
and U17152 (N_17152,N_15072,N_15443);
or U17153 (N_17153,N_15654,N_14811);
or U17154 (N_17154,N_14096,N_15039);
and U17155 (N_17155,N_14533,N_15150);
or U17156 (N_17156,N_14541,N_15463);
and U17157 (N_17157,N_15114,N_14012);
nand U17158 (N_17158,N_14291,N_14451);
and U17159 (N_17159,N_15177,N_14031);
xnor U17160 (N_17160,N_15819,N_14540);
or U17161 (N_17161,N_14428,N_15182);
and U17162 (N_17162,N_15142,N_15739);
xor U17163 (N_17163,N_15119,N_15080);
and U17164 (N_17164,N_15257,N_15354);
nand U17165 (N_17165,N_14775,N_14455);
nor U17166 (N_17166,N_15180,N_15661);
xor U17167 (N_17167,N_14416,N_15716);
xnor U17168 (N_17168,N_15330,N_15308);
or U17169 (N_17169,N_14207,N_15194);
and U17170 (N_17170,N_14978,N_14252);
nor U17171 (N_17171,N_15775,N_14563);
and U17172 (N_17172,N_14977,N_15506);
xnor U17173 (N_17173,N_15083,N_15455);
or U17174 (N_17174,N_15871,N_14715);
xnor U17175 (N_17175,N_14370,N_14131);
nand U17176 (N_17176,N_14641,N_15399);
and U17177 (N_17177,N_14456,N_14771);
and U17178 (N_17178,N_15424,N_14885);
nand U17179 (N_17179,N_15992,N_14189);
or U17180 (N_17180,N_14198,N_14674);
and U17181 (N_17181,N_15148,N_15811);
nor U17182 (N_17182,N_14029,N_14396);
nor U17183 (N_17183,N_15139,N_15845);
or U17184 (N_17184,N_15118,N_15485);
xnor U17185 (N_17185,N_14156,N_14917);
nand U17186 (N_17186,N_15865,N_14180);
nor U17187 (N_17187,N_14661,N_15902);
nand U17188 (N_17188,N_14678,N_14555);
nor U17189 (N_17189,N_14898,N_14081);
nand U17190 (N_17190,N_15383,N_15312);
xor U17191 (N_17191,N_15983,N_15493);
or U17192 (N_17192,N_15025,N_14556);
xor U17193 (N_17193,N_14489,N_15473);
nand U17194 (N_17194,N_15946,N_14254);
and U17195 (N_17195,N_14743,N_14548);
and U17196 (N_17196,N_15982,N_14882);
or U17197 (N_17197,N_15306,N_15350);
and U17198 (N_17198,N_14920,N_15056);
xnor U17199 (N_17199,N_15962,N_14403);
or U17200 (N_17200,N_15617,N_15090);
nand U17201 (N_17201,N_14573,N_14785);
nand U17202 (N_17202,N_14244,N_15847);
nand U17203 (N_17203,N_14402,N_14954);
nand U17204 (N_17204,N_14445,N_15087);
nand U17205 (N_17205,N_15059,N_14778);
and U17206 (N_17206,N_14896,N_14528);
nor U17207 (N_17207,N_14888,N_15515);
nand U17208 (N_17208,N_14126,N_15027);
xnor U17209 (N_17209,N_15741,N_15546);
nor U17210 (N_17210,N_14541,N_15908);
nor U17211 (N_17211,N_14754,N_15914);
nand U17212 (N_17212,N_15908,N_15296);
and U17213 (N_17213,N_14886,N_14087);
nand U17214 (N_17214,N_15634,N_14693);
and U17215 (N_17215,N_15221,N_15451);
nand U17216 (N_17216,N_15276,N_14652);
xnor U17217 (N_17217,N_14324,N_15603);
nor U17218 (N_17218,N_15293,N_14243);
nor U17219 (N_17219,N_15857,N_14577);
xnor U17220 (N_17220,N_15281,N_15905);
or U17221 (N_17221,N_15435,N_15334);
or U17222 (N_17222,N_15613,N_15419);
xor U17223 (N_17223,N_14754,N_14542);
and U17224 (N_17224,N_15561,N_15544);
nor U17225 (N_17225,N_15198,N_15719);
xor U17226 (N_17226,N_14454,N_15771);
or U17227 (N_17227,N_15999,N_14902);
xor U17228 (N_17228,N_14912,N_14007);
and U17229 (N_17229,N_15914,N_15232);
and U17230 (N_17230,N_15147,N_14373);
nand U17231 (N_17231,N_14621,N_15393);
nor U17232 (N_17232,N_15876,N_14936);
and U17233 (N_17233,N_14990,N_14471);
nor U17234 (N_17234,N_14494,N_15790);
and U17235 (N_17235,N_14623,N_15034);
nand U17236 (N_17236,N_15916,N_15191);
nor U17237 (N_17237,N_15165,N_14854);
nand U17238 (N_17238,N_15279,N_14899);
xnor U17239 (N_17239,N_15070,N_14656);
nor U17240 (N_17240,N_14459,N_15276);
nand U17241 (N_17241,N_15601,N_15941);
xnor U17242 (N_17242,N_14505,N_14600);
nand U17243 (N_17243,N_14655,N_15748);
nand U17244 (N_17244,N_15100,N_15482);
nand U17245 (N_17245,N_15345,N_15996);
xnor U17246 (N_17246,N_15137,N_14558);
xor U17247 (N_17247,N_14747,N_15454);
xnor U17248 (N_17248,N_15895,N_14784);
nor U17249 (N_17249,N_14939,N_15486);
xor U17250 (N_17250,N_15037,N_15714);
nor U17251 (N_17251,N_14959,N_14639);
nor U17252 (N_17252,N_14356,N_15043);
nand U17253 (N_17253,N_14276,N_14947);
or U17254 (N_17254,N_14266,N_14897);
xnor U17255 (N_17255,N_15788,N_15792);
and U17256 (N_17256,N_14487,N_15355);
or U17257 (N_17257,N_14038,N_14699);
nand U17258 (N_17258,N_14750,N_15959);
and U17259 (N_17259,N_14509,N_15942);
nor U17260 (N_17260,N_14964,N_15898);
nand U17261 (N_17261,N_14128,N_15519);
and U17262 (N_17262,N_14947,N_15467);
or U17263 (N_17263,N_15193,N_14056);
and U17264 (N_17264,N_15416,N_14291);
and U17265 (N_17265,N_15120,N_14474);
and U17266 (N_17266,N_14143,N_14954);
or U17267 (N_17267,N_15506,N_15654);
or U17268 (N_17268,N_14767,N_14742);
xnor U17269 (N_17269,N_14158,N_15358);
nor U17270 (N_17270,N_14041,N_14328);
xor U17271 (N_17271,N_14473,N_14878);
nor U17272 (N_17272,N_14350,N_15406);
and U17273 (N_17273,N_15656,N_14156);
nand U17274 (N_17274,N_15106,N_15917);
nand U17275 (N_17275,N_15928,N_15903);
xor U17276 (N_17276,N_14640,N_14536);
nor U17277 (N_17277,N_14970,N_15869);
and U17278 (N_17278,N_14016,N_15066);
and U17279 (N_17279,N_14954,N_15513);
xor U17280 (N_17280,N_15830,N_15112);
or U17281 (N_17281,N_15226,N_15274);
nor U17282 (N_17282,N_15910,N_14207);
xor U17283 (N_17283,N_15664,N_15697);
xnor U17284 (N_17284,N_14112,N_14477);
and U17285 (N_17285,N_15349,N_15286);
nand U17286 (N_17286,N_15701,N_15997);
nor U17287 (N_17287,N_14619,N_15699);
xnor U17288 (N_17288,N_15237,N_15552);
xor U17289 (N_17289,N_15638,N_14765);
nand U17290 (N_17290,N_15784,N_14378);
or U17291 (N_17291,N_14848,N_14253);
or U17292 (N_17292,N_14549,N_15583);
or U17293 (N_17293,N_15013,N_14662);
nand U17294 (N_17294,N_15929,N_14707);
xor U17295 (N_17295,N_14113,N_14268);
nand U17296 (N_17296,N_14047,N_14044);
nand U17297 (N_17297,N_14877,N_15910);
or U17298 (N_17298,N_15968,N_15752);
nand U17299 (N_17299,N_15747,N_14717);
and U17300 (N_17300,N_14196,N_15458);
xor U17301 (N_17301,N_15968,N_14685);
nor U17302 (N_17302,N_15719,N_14357);
nor U17303 (N_17303,N_15992,N_15743);
xnor U17304 (N_17304,N_14635,N_15949);
nand U17305 (N_17305,N_15475,N_15654);
or U17306 (N_17306,N_15689,N_15363);
xor U17307 (N_17307,N_15489,N_14349);
nand U17308 (N_17308,N_15764,N_15263);
xor U17309 (N_17309,N_15152,N_14487);
nor U17310 (N_17310,N_15123,N_14450);
nor U17311 (N_17311,N_14342,N_14459);
and U17312 (N_17312,N_15628,N_14213);
nand U17313 (N_17313,N_15489,N_15944);
xnor U17314 (N_17314,N_15401,N_15176);
or U17315 (N_17315,N_14099,N_15485);
or U17316 (N_17316,N_14531,N_15280);
and U17317 (N_17317,N_15102,N_15915);
or U17318 (N_17318,N_14172,N_14620);
or U17319 (N_17319,N_15913,N_14979);
or U17320 (N_17320,N_14037,N_15684);
or U17321 (N_17321,N_15970,N_15429);
nor U17322 (N_17322,N_15006,N_14724);
or U17323 (N_17323,N_14659,N_14229);
nor U17324 (N_17324,N_15461,N_15042);
nand U17325 (N_17325,N_14986,N_14356);
xnor U17326 (N_17326,N_15783,N_15554);
or U17327 (N_17327,N_15863,N_14656);
nand U17328 (N_17328,N_14505,N_14185);
and U17329 (N_17329,N_14972,N_15433);
and U17330 (N_17330,N_14855,N_14628);
nor U17331 (N_17331,N_15395,N_14286);
or U17332 (N_17332,N_15942,N_15932);
xnor U17333 (N_17333,N_15839,N_15224);
and U17334 (N_17334,N_14921,N_15094);
and U17335 (N_17335,N_14751,N_14844);
or U17336 (N_17336,N_14284,N_14298);
or U17337 (N_17337,N_14852,N_15184);
xnor U17338 (N_17338,N_14830,N_14092);
nand U17339 (N_17339,N_15090,N_14776);
or U17340 (N_17340,N_15346,N_15776);
nor U17341 (N_17341,N_14961,N_14252);
or U17342 (N_17342,N_14716,N_15750);
nor U17343 (N_17343,N_15366,N_15081);
nand U17344 (N_17344,N_14246,N_14901);
xnor U17345 (N_17345,N_15435,N_15607);
nor U17346 (N_17346,N_15175,N_15233);
or U17347 (N_17347,N_15586,N_14645);
nand U17348 (N_17348,N_15111,N_15066);
and U17349 (N_17349,N_15886,N_14686);
xnor U17350 (N_17350,N_15097,N_14518);
or U17351 (N_17351,N_14751,N_14342);
nor U17352 (N_17352,N_14986,N_14867);
or U17353 (N_17353,N_14882,N_14071);
nand U17354 (N_17354,N_15866,N_15429);
nor U17355 (N_17355,N_14127,N_15787);
nand U17356 (N_17356,N_14993,N_15357);
or U17357 (N_17357,N_14200,N_15664);
or U17358 (N_17358,N_15731,N_15900);
or U17359 (N_17359,N_14765,N_14129);
or U17360 (N_17360,N_14988,N_15768);
or U17361 (N_17361,N_15070,N_15612);
nor U17362 (N_17362,N_14959,N_14568);
and U17363 (N_17363,N_14705,N_14025);
and U17364 (N_17364,N_15613,N_15973);
xor U17365 (N_17365,N_15866,N_14020);
xnor U17366 (N_17366,N_15330,N_15434);
or U17367 (N_17367,N_14539,N_14452);
or U17368 (N_17368,N_14636,N_15084);
or U17369 (N_17369,N_14172,N_14858);
nor U17370 (N_17370,N_15568,N_15261);
or U17371 (N_17371,N_15057,N_14054);
nand U17372 (N_17372,N_14695,N_15494);
nor U17373 (N_17373,N_14944,N_14325);
or U17374 (N_17374,N_14516,N_15015);
xor U17375 (N_17375,N_15155,N_14735);
and U17376 (N_17376,N_15145,N_15321);
xnor U17377 (N_17377,N_15645,N_15884);
nor U17378 (N_17378,N_15360,N_15365);
nand U17379 (N_17379,N_14332,N_15753);
xnor U17380 (N_17380,N_15109,N_14374);
nor U17381 (N_17381,N_14029,N_14030);
and U17382 (N_17382,N_14900,N_15956);
xor U17383 (N_17383,N_15647,N_15591);
nor U17384 (N_17384,N_14023,N_15718);
and U17385 (N_17385,N_14242,N_15077);
xor U17386 (N_17386,N_14752,N_15609);
nand U17387 (N_17387,N_14674,N_14214);
or U17388 (N_17388,N_15609,N_14758);
nand U17389 (N_17389,N_15836,N_14742);
xnor U17390 (N_17390,N_15670,N_14467);
xnor U17391 (N_17391,N_15218,N_15345);
xor U17392 (N_17392,N_15000,N_15880);
or U17393 (N_17393,N_15084,N_15992);
xnor U17394 (N_17394,N_15303,N_14196);
or U17395 (N_17395,N_15462,N_15187);
nor U17396 (N_17396,N_15408,N_14071);
or U17397 (N_17397,N_15623,N_14577);
xor U17398 (N_17398,N_14267,N_14439);
or U17399 (N_17399,N_15041,N_15164);
xor U17400 (N_17400,N_15774,N_14071);
and U17401 (N_17401,N_14117,N_15659);
and U17402 (N_17402,N_14445,N_15656);
nor U17403 (N_17403,N_15622,N_14039);
and U17404 (N_17404,N_14016,N_14056);
or U17405 (N_17405,N_14242,N_14668);
or U17406 (N_17406,N_15209,N_15997);
and U17407 (N_17407,N_14044,N_15804);
or U17408 (N_17408,N_14130,N_14237);
and U17409 (N_17409,N_15206,N_14923);
nand U17410 (N_17410,N_14907,N_14409);
nand U17411 (N_17411,N_14203,N_14031);
nand U17412 (N_17412,N_15295,N_14918);
nor U17413 (N_17413,N_15374,N_15119);
or U17414 (N_17414,N_14702,N_15009);
and U17415 (N_17415,N_15998,N_15820);
or U17416 (N_17416,N_15110,N_14685);
nor U17417 (N_17417,N_14461,N_15963);
nand U17418 (N_17418,N_15603,N_14434);
nand U17419 (N_17419,N_14394,N_15087);
xnor U17420 (N_17420,N_14076,N_15619);
nor U17421 (N_17421,N_14718,N_15538);
nor U17422 (N_17422,N_15397,N_14729);
and U17423 (N_17423,N_14367,N_14887);
or U17424 (N_17424,N_14006,N_15172);
nor U17425 (N_17425,N_14189,N_15498);
or U17426 (N_17426,N_15951,N_15238);
nor U17427 (N_17427,N_14152,N_15179);
nor U17428 (N_17428,N_14936,N_14741);
or U17429 (N_17429,N_15122,N_14216);
or U17430 (N_17430,N_14280,N_15156);
xnor U17431 (N_17431,N_14284,N_15645);
and U17432 (N_17432,N_15762,N_15784);
and U17433 (N_17433,N_15114,N_15800);
nand U17434 (N_17434,N_14699,N_15144);
nand U17435 (N_17435,N_14294,N_15927);
nor U17436 (N_17436,N_14795,N_15346);
nor U17437 (N_17437,N_14134,N_15775);
and U17438 (N_17438,N_15032,N_14209);
or U17439 (N_17439,N_14444,N_14736);
nand U17440 (N_17440,N_15911,N_15868);
nor U17441 (N_17441,N_15826,N_14351);
and U17442 (N_17442,N_15460,N_14661);
nand U17443 (N_17443,N_14819,N_14735);
nand U17444 (N_17444,N_15836,N_15979);
nor U17445 (N_17445,N_14047,N_14491);
and U17446 (N_17446,N_15141,N_14803);
xor U17447 (N_17447,N_15303,N_15908);
nor U17448 (N_17448,N_14289,N_15941);
or U17449 (N_17449,N_15155,N_14613);
xor U17450 (N_17450,N_14221,N_15429);
or U17451 (N_17451,N_15734,N_14464);
or U17452 (N_17452,N_14691,N_14980);
nand U17453 (N_17453,N_15434,N_15361);
xor U17454 (N_17454,N_14313,N_14188);
nor U17455 (N_17455,N_15644,N_15940);
and U17456 (N_17456,N_14311,N_15609);
xnor U17457 (N_17457,N_14646,N_14044);
or U17458 (N_17458,N_14547,N_14382);
or U17459 (N_17459,N_15136,N_15114);
xnor U17460 (N_17460,N_15904,N_15999);
nand U17461 (N_17461,N_14157,N_15434);
or U17462 (N_17462,N_14026,N_15014);
or U17463 (N_17463,N_14734,N_14669);
or U17464 (N_17464,N_14950,N_14290);
or U17465 (N_17465,N_15381,N_15076);
or U17466 (N_17466,N_15889,N_14610);
or U17467 (N_17467,N_14513,N_15484);
nor U17468 (N_17468,N_14871,N_15468);
nand U17469 (N_17469,N_15136,N_14967);
nand U17470 (N_17470,N_15983,N_14435);
or U17471 (N_17471,N_14097,N_14915);
nand U17472 (N_17472,N_14729,N_15477);
or U17473 (N_17473,N_15691,N_15051);
nor U17474 (N_17474,N_15884,N_14275);
and U17475 (N_17475,N_15133,N_15290);
and U17476 (N_17476,N_14452,N_15445);
or U17477 (N_17477,N_14384,N_15582);
xor U17478 (N_17478,N_14823,N_15121);
or U17479 (N_17479,N_15048,N_15289);
nand U17480 (N_17480,N_14682,N_15493);
and U17481 (N_17481,N_15407,N_14566);
or U17482 (N_17482,N_15403,N_14230);
and U17483 (N_17483,N_14180,N_15923);
or U17484 (N_17484,N_15745,N_14571);
xor U17485 (N_17485,N_15973,N_14636);
nand U17486 (N_17486,N_14093,N_15435);
xnor U17487 (N_17487,N_15051,N_15034);
nand U17488 (N_17488,N_14914,N_15852);
or U17489 (N_17489,N_14899,N_15907);
or U17490 (N_17490,N_15116,N_15614);
and U17491 (N_17491,N_15284,N_14456);
nor U17492 (N_17492,N_15122,N_15452);
or U17493 (N_17493,N_14071,N_14360);
xnor U17494 (N_17494,N_15258,N_15458);
nand U17495 (N_17495,N_14340,N_15010);
xor U17496 (N_17496,N_15735,N_15215);
and U17497 (N_17497,N_15295,N_14575);
xor U17498 (N_17498,N_15649,N_14749);
and U17499 (N_17499,N_14216,N_15698);
xnor U17500 (N_17500,N_14995,N_14521);
nor U17501 (N_17501,N_15172,N_14266);
nand U17502 (N_17502,N_14074,N_14823);
nor U17503 (N_17503,N_14803,N_15536);
and U17504 (N_17504,N_14508,N_14538);
or U17505 (N_17505,N_14990,N_14608);
nand U17506 (N_17506,N_14201,N_15544);
nor U17507 (N_17507,N_15392,N_14492);
nand U17508 (N_17508,N_14638,N_15270);
nand U17509 (N_17509,N_14589,N_14739);
xnor U17510 (N_17510,N_14709,N_14376);
nand U17511 (N_17511,N_15927,N_15947);
nand U17512 (N_17512,N_15790,N_14649);
nor U17513 (N_17513,N_14208,N_15941);
and U17514 (N_17514,N_15810,N_15557);
or U17515 (N_17515,N_14158,N_15893);
or U17516 (N_17516,N_15583,N_14213);
and U17517 (N_17517,N_15217,N_14166);
xnor U17518 (N_17518,N_14776,N_15134);
nor U17519 (N_17519,N_15184,N_15362);
or U17520 (N_17520,N_15521,N_14680);
and U17521 (N_17521,N_15939,N_15880);
xnor U17522 (N_17522,N_15414,N_15588);
nor U17523 (N_17523,N_15275,N_15790);
and U17524 (N_17524,N_14950,N_15532);
xnor U17525 (N_17525,N_14838,N_15033);
nor U17526 (N_17526,N_14678,N_15099);
xnor U17527 (N_17527,N_14748,N_15186);
nor U17528 (N_17528,N_15166,N_14433);
nor U17529 (N_17529,N_15318,N_15856);
or U17530 (N_17530,N_15587,N_14155);
nor U17531 (N_17531,N_14452,N_15544);
and U17532 (N_17532,N_15865,N_14976);
nand U17533 (N_17533,N_14493,N_14542);
xnor U17534 (N_17534,N_15963,N_14278);
xor U17535 (N_17535,N_15119,N_14003);
xor U17536 (N_17536,N_14040,N_15091);
nor U17537 (N_17537,N_14757,N_15307);
xor U17538 (N_17538,N_14064,N_15237);
nand U17539 (N_17539,N_14050,N_14213);
or U17540 (N_17540,N_15117,N_14685);
or U17541 (N_17541,N_15955,N_15360);
and U17542 (N_17542,N_15668,N_14079);
or U17543 (N_17543,N_15587,N_15252);
nand U17544 (N_17544,N_14134,N_15121);
nand U17545 (N_17545,N_14804,N_15416);
nor U17546 (N_17546,N_14459,N_15566);
or U17547 (N_17547,N_14874,N_15432);
nand U17548 (N_17548,N_14592,N_14583);
xor U17549 (N_17549,N_14587,N_14623);
and U17550 (N_17550,N_15435,N_15708);
xnor U17551 (N_17551,N_15137,N_15921);
nand U17552 (N_17552,N_14100,N_15941);
xor U17553 (N_17553,N_15244,N_15298);
or U17554 (N_17554,N_14584,N_15666);
nor U17555 (N_17555,N_14208,N_14533);
xnor U17556 (N_17556,N_15423,N_15114);
nor U17557 (N_17557,N_14399,N_14313);
nor U17558 (N_17558,N_14068,N_15507);
xnor U17559 (N_17559,N_14212,N_15766);
and U17560 (N_17560,N_14046,N_15993);
and U17561 (N_17561,N_14075,N_14669);
nand U17562 (N_17562,N_14822,N_15683);
xor U17563 (N_17563,N_14109,N_15875);
and U17564 (N_17564,N_15068,N_14162);
nor U17565 (N_17565,N_14497,N_15515);
xor U17566 (N_17566,N_14132,N_15987);
or U17567 (N_17567,N_14995,N_14179);
and U17568 (N_17568,N_14568,N_15380);
xnor U17569 (N_17569,N_14404,N_14400);
and U17570 (N_17570,N_15389,N_15948);
or U17571 (N_17571,N_15907,N_14260);
nor U17572 (N_17572,N_14887,N_14567);
xnor U17573 (N_17573,N_14996,N_14745);
xor U17574 (N_17574,N_14585,N_15813);
nand U17575 (N_17575,N_14575,N_14504);
nor U17576 (N_17576,N_15563,N_14646);
nand U17577 (N_17577,N_15614,N_14145);
and U17578 (N_17578,N_15490,N_15612);
and U17579 (N_17579,N_15885,N_15474);
and U17580 (N_17580,N_15411,N_14717);
or U17581 (N_17581,N_15168,N_14922);
or U17582 (N_17582,N_15872,N_15090);
and U17583 (N_17583,N_15369,N_15615);
nor U17584 (N_17584,N_15264,N_15292);
and U17585 (N_17585,N_14460,N_15225);
nor U17586 (N_17586,N_14045,N_15917);
xnor U17587 (N_17587,N_15007,N_15398);
and U17588 (N_17588,N_15611,N_14407);
or U17589 (N_17589,N_14705,N_15726);
and U17590 (N_17590,N_14691,N_15163);
or U17591 (N_17591,N_15290,N_14420);
xor U17592 (N_17592,N_15886,N_15810);
nor U17593 (N_17593,N_15777,N_15804);
or U17594 (N_17594,N_15431,N_14191);
and U17595 (N_17595,N_15705,N_15016);
nand U17596 (N_17596,N_14050,N_15013);
xor U17597 (N_17597,N_15604,N_15480);
xnor U17598 (N_17598,N_14666,N_14908);
nand U17599 (N_17599,N_15711,N_15035);
nor U17600 (N_17600,N_14683,N_14830);
nand U17601 (N_17601,N_14152,N_14871);
nor U17602 (N_17602,N_15088,N_15414);
and U17603 (N_17603,N_15103,N_15272);
xor U17604 (N_17604,N_14339,N_15107);
and U17605 (N_17605,N_14342,N_14585);
and U17606 (N_17606,N_14602,N_15443);
or U17607 (N_17607,N_14553,N_14038);
nor U17608 (N_17608,N_14459,N_15000);
xor U17609 (N_17609,N_15052,N_14253);
nand U17610 (N_17610,N_15679,N_15106);
or U17611 (N_17611,N_14353,N_14808);
nand U17612 (N_17612,N_15964,N_14760);
and U17613 (N_17613,N_15168,N_15667);
nand U17614 (N_17614,N_14821,N_15443);
xnor U17615 (N_17615,N_14372,N_15745);
and U17616 (N_17616,N_14546,N_15597);
and U17617 (N_17617,N_15615,N_15051);
nor U17618 (N_17618,N_14697,N_15516);
nand U17619 (N_17619,N_14477,N_15720);
or U17620 (N_17620,N_14887,N_15164);
xor U17621 (N_17621,N_14792,N_14407);
and U17622 (N_17622,N_15494,N_14042);
and U17623 (N_17623,N_14773,N_15273);
nor U17624 (N_17624,N_15010,N_15960);
or U17625 (N_17625,N_15928,N_14421);
or U17626 (N_17626,N_14769,N_15393);
or U17627 (N_17627,N_15367,N_15756);
and U17628 (N_17628,N_15987,N_15645);
nand U17629 (N_17629,N_15725,N_15219);
or U17630 (N_17630,N_15753,N_15784);
xor U17631 (N_17631,N_14999,N_15595);
or U17632 (N_17632,N_14506,N_15181);
and U17633 (N_17633,N_15741,N_15125);
nor U17634 (N_17634,N_14192,N_14014);
nand U17635 (N_17635,N_14313,N_15099);
and U17636 (N_17636,N_14021,N_14050);
or U17637 (N_17637,N_15887,N_15689);
nor U17638 (N_17638,N_14819,N_15187);
nor U17639 (N_17639,N_14526,N_15157);
nand U17640 (N_17640,N_14140,N_14936);
nor U17641 (N_17641,N_15175,N_14981);
xnor U17642 (N_17642,N_14750,N_15736);
or U17643 (N_17643,N_14886,N_14677);
nor U17644 (N_17644,N_14869,N_15810);
nand U17645 (N_17645,N_14528,N_14997);
or U17646 (N_17646,N_14473,N_15897);
xor U17647 (N_17647,N_14605,N_14442);
nor U17648 (N_17648,N_15715,N_15916);
or U17649 (N_17649,N_15558,N_15148);
nor U17650 (N_17650,N_14591,N_14414);
and U17651 (N_17651,N_15188,N_14746);
or U17652 (N_17652,N_14079,N_14456);
or U17653 (N_17653,N_14008,N_15208);
nand U17654 (N_17654,N_15732,N_15153);
nor U17655 (N_17655,N_15696,N_14367);
nand U17656 (N_17656,N_15968,N_15702);
xor U17657 (N_17657,N_15447,N_15420);
nand U17658 (N_17658,N_15652,N_15075);
nand U17659 (N_17659,N_14450,N_14763);
nand U17660 (N_17660,N_15908,N_14403);
nand U17661 (N_17661,N_15480,N_15857);
nor U17662 (N_17662,N_15383,N_14561);
xnor U17663 (N_17663,N_15798,N_14124);
or U17664 (N_17664,N_14360,N_14830);
nand U17665 (N_17665,N_15361,N_14374);
and U17666 (N_17666,N_14599,N_14777);
nor U17667 (N_17667,N_14122,N_14469);
xor U17668 (N_17668,N_15330,N_14564);
and U17669 (N_17669,N_14393,N_14791);
xnor U17670 (N_17670,N_14930,N_15512);
nand U17671 (N_17671,N_14488,N_15182);
nand U17672 (N_17672,N_15113,N_15045);
and U17673 (N_17673,N_15403,N_14994);
nand U17674 (N_17674,N_14565,N_15624);
or U17675 (N_17675,N_14007,N_14828);
nor U17676 (N_17676,N_15130,N_14200);
and U17677 (N_17677,N_14291,N_15858);
xor U17678 (N_17678,N_14472,N_15126);
and U17679 (N_17679,N_15778,N_14241);
xnor U17680 (N_17680,N_14571,N_15382);
nor U17681 (N_17681,N_15801,N_14246);
nor U17682 (N_17682,N_15789,N_14911);
and U17683 (N_17683,N_15453,N_15439);
and U17684 (N_17684,N_14454,N_14382);
nand U17685 (N_17685,N_15214,N_15535);
or U17686 (N_17686,N_15262,N_15411);
nand U17687 (N_17687,N_15615,N_14190);
xnor U17688 (N_17688,N_15140,N_15858);
nand U17689 (N_17689,N_14466,N_14818);
nor U17690 (N_17690,N_15855,N_14596);
xor U17691 (N_17691,N_14029,N_14637);
and U17692 (N_17692,N_15879,N_15000);
nor U17693 (N_17693,N_14686,N_15114);
xnor U17694 (N_17694,N_15803,N_15457);
or U17695 (N_17695,N_15286,N_14458);
nor U17696 (N_17696,N_14564,N_14714);
or U17697 (N_17697,N_14322,N_15034);
or U17698 (N_17698,N_15179,N_14164);
and U17699 (N_17699,N_15320,N_15696);
and U17700 (N_17700,N_15732,N_15563);
nor U17701 (N_17701,N_15906,N_15339);
and U17702 (N_17702,N_15246,N_15890);
nor U17703 (N_17703,N_14389,N_15861);
and U17704 (N_17704,N_14537,N_14583);
nand U17705 (N_17705,N_15389,N_15056);
nand U17706 (N_17706,N_15530,N_14289);
or U17707 (N_17707,N_15365,N_15636);
and U17708 (N_17708,N_14907,N_15035);
nor U17709 (N_17709,N_14337,N_15982);
nand U17710 (N_17710,N_15400,N_14800);
xnor U17711 (N_17711,N_14235,N_15448);
or U17712 (N_17712,N_14941,N_15436);
nand U17713 (N_17713,N_15407,N_15897);
and U17714 (N_17714,N_15242,N_15785);
or U17715 (N_17715,N_14566,N_14532);
nor U17716 (N_17716,N_15034,N_15258);
nor U17717 (N_17717,N_15882,N_14074);
nor U17718 (N_17718,N_14929,N_14525);
xor U17719 (N_17719,N_15352,N_14532);
nand U17720 (N_17720,N_15748,N_15878);
xor U17721 (N_17721,N_15705,N_14846);
nor U17722 (N_17722,N_15535,N_14023);
nand U17723 (N_17723,N_14648,N_14074);
or U17724 (N_17724,N_14777,N_15381);
and U17725 (N_17725,N_14615,N_14814);
and U17726 (N_17726,N_14215,N_15045);
xnor U17727 (N_17727,N_15764,N_15980);
or U17728 (N_17728,N_15794,N_14984);
nor U17729 (N_17729,N_15789,N_14278);
xnor U17730 (N_17730,N_14897,N_15270);
or U17731 (N_17731,N_14375,N_14137);
and U17732 (N_17732,N_14965,N_14987);
and U17733 (N_17733,N_15930,N_14688);
and U17734 (N_17734,N_15303,N_14825);
xor U17735 (N_17735,N_15328,N_14359);
nor U17736 (N_17736,N_14378,N_14089);
and U17737 (N_17737,N_15229,N_15209);
or U17738 (N_17738,N_14174,N_14807);
xor U17739 (N_17739,N_15999,N_15931);
xnor U17740 (N_17740,N_14106,N_14395);
nand U17741 (N_17741,N_15173,N_15226);
xor U17742 (N_17742,N_15495,N_15167);
or U17743 (N_17743,N_14648,N_14354);
xor U17744 (N_17744,N_15180,N_14021);
and U17745 (N_17745,N_15896,N_15080);
nor U17746 (N_17746,N_15656,N_14166);
nand U17747 (N_17747,N_15197,N_15804);
nor U17748 (N_17748,N_15026,N_15971);
xor U17749 (N_17749,N_15709,N_15222);
xnor U17750 (N_17750,N_15478,N_14051);
xor U17751 (N_17751,N_14027,N_14252);
and U17752 (N_17752,N_15284,N_15130);
nand U17753 (N_17753,N_14005,N_15278);
and U17754 (N_17754,N_15771,N_14982);
or U17755 (N_17755,N_14607,N_14517);
nand U17756 (N_17756,N_14011,N_14844);
xnor U17757 (N_17757,N_15290,N_15429);
nand U17758 (N_17758,N_14581,N_15234);
xor U17759 (N_17759,N_14722,N_15185);
xor U17760 (N_17760,N_15566,N_15363);
nor U17761 (N_17761,N_14627,N_15873);
nor U17762 (N_17762,N_15332,N_14327);
nand U17763 (N_17763,N_15629,N_15587);
nand U17764 (N_17764,N_14643,N_14300);
and U17765 (N_17765,N_15486,N_15846);
nand U17766 (N_17766,N_14439,N_15983);
or U17767 (N_17767,N_15394,N_15261);
nor U17768 (N_17768,N_14425,N_14680);
nand U17769 (N_17769,N_14996,N_15893);
xor U17770 (N_17770,N_15062,N_15646);
xnor U17771 (N_17771,N_14803,N_15321);
or U17772 (N_17772,N_15902,N_14449);
nor U17773 (N_17773,N_15249,N_15151);
xor U17774 (N_17774,N_14043,N_14437);
or U17775 (N_17775,N_15266,N_15073);
nand U17776 (N_17776,N_14771,N_14440);
xor U17777 (N_17777,N_14777,N_14436);
nor U17778 (N_17778,N_14481,N_14688);
and U17779 (N_17779,N_15582,N_15219);
or U17780 (N_17780,N_15372,N_14924);
nor U17781 (N_17781,N_14539,N_15597);
xnor U17782 (N_17782,N_14484,N_15239);
nor U17783 (N_17783,N_14800,N_14724);
xnor U17784 (N_17784,N_15516,N_15239);
nor U17785 (N_17785,N_14254,N_14578);
nand U17786 (N_17786,N_15759,N_15956);
nor U17787 (N_17787,N_14443,N_15976);
nor U17788 (N_17788,N_15355,N_15947);
or U17789 (N_17789,N_15426,N_14193);
nand U17790 (N_17790,N_14157,N_15138);
xnor U17791 (N_17791,N_14627,N_15272);
or U17792 (N_17792,N_14961,N_14989);
or U17793 (N_17793,N_14998,N_15444);
or U17794 (N_17794,N_14774,N_15871);
xnor U17795 (N_17795,N_15330,N_14465);
nand U17796 (N_17796,N_15574,N_15082);
or U17797 (N_17797,N_14979,N_14331);
or U17798 (N_17798,N_14272,N_15192);
and U17799 (N_17799,N_14933,N_15236);
xnor U17800 (N_17800,N_14529,N_15107);
and U17801 (N_17801,N_15305,N_15837);
and U17802 (N_17802,N_14182,N_14404);
nor U17803 (N_17803,N_14733,N_15033);
and U17804 (N_17804,N_14280,N_14486);
nor U17805 (N_17805,N_15475,N_14194);
or U17806 (N_17806,N_14943,N_15726);
nand U17807 (N_17807,N_15021,N_14552);
or U17808 (N_17808,N_15312,N_14878);
xnor U17809 (N_17809,N_15140,N_15605);
nor U17810 (N_17810,N_15850,N_14827);
nor U17811 (N_17811,N_15237,N_15315);
or U17812 (N_17812,N_14089,N_15018);
and U17813 (N_17813,N_14394,N_15302);
or U17814 (N_17814,N_15849,N_14313);
xnor U17815 (N_17815,N_14191,N_14115);
xnor U17816 (N_17816,N_14477,N_15177);
or U17817 (N_17817,N_14970,N_14550);
nand U17818 (N_17818,N_14508,N_15125);
and U17819 (N_17819,N_14593,N_15451);
xor U17820 (N_17820,N_15935,N_15801);
nand U17821 (N_17821,N_14907,N_15931);
xnor U17822 (N_17822,N_15691,N_15005);
nor U17823 (N_17823,N_15534,N_15124);
xnor U17824 (N_17824,N_14213,N_14501);
xnor U17825 (N_17825,N_15868,N_15934);
xnor U17826 (N_17826,N_14868,N_15373);
nand U17827 (N_17827,N_15128,N_14342);
or U17828 (N_17828,N_14547,N_14475);
nor U17829 (N_17829,N_14465,N_14649);
nor U17830 (N_17830,N_14266,N_14888);
xnor U17831 (N_17831,N_14365,N_15912);
xnor U17832 (N_17832,N_14915,N_14559);
xor U17833 (N_17833,N_14130,N_14524);
xnor U17834 (N_17834,N_15775,N_15064);
or U17835 (N_17835,N_14528,N_15292);
xnor U17836 (N_17836,N_15016,N_15120);
xor U17837 (N_17837,N_14590,N_14675);
nor U17838 (N_17838,N_15903,N_14290);
and U17839 (N_17839,N_14995,N_14347);
or U17840 (N_17840,N_14660,N_15500);
and U17841 (N_17841,N_15133,N_15247);
xnor U17842 (N_17842,N_14929,N_14347);
or U17843 (N_17843,N_15321,N_14111);
nand U17844 (N_17844,N_14756,N_15409);
or U17845 (N_17845,N_14175,N_15275);
nor U17846 (N_17846,N_15336,N_14010);
or U17847 (N_17847,N_14544,N_15313);
nand U17848 (N_17848,N_14097,N_15391);
nand U17849 (N_17849,N_15894,N_15717);
nor U17850 (N_17850,N_15976,N_14827);
and U17851 (N_17851,N_15969,N_15468);
xnor U17852 (N_17852,N_14956,N_14685);
nor U17853 (N_17853,N_15346,N_14754);
or U17854 (N_17854,N_14656,N_15051);
and U17855 (N_17855,N_14722,N_15361);
and U17856 (N_17856,N_14879,N_15672);
xor U17857 (N_17857,N_15958,N_15638);
xor U17858 (N_17858,N_14396,N_15365);
and U17859 (N_17859,N_15778,N_15839);
and U17860 (N_17860,N_14267,N_15145);
nand U17861 (N_17861,N_14827,N_14806);
and U17862 (N_17862,N_14863,N_15601);
xnor U17863 (N_17863,N_14560,N_15840);
xnor U17864 (N_17864,N_14897,N_15287);
and U17865 (N_17865,N_15023,N_15983);
nand U17866 (N_17866,N_14423,N_15116);
or U17867 (N_17867,N_15303,N_15601);
or U17868 (N_17868,N_15554,N_15828);
or U17869 (N_17869,N_15970,N_14515);
and U17870 (N_17870,N_14831,N_14854);
xnor U17871 (N_17871,N_14934,N_15912);
or U17872 (N_17872,N_14664,N_15891);
nor U17873 (N_17873,N_14032,N_14797);
xnor U17874 (N_17874,N_15106,N_15546);
nand U17875 (N_17875,N_15176,N_14467);
or U17876 (N_17876,N_15294,N_15002);
nand U17877 (N_17877,N_14647,N_15635);
or U17878 (N_17878,N_15423,N_14105);
xor U17879 (N_17879,N_14863,N_15213);
or U17880 (N_17880,N_14868,N_14025);
or U17881 (N_17881,N_15278,N_14496);
nor U17882 (N_17882,N_15071,N_14366);
or U17883 (N_17883,N_15255,N_14289);
and U17884 (N_17884,N_15445,N_14090);
nor U17885 (N_17885,N_15190,N_15346);
xor U17886 (N_17886,N_15297,N_14601);
or U17887 (N_17887,N_14845,N_15621);
and U17888 (N_17888,N_15168,N_14136);
nor U17889 (N_17889,N_14228,N_14436);
and U17890 (N_17890,N_15683,N_14916);
or U17891 (N_17891,N_15252,N_15766);
nand U17892 (N_17892,N_14465,N_15868);
or U17893 (N_17893,N_14316,N_14380);
and U17894 (N_17894,N_15931,N_14882);
nand U17895 (N_17895,N_14890,N_15023);
and U17896 (N_17896,N_14610,N_14551);
nor U17897 (N_17897,N_15889,N_15376);
nand U17898 (N_17898,N_15464,N_15217);
nand U17899 (N_17899,N_15604,N_15767);
nand U17900 (N_17900,N_14565,N_15660);
and U17901 (N_17901,N_15946,N_14484);
nand U17902 (N_17902,N_14143,N_15053);
xnor U17903 (N_17903,N_15615,N_15056);
or U17904 (N_17904,N_15481,N_15131);
xnor U17905 (N_17905,N_15526,N_15767);
xnor U17906 (N_17906,N_14711,N_14227);
and U17907 (N_17907,N_15645,N_14463);
and U17908 (N_17908,N_15495,N_14420);
and U17909 (N_17909,N_15880,N_15760);
or U17910 (N_17910,N_15562,N_14004);
nor U17911 (N_17911,N_15665,N_14021);
and U17912 (N_17912,N_14387,N_15067);
nor U17913 (N_17913,N_14059,N_15349);
nand U17914 (N_17914,N_15732,N_14109);
and U17915 (N_17915,N_14933,N_14428);
nand U17916 (N_17916,N_15856,N_14707);
or U17917 (N_17917,N_14596,N_14137);
and U17918 (N_17918,N_15586,N_15177);
or U17919 (N_17919,N_15000,N_15727);
nor U17920 (N_17920,N_15910,N_14989);
or U17921 (N_17921,N_14033,N_15967);
or U17922 (N_17922,N_15968,N_15296);
and U17923 (N_17923,N_15325,N_14246);
or U17924 (N_17924,N_14022,N_15990);
or U17925 (N_17925,N_14791,N_15149);
xor U17926 (N_17926,N_15202,N_14853);
and U17927 (N_17927,N_15861,N_14109);
nor U17928 (N_17928,N_14732,N_15783);
and U17929 (N_17929,N_14430,N_14435);
or U17930 (N_17930,N_15666,N_14360);
xnor U17931 (N_17931,N_15958,N_14497);
nand U17932 (N_17932,N_14981,N_14933);
xnor U17933 (N_17933,N_15202,N_15177);
nor U17934 (N_17934,N_15398,N_15227);
nand U17935 (N_17935,N_14938,N_15190);
and U17936 (N_17936,N_15784,N_14471);
nor U17937 (N_17937,N_14585,N_15152);
nand U17938 (N_17938,N_14955,N_15400);
nand U17939 (N_17939,N_14284,N_15640);
xnor U17940 (N_17940,N_15295,N_15704);
nor U17941 (N_17941,N_14963,N_14394);
nor U17942 (N_17942,N_14956,N_14073);
nor U17943 (N_17943,N_15974,N_14882);
nor U17944 (N_17944,N_14445,N_15010);
nand U17945 (N_17945,N_15450,N_14417);
nand U17946 (N_17946,N_14437,N_15950);
xor U17947 (N_17947,N_14036,N_15025);
xnor U17948 (N_17948,N_14345,N_15601);
and U17949 (N_17949,N_14695,N_14602);
nor U17950 (N_17950,N_15177,N_15745);
and U17951 (N_17951,N_15149,N_14091);
nor U17952 (N_17952,N_14076,N_15139);
xnor U17953 (N_17953,N_14133,N_14874);
and U17954 (N_17954,N_15962,N_14803);
and U17955 (N_17955,N_15255,N_15448);
and U17956 (N_17956,N_15312,N_14272);
nor U17957 (N_17957,N_15238,N_15713);
nand U17958 (N_17958,N_15205,N_14415);
nor U17959 (N_17959,N_14045,N_14027);
and U17960 (N_17960,N_15133,N_14939);
nor U17961 (N_17961,N_15778,N_14059);
and U17962 (N_17962,N_14994,N_14576);
nor U17963 (N_17963,N_15007,N_14539);
nand U17964 (N_17964,N_15181,N_15249);
xnor U17965 (N_17965,N_15430,N_15814);
nor U17966 (N_17966,N_14703,N_14502);
or U17967 (N_17967,N_15133,N_15551);
or U17968 (N_17968,N_14936,N_14763);
xor U17969 (N_17969,N_15422,N_14202);
xnor U17970 (N_17970,N_15804,N_15605);
and U17971 (N_17971,N_14830,N_14341);
nor U17972 (N_17972,N_14656,N_14731);
xor U17973 (N_17973,N_15576,N_14850);
nor U17974 (N_17974,N_14201,N_14227);
or U17975 (N_17975,N_15480,N_15643);
or U17976 (N_17976,N_15909,N_14447);
nand U17977 (N_17977,N_14444,N_15781);
xor U17978 (N_17978,N_15790,N_14980);
nand U17979 (N_17979,N_15293,N_15466);
nand U17980 (N_17980,N_15824,N_15097);
or U17981 (N_17981,N_15063,N_15387);
xor U17982 (N_17982,N_15390,N_15999);
nor U17983 (N_17983,N_14123,N_15002);
xor U17984 (N_17984,N_15759,N_15921);
nand U17985 (N_17985,N_15150,N_15225);
and U17986 (N_17986,N_15933,N_15069);
nor U17987 (N_17987,N_14847,N_15351);
xnor U17988 (N_17988,N_14130,N_14699);
and U17989 (N_17989,N_14118,N_14106);
nand U17990 (N_17990,N_15744,N_15953);
xnor U17991 (N_17991,N_15370,N_15180);
and U17992 (N_17992,N_14000,N_14240);
and U17993 (N_17993,N_15107,N_15996);
and U17994 (N_17994,N_15541,N_14915);
or U17995 (N_17995,N_14698,N_14334);
nor U17996 (N_17996,N_14203,N_14519);
and U17997 (N_17997,N_15475,N_15180);
and U17998 (N_17998,N_15929,N_15590);
nor U17999 (N_17999,N_15714,N_14254);
and U18000 (N_18000,N_16856,N_16880);
or U18001 (N_18001,N_16310,N_17743);
xnor U18002 (N_18002,N_16592,N_17288);
xor U18003 (N_18003,N_16632,N_17494);
or U18004 (N_18004,N_16874,N_17291);
nor U18005 (N_18005,N_16468,N_17292);
xnor U18006 (N_18006,N_16922,N_17980);
and U18007 (N_18007,N_17495,N_17393);
nor U18008 (N_18008,N_17848,N_16697);
or U18009 (N_18009,N_16802,N_16510);
and U18010 (N_18010,N_17294,N_17186);
nand U18011 (N_18011,N_17118,N_16025);
nand U18012 (N_18012,N_16463,N_17509);
nor U18013 (N_18013,N_17303,N_16116);
nor U18014 (N_18014,N_16607,N_16621);
xnor U18015 (N_18015,N_17085,N_17939);
nand U18016 (N_18016,N_17368,N_16040);
and U18017 (N_18017,N_16174,N_17219);
nor U18018 (N_18018,N_16909,N_16213);
nand U18019 (N_18019,N_16228,N_17811);
nor U18020 (N_18020,N_17719,N_16866);
nor U18021 (N_18021,N_17262,N_17735);
and U18022 (N_18022,N_17637,N_16104);
xnor U18023 (N_18023,N_17856,N_17968);
or U18024 (N_18024,N_17401,N_16290);
or U18025 (N_18025,N_16636,N_17164);
xor U18026 (N_18026,N_16059,N_17499);
xnor U18027 (N_18027,N_16189,N_17756);
nor U18028 (N_18028,N_17093,N_16335);
nand U18029 (N_18029,N_16926,N_16186);
nand U18030 (N_18030,N_16937,N_16549);
nor U18031 (N_18031,N_17124,N_16606);
or U18032 (N_18032,N_16226,N_16391);
or U18033 (N_18033,N_17923,N_16865);
nor U18034 (N_18034,N_17363,N_16265);
and U18035 (N_18035,N_16207,N_17297);
xor U18036 (N_18036,N_17145,N_17695);
nand U18037 (N_18037,N_17688,N_16431);
nand U18038 (N_18038,N_17081,N_17705);
nor U18039 (N_18039,N_17628,N_17766);
nor U18040 (N_18040,N_17448,N_17862);
xor U18041 (N_18041,N_17112,N_17526);
and U18042 (N_18042,N_17426,N_16884);
xor U18043 (N_18043,N_16185,N_16959);
nand U18044 (N_18044,N_16602,N_16058);
and U18045 (N_18045,N_16850,N_17801);
nor U18046 (N_18046,N_17813,N_17435);
and U18047 (N_18047,N_17308,N_17272);
nor U18048 (N_18048,N_17890,N_17563);
xor U18049 (N_18049,N_17236,N_16048);
and U18050 (N_18050,N_17534,N_16181);
and U18051 (N_18051,N_17892,N_16947);
or U18052 (N_18052,N_17433,N_16542);
and U18053 (N_18053,N_17804,N_16485);
and U18054 (N_18054,N_17920,N_17834);
nand U18055 (N_18055,N_17972,N_17136);
and U18056 (N_18056,N_16599,N_16410);
xnor U18057 (N_18057,N_16751,N_17720);
nor U18058 (N_18058,N_16656,N_17781);
or U18059 (N_18059,N_17990,N_17907);
xnor U18060 (N_18060,N_17046,N_16035);
nor U18061 (N_18061,N_17427,N_16872);
xnor U18062 (N_18062,N_16562,N_17127);
or U18063 (N_18063,N_16669,N_17226);
and U18064 (N_18064,N_17455,N_16683);
xor U18065 (N_18065,N_16440,N_16852);
and U18066 (N_18066,N_16948,N_17643);
xor U18067 (N_18067,N_17020,N_16543);
nor U18068 (N_18068,N_16408,N_17174);
and U18069 (N_18069,N_16445,N_17881);
and U18070 (N_18070,N_17784,N_17759);
and U18071 (N_18071,N_17536,N_16817);
nand U18072 (N_18072,N_17828,N_17649);
nor U18073 (N_18073,N_16140,N_16955);
xnor U18074 (N_18074,N_17909,N_17931);
and U18075 (N_18075,N_16101,N_16826);
xnor U18076 (N_18076,N_16438,N_17454);
nand U18077 (N_18077,N_17449,N_17380);
nor U18078 (N_18078,N_16509,N_17281);
xnor U18079 (N_18079,N_17561,N_16582);
or U18080 (N_18080,N_16991,N_17018);
and U18081 (N_18081,N_16105,N_17691);
xnor U18082 (N_18082,N_16491,N_16862);
nand U18083 (N_18083,N_16687,N_17717);
nor U18084 (N_18084,N_17780,N_16647);
xor U18085 (N_18085,N_16833,N_16779);
or U18086 (N_18086,N_17192,N_16306);
nor U18087 (N_18087,N_17234,N_17230);
xnor U18088 (N_18088,N_17535,N_16120);
nor U18089 (N_18089,N_17604,N_16529);
xnor U18090 (N_18090,N_16453,N_16029);
and U18091 (N_18091,N_16601,N_16635);
nand U18092 (N_18092,N_16313,N_17932);
nor U18093 (N_18093,N_16329,N_16027);
nand U18094 (N_18094,N_17423,N_16848);
nor U18095 (N_18095,N_16286,N_17581);
and U18096 (N_18096,N_17102,N_17988);
or U18097 (N_18097,N_17753,N_17876);
nand U18098 (N_18098,N_16489,N_16768);
nor U18099 (N_18099,N_16405,N_16616);
or U18100 (N_18100,N_16983,N_16237);
or U18101 (N_18101,N_17944,N_16071);
or U18102 (N_18102,N_17520,N_17082);
or U18103 (N_18103,N_17502,N_17524);
xor U18104 (N_18104,N_17383,N_17598);
and U18105 (N_18105,N_16704,N_17098);
nor U18106 (N_18106,N_17023,N_17579);
nor U18107 (N_18107,N_16421,N_16209);
nand U18108 (N_18108,N_16744,N_16422);
xnor U18109 (N_18109,N_17077,N_17349);
nand U18110 (N_18110,N_17653,N_17319);
or U18111 (N_18111,N_17715,N_16590);
nor U18112 (N_18112,N_17739,N_17338);
nor U18113 (N_18113,N_16674,N_16091);
and U18114 (N_18114,N_17417,N_16586);
nand U18115 (N_18115,N_16709,N_16062);
and U18116 (N_18116,N_16426,N_16544);
nand U18117 (N_18117,N_17721,N_16096);
or U18118 (N_18118,N_17877,N_17012);
and U18119 (N_18119,N_17964,N_16749);
nand U18120 (N_18120,N_17318,N_16578);
nor U18121 (N_18121,N_16006,N_16844);
xor U18122 (N_18122,N_16811,N_16508);
nand U18123 (N_18123,N_16386,N_17492);
and U18124 (N_18124,N_16712,N_16879);
and U18125 (N_18125,N_17440,N_16974);
xnor U18126 (N_18126,N_16016,N_17062);
nand U18127 (N_18127,N_17031,N_16137);
and U18128 (N_18128,N_17962,N_17976);
nor U18129 (N_18129,N_17960,N_16256);
or U18130 (N_18130,N_16436,N_17884);
xnor U18131 (N_18131,N_17723,N_16383);
nor U18132 (N_18132,N_16156,N_17092);
nor U18133 (N_18133,N_17341,N_17106);
nor U18134 (N_18134,N_17444,N_17107);
or U18135 (N_18135,N_16633,N_17882);
nand U18136 (N_18136,N_17463,N_16328);
or U18137 (N_18137,N_17704,N_17070);
nor U18138 (N_18138,N_17994,N_17914);
or U18139 (N_18139,N_16278,N_16846);
xor U18140 (N_18140,N_17625,N_17546);
nor U18141 (N_18141,N_16017,N_17282);
xor U18142 (N_18142,N_17360,N_17168);
xor U18143 (N_18143,N_16610,N_16989);
nand U18144 (N_18144,N_17618,N_16611);
xor U18145 (N_18145,N_16694,N_17908);
xnor U18146 (N_18146,N_16793,N_17453);
nand U18147 (N_18147,N_16452,N_17068);
nor U18148 (N_18148,N_16681,N_16138);
nand U18149 (N_18149,N_16663,N_16293);
nor U18150 (N_18150,N_16679,N_16796);
nand U18151 (N_18151,N_16492,N_17396);
or U18152 (N_18152,N_17539,N_17952);
or U18153 (N_18153,N_17104,N_17767);
xnor U18154 (N_18154,N_16588,N_17265);
and U18155 (N_18155,N_16081,N_16842);
or U18156 (N_18156,N_17725,N_17777);
xnor U18157 (N_18157,N_16579,N_16362);
or U18158 (N_18158,N_17842,N_16248);
or U18159 (N_18159,N_17824,N_17967);
xnor U18160 (N_18160,N_17608,N_16394);
or U18161 (N_18161,N_16314,N_16855);
nand U18162 (N_18162,N_16953,N_17622);
and U18163 (N_18163,N_16118,N_16942);
nand U18164 (N_18164,N_16200,N_16164);
or U18165 (N_18165,N_17017,N_17010);
xnor U18166 (N_18166,N_17026,N_17627);
and U18167 (N_18167,N_17574,N_16132);
nor U18168 (N_18168,N_17763,N_16502);
nor U18169 (N_18169,N_17887,N_17633);
or U18170 (N_18170,N_16057,N_16785);
and U18171 (N_18171,N_17241,N_16242);
xor U18172 (N_18172,N_17209,N_16399);
xnor U18173 (N_18173,N_16157,N_17126);
nand U18174 (N_18174,N_17754,N_17501);
nand U18175 (N_18175,N_17436,N_17312);
xor U18176 (N_18176,N_17771,N_16659);
nor U18177 (N_18177,N_17762,N_17961);
or U18178 (N_18178,N_16678,N_16158);
and U18179 (N_18179,N_17225,N_16318);
or U18180 (N_18180,N_16475,N_17530);
and U18181 (N_18181,N_17442,N_17403);
or U18182 (N_18182,N_17275,N_16946);
xor U18183 (N_18183,N_17028,N_16945);
nor U18184 (N_18184,N_16890,N_17395);
nand U18185 (N_18185,N_17242,N_17858);
or U18186 (N_18186,N_16642,N_17567);
nand U18187 (N_18187,N_16370,N_17337);
or U18188 (N_18188,N_17505,N_16086);
nand U18189 (N_18189,N_17684,N_16925);
nand U18190 (N_18190,N_17222,N_17518);
and U18191 (N_18191,N_16134,N_16756);
or U18192 (N_18192,N_17795,N_16790);
xor U18193 (N_18193,N_17983,N_17918);
or U18194 (N_18194,N_16834,N_16653);
and U18195 (N_18195,N_17666,N_17532);
nand U18196 (N_18196,N_17991,N_17954);
xor U18197 (N_18197,N_17016,N_17064);
or U18198 (N_18198,N_17184,N_16446);
xor U18199 (N_18199,N_16280,N_16652);
xnor U18200 (N_18200,N_16353,N_16645);
and U18201 (N_18201,N_16604,N_17090);
nand U18202 (N_18202,N_16486,N_17354);
xnor U18203 (N_18203,N_16902,N_17927);
nand U18204 (N_18204,N_16295,N_16513);
xor U18205 (N_18205,N_16819,N_16803);
nand U18206 (N_18206,N_16605,N_17531);
and U18207 (N_18207,N_16364,N_16589);
and U18208 (N_18208,N_17747,N_16994);
and U18209 (N_18209,N_17897,N_16985);
and U18210 (N_18210,N_16236,N_17768);
and U18211 (N_18211,N_16932,N_16342);
nor U18212 (N_18212,N_16375,N_17317);
and U18213 (N_18213,N_17080,N_17021);
or U18214 (N_18214,N_17676,N_16480);
or U18215 (N_18215,N_16730,N_17218);
nand U18216 (N_18216,N_17979,N_17738);
nand U18217 (N_18217,N_16461,N_16069);
or U18218 (N_18218,N_16352,N_17537);
nor U18219 (N_18219,N_16312,N_16095);
nor U18220 (N_18220,N_16759,N_16193);
or U18221 (N_18221,N_16943,N_17592);
or U18222 (N_18222,N_16877,N_17468);
or U18223 (N_18223,N_16952,N_16056);
xnor U18224 (N_18224,N_16054,N_16690);
nor U18225 (N_18225,N_17036,N_16684);
nor U18226 (N_18226,N_17957,N_17141);
xnor U18227 (N_18227,N_17330,N_16246);
nand U18228 (N_18228,N_17500,N_17549);
xor U18229 (N_18229,N_17573,N_16051);
or U18230 (N_18230,N_16011,N_16417);
nand U18231 (N_18231,N_16359,N_17673);
xor U18232 (N_18232,N_17840,N_16028);
nand U18233 (N_18233,N_16222,N_16668);
xnor U18234 (N_18234,N_16532,N_17470);
or U18235 (N_18235,N_16389,N_16563);
xnor U18236 (N_18236,N_16619,N_17818);
nor U18237 (N_18237,N_17517,N_16007);
xnor U18238 (N_18238,N_17378,N_17353);
or U18239 (N_18239,N_17034,N_16454);
nand U18240 (N_18240,N_16045,N_17324);
nor U18241 (N_18241,N_17343,N_16487);
nand U18242 (N_18242,N_17415,N_17243);
and U18243 (N_18243,N_16337,N_16765);
xnor U18244 (N_18244,N_17488,N_16898);
nand U18245 (N_18245,N_16908,N_16240);
and U18246 (N_18246,N_16341,N_16176);
nor U18247 (N_18247,N_17091,N_16559);
and U18248 (N_18248,N_17389,N_16581);
nor U18249 (N_18249,N_16249,N_17414);
or U18250 (N_18250,N_17646,N_16757);
xnor U18251 (N_18251,N_17256,N_16212);
nand U18252 (N_18252,N_17372,N_17235);
or U18253 (N_18253,N_16476,N_17086);
xnor U18254 (N_18254,N_16807,N_17726);
xnor U18255 (N_18255,N_16205,N_16919);
and U18256 (N_18256,N_17659,N_16488);
nor U18257 (N_18257,N_17003,N_16307);
nand U18258 (N_18258,N_16875,N_17366);
xor U18259 (N_18259,N_16015,N_17683);
nand U18260 (N_18260,N_16350,N_16130);
xnor U18261 (N_18261,N_16651,N_16064);
nor U18262 (N_18262,N_16360,N_16847);
or U18263 (N_18263,N_16407,N_17589);
nand U18264 (N_18264,N_17689,N_16971);
and U18265 (N_18265,N_16496,N_17156);
and U18266 (N_18266,N_17279,N_17461);
and U18267 (N_18267,N_17117,N_17004);
nand U18268 (N_18268,N_17129,N_16764);
nor U18269 (N_18269,N_17806,N_17079);
nand U18270 (N_18270,N_16675,N_16172);
or U18271 (N_18271,N_17377,N_17571);
nand U18272 (N_18272,N_17917,N_16477);
or U18273 (N_18273,N_16973,N_16799);
nand U18274 (N_18274,N_16152,N_17072);
nor U18275 (N_18275,N_16747,N_16354);
nor U18276 (N_18276,N_16680,N_17822);
nand U18277 (N_18277,N_16878,N_17859);
nor U18278 (N_18278,N_16813,N_16624);
nor U18279 (N_18279,N_16433,N_17493);
or U18280 (N_18280,N_16899,N_16385);
nor U18281 (N_18281,N_17166,N_16661);
nand U18282 (N_18282,N_17221,N_17042);
or U18283 (N_18283,N_17560,N_17307);
xor U18284 (N_18284,N_16083,N_17247);
xnor U18285 (N_18285,N_17327,N_16725);
xor U18286 (N_18286,N_16886,N_16494);
nand U18287 (N_18287,N_16264,N_16424);
nor U18288 (N_18288,N_16892,N_16639);
and U18289 (N_18289,N_16821,N_17176);
nand U18290 (N_18290,N_16416,N_16810);
nand U18291 (N_18291,N_16522,N_16202);
and U18292 (N_18292,N_16311,N_17253);
nor U18293 (N_18293,N_16792,N_17421);
or U18294 (N_18294,N_17621,N_16349);
nor U18295 (N_18295,N_16267,N_17938);
nand U18296 (N_18296,N_16055,N_17992);
xnor U18297 (N_18297,N_17496,N_17473);
or U18298 (N_18298,N_16568,N_17728);
and U18299 (N_18299,N_16148,N_17466);
nor U18300 (N_18300,N_16478,N_17851);
nor U18301 (N_18301,N_17748,N_17749);
nor U18302 (N_18302,N_17438,N_17044);
nand U18303 (N_18303,N_17981,N_17159);
nand U18304 (N_18304,N_17147,N_16037);
and U18305 (N_18305,N_17973,N_16646);
or U18306 (N_18306,N_17119,N_16975);
or U18307 (N_18307,N_17609,N_16501);
or U18308 (N_18308,N_17541,N_17151);
nand U18309 (N_18309,N_16672,N_17565);
xor U18310 (N_18310,N_16517,N_16851);
or U18311 (N_18311,N_16020,N_17919);
nor U18312 (N_18312,N_17788,N_17173);
nand U18313 (N_18313,N_17569,N_16565);
nand U18314 (N_18314,N_16644,N_17706);
and U18315 (N_18315,N_17032,N_17479);
or U18316 (N_18316,N_16634,N_16882);
nand U18317 (N_18317,N_17975,N_16887);
nand U18318 (N_18318,N_16187,N_16753);
or U18319 (N_18319,N_17290,N_16182);
xnor U18320 (N_18320,N_16603,N_17358);
nor U18321 (N_18321,N_17266,N_17911);
or U18322 (N_18322,N_16251,N_16357);
nand U18323 (N_18323,N_17740,N_16178);
or U18324 (N_18324,N_16963,N_17451);
nor U18325 (N_18325,N_16239,N_16085);
xor U18326 (N_18326,N_16993,N_17103);
xor U18327 (N_18327,N_17200,N_16155);
or U18328 (N_18328,N_16881,N_17629);
or U18329 (N_18329,N_16888,N_17602);
nand U18330 (N_18330,N_17915,N_16854);
nor U18331 (N_18331,N_17867,N_17736);
or U18332 (N_18332,N_17644,N_16470);
nor U18333 (N_18333,N_17286,N_17323);
or U18334 (N_18334,N_16863,N_17654);
and U18335 (N_18335,N_16752,N_16358);
nand U18336 (N_18336,N_17175,N_16458);
nand U18337 (N_18337,N_16308,N_17464);
or U18338 (N_18338,N_16270,N_16840);
nand U18339 (N_18339,N_17478,N_17902);
or U18340 (N_18340,N_17959,N_16710);
nand U18341 (N_18341,N_16112,N_17237);
xor U18342 (N_18342,N_17424,N_17187);
xor U18343 (N_18343,N_17154,N_17316);
or U18344 (N_18344,N_16664,N_16536);
nand U18345 (N_18345,N_16225,N_16783);
nand U18346 (N_18346,N_16995,N_16596);
and U18347 (N_18347,N_17277,N_17658);
nor U18348 (N_18348,N_17065,N_17583);
or U18349 (N_18349,N_16595,N_16805);
or U18350 (N_18350,N_17808,N_16727);
nand U18351 (N_18351,N_16419,N_16272);
xor U18352 (N_18352,N_16940,N_17146);
xnor U18353 (N_18353,N_17181,N_16654);
or U18354 (N_18354,N_17190,N_16093);
or U18355 (N_18355,N_17336,N_16514);
xnor U18356 (N_18356,N_17447,N_17697);
or U18357 (N_18357,N_16982,N_16450);
and U18358 (N_18358,N_16292,N_17727);
and U18359 (N_18359,N_17309,N_17109);
or U18360 (N_18360,N_17203,N_16073);
nor U18361 (N_18361,N_17678,N_16666);
xor U18362 (N_18362,N_17572,N_16122);
and U18363 (N_18363,N_16920,N_17205);
nand U18364 (N_18364,N_16766,N_17969);
xnor U18365 (N_18365,N_16526,N_16080);
nand U18366 (N_18366,N_17165,N_17669);
and U18367 (N_18367,N_16493,N_16170);
or U18368 (N_18368,N_16570,N_17467);
xor U18369 (N_18369,N_16662,N_16466);
nand U18370 (N_18370,N_17320,N_16692);
or U18371 (N_18371,N_16079,N_17095);
xor U18372 (N_18372,N_17367,N_17460);
and U18373 (N_18373,N_17667,N_16021);
nand U18374 (N_18374,N_17278,N_17681);
xnor U18375 (N_18375,N_16797,N_16125);
nand U18376 (N_18376,N_16530,N_17638);
nor U18377 (N_18377,N_16685,N_16490);
nor U18378 (N_18378,N_17935,N_16503);
nand U18379 (N_18379,N_17830,N_16323);
nor U18380 (N_18380,N_17562,N_17364);
and U18381 (N_18381,N_17158,N_16572);
nor U18382 (N_18382,N_16716,N_17038);
nor U18383 (N_18383,N_17742,N_16627);
nor U18384 (N_18384,N_17326,N_17099);
or U18385 (N_18385,N_17543,N_17100);
nand U18386 (N_18386,N_16771,N_16822);
or U18387 (N_18387,N_17069,N_17160);
xnor U18388 (N_18388,N_17547,N_17239);
nor U18389 (N_18389,N_16388,N_16906);
nand U18390 (N_18390,N_16343,N_16441);
nor U18391 (N_18391,N_17829,N_16184);
or U18392 (N_18392,N_17770,N_16124);
or U18393 (N_18393,N_16188,N_16074);
nand U18394 (N_18394,N_17937,N_16520);
xor U18395 (N_18395,N_17556,N_17115);
xor U18396 (N_18396,N_16843,N_16696);
xor U18397 (N_18397,N_17694,N_17839);
nor U18398 (N_18398,N_17873,N_16327);
and U18399 (N_18399,N_17752,N_17554);
nand U18400 (N_18400,N_16857,N_16050);
xnor U18401 (N_18401,N_17246,N_16257);
and U18402 (N_18402,N_17402,N_17198);
nor U18403 (N_18403,N_16469,N_16097);
xor U18404 (N_18404,N_16179,N_16333);
xor U18405 (N_18405,N_16827,N_17861);
nor U18406 (N_18406,N_16474,N_17287);
or U18407 (N_18407,N_16598,N_16317);
nor U18408 (N_18408,N_17514,N_16889);
nor U18409 (N_18409,N_17207,N_16760);
nor U18410 (N_18410,N_17305,N_16141);
nand U18411 (N_18411,N_16110,N_16550);
nor U18412 (N_18412,N_16976,N_16845);
nand U18413 (N_18413,N_16700,N_17950);
xnor U18414 (N_18414,N_17899,N_17180);
nand U18415 (N_18415,N_16065,N_17280);
nand U18416 (N_18416,N_17685,N_16558);
or U18417 (N_18417,N_17452,N_16289);
nand U18418 (N_18418,N_16557,N_17974);
nor U18419 (N_18419,N_16398,N_16401);
and U18420 (N_18420,N_17816,N_17929);
and U18421 (N_18421,N_16540,N_16484);
nor U18422 (N_18422,N_16935,N_17465);
nand U18423 (N_18423,N_16832,N_17716);
nand U18424 (N_18424,N_17564,N_17626);
or U18425 (N_18425,N_17984,N_17648);
and U18426 (N_18426,N_17388,N_16263);
nand U18427 (N_18427,N_16835,N_17373);
xor U18428 (N_18428,N_17963,N_16192);
and U18429 (N_18429,N_17379,N_16523);
or U18430 (N_18430,N_17111,N_17369);
and U18431 (N_18431,N_17789,N_16098);
and U18432 (N_18432,N_16271,N_16334);
and U18433 (N_18433,N_16916,N_16411);
xor U18434 (N_18434,N_16658,N_17037);
xnor U18435 (N_18435,N_16511,N_16736);
and U18436 (N_18436,N_16117,N_17613);
xor U18437 (N_18437,N_16036,N_16600);
and U18438 (N_18438,N_17672,N_17157);
xnor U18439 (N_18439,N_17989,N_17477);
and U18440 (N_18440,N_17596,N_17712);
nand U18441 (N_18441,N_17482,N_16699);
nor U18442 (N_18442,N_16076,N_17866);
nand U18443 (N_18443,N_16698,N_16229);
or U18444 (N_18444,N_16622,N_17067);
nor U18445 (N_18445,N_17193,N_16052);
xnor U18446 (N_18446,N_16153,N_16042);
and U18447 (N_18447,N_16163,N_17522);
or U18448 (N_18448,N_17122,N_17844);
nor U18449 (N_18449,N_16135,N_17506);
or U18450 (N_18450,N_17891,N_17610);
and U18451 (N_18451,N_17630,N_16527);
xor U18452 (N_18452,N_17179,N_16034);
or U18453 (N_18453,N_17833,N_17250);
or U18454 (N_18454,N_17051,N_17843);
or U18455 (N_18455,N_16113,N_17584);
or U18456 (N_18456,N_16738,N_17521);
xnor U18457 (N_18457,N_17878,N_17139);
nand U18458 (N_18458,N_16418,N_17285);
nand U18459 (N_18459,N_16957,N_17778);
xnor U18460 (N_18460,N_16238,N_16321);
or U18461 (N_18461,N_16951,N_16719);
and U18462 (N_18462,N_16537,N_16183);
xor U18463 (N_18463,N_17276,N_17013);
and U18464 (N_18464,N_17298,N_16960);
xnor U18465 (N_18465,N_16954,N_16439);
or U18466 (N_18466,N_16631,N_16820);
nand U18467 (N_18467,N_16936,N_16024);
xor U18468 (N_18468,N_17487,N_16740);
nor U18469 (N_18469,N_17568,N_16714);
nor U18470 (N_18470,N_17893,N_16689);
and U18471 (N_18471,N_17619,N_17390);
and U18472 (N_18472,N_17167,N_16460);
or U18473 (N_18473,N_16302,N_17000);
and U18474 (N_18474,N_17734,N_16497);
nor U18475 (N_18475,N_16201,N_17879);
xor U18476 (N_18476,N_17043,N_17605);
nor U18477 (N_18477,N_16442,N_17922);
or U18478 (N_18478,N_16836,N_17008);
or U18479 (N_18479,N_17394,N_17847);
or U18480 (N_18480,N_17814,N_17998);
xnor U18481 (N_18481,N_16941,N_17651);
and U18482 (N_18482,N_17404,N_16591);
and U18483 (N_18483,N_16555,N_17310);
or U18484 (N_18484,N_16506,N_16220);
xor U18485 (N_18485,N_17951,N_16231);
or U18486 (N_18486,N_17212,N_17790);
and U18487 (N_18487,N_17730,N_17284);
nand U18488 (N_18488,N_16758,N_16428);
xor U18489 (N_18489,N_16355,N_16958);
nand U18490 (N_18490,N_17413,N_16472);
nor U18491 (N_18491,N_17429,N_17339);
or U18492 (N_18492,N_16962,N_16724);
xor U18493 (N_18493,N_16483,N_16929);
nor U18494 (N_18494,N_17798,N_16978);
nor U18495 (N_18495,N_16315,N_17821);
xor U18496 (N_18496,N_16344,N_17640);
and U18497 (N_18497,N_16640,N_17978);
and U18498 (N_18498,N_17599,N_16984);
xnor U18499 (N_18499,N_17328,N_17196);
nand U18500 (N_18500,N_17114,N_16038);
xor U18501 (N_18501,N_16049,N_16626);
nor U18502 (N_18502,N_17346,N_16703);
nand U18503 (N_18503,N_17933,N_17591);
nand U18504 (N_18504,N_17614,N_17329);
and U18505 (N_18505,N_16637,N_17993);
nor U18506 (N_18506,N_17955,N_17875);
and U18507 (N_18507,N_17475,N_17428);
nand U18508 (N_18508,N_17215,N_16791);
nor U18509 (N_18509,N_17335,N_16814);
nand U18510 (N_18510,N_16707,N_16623);
nand U18511 (N_18511,N_16284,N_17296);
xor U18512 (N_18512,N_16078,N_17977);
or U18513 (N_18513,N_17321,N_17836);
nor U18514 (N_18514,N_16241,N_17486);
or U18515 (N_18515,N_17718,N_17772);
nand U18516 (N_18516,N_16650,N_16883);
or U18517 (N_18517,N_17024,N_16717);
nand U18518 (N_18518,N_16384,N_17662);
or U18519 (N_18519,N_16131,N_16014);
and U18520 (N_18520,N_17116,N_17137);
xnor U18521 (N_18521,N_16000,N_17513);
nand U18522 (N_18522,N_16425,N_16244);
nand U18523 (N_18523,N_16869,N_17430);
and U18524 (N_18524,N_16197,N_16026);
nand U18525 (N_18525,N_17457,N_16504);
and U18526 (N_18526,N_16608,N_17131);
nor U18527 (N_18527,N_16789,N_17817);
and U18528 (N_18528,N_16210,N_16949);
or U18529 (N_18529,N_16177,N_16964);
or U18530 (N_18530,N_17002,N_16566);
nor U18531 (N_18531,N_16554,N_17642);
xor U18532 (N_18532,N_16322,N_17557);
xnor U18533 (N_18533,N_16005,N_16427);
and U18534 (N_18534,N_16139,N_16535);
nand U18535 (N_18535,N_16597,N_16227);
xnor U18536 (N_18536,N_16044,N_16126);
xor U18537 (N_18537,N_16722,N_17886);
and U18538 (N_18538,N_16546,N_16551);
and U18539 (N_18539,N_16781,N_17304);
nor U18540 (N_18540,N_17060,N_17785);
xor U18541 (N_18541,N_16216,N_16194);
and U18542 (N_18542,N_17576,N_16002);
and U18543 (N_18543,N_16515,N_17233);
xor U18544 (N_18544,N_17677,N_16090);
nor U18545 (N_18545,N_16376,N_16828);
and U18546 (N_18546,N_17566,N_17050);
or U18547 (N_18547,N_16731,N_16136);
and U18548 (N_18548,N_17511,N_16728);
or U18549 (N_18549,N_16885,N_16777);
nand U18550 (N_18550,N_16547,N_16977);
nand U18551 (N_18551,N_17342,N_16516);
and U18552 (N_18552,N_16649,N_16396);
nand U18553 (N_18553,N_16761,N_17340);
and U18554 (N_18554,N_16742,N_17652);
and U18555 (N_18555,N_17283,N_16109);
or U18556 (N_18556,N_16464,N_16915);
and U18557 (N_18557,N_17503,N_16617);
xor U18558 (N_18558,N_16009,N_16587);
nand U18559 (N_18559,N_16939,N_16143);
and U18560 (N_18560,N_16390,N_17860);
and U18561 (N_18561,N_17650,N_16077);
xnor U18562 (N_18562,N_17510,N_17073);
and U18563 (N_18563,N_16356,N_16512);
xnor U18564 (N_18564,N_16950,N_17906);
xnor U18565 (N_18565,N_16304,N_17311);
nor U18566 (N_18566,N_16999,N_16552);
nor U18567 (N_18567,N_16723,N_17940);
and U18568 (N_18568,N_17900,N_16648);
or U18569 (N_18569,N_16070,N_16734);
nor U18570 (N_18570,N_16775,N_16392);
nand U18571 (N_18571,N_16412,N_17699);
or U18572 (N_18572,N_16961,N_17660);
nand U18573 (N_18573,N_16615,N_17052);
xnor U18574 (N_18574,N_17387,N_16981);
or U18575 (N_18575,N_17223,N_16701);
xnor U18576 (N_18576,N_16379,N_17529);
nor U18577 (N_18577,N_17805,N_16144);
nor U18578 (N_18578,N_17665,N_16467);
xnor U18579 (N_18579,N_16825,N_16917);
and U18580 (N_18580,N_16987,N_17515);
and U18581 (N_18581,N_17035,N_17425);
and U18582 (N_18582,N_16498,N_16128);
and U18583 (N_18583,N_16901,N_16992);
xnor U18584 (N_18584,N_16196,N_17189);
nor U18585 (N_18585,N_16574,N_17409);
and U18586 (N_18586,N_16990,N_16223);
or U18587 (N_18587,N_16667,N_16094);
nand U18588 (N_18588,N_16708,N_17140);
nand U18589 (N_18589,N_16691,N_17894);
xnor U18590 (N_18590,N_16594,N_17153);
nand U18591 (N_18591,N_17224,N_16348);
and U18592 (N_18592,N_16087,N_17231);
nor U18593 (N_18593,N_17631,N_17306);
or U18594 (N_18594,N_16413,N_17516);
and U18595 (N_18595,N_17220,N_16199);
and U18596 (N_18596,N_17987,N_17835);
and U18597 (N_18597,N_17348,N_17471);
or U18598 (N_18598,N_17001,N_17985);
and U18599 (N_18599,N_16931,N_17259);
and U18600 (N_18600,N_16573,N_16457);
or U18601 (N_18601,N_17820,N_16746);
nor U18602 (N_18602,N_17407,N_17601);
xnor U18603 (N_18603,N_16870,N_17982);
and U18604 (N_18604,N_16613,N_17120);
nor U18605 (N_18605,N_16230,N_16831);
or U18606 (N_18606,N_17251,N_17611);
xor U18607 (N_18607,N_17392,N_16853);
or U18608 (N_18608,N_16151,N_16518);
nand U18609 (N_18609,N_16612,N_17645);
nor U18610 (N_18610,N_17443,N_16320);
nor U18611 (N_18611,N_16218,N_17027);
or U18612 (N_18612,N_17199,N_16965);
nand U18613 (N_18613,N_17995,N_17313);
nor U18614 (N_18614,N_16670,N_16754);
and U18615 (N_18615,N_17228,N_16001);
nor U18616 (N_18616,N_17101,N_17585);
nand U18617 (N_18617,N_17398,N_17773);
nor U18618 (N_18618,N_16720,N_17213);
nand U18619 (N_18619,N_17533,N_16471);
nand U18620 (N_18620,N_16169,N_17508);
nor U18621 (N_18621,N_16068,N_16339);
and U18622 (N_18622,N_16247,N_16913);
nand U18623 (N_18623,N_17958,N_17765);
nor U18624 (N_18624,N_16432,N_16655);
or U18625 (N_18625,N_16778,N_16695);
xnor U18626 (N_18626,N_16970,N_16437);
and U18627 (N_18627,N_17930,N_17132);
or U18628 (N_18628,N_16895,N_17255);
or U18629 (N_18629,N_16309,N_16657);
nand U18630 (N_18630,N_17045,N_17289);
nor U18631 (N_18631,N_17883,N_17733);
nand U18632 (N_18632,N_17481,N_17603);
xnor U18633 (N_18633,N_17744,N_16274);
nor U18634 (N_18634,N_16400,N_17362);
or U18635 (N_18635,N_16548,N_17863);
nand U18636 (N_18636,N_16326,N_16676);
or U18637 (N_18637,N_16780,N_16146);
nand U18638 (N_18638,N_17361,N_17701);
xor U18639 (N_18639,N_16013,N_16907);
xnor U18640 (N_18640,N_16868,N_16837);
or U18641 (N_18641,N_17097,N_16167);
or U18642 (N_18642,N_16767,N_16618);
and U18643 (N_18643,N_17901,N_16129);
xnor U18644 (N_18644,N_16748,N_17956);
nand U18645 (N_18645,N_16861,N_17047);
nor U18646 (N_18646,N_17552,N_17831);
nand U18647 (N_18647,N_16688,N_17087);
and U18648 (N_18648,N_16367,N_17210);
nor U18649 (N_18649,N_17582,N_17033);
nand U18650 (N_18650,N_16927,N_16319);
nand U18651 (N_18651,N_17698,N_17022);
or U18652 (N_18652,N_16031,N_16368);
and U18653 (N_18653,N_16397,N_16296);
or U18654 (N_18654,N_16923,N_16347);
nand U18655 (N_18655,N_17076,N_17670);
xnor U18656 (N_18656,N_17615,N_17201);
nand U18657 (N_18657,N_17009,N_17947);
nor U18658 (N_18658,N_17011,N_17257);
xnor U18659 (N_18659,N_17053,N_17094);
nor U18660 (N_18660,N_16338,N_17846);
xnor U18661 (N_18661,N_17544,N_17439);
xor U18662 (N_18662,N_17161,N_16108);
nand U18663 (N_18663,N_16733,N_16369);
or U18664 (N_18664,N_17793,N_16403);
and U18665 (N_18665,N_16171,N_16456);
and U18666 (N_18666,N_17476,N_16106);
nor U18667 (N_18667,N_17268,N_17724);
xnor U18668 (N_18668,N_16114,N_16279);
nand U18669 (N_18669,N_17745,N_16829);
and U18670 (N_18670,N_17782,N_16673);
or U18671 (N_18671,N_16904,N_17708);
nor U18672 (N_18672,N_17800,N_17270);
and U18673 (N_18673,N_17163,N_17204);
nor U18674 (N_18674,N_17921,N_17345);
nor U18675 (N_18675,N_17397,N_16715);
and U18676 (N_18676,N_17125,N_16531);
and U18677 (N_18677,N_17825,N_16297);
nor U18678 (N_18678,N_17791,N_17133);
xor U18679 (N_18679,N_17227,N_17177);
or U18680 (N_18680,N_16147,N_17084);
nor U18681 (N_18681,N_17459,N_16776);
nand U18682 (N_18682,N_16660,N_16564);
and U18683 (N_18683,N_16273,N_17434);
nor U18684 (N_18684,N_16258,N_17244);
xor U18685 (N_18685,N_17709,N_16060);
nand U18686 (N_18686,N_17807,N_16142);
nand U18687 (N_18687,N_17657,N_17252);
nor U18688 (N_18688,N_17871,N_16891);
xor U18689 (N_18689,N_17216,N_16849);
xor U18690 (N_18690,N_17138,N_17550);
nand U18691 (N_18691,N_17134,N_17469);
nand U18692 (N_18692,N_17350,N_16250);
nand U18693 (N_18693,N_17191,N_16815);
nand U18694 (N_18694,N_17089,N_16232);
nor U18695 (N_18695,N_16262,N_16897);
or U18696 (N_18696,N_17593,N_16944);
xor U18697 (N_18697,N_17110,N_17617);
nor U18698 (N_18698,N_17355,N_17142);
and U18699 (N_18699,N_17751,N_16119);
nand U18700 (N_18700,N_16561,N_16545);
and U18701 (N_18701,N_17005,N_16772);
nor U18702 (N_18702,N_16839,N_17663);
nor U18703 (N_18703,N_17295,N_17600);
and U18704 (N_18704,N_16161,N_16305);
nand U18705 (N_18705,N_16235,N_17456);
nand U18706 (N_18706,N_17410,N_16481);
xor U18707 (N_18707,N_16190,N_17374);
xor U18708 (N_18708,N_16903,N_16374);
xor U18709 (N_18709,N_16180,N_16905);
or U18710 (N_18710,N_16168,N_17540);
or U18711 (N_18711,N_17484,N_17616);
or U18712 (N_18712,N_16682,N_16084);
xnor U18713 (N_18713,N_17412,N_16500);
and U18714 (N_18714,N_16809,N_17570);
nand U18715 (N_18715,N_17108,N_17325);
and U18716 (N_18716,N_17686,N_17182);
nor U18717 (N_18717,N_17057,N_17019);
nand U18718 (N_18718,N_17420,N_16787);
or U18719 (N_18719,N_17597,N_17674);
or U18720 (N_18720,N_16206,N_16115);
nand U18721 (N_18721,N_17872,N_16763);
and U18722 (N_18722,N_17587,N_16795);
nor U18723 (N_18723,N_17014,N_16806);
nor U18724 (N_18724,N_16043,N_16414);
or U18725 (N_18725,N_17722,N_17620);
or U18726 (N_18726,N_16745,N_17128);
or U18727 (N_18727,N_17267,N_17910);
and U18728 (N_18728,N_16871,N_17121);
nand U18729 (N_18729,N_17185,N_16912);
nor U18730 (N_18730,N_17039,N_17480);
and U18731 (N_18731,N_16195,N_17171);
and U18732 (N_18732,N_17888,N_17078);
nand U18733 (N_18733,N_16204,N_16630);
nand U18734 (N_18734,N_16217,N_17183);
nand U18735 (N_18735,N_17696,N_16864);
nand U18736 (N_18736,N_17852,N_17577);
nor U18737 (N_18737,N_17607,N_16585);
nand U18738 (N_18738,N_16911,N_17776);
and U18739 (N_18739,N_16041,N_16291);
xnor U18740 (N_18740,N_17692,N_16525);
and U18741 (N_18741,N_16986,N_17055);
nand U18742 (N_18742,N_17483,N_16528);
xor U18743 (N_18743,N_17647,N_17764);
xnor U18744 (N_18744,N_16539,N_16451);
and U18745 (N_18745,N_17432,N_17999);
nand U18746 (N_18746,N_16324,N_17314);
nor U18747 (N_18747,N_16641,N_16507);
or U18748 (N_18748,N_16162,N_17713);
or U18749 (N_18749,N_16867,N_16102);
xnor U18750 (N_18750,N_16894,N_17334);
xnor U18751 (N_18751,N_17913,N_16283);
nand U18752 (N_18752,N_16996,N_17217);
nor U18753 (N_18753,N_16066,N_16429);
or U18754 (N_18754,N_17575,N_17693);
xnor U18755 (N_18755,N_16533,N_17061);
and U18756 (N_18756,N_17152,N_16099);
nor U18757 (N_18757,N_17905,N_17924);
or U18758 (N_18758,N_16253,N_16219);
nor U18759 (N_18759,N_17525,N_17331);
xnor U18760 (N_18760,N_16316,N_17870);
nor U18761 (N_18761,N_17703,N_16010);
nor U18762 (N_18762,N_16127,N_16243);
or U18763 (N_18763,N_17315,N_17761);
xnor U18764 (N_18764,N_17559,N_17301);
and U18765 (N_18765,N_16215,N_17849);
nand U18766 (N_18766,N_17385,N_17162);
xor U18767 (N_18767,N_17365,N_16149);
xnor U18768 (N_18768,N_16713,N_16928);
nand U18769 (N_18769,N_16393,N_17661);
nand U18770 (N_18770,N_16569,N_16294);
and U18771 (N_18771,N_17135,N_17071);
or U18772 (N_18772,N_16794,N_17006);
nor U18773 (N_18773,N_17075,N_16750);
xor U18774 (N_18774,N_17934,N_17750);
nor U18775 (N_18775,N_16377,N_17273);
xnor U18776 (N_18776,N_16479,N_17155);
nor U18777 (N_18777,N_16718,N_17431);
or U18778 (N_18778,N_17399,N_17953);
nor U18779 (N_18779,N_16381,N_16303);
or U18780 (N_18780,N_17490,N_17810);
nand U18781 (N_18781,N_16150,N_17015);
nor U18782 (N_18782,N_16741,N_17232);
or U18783 (N_18783,N_17519,N_16449);
xnor U18784 (N_18784,N_17446,N_16160);
or U18785 (N_18785,N_17769,N_16277);
nor U18786 (N_18786,N_16266,N_17837);
xor U18787 (N_18787,N_16739,N_17815);
or U18788 (N_18788,N_17357,N_16175);
nand U18789 (N_18789,N_16395,N_17056);
and U18790 (N_18790,N_17498,N_17376);
or U18791 (N_18791,N_16997,N_16643);
nor U18792 (N_18792,N_17254,N_16123);
or U18793 (N_18793,N_16576,N_17945);
nor U18794 (N_18794,N_16351,N_17904);
nand U18795 (N_18795,N_17635,N_16406);
nand U18796 (N_18796,N_17707,N_16801);
xor U18797 (N_18797,N_17245,N_17406);
and U18798 (N_18798,N_16245,N_17623);
or U18799 (N_18799,N_17149,N_17194);
or U18800 (N_18800,N_17007,N_17450);
and U18801 (N_18801,N_16583,N_16159);
xor U18802 (N_18802,N_16018,N_17548);
or U18803 (N_18803,N_16567,N_17437);
or U18804 (N_18804,N_17606,N_17664);
or U18805 (N_18805,N_17344,N_16541);
and U18806 (N_18806,N_17523,N_16782);
nor U18807 (N_18807,N_16841,N_16030);
and U18808 (N_18808,N_17812,N_16300);
and U18809 (N_18809,N_16287,N_17711);
or U18810 (N_18810,N_17150,N_16234);
or U18811 (N_18811,N_16082,N_17580);
nand U18812 (N_18812,N_17489,N_17997);
nand U18813 (N_18813,N_16628,N_16121);
nand U18814 (N_18814,N_16743,N_16268);
and U18815 (N_18815,N_16067,N_17803);
and U18816 (N_18816,N_17375,N_17594);
xor U18817 (N_18817,N_17528,N_16387);
nor U18818 (N_18818,N_16702,N_17841);
or U18819 (N_18819,N_17096,N_16145);
nor U18820 (N_18820,N_16133,N_17838);
nand U18821 (N_18821,N_17083,N_16956);
nand U18822 (N_18822,N_16473,N_16830);
nand U18823 (N_18823,N_16019,N_17391);
nand U18824 (N_18824,N_16361,N_16415);
nor U18825 (N_18825,N_17458,N_16047);
and U18826 (N_18826,N_16773,N_17986);
xor U18827 (N_18827,N_17624,N_17578);
and U18828 (N_18828,N_16366,N_17639);
nor U18829 (N_18829,N_17041,N_17300);
nor U18830 (N_18830,N_16770,N_17170);
and U18831 (N_18831,N_17588,N_17208);
and U18832 (N_18832,N_16914,N_16443);
or U18833 (N_18833,N_16211,N_16039);
and U18834 (N_18834,N_16495,N_17551);
xnor U18835 (N_18835,N_17491,N_17971);
nor U18836 (N_18836,N_16332,N_16988);
and U18837 (N_18837,N_17868,N_17702);
and U18838 (N_18838,N_16571,N_17869);
and U18839 (N_18839,N_16966,N_16046);
nand U18840 (N_18840,N_17823,N_16967);
and U18841 (N_18841,N_17943,N_16638);
xor U18842 (N_18842,N_16053,N_16896);
xor U18843 (N_18843,N_17774,N_16910);
xnor U18844 (N_18844,N_17936,N_17775);
xor U18845 (N_18845,N_17731,N_16252);
nor U18846 (N_18846,N_16340,N_16938);
xor U18847 (N_18847,N_17418,N_16198);
and U18848 (N_18848,N_16577,N_17729);
and U18849 (N_18849,N_17949,N_16972);
nand U18850 (N_18850,N_17400,N_17386);
xor U18851 (N_18851,N_16382,N_17786);
nand U18852 (N_18852,N_17966,N_17819);
nor U18853 (N_18853,N_16301,N_16732);
xnor U18854 (N_18854,N_17916,N_17419);
xor U18855 (N_18855,N_17710,N_17264);
nor U18856 (N_18856,N_17030,N_16430);
or U18857 (N_18857,N_17679,N_16524);
or U18858 (N_18858,N_17202,N_17928);
and U18859 (N_18859,N_17123,N_16804);
xor U18860 (N_18860,N_17755,N_17545);
nand U18861 (N_18861,N_17680,N_17970);
xnor U18862 (N_18862,N_17178,N_17485);
nand U18863 (N_18863,N_17248,N_16092);
nand U18864 (N_18864,N_16404,N_17799);
nand U18865 (N_18865,N_17802,N_16499);
xnor U18866 (N_18866,N_17854,N_16824);
nand U18867 (N_18867,N_16762,N_16575);
and U18868 (N_18868,N_17527,N_17880);
nand U18869 (N_18869,N_17632,N_16402);
or U18870 (N_18870,N_16075,N_16726);
nor U18871 (N_18871,N_16584,N_16103);
nor U18872 (N_18872,N_17903,N_17553);
xor U18873 (N_18873,N_16380,N_16553);
xor U18874 (N_18874,N_17668,N_16462);
and U18875 (N_18875,N_17634,N_17347);
and U18876 (N_18876,N_16808,N_16816);
or U18877 (N_18877,N_17612,N_17794);
nand U18878 (N_18878,N_17732,N_17700);
nor U18879 (N_18879,N_17371,N_16519);
or U18880 (N_18880,N_17066,N_16858);
or U18881 (N_18881,N_16345,N_16505);
or U18882 (N_18882,N_16784,N_17260);
and U18883 (N_18883,N_17853,N_17797);
nor U18884 (N_18884,N_17671,N_17512);
xor U18885 (N_18885,N_16372,N_16325);
xor U18886 (N_18886,N_17172,N_16022);
nor U18887 (N_18887,N_17885,N_17655);
and U18888 (N_18888,N_17411,N_17946);
or U18889 (N_18889,N_16693,N_17783);
and U18890 (N_18890,N_17356,N_16448);
nor U18891 (N_18891,N_17641,N_17405);
nor U18892 (N_18892,N_17063,N_16979);
or U18893 (N_18893,N_16346,N_17322);
and U18894 (N_18894,N_16921,N_16900);
or U18895 (N_18895,N_17826,N_16671);
nand U18896 (N_18896,N_16459,N_16434);
nor U18897 (N_18897,N_17238,N_16224);
nor U18898 (N_18898,N_17240,N_16378);
and U18899 (N_18899,N_16800,N_17675);
nand U18900 (N_18900,N_16033,N_17865);
or U18901 (N_18901,N_16004,N_16208);
nand U18902 (N_18902,N_17130,N_16860);
nand U18903 (N_18903,N_16924,N_17195);
xnor U18904 (N_18904,N_16893,N_16755);
or U18905 (N_18905,N_17542,N_17737);
nor U18906 (N_18906,N_17332,N_17211);
nor U18907 (N_18907,N_16788,N_16521);
nor U18908 (N_18908,N_16299,N_17714);
and U18909 (N_18909,N_17105,N_16444);
nor U18910 (N_18910,N_16930,N_17474);
xnor U18911 (N_18911,N_16214,N_17058);
nand U18912 (N_18912,N_17792,N_17809);
nor U18913 (N_18913,N_17293,N_17263);
and U18914 (N_18914,N_16838,N_16173);
xnor U18915 (N_18915,N_17996,N_16330);
nor U18916 (N_18916,N_17359,N_17538);
or U18917 (N_18917,N_17965,N_16998);
and U18918 (N_18918,N_16735,N_17214);
and U18919 (N_18919,N_17942,N_17948);
xnor U18920 (N_18920,N_16729,N_16111);
or U18921 (N_18921,N_16365,N_17636);
and U18922 (N_18922,N_16482,N_16968);
nand U18923 (N_18923,N_16859,N_16934);
xnor U18924 (N_18924,N_16003,N_17558);
and U18925 (N_18925,N_16969,N_16706);
xnor U18926 (N_18926,N_17925,N_16166);
nor U18927 (N_18927,N_17895,N_16593);
and U18928 (N_18928,N_16665,N_17855);
xnor U18929 (N_18929,N_16100,N_16288);
nand U18930 (N_18930,N_17926,N_16373);
xnor U18931 (N_18931,N_17586,N_17333);
or U18932 (N_18932,N_17048,N_16465);
or U18933 (N_18933,N_17787,N_17590);
xor U18934 (N_18934,N_17148,N_16686);
xor U18935 (N_18935,N_17595,N_16088);
or U18936 (N_18936,N_16677,N_16812);
and U18937 (N_18937,N_16298,N_16203);
xor U18938 (N_18938,N_16534,N_16625);
or U18939 (N_18939,N_16580,N_16072);
or U18940 (N_18940,N_16409,N_17845);
and U18941 (N_18941,N_17274,N_17682);
or U18942 (N_18942,N_16933,N_16455);
nor U18943 (N_18943,N_17555,N_16331);
xnor U18944 (N_18944,N_17422,N_16435);
nand U18945 (N_18945,N_17796,N_17758);
nand U18946 (N_18946,N_16255,N_17249);
nor U18947 (N_18947,N_16012,N_16089);
nor U18948 (N_18948,N_17258,N_17687);
nand U18949 (N_18949,N_16269,N_16282);
nor U18950 (N_18950,N_17850,N_17088);
or U18951 (N_18951,N_16609,N_16259);
or U18952 (N_18952,N_16107,N_16447);
xnor U18953 (N_18953,N_17113,N_17779);
xnor U18954 (N_18954,N_16363,N_17757);
nor U18955 (N_18955,N_16918,N_16154);
nor U18956 (N_18956,N_17384,N_16614);
xor U18957 (N_18957,N_17351,N_17741);
or U18958 (N_18958,N_16737,N_17656);
nand U18959 (N_18959,N_17874,N_17827);
xnor U18960 (N_18960,N_17445,N_17271);
and U18961 (N_18961,N_17269,N_17261);
xor U18962 (N_18962,N_17025,N_17302);
nor U18963 (N_18963,N_16260,N_17507);
or U18964 (N_18964,N_17382,N_16774);
xor U18965 (N_18965,N_16276,N_16281);
nand U18966 (N_18966,N_16275,N_16261);
and U18967 (N_18967,N_17472,N_17889);
and U18968 (N_18968,N_17864,N_16556);
nor U18969 (N_18969,N_17143,N_17441);
and U18970 (N_18970,N_16620,N_16786);
or U18971 (N_18971,N_17416,N_17040);
or U18972 (N_18972,N_17074,N_17197);
nand U18973 (N_18973,N_16980,N_17229);
nor U18974 (N_18974,N_17832,N_17352);
nand U18975 (N_18975,N_16191,N_16876);
xnor U18976 (N_18976,N_17912,N_16818);
xor U18977 (N_18977,N_16032,N_17029);
nor U18978 (N_18978,N_17896,N_17504);
xnor U18979 (N_18979,N_16423,N_17462);
and U18980 (N_18980,N_16823,N_16769);
xnor U18981 (N_18981,N_17370,N_16538);
xor U18982 (N_18982,N_17898,N_16873);
xnor U18983 (N_18983,N_17746,N_16371);
and U18984 (N_18984,N_17169,N_16711);
xnor U18985 (N_18985,N_17408,N_17206);
nand U18986 (N_18986,N_16285,N_16008);
or U18987 (N_18987,N_16254,N_16023);
nor U18988 (N_18988,N_16420,N_16063);
and U18989 (N_18989,N_17049,N_16705);
nand U18990 (N_18990,N_17144,N_16061);
xor U18991 (N_18991,N_17299,N_17059);
and U18992 (N_18992,N_16721,N_17497);
nand U18993 (N_18993,N_17760,N_17690);
nand U18994 (N_18994,N_17381,N_16560);
or U18995 (N_18995,N_16233,N_16336);
nor U18996 (N_18996,N_17941,N_17188);
or U18997 (N_18997,N_17857,N_16798);
nand U18998 (N_18998,N_17054,N_16221);
nand U18999 (N_18999,N_16165,N_16629);
and U19000 (N_19000,N_16468,N_16201);
and U19001 (N_19001,N_17802,N_16145);
nor U19002 (N_19002,N_17689,N_16230);
and U19003 (N_19003,N_16480,N_16845);
nor U19004 (N_19004,N_16632,N_17969);
xnor U19005 (N_19005,N_16026,N_16224);
nor U19006 (N_19006,N_17338,N_17649);
or U19007 (N_19007,N_17251,N_16232);
xnor U19008 (N_19008,N_17029,N_16475);
nand U19009 (N_19009,N_17691,N_16966);
nand U19010 (N_19010,N_17256,N_17119);
and U19011 (N_19011,N_16061,N_17209);
nand U19012 (N_19012,N_16478,N_17866);
and U19013 (N_19013,N_17490,N_16039);
and U19014 (N_19014,N_17229,N_17734);
and U19015 (N_19015,N_16941,N_17147);
nand U19016 (N_19016,N_17738,N_17560);
nor U19017 (N_19017,N_16120,N_16924);
and U19018 (N_19018,N_16872,N_17966);
nor U19019 (N_19019,N_17352,N_17620);
nor U19020 (N_19020,N_17289,N_17414);
and U19021 (N_19021,N_16520,N_16908);
or U19022 (N_19022,N_17839,N_16084);
xnor U19023 (N_19023,N_16482,N_16534);
and U19024 (N_19024,N_16430,N_17244);
or U19025 (N_19025,N_16698,N_17587);
and U19026 (N_19026,N_17686,N_17133);
xor U19027 (N_19027,N_16236,N_17552);
and U19028 (N_19028,N_16279,N_17473);
or U19029 (N_19029,N_16541,N_16724);
nor U19030 (N_19030,N_17949,N_17484);
nor U19031 (N_19031,N_17514,N_17241);
nor U19032 (N_19032,N_17082,N_17617);
nor U19033 (N_19033,N_17023,N_17772);
and U19034 (N_19034,N_16195,N_16597);
xor U19035 (N_19035,N_16232,N_17849);
nor U19036 (N_19036,N_17599,N_17324);
or U19037 (N_19037,N_17207,N_17032);
nor U19038 (N_19038,N_17483,N_17491);
xor U19039 (N_19039,N_16585,N_17867);
or U19040 (N_19040,N_17879,N_16935);
and U19041 (N_19041,N_16893,N_17971);
nand U19042 (N_19042,N_17416,N_16389);
or U19043 (N_19043,N_17686,N_17015);
and U19044 (N_19044,N_16077,N_16094);
nand U19045 (N_19045,N_17127,N_16993);
nor U19046 (N_19046,N_16360,N_16898);
or U19047 (N_19047,N_17243,N_16547);
and U19048 (N_19048,N_17363,N_16496);
and U19049 (N_19049,N_16472,N_17135);
nand U19050 (N_19050,N_16324,N_16472);
nor U19051 (N_19051,N_16649,N_17438);
xor U19052 (N_19052,N_17030,N_17417);
or U19053 (N_19053,N_17456,N_16812);
and U19054 (N_19054,N_16399,N_17361);
and U19055 (N_19055,N_16410,N_17782);
nand U19056 (N_19056,N_17571,N_16306);
or U19057 (N_19057,N_17162,N_17882);
nor U19058 (N_19058,N_16314,N_17525);
and U19059 (N_19059,N_16526,N_17672);
nand U19060 (N_19060,N_16021,N_16600);
or U19061 (N_19061,N_17736,N_16724);
and U19062 (N_19062,N_17953,N_16546);
nand U19063 (N_19063,N_16865,N_17260);
xnor U19064 (N_19064,N_16394,N_17805);
xor U19065 (N_19065,N_17964,N_16474);
xnor U19066 (N_19066,N_17657,N_16024);
or U19067 (N_19067,N_16893,N_17141);
nor U19068 (N_19068,N_16979,N_16779);
or U19069 (N_19069,N_17237,N_17575);
xnor U19070 (N_19070,N_17649,N_16011);
and U19071 (N_19071,N_17757,N_16349);
nand U19072 (N_19072,N_17843,N_16799);
nor U19073 (N_19073,N_16283,N_17217);
nand U19074 (N_19074,N_16014,N_17342);
xnor U19075 (N_19075,N_16733,N_16940);
nor U19076 (N_19076,N_16904,N_16071);
xnor U19077 (N_19077,N_17022,N_17435);
nand U19078 (N_19078,N_16739,N_17157);
or U19079 (N_19079,N_17189,N_17672);
nor U19080 (N_19080,N_17787,N_16899);
xor U19081 (N_19081,N_17176,N_17121);
xnor U19082 (N_19082,N_17610,N_16554);
xor U19083 (N_19083,N_17504,N_16933);
nand U19084 (N_19084,N_16778,N_17226);
nor U19085 (N_19085,N_16139,N_16220);
and U19086 (N_19086,N_17407,N_16246);
xor U19087 (N_19087,N_16237,N_16624);
xnor U19088 (N_19088,N_17651,N_17390);
nor U19089 (N_19089,N_16178,N_17847);
nand U19090 (N_19090,N_17466,N_17622);
and U19091 (N_19091,N_16347,N_17802);
and U19092 (N_19092,N_16470,N_16031);
nor U19093 (N_19093,N_17048,N_17894);
nor U19094 (N_19094,N_16676,N_17724);
nor U19095 (N_19095,N_17921,N_17531);
or U19096 (N_19096,N_17053,N_17830);
xnor U19097 (N_19097,N_17489,N_16918);
and U19098 (N_19098,N_17683,N_17486);
and U19099 (N_19099,N_17806,N_16548);
xnor U19100 (N_19100,N_17015,N_17637);
nand U19101 (N_19101,N_17915,N_16069);
nor U19102 (N_19102,N_16616,N_17467);
nor U19103 (N_19103,N_16428,N_17191);
xnor U19104 (N_19104,N_16542,N_17941);
nand U19105 (N_19105,N_16561,N_17446);
xor U19106 (N_19106,N_17685,N_17974);
nand U19107 (N_19107,N_17806,N_16273);
and U19108 (N_19108,N_16485,N_17842);
xor U19109 (N_19109,N_17819,N_16500);
or U19110 (N_19110,N_17892,N_17964);
nor U19111 (N_19111,N_17712,N_16254);
xor U19112 (N_19112,N_16926,N_16019);
nor U19113 (N_19113,N_16864,N_17049);
nand U19114 (N_19114,N_17633,N_17475);
and U19115 (N_19115,N_16420,N_17550);
nand U19116 (N_19116,N_16253,N_17627);
nand U19117 (N_19117,N_17330,N_16647);
and U19118 (N_19118,N_16556,N_17432);
and U19119 (N_19119,N_17967,N_16458);
or U19120 (N_19120,N_16944,N_17362);
or U19121 (N_19121,N_16780,N_17126);
xor U19122 (N_19122,N_16989,N_17915);
nor U19123 (N_19123,N_16009,N_16241);
nor U19124 (N_19124,N_16606,N_17706);
nor U19125 (N_19125,N_17242,N_17499);
or U19126 (N_19126,N_16680,N_17018);
nand U19127 (N_19127,N_16927,N_17625);
nor U19128 (N_19128,N_16230,N_16439);
xnor U19129 (N_19129,N_17180,N_16191);
and U19130 (N_19130,N_16520,N_16229);
nand U19131 (N_19131,N_17490,N_16849);
nand U19132 (N_19132,N_16024,N_16506);
xor U19133 (N_19133,N_17628,N_17926);
or U19134 (N_19134,N_16579,N_16587);
and U19135 (N_19135,N_17876,N_16930);
nand U19136 (N_19136,N_16172,N_17098);
and U19137 (N_19137,N_16495,N_17654);
xnor U19138 (N_19138,N_17086,N_17000);
nand U19139 (N_19139,N_16984,N_17334);
nand U19140 (N_19140,N_16820,N_17713);
xnor U19141 (N_19141,N_17817,N_16673);
xnor U19142 (N_19142,N_17364,N_16196);
nand U19143 (N_19143,N_16960,N_17206);
nand U19144 (N_19144,N_17300,N_17657);
xor U19145 (N_19145,N_16879,N_16625);
and U19146 (N_19146,N_16284,N_17365);
xor U19147 (N_19147,N_16439,N_17421);
nand U19148 (N_19148,N_16690,N_16817);
or U19149 (N_19149,N_16894,N_17867);
or U19150 (N_19150,N_17488,N_16219);
and U19151 (N_19151,N_16878,N_16600);
nor U19152 (N_19152,N_17628,N_17760);
nor U19153 (N_19153,N_16121,N_17347);
xor U19154 (N_19154,N_16725,N_16165);
nor U19155 (N_19155,N_16877,N_16867);
and U19156 (N_19156,N_16949,N_17849);
or U19157 (N_19157,N_16906,N_16015);
or U19158 (N_19158,N_16337,N_17630);
xnor U19159 (N_19159,N_16722,N_16703);
or U19160 (N_19160,N_17176,N_17112);
or U19161 (N_19161,N_17717,N_16347);
nor U19162 (N_19162,N_17788,N_16776);
nor U19163 (N_19163,N_16226,N_17089);
nand U19164 (N_19164,N_17758,N_17723);
and U19165 (N_19165,N_17114,N_16801);
or U19166 (N_19166,N_17445,N_16808);
xor U19167 (N_19167,N_16078,N_17619);
xnor U19168 (N_19168,N_17275,N_16479);
and U19169 (N_19169,N_16476,N_17867);
and U19170 (N_19170,N_17874,N_17913);
nor U19171 (N_19171,N_17764,N_16395);
nor U19172 (N_19172,N_16208,N_17720);
xor U19173 (N_19173,N_16527,N_16416);
nand U19174 (N_19174,N_16369,N_17286);
and U19175 (N_19175,N_17330,N_16630);
nand U19176 (N_19176,N_16749,N_17626);
or U19177 (N_19177,N_16283,N_16988);
xor U19178 (N_19178,N_16543,N_17472);
nand U19179 (N_19179,N_17105,N_17632);
and U19180 (N_19180,N_16477,N_17969);
nand U19181 (N_19181,N_17400,N_17394);
nor U19182 (N_19182,N_17154,N_17537);
and U19183 (N_19183,N_16444,N_17545);
nor U19184 (N_19184,N_17615,N_16193);
nand U19185 (N_19185,N_17248,N_17800);
or U19186 (N_19186,N_17515,N_17334);
nor U19187 (N_19187,N_16936,N_17895);
nor U19188 (N_19188,N_17863,N_17557);
and U19189 (N_19189,N_16886,N_16169);
or U19190 (N_19190,N_16961,N_17236);
and U19191 (N_19191,N_16227,N_16941);
xnor U19192 (N_19192,N_17602,N_17716);
xor U19193 (N_19193,N_17671,N_17539);
or U19194 (N_19194,N_17340,N_16139);
nor U19195 (N_19195,N_16058,N_17565);
nand U19196 (N_19196,N_17206,N_16014);
or U19197 (N_19197,N_17066,N_17575);
or U19198 (N_19198,N_16804,N_17431);
nor U19199 (N_19199,N_17064,N_17528);
xnor U19200 (N_19200,N_17245,N_16939);
nor U19201 (N_19201,N_16837,N_16157);
xor U19202 (N_19202,N_17309,N_17679);
or U19203 (N_19203,N_16590,N_17381);
xor U19204 (N_19204,N_17007,N_17473);
nor U19205 (N_19205,N_17228,N_17132);
or U19206 (N_19206,N_16378,N_17364);
nor U19207 (N_19207,N_16430,N_16562);
and U19208 (N_19208,N_17783,N_17829);
nand U19209 (N_19209,N_17942,N_17093);
and U19210 (N_19210,N_17034,N_17227);
nor U19211 (N_19211,N_16538,N_16449);
nor U19212 (N_19212,N_17314,N_17317);
nand U19213 (N_19213,N_17663,N_17161);
and U19214 (N_19214,N_17267,N_17196);
nand U19215 (N_19215,N_16444,N_17241);
nor U19216 (N_19216,N_16502,N_17172);
nor U19217 (N_19217,N_16238,N_16773);
and U19218 (N_19218,N_16851,N_17228);
xnor U19219 (N_19219,N_16193,N_17469);
or U19220 (N_19220,N_17039,N_17988);
nand U19221 (N_19221,N_16442,N_16982);
and U19222 (N_19222,N_16933,N_16827);
or U19223 (N_19223,N_17585,N_16953);
or U19224 (N_19224,N_17080,N_17496);
nor U19225 (N_19225,N_17042,N_17100);
xnor U19226 (N_19226,N_16266,N_17036);
nor U19227 (N_19227,N_16884,N_17088);
nand U19228 (N_19228,N_17331,N_16470);
and U19229 (N_19229,N_17904,N_17304);
and U19230 (N_19230,N_16676,N_17142);
nand U19231 (N_19231,N_17774,N_16943);
nand U19232 (N_19232,N_16951,N_17571);
and U19233 (N_19233,N_16129,N_17223);
and U19234 (N_19234,N_17218,N_17318);
nand U19235 (N_19235,N_16828,N_17845);
nand U19236 (N_19236,N_16760,N_17007);
xnor U19237 (N_19237,N_16959,N_16540);
or U19238 (N_19238,N_16845,N_17201);
nor U19239 (N_19239,N_16801,N_17467);
xor U19240 (N_19240,N_17985,N_17796);
nor U19241 (N_19241,N_17281,N_16426);
and U19242 (N_19242,N_16500,N_17234);
and U19243 (N_19243,N_16926,N_17953);
and U19244 (N_19244,N_16977,N_16067);
nand U19245 (N_19245,N_17973,N_16504);
and U19246 (N_19246,N_17067,N_17043);
xnor U19247 (N_19247,N_16116,N_17187);
nand U19248 (N_19248,N_17946,N_17785);
and U19249 (N_19249,N_17304,N_17358);
or U19250 (N_19250,N_17319,N_16196);
nor U19251 (N_19251,N_16596,N_16093);
and U19252 (N_19252,N_17019,N_16559);
or U19253 (N_19253,N_17112,N_16831);
and U19254 (N_19254,N_17757,N_17519);
xor U19255 (N_19255,N_17473,N_17304);
or U19256 (N_19256,N_17541,N_16520);
xnor U19257 (N_19257,N_16799,N_16365);
or U19258 (N_19258,N_16568,N_17215);
xor U19259 (N_19259,N_17641,N_17976);
and U19260 (N_19260,N_17791,N_17053);
or U19261 (N_19261,N_16286,N_16761);
nor U19262 (N_19262,N_17897,N_16222);
nand U19263 (N_19263,N_17322,N_17931);
nor U19264 (N_19264,N_17591,N_17460);
or U19265 (N_19265,N_17919,N_16241);
or U19266 (N_19266,N_17393,N_17731);
or U19267 (N_19267,N_17699,N_17443);
nand U19268 (N_19268,N_17789,N_17537);
and U19269 (N_19269,N_17609,N_17754);
nor U19270 (N_19270,N_16778,N_16523);
nor U19271 (N_19271,N_17104,N_17318);
xor U19272 (N_19272,N_17468,N_17149);
nand U19273 (N_19273,N_16941,N_17982);
or U19274 (N_19274,N_16137,N_17699);
xnor U19275 (N_19275,N_17837,N_17325);
or U19276 (N_19276,N_17003,N_16375);
xnor U19277 (N_19277,N_16648,N_16738);
or U19278 (N_19278,N_17229,N_17808);
xnor U19279 (N_19279,N_17538,N_16792);
xor U19280 (N_19280,N_17943,N_16015);
nor U19281 (N_19281,N_16912,N_17198);
and U19282 (N_19282,N_16869,N_17136);
or U19283 (N_19283,N_16414,N_16371);
or U19284 (N_19284,N_16098,N_17285);
nor U19285 (N_19285,N_16217,N_16455);
xor U19286 (N_19286,N_17379,N_16144);
nor U19287 (N_19287,N_17517,N_16017);
or U19288 (N_19288,N_17258,N_16309);
nor U19289 (N_19289,N_16454,N_17671);
nand U19290 (N_19290,N_16528,N_16413);
nand U19291 (N_19291,N_17748,N_16876);
and U19292 (N_19292,N_16428,N_16821);
and U19293 (N_19293,N_17921,N_16285);
nor U19294 (N_19294,N_16386,N_16129);
and U19295 (N_19295,N_17135,N_16409);
and U19296 (N_19296,N_17011,N_17240);
xor U19297 (N_19297,N_17990,N_17570);
or U19298 (N_19298,N_16633,N_16276);
xor U19299 (N_19299,N_16622,N_17979);
nand U19300 (N_19300,N_16211,N_16122);
and U19301 (N_19301,N_16530,N_17966);
and U19302 (N_19302,N_17752,N_16319);
or U19303 (N_19303,N_17474,N_17072);
nor U19304 (N_19304,N_16350,N_17549);
or U19305 (N_19305,N_17803,N_17875);
xor U19306 (N_19306,N_16824,N_16881);
nand U19307 (N_19307,N_16199,N_17433);
nor U19308 (N_19308,N_17353,N_17568);
and U19309 (N_19309,N_16972,N_17865);
nand U19310 (N_19310,N_17920,N_17720);
nand U19311 (N_19311,N_16535,N_17429);
or U19312 (N_19312,N_16151,N_16866);
nand U19313 (N_19313,N_17470,N_17468);
or U19314 (N_19314,N_16365,N_17241);
xnor U19315 (N_19315,N_17431,N_16541);
or U19316 (N_19316,N_16073,N_17298);
nor U19317 (N_19317,N_16718,N_17365);
xor U19318 (N_19318,N_16196,N_17581);
xor U19319 (N_19319,N_17137,N_17633);
nor U19320 (N_19320,N_16114,N_16834);
nor U19321 (N_19321,N_16089,N_16990);
xor U19322 (N_19322,N_17972,N_17867);
xor U19323 (N_19323,N_17608,N_17427);
or U19324 (N_19324,N_17409,N_17746);
nor U19325 (N_19325,N_17194,N_17862);
or U19326 (N_19326,N_16813,N_16200);
and U19327 (N_19327,N_17332,N_17619);
and U19328 (N_19328,N_16963,N_17062);
and U19329 (N_19329,N_17608,N_17283);
nand U19330 (N_19330,N_17252,N_17411);
and U19331 (N_19331,N_16665,N_17359);
nand U19332 (N_19332,N_16113,N_17972);
or U19333 (N_19333,N_17552,N_17533);
or U19334 (N_19334,N_17600,N_17361);
and U19335 (N_19335,N_17985,N_17978);
or U19336 (N_19336,N_16656,N_17597);
and U19337 (N_19337,N_16528,N_16517);
and U19338 (N_19338,N_16912,N_17160);
nor U19339 (N_19339,N_16348,N_16346);
or U19340 (N_19340,N_17048,N_17366);
xnor U19341 (N_19341,N_17820,N_16332);
and U19342 (N_19342,N_16454,N_16020);
or U19343 (N_19343,N_16193,N_17913);
nor U19344 (N_19344,N_16162,N_17035);
nor U19345 (N_19345,N_16484,N_17025);
xor U19346 (N_19346,N_16963,N_16043);
and U19347 (N_19347,N_16554,N_17560);
xor U19348 (N_19348,N_16721,N_17638);
xor U19349 (N_19349,N_17217,N_17205);
or U19350 (N_19350,N_17763,N_16518);
xnor U19351 (N_19351,N_16387,N_17036);
nor U19352 (N_19352,N_16091,N_16088);
nor U19353 (N_19353,N_17550,N_17140);
or U19354 (N_19354,N_17708,N_16418);
nor U19355 (N_19355,N_16556,N_16526);
nor U19356 (N_19356,N_16579,N_16239);
nor U19357 (N_19357,N_17596,N_16231);
nand U19358 (N_19358,N_16415,N_16255);
nand U19359 (N_19359,N_17653,N_16869);
xor U19360 (N_19360,N_17950,N_16203);
or U19361 (N_19361,N_16304,N_16323);
and U19362 (N_19362,N_16708,N_16216);
nand U19363 (N_19363,N_16938,N_17774);
and U19364 (N_19364,N_17416,N_17418);
or U19365 (N_19365,N_17626,N_17657);
nand U19366 (N_19366,N_17236,N_16127);
nor U19367 (N_19367,N_17417,N_16270);
nor U19368 (N_19368,N_16378,N_16479);
or U19369 (N_19369,N_17675,N_16175);
nand U19370 (N_19370,N_17880,N_16356);
xor U19371 (N_19371,N_16154,N_17603);
or U19372 (N_19372,N_16602,N_16383);
xnor U19373 (N_19373,N_17855,N_16560);
nor U19374 (N_19374,N_17503,N_17322);
xnor U19375 (N_19375,N_16855,N_17483);
or U19376 (N_19376,N_16763,N_16043);
and U19377 (N_19377,N_17170,N_17749);
or U19378 (N_19378,N_17072,N_17297);
and U19379 (N_19379,N_17958,N_16761);
or U19380 (N_19380,N_16274,N_17739);
or U19381 (N_19381,N_16162,N_17604);
nand U19382 (N_19382,N_16300,N_16026);
xnor U19383 (N_19383,N_17098,N_17778);
xnor U19384 (N_19384,N_17041,N_17572);
nor U19385 (N_19385,N_17482,N_17604);
nand U19386 (N_19386,N_17587,N_16596);
nand U19387 (N_19387,N_16736,N_17441);
nand U19388 (N_19388,N_17237,N_16163);
xnor U19389 (N_19389,N_17271,N_16590);
xnor U19390 (N_19390,N_17945,N_17040);
or U19391 (N_19391,N_17066,N_17752);
nand U19392 (N_19392,N_16469,N_17969);
nor U19393 (N_19393,N_16300,N_16246);
xor U19394 (N_19394,N_16612,N_16402);
nor U19395 (N_19395,N_17854,N_16086);
and U19396 (N_19396,N_16261,N_17601);
nand U19397 (N_19397,N_16966,N_17187);
xor U19398 (N_19398,N_16483,N_17783);
nand U19399 (N_19399,N_16597,N_16053);
xor U19400 (N_19400,N_16339,N_16713);
or U19401 (N_19401,N_16040,N_16457);
or U19402 (N_19402,N_16996,N_16997);
xnor U19403 (N_19403,N_17788,N_17933);
nor U19404 (N_19404,N_17740,N_16974);
xor U19405 (N_19405,N_16960,N_16313);
nand U19406 (N_19406,N_17258,N_16515);
xnor U19407 (N_19407,N_16146,N_16282);
nor U19408 (N_19408,N_16887,N_17208);
xnor U19409 (N_19409,N_16511,N_16036);
xnor U19410 (N_19410,N_16829,N_16081);
and U19411 (N_19411,N_17607,N_17486);
xnor U19412 (N_19412,N_16598,N_16922);
or U19413 (N_19413,N_17025,N_17326);
or U19414 (N_19414,N_16837,N_16305);
xor U19415 (N_19415,N_17211,N_16888);
or U19416 (N_19416,N_17071,N_17570);
or U19417 (N_19417,N_17607,N_16754);
xor U19418 (N_19418,N_16341,N_17737);
xnor U19419 (N_19419,N_17872,N_17294);
and U19420 (N_19420,N_17917,N_17447);
and U19421 (N_19421,N_16751,N_16976);
nor U19422 (N_19422,N_16319,N_17546);
or U19423 (N_19423,N_17566,N_17325);
and U19424 (N_19424,N_16706,N_17418);
and U19425 (N_19425,N_16257,N_17071);
xnor U19426 (N_19426,N_17178,N_17936);
or U19427 (N_19427,N_16015,N_16980);
nor U19428 (N_19428,N_16167,N_16703);
and U19429 (N_19429,N_17861,N_17918);
xnor U19430 (N_19430,N_17833,N_17913);
or U19431 (N_19431,N_16186,N_16221);
and U19432 (N_19432,N_16774,N_17015);
or U19433 (N_19433,N_16385,N_17211);
nor U19434 (N_19434,N_16040,N_17459);
nor U19435 (N_19435,N_17465,N_16668);
and U19436 (N_19436,N_17861,N_17547);
xnor U19437 (N_19437,N_16755,N_16433);
xor U19438 (N_19438,N_17306,N_16171);
or U19439 (N_19439,N_17802,N_17751);
or U19440 (N_19440,N_17207,N_16470);
xor U19441 (N_19441,N_17194,N_17711);
xor U19442 (N_19442,N_16680,N_17240);
nand U19443 (N_19443,N_17426,N_16034);
xor U19444 (N_19444,N_17474,N_17141);
and U19445 (N_19445,N_16767,N_16270);
and U19446 (N_19446,N_16904,N_16321);
nand U19447 (N_19447,N_16134,N_17537);
or U19448 (N_19448,N_16720,N_16515);
and U19449 (N_19449,N_16321,N_16540);
nor U19450 (N_19450,N_16909,N_17877);
xor U19451 (N_19451,N_16391,N_16239);
nand U19452 (N_19452,N_16841,N_17339);
nand U19453 (N_19453,N_17779,N_17316);
nand U19454 (N_19454,N_16052,N_16112);
and U19455 (N_19455,N_16997,N_17121);
nor U19456 (N_19456,N_17122,N_17339);
nor U19457 (N_19457,N_16993,N_17999);
or U19458 (N_19458,N_16195,N_16665);
or U19459 (N_19459,N_16484,N_17788);
or U19460 (N_19460,N_16374,N_16682);
nand U19461 (N_19461,N_17780,N_17465);
and U19462 (N_19462,N_17254,N_16204);
xnor U19463 (N_19463,N_17951,N_17675);
and U19464 (N_19464,N_16192,N_16821);
nor U19465 (N_19465,N_16470,N_16772);
nor U19466 (N_19466,N_16132,N_16554);
or U19467 (N_19467,N_16166,N_17742);
and U19468 (N_19468,N_17198,N_17337);
or U19469 (N_19469,N_17019,N_16421);
nand U19470 (N_19470,N_17444,N_16976);
and U19471 (N_19471,N_16201,N_17450);
xnor U19472 (N_19472,N_16315,N_17358);
and U19473 (N_19473,N_17443,N_17821);
nand U19474 (N_19474,N_17047,N_16036);
and U19475 (N_19475,N_17057,N_17592);
and U19476 (N_19476,N_16662,N_17421);
xnor U19477 (N_19477,N_16627,N_16746);
and U19478 (N_19478,N_17938,N_16037);
xor U19479 (N_19479,N_17693,N_16025);
nor U19480 (N_19480,N_17040,N_17171);
xnor U19481 (N_19481,N_17706,N_17041);
and U19482 (N_19482,N_17763,N_16641);
and U19483 (N_19483,N_17152,N_17485);
nor U19484 (N_19484,N_16649,N_16228);
xor U19485 (N_19485,N_16692,N_17650);
and U19486 (N_19486,N_17305,N_17411);
xnor U19487 (N_19487,N_17538,N_17366);
or U19488 (N_19488,N_17646,N_16116);
and U19489 (N_19489,N_17407,N_16085);
or U19490 (N_19490,N_16348,N_16400);
or U19491 (N_19491,N_17470,N_17191);
and U19492 (N_19492,N_17618,N_16646);
or U19493 (N_19493,N_16236,N_16790);
xnor U19494 (N_19494,N_16802,N_16176);
and U19495 (N_19495,N_16357,N_17747);
nor U19496 (N_19496,N_16310,N_16694);
or U19497 (N_19497,N_17976,N_17610);
xnor U19498 (N_19498,N_17472,N_17482);
xnor U19499 (N_19499,N_16429,N_17595);
or U19500 (N_19500,N_17847,N_16144);
nand U19501 (N_19501,N_17444,N_16913);
or U19502 (N_19502,N_17380,N_16882);
nor U19503 (N_19503,N_16871,N_17034);
nor U19504 (N_19504,N_16047,N_17214);
nand U19505 (N_19505,N_16588,N_16428);
nor U19506 (N_19506,N_16962,N_16839);
or U19507 (N_19507,N_16231,N_17277);
nand U19508 (N_19508,N_17825,N_17739);
xor U19509 (N_19509,N_17131,N_16544);
nand U19510 (N_19510,N_16658,N_17234);
nand U19511 (N_19511,N_17947,N_16663);
nor U19512 (N_19512,N_16277,N_17408);
xor U19513 (N_19513,N_17353,N_17003);
or U19514 (N_19514,N_17213,N_17063);
or U19515 (N_19515,N_16011,N_16422);
nand U19516 (N_19516,N_17749,N_16969);
and U19517 (N_19517,N_16046,N_16073);
xnor U19518 (N_19518,N_17397,N_16246);
xnor U19519 (N_19519,N_17691,N_17179);
and U19520 (N_19520,N_16598,N_17248);
and U19521 (N_19521,N_17565,N_16561);
nor U19522 (N_19522,N_16037,N_17149);
xor U19523 (N_19523,N_16637,N_17767);
or U19524 (N_19524,N_17525,N_17730);
nand U19525 (N_19525,N_17837,N_17105);
or U19526 (N_19526,N_17404,N_17342);
xor U19527 (N_19527,N_17023,N_16062);
or U19528 (N_19528,N_16309,N_16628);
or U19529 (N_19529,N_17830,N_17162);
nor U19530 (N_19530,N_16504,N_16709);
or U19531 (N_19531,N_16516,N_16540);
and U19532 (N_19532,N_17713,N_17164);
nand U19533 (N_19533,N_16500,N_16738);
or U19534 (N_19534,N_17273,N_17002);
xor U19535 (N_19535,N_16550,N_17973);
and U19536 (N_19536,N_16809,N_17937);
and U19537 (N_19537,N_17507,N_17729);
and U19538 (N_19538,N_17880,N_17006);
or U19539 (N_19539,N_16428,N_17532);
xnor U19540 (N_19540,N_17747,N_16744);
nor U19541 (N_19541,N_16305,N_16375);
nor U19542 (N_19542,N_16846,N_16848);
nand U19543 (N_19543,N_16382,N_16223);
nand U19544 (N_19544,N_16023,N_16770);
xnor U19545 (N_19545,N_17604,N_17980);
or U19546 (N_19546,N_16811,N_16776);
nor U19547 (N_19547,N_16412,N_16530);
xnor U19548 (N_19548,N_17123,N_16113);
nand U19549 (N_19549,N_16052,N_16626);
xnor U19550 (N_19550,N_16672,N_17461);
or U19551 (N_19551,N_16644,N_16788);
nand U19552 (N_19552,N_16264,N_16835);
and U19553 (N_19553,N_16677,N_17680);
or U19554 (N_19554,N_17073,N_16313);
xnor U19555 (N_19555,N_17871,N_17855);
xnor U19556 (N_19556,N_16660,N_16850);
or U19557 (N_19557,N_17708,N_16423);
xor U19558 (N_19558,N_16473,N_17642);
xnor U19559 (N_19559,N_17572,N_17052);
and U19560 (N_19560,N_16851,N_17342);
nand U19561 (N_19561,N_16839,N_16657);
and U19562 (N_19562,N_16028,N_17524);
and U19563 (N_19563,N_17395,N_16913);
and U19564 (N_19564,N_17506,N_17216);
nand U19565 (N_19565,N_17497,N_16967);
xor U19566 (N_19566,N_17632,N_16268);
and U19567 (N_19567,N_17585,N_16199);
or U19568 (N_19568,N_16308,N_16850);
nor U19569 (N_19569,N_17794,N_17390);
or U19570 (N_19570,N_16419,N_17409);
and U19571 (N_19571,N_17535,N_17974);
nand U19572 (N_19572,N_16375,N_17614);
nand U19573 (N_19573,N_17348,N_17332);
or U19574 (N_19574,N_17528,N_17029);
xor U19575 (N_19575,N_16363,N_16695);
or U19576 (N_19576,N_17261,N_17192);
and U19577 (N_19577,N_17137,N_17713);
or U19578 (N_19578,N_17108,N_17148);
nand U19579 (N_19579,N_17343,N_17619);
nor U19580 (N_19580,N_16388,N_16328);
nand U19581 (N_19581,N_17164,N_17252);
or U19582 (N_19582,N_17755,N_17895);
xnor U19583 (N_19583,N_16239,N_17701);
and U19584 (N_19584,N_17484,N_16664);
nand U19585 (N_19585,N_16687,N_17573);
nor U19586 (N_19586,N_16726,N_16667);
and U19587 (N_19587,N_17955,N_16788);
nand U19588 (N_19588,N_16603,N_16229);
xor U19589 (N_19589,N_17463,N_16981);
xnor U19590 (N_19590,N_17931,N_16889);
nand U19591 (N_19591,N_17903,N_16367);
nand U19592 (N_19592,N_16107,N_16891);
nand U19593 (N_19593,N_17753,N_17890);
or U19594 (N_19594,N_17357,N_17350);
and U19595 (N_19595,N_17218,N_17407);
or U19596 (N_19596,N_16276,N_17159);
or U19597 (N_19597,N_16656,N_16500);
or U19598 (N_19598,N_16581,N_17859);
xor U19599 (N_19599,N_17959,N_17819);
xor U19600 (N_19600,N_16033,N_16119);
nand U19601 (N_19601,N_17959,N_17856);
nor U19602 (N_19602,N_16417,N_17140);
nor U19603 (N_19603,N_17436,N_17939);
xnor U19604 (N_19604,N_17528,N_17530);
and U19605 (N_19605,N_16928,N_16730);
nor U19606 (N_19606,N_16595,N_17713);
nor U19607 (N_19607,N_17864,N_17166);
nor U19608 (N_19608,N_17894,N_17018);
xor U19609 (N_19609,N_17312,N_17785);
and U19610 (N_19610,N_17956,N_16812);
nor U19611 (N_19611,N_17888,N_16459);
nand U19612 (N_19612,N_16044,N_16611);
xor U19613 (N_19613,N_16316,N_17530);
xnor U19614 (N_19614,N_17495,N_17768);
or U19615 (N_19615,N_17158,N_17977);
nand U19616 (N_19616,N_17595,N_16933);
nand U19617 (N_19617,N_17911,N_17647);
nand U19618 (N_19618,N_16764,N_17197);
nand U19619 (N_19619,N_17817,N_17736);
nor U19620 (N_19620,N_16560,N_17634);
and U19621 (N_19621,N_16615,N_16841);
nand U19622 (N_19622,N_17707,N_16152);
or U19623 (N_19623,N_16938,N_16941);
xor U19624 (N_19624,N_17236,N_17505);
nor U19625 (N_19625,N_16646,N_17430);
nor U19626 (N_19626,N_16529,N_17460);
xor U19627 (N_19627,N_16795,N_16847);
xnor U19628 (N_19628,N_16143,N_16177);
nand U19629 (N_19629,N_16690,N_16501);
xnor U19630 (N_19630,N_16292,N_16945);
or U19631 (N_19631,N_16816,N_17146);
or U19632 (N_19632,N_16239,N_16939);
nor U19633 (N_19633,N_16473,N_16153);
and U19634 (N_19634,N_16130,N_16878);
nand U19635 (N_19635,N_16501,N_16071);
nand U19636 (N_19636,N_16710,N_16683);
nor U19637 (N_19637,N_16985,N_17269);
or U19638 (N_19638,N_17953,N_16868);
nor U19639 (N_19639,N_17800,N_17000);
nor U19640 (N_19640,N_16251,N_17830);
nand U19641 (N_19641,N_16121,N_17736);
nor U19642 (N_19642,N_17617,N_17481);
nor U19643 (N_19643,N_16383,N_17481);
xor U19644 (N_19644,N_17263,N_17834);
and U19645 (N_19645,N_17925,N_17401);
nor U19646 (N_19646,N_16281,N_16348);
nand U19647 (N_19647,N_16663,N_16909);
xor U19648 (N_19648,N_17382,N_17682);
and U19649 (N_19649,N_17199,N_16586);
xor U19650 (N_19650,N_16569,N_16564);
xor U19651 (N_19651,N_17201,N_17721);
and U19652 (N_19652,N_17984,N_17591);
nand U19653 (N_19653,N_17872,N_17513);
xnor U19654 (N_19654,N_16460,N_17315);
or U19655 (N_19655,N_17539,N_16751);
or U19656 (N_19656,N_17373,N_17355);
nor U19657 (N_19657,N_16019,N_16436);
nor U19658 (N_19658,N_17368,N_17096);
nand U19659 (N_19659,N_17714,N_17992);
and U19660 (N_19660,N_16008,N_17559);
and U19661 (N_19661,N_16221,N_17699);
nand U19662 (N_19662,N_17462,N_16401);
nand U19663 (N_19663,N_16879,N_16716);
or U19664 (N_19664,N_17652,N_17982);
and U19665 (N_19665,N_17737,N_17832);
and U19666 (N_19666,N_17414,N_16845);
nand U19667 (N_19667,N_16959,N_17798);
nand U19668 (N_19668,N_17975,N_17250);
nand U19669 (N_19669,N_17474,N_17235);
and U19670 (N_19670,N_17919,N_17149);
or U19671 (N_19671,N_17947,N_16174);
and U19672 (N_19672,N_16667,N_16093);
nand U19673 (N_19673,N_16992,N_17585);
nand U19674 (N_19674,N_17358,N_16889);
and U19675 (N_19675,N_16639,N_17497);
xor U19676 (N_19676,N_16948,N_16980);
nand U19677 (N_19677,N_17558,N_17357);
nor U19678 (N_19678,N_16463,N_17458);
or U19679 (N_19679,N_17426,N_17191);
xnor U19680 (N_19680,N_16138,N_16349);
xor U19681 (N_19681,N_17759,N_17103);
xor U19682 (N_19682,N_16761,N_17567);
or U19683 (N_19683,N_17518,N_17529);
nand U19684 (N_19684,N_16577,N_17521);
and U19685 (N_19685,N_16570,N_16056);
nand U19686 (N_19686,N_16286,N_16369);
and U19687 (N_19687,N_16443,N_17934);
and U19688 (N_19688,N_16368,N_17876);
and U19689 (N_19689,N_17794,N_17821);
and U19690 (N_19690,N_17553,N_16946);
xnor U19691 (N_19691,N_16133,N_16841);
nand U19692 (N_19692,N_16329,N_17609);
and U19693 (N_19693,N_16782,N_16384);
nand U19694 (N_19694,N_17612,N_16422);
nor U19695 (N_19695,N_17515,N_17705);
or U19696 (N_19696,N_16798,N_17813);
nand U19697 (N_19697,N_17440,N_16194);
nand U19698 (N_19698,N_17504,N_17201);
and U19699 (N_19699,N_17615,N_17761);
and U19700 (N_19700,N_17352,N_17781);
xnor U19701 (N_19701,N_16286,N_17004);
nor U19702 (N_19702,N_17497,N_16485);
nor U19703 (N_19703,N_17606,N_16969);
nor U19704 (N_19704,N_16759,N_17797);
xor U19705 (N_19705,N_16408,N_17081);
nor U19706 (N_19706,N_17006,N_16298);
and U19707 (N_19707,N_17237,N_16279);
nand U19708 (N_19708,N_16315,N_16399);
nor U19709 (N_19709,N_17890,N_17387);
and U19710 (N_19710,N_16211,N_17270);
nor U19711 (N_19711,N_17392,N_16128);
and U19712 (N_19712,N_17168,N_16107);
or U19713 (N_19713,N_16657,N_17762);
nor U19714 (N_19714,N_17810,N_16737);
or U19715 (N_19715,N_16734,N_16991);
xnor U19716 (N_19716,N_17920,N_16173);
nand U19717 (N_19717,N_16825,N_16813);
or U19718 (N_19718,N_17355,N_17622);
nor U19719 (N_19719,N_16415,N_16822);
and U19720 (N_19720,N_16348,N_16300);
nor U19721 (N_19721,N_16884,N_17385);
nand U19722 (N_19722,N_17738,N_17880);
and U19723 (N_19723,N_16181,N_17845);
and U19724 (N_19724,N_17257,N_16211);
nor U19725 (N_19725,N_17510,N_17226);
nor U19726 (N_19726,N_17820,N_16408);
or U19727 (N_19727,N_17964,N_16975);
and U19728 (N_19728,N_17794,N_17871);
nor U19729 (N_19729,N_16279,N_16614);
and U19730 (N_19730,N_17762,N_16278);
xor U19731 (N_19731,N_17434,N_16783);
and U19732 (N_19732,N_17436,N_16422);
or U19733 (N_19733,N_17792,N_17320);
nand U19734 (N_19734,N_16302,N_17607);
and U19735 (N_19735,N_16915,N_16230);
or U19736 (N_19736,N_17799,N_17902);
nand U19737 (N_19737,N_17742,N_17883);
or U19738 (N_19738,N_17718,N_17849);
nor U19739 (N_19739,N_16678,N_17610);
nand U19740 (N_19740,N_17397,N_17294);
and U19741 (N_19741,N_17938,N_17153);
nand U19742 (N_19742,N_16420,N_17206);
nand U19743 (N_19743,N_17857,N_17203);
and U19744 (N_19744,N_17512,N_16448);
nand U19745 (N_19745,N_16471,N_16938);
nand U19746 (N_19746,N_16863,N_17375);
nand U19747 (N_19747,N_17509,N_17504);
xnor U19748 (N_19748,N_17688,N_17285);
nand U19749 (N_19749,N_17589,N_16578);
nand U19750 (N_19750,N_16636,N_16294);
xor U19751 (N_19751,N_17936,N_16231);
nor U19752 (N_19752,N_17027,N_16722);
nand U19753 (N_19753,N_16082,N_16713);
nor U19754 (N_19754,N_17380,N_16251);
and U19755 (N_19755,N_16903,N_16695);
or U19756 (N_19756,N_16982,N_16685);
and U19757 (N_19757,N_16270,N_16942);
xor U19758 (N_19758,N_16408,N_17059);
and U19759 (N_19759,N_16130,N_16067);
nor U19760 (N_19760,N_17924,N_17373);
or U19761 (N_19761,N_17184,N_17036);
nand U19762 (N_19762,N_16361,N_16952);
and U19763 (N_19763,N_17965,N_16422);
or U19764 (N_19764,N_17283,N_17352);
and U19765 (N_19765,N_17440,N_17868);
nor U19766 (N_19766,N_16223,N_16662);
nor U19767 (N_19767,N_17754,N_17108);
nor U19768 (N_19768,N_16490,N_16423);
nor U19769 (N_19769,N_16860,N_16203);
nand U19770 (N_19770,N_16716,N_16020);
or U19771 (N_19771,N_16888,N_17944);
nand U19772 (N_19772,N_16936,N_16901);
xnor U19773 (N_19773,N_16007,N_16832);
nand U19774 (N_19774,N_16246,N_17343);
nand U19775 (N_19775,N_17235,N_16335);
nand U19776 (N_19776,N_17438,N_16977);
or U19777 (N_19777,N_17624,N_17436);
and U19778 (N_19778,N_17194,N_16370);
and U19779 (N_19779,N_16457,N_16135);
and U19780 (N_19780,N_16969,N_16676);
nand U19781 (N_19781,N_16269,N_16486);
xnor U19782 (N_19782,N_16461,N_16066);
nand U19783 (N_19783,N_17822,N_16829);
xnor U19784 (N_19784,N_17674,N_17315);
and U19785 (N_19785,N_17995,N_17336);
nor U19786 (N_19786,N_16993,N_17261);
nor U19787 (N_19787,N_16518,N_16788);
or U19788 (N_19788,N_16322,N_16264);
or U19789 (N_19789,N_17987,N_17705);
or U19790 (N_19790,N_16740,N_17501);
xnor U19791 (N_19791,N_17419,N_17094);
xor U19792 (N_19792,N_16165,N_17256);
nand U19793 (N_19793,N_16124,N_17347);
and U19794 (N_19794,N_17693,N_17994);
xnor U19795 (N_19795,N_17679,N_16636);
xor U19796 (N_19796,N_17351,N_17772);
nand U19797 (N_19797,N_17663,N_17670);
nand U19798 (N_19798,N_16566,N_16850);
nand U19799 (N_19799,N_17340,N_16788);
and U19800 (N_19800,N_17517,N_16418);
nor U19801 (N_19801,N_17292,N_16751);
or U19802 (N_19802,N_17640,N_16463);
or U19803 (N_19803,N_16161,N_16279);
and U19804 (N_19804,N_17620,N_17306);
nand U19805 (N_19805,N_17664,N_17317);
and U19806 (N_19806,N_17362,N_17506);
nor U19807 (N_19807,N_16866,N_17011);
nor U19808 (N_19808,N_17616,N_17124);
and U19809 (N_19809,N_16674,N_17119);
nand U19810 (N_19810,N_16925,N_17524);
nand U19811 (N_19811,N_17227,N_16053);
nor U19812 (N_19812,N_17903,N_17023);
nor U19813 (N_19813,N_16649,N_17235);
xor U19814 (N_19814,N_16829,N_17362);
nand U19815 (N_19815,N_16613,N_17606);
nand U19816 (N_19816,N_16029,N_17120);
xor U19817 (N_19817,N_16254,N_16847);
nor U19818 (N_19818,N_16372,N_17139);
nor U19819 (N_19819,N_17926,N_16121);
nor U19820 (N_19820,N_17298,N_16473);
nor U19821 (N_19821,N_16468,N_17672);
or U19822 (N_19822,N_16040,N_17920);
nand U19823 (N_19823,N_16061,N_17828);
nand U19824 (N_19824,N_16266,N_17841);
or U19825 (N_19825,N_16735,N_17338);
nand U19826 (N_19826,N_16583,N_16783);
and U19827 (N_19827,N_16354,N_16308);
xor U19828 (N_19828,N_17050,N_16388);
xor U19829 (N_19829,N_17936,N_17748);
nand U19830 (N_19830,N_17456,N_16727);
or U19831 (N_19831,N_16906,N_17267);
nand U19832 (N_19832,N_16983,N_16266);
nand U19833 (N_19833,N_16716,N_17500);
nand U19834 (N_19834,N_17510,N_17694);
and U19835 (N_19835,N_16935,N_17392);
xnor U19836 (N_19836,N_17159,N_16183);
nor U19837 (N_19837,N_17531,N_17847);
nor U19838 (N_19838,N_17026,N_17181);
nand U19839 (N_19839,N_17239,N_17707);
nor U19840 (N_19840,N_17903,N_16599);
nor U19841 (N_19841,N_17726,N_17572);
and U19842 (N_19842,N_17973,N_17459);
or U19843 (N_19843,N_16422,N_17523);
xnor U19844 (N_19844,N_16910,N_16859);
and U19845 (N_19845,N_16435,N_16114);
xnor U19846 (N_19846,N_16099,N_16326);
and U19847 (N_19847,N_16607,N_16394);
and U19848 (N_19848,N_16317,N_16851);
nand U19849 (N_19849,N_16520,N_16349);
and U19850 (N_19850,N_17948,N_17292);
nand U19851 (N_19851,N_17680,N_16949);
nand U19852 (N_19852,N_17108,N_16906);
nand U19853 (N_19853,N_16205,N_17109);
nand U19854 (N_19854,N_17892,N_16250);
and U19855 (N_19855,N_17110,N_16574);
xnor U19856 (N_19856,N_16640,N_17396);
xnor U19857 (N_19857,N_17692,N_17190);
nor U19858 (N_19858,N_16364,N_16719);
nor U19859 (N_19859,N_17071,N_17567);
nor U19860 (N_19860,N_17373,N_17088);
xor U19861 (N_19861,N_16342,N_17607);
and U19862 (N_19862,N_16502,N_17863);
nor U19863 (N_19863,N_16850,N_16588);
or U19864 (N_19864,N_17786,N_17147);
nand U19865 (N_19865,N_16796,N_16755);
or U19866 (N_19866,N_17740,N_16340);
xnor U19867 (N_19867,N_16201,N_16517);
nand U19868 (N_19868,N_17039,N_17416);
nand U19869 (N_19869,N_17676,N_16110);
xnor U19870 (N_19870,N_16468,N_16989);
nor U19871 (N_19871,N_16678,N_17689);
nand U19872 (N_19872,N_16400,N_16299);
or U19873 (N_19873,N_17047,N_16745);
nor U19874 (N_19874,N_16605,N_17124);
nand U19875 (N_19875,N_17685,N_16366);
xnor U19876 (N_19876,N_16753,N_17307);
xnor U19877 (N_19877,N_16720,N_16438);
nand U19878 (N_19878,N_16387,N_16156);
xor U19879 (N_19879,N_17276,N_16111);
xor U19880 (N_19880,N_17583,N_17325);
nor U19881 (N_19881,N_16494,N_17205);
nor U19882 (N_19882,N_16765,N_17700);
nor U19883 (N_19883,N_16851,N_16670);
or U19884 (N_19884,N_16605,N_16733);
nor U19885 (N_19885,N_16492,N_17609);
xor U19886 (N_19886,N_16252,N_16664);
or U19887 (N_19887,N_17539,N_17883);
or U19888 (N_19888,N_17552,N_16887);
nor U19889 (N_19889,N_17788,N_16045);
or U19890 (N_19890,N_16620,N_17188);
nand U19891 (N_19891,N_17871,N_16758);
xnor U19892 (N_19892,N_16317,N_17647);
nor U19893 (N_19893,N_16488,N_16691);
or U19894 (N_19894,N_17104,N_16441);
xnor U19895 (N_19895,N_16404,N_17540);
nand U19896 (N_19896,N_16477,N_16447);
xor U19897 (N_19897,N_17359,N_16145);
and U19898 (N_19898,N_16323,N_16349);
nor U19899 (N_19899,N_16442,N_16500);
xor U19900 (N_19900,N_16575,N_16472);
nor U19901 (N_19901,N_16732,N_17852);
and U19902 (N_19902,N_16897,N_17378);
and U19903 (N_19903,N_17275,N_16077);
xor U19904 (N_19904,N_16434,N_16335);
nand U19905 (N_19905,N_16953,N_16454);
or U19906 (N_19906,N_16126,N_16114);
and U19907 (N_19907,N_16928,N_17114);
nor U19908 (N_19908,N_16633,N_17878);
nand U19909 (N_19909,N_16228,N_17003);
nor U19910 (N_19910,N_16642,N_16338);
nor U19911 (N_19911,N_17989,N_17916);
or U19912 (N_19912,N_17369,N_17869);
and U19913 (N_19913,N_16477,N_16294);
and U19914 (N_19914,N_16110,N_16371);
and U19915 (N_19915,N_16503,N_16026);
nor U19916 (N_19916,N_17458,N_16974);
nand U19917 (N_19917,N_16618,N_16993);
or U19918 (N_19918,N_16067,N_16139);
and U19919 (N_19919,N_16743,N_17838);
xnor U19920 (N_19920,N_16084,N_16008);
and U19921 (N_19921,N_17341,N_17347);
xnor U19922 (N_19922,N_17748,N_17863);
nand U19923 (N_19923,N_16548,N_17221);
nand U19924 (N_19924,N_16566,N_17166);
or U19925 (N_19925,N_17393,N_17362);
and U19926 (N_19926,N_16572,N_17116);
or U19927 (N_19927,N_17999,N_17753);
nor U19928 (N_19928,N_17476,N_17919);
xnor U19929 (N_19929,N_17009,N_16912);
nor U19930 (N_19930,N_16476,N_16116);
nand U19931 (N_19931,N_16914,N_16704);
xor U19932 (N_19932,N_17551,N_17991);
or U19933 (N_19933,N_16204,N_16566);
and U19934 (N_19934,N_17258,N_16358);
and U19935 (N_19935,N_16488,N_17477);
nor U19936 (N_19936,N_16839,N_17072);
xor U19937 (N_19937,N_16607,N_17394);
nand U19938 (N_19938,N_16593,N_17606);
and U19939 (N_19939,N_17647,N_16434);
xor U19940 (N_19940,N_17190,N_17120);
nor U19941 (N_19941,N_17666,N_16041);
nor U19942 (N_19942,N_16805,N_16166);
and U19943 (N_19943,N_16349,N_16629);
or U19944 (N_19944,N_16104,N_17265);
xor U19945 (N_19945,N_17019,N_17358);
and U19946 (N_19946,N_17503,N_16463);
nor U19947 (N_19947,N_16197,N_16539);
or U19948 (N_19948,N_16894,N_17197);
nand U19949 (N_19949,N_16051,N_16032);
and U19950 (N_19950,N_17859,N_16815);
nor U19951 (N_19951,N_16255,N_16884);
nand U19952 (N_19952,N_17179,N_17601);
or U19953 (N_19953,N_17154,N_17443);
xnor U19954 (N_19954,N_17561,N_17018);
or U19955 (N_19955,N_17552,N_16747);
nand U19956 (N_19956,N_17435,N_16631);
xor U19957 (N_19957,N_17581,N_17127);
nor U19958 (N_19958,N_16976,N_17777);
xnor U19959 (N_19959,N_17276,N_16762);
and U19960 (N_19960,N_17240,N_16687);
xor U19961 (N_19961,N_16477,N_17350);
or U19962 (N_19962,N_17549,N_16483);
and U19963 (N_19963,N_17233,N_17068);
nand U19964 (N_19964,N_17228,N_16588);
nor U19965 (N_19965,N_17946,N_17600);
and U19966 (N_19966,N_16430,N_16594);
xnor U19967 (N_19967,N_17503,N_17752);
xnor U19968 (N_19968,N_17195,N_17723);
nor U19969 (N_19969,N_17502,N_17038);
nor U19970 (N_19970,N_16770,N_16645);
and U19971 (N_19971,N_16562,N_17297);
nand U19972 (N_19972,N_16234,N_16520);
and U19973 (N_19973,N_16559,N_17903);
nor U19974 (N_19974,N_17964,N_17045);
or U19975 (N_19975,N_17681,N_17151);
and U19976 (N_19976,N_17888,N_16465);
and U19977 (N_19977,N_17149,N_16846);
nand U19978 (N_19978,N_17209,N_17189);
and U19979 (N_19979,N_17164,N_16650);
nand U19980 (N_19980,N_16002,N_17548);
nand U19981 (N_19981,N_17939,N_16903);
xor U19982 (N_19982,N_16960,N_17269);
nor U19983 (N_19983,N_16278,N_16612);
or U19984 (N_19984,N_17868,N_17865);
nor U19985 (N_19985,N_17582,N_17692);
nor U19986 (N_19986,N_17695,N_16799);
xnor U19987 (N_19987,N_16211,N_16709);
nand U19988 (N_19988,N_17766,N_16221);
and U19989 (N_19989,N_16167,N_17014);
nor U19990 (N_19990,N_17454,N_16342);
and U19991 (N_19991,N_16129,N_17201);
xor U19992 (N_19992,N_17736,N_17358);
or U19993 (N_19993,N_16828,N_17862);
and U19994 (N_19994,N_17649,N_16502);
nand U19995 (N_19995,N_17472,N_17512);
or U19996 (N_19996,N_16844,N_17058);
and U19997 (N_19997,N_17018,N_16453);
or U19998 (N_19998,N_17723,N_17255);
nand U19999 (N_19999,N_16198,N_16501);
nand U20000 (N_20000,N_18633,N_19047);
nor U20001 (N_20001,N_19918,N_18226);
xor U20002 (N_20002,N_19692,N_19401);
nand U20003 (N_20003,N_18130,N_19435);
or U20004 (N_20004,N_19619,N_19444);
nor U20005 (N_20005,N_18474,N_19792);
nor U20006 (N_20006,N_19524,N_19715);
and U20007 (N_20007,N_18879,N_19756);
xor U20008 (N_20008,N_18017,N_18685);
and U20009 (N_20009,N_19812,N_18638);
nor U20010 (N_20010,N_18236,N_18037);
xnor U20011 (N_20011,N_18352,N_19602);
xor U20012 (N_20012,N_19656,N_19098);
and U20013 (N_20013,N_18794,N_18376);
or U20014 (N_20014,N_18332,N_18217);
xor U20015 (N_20015,N_19860,N_18787);
and U20016 (N_20016,N_18694,N_18378);
xor U20017 (N_20017,N_18229,N_19407);
nor U20018 (N_20018,N_19273,N_18262);
and U20019 (N_20019,N_19445,N_18979);
xnor U20020 (N_20020,N_18359,N_18180);
and U20021 (N_20021,N_18254,N_19381);
nand U20022 (N_20022,N_19202,N_19084);
and U20023 (N_20023,N_19873,N_18384);
nor U20024 (N_20024,N_18123,N_18019);
nand U20025 (N_20025,N_19997,N_19956);
xor U20026 (N_20026,N_19932,N_18839);
xor U20027 (N_20027,N_19388,N_18976);
nor U20028 (N_20028,N_19744,N_19820);
nor U20029 (N_20029,N_19788,N_19944);
or U20030 (N_20030,N_18868,N_18422);
and U20031 (N_20031,N_18552,N_19746);
nand U20032 (N_20032,N_18972,N_19092);
or U20033 (N_20033,N_18690,N_19433);
nand U20034 (N_20034,N_19802,N_18780);
xnor U20035 (N_20035,N_19907,N_18782);
and U20036 (N_20036,N_19431,N_19199);
nand U20037 (N_20037,N_18047,N_19420);
or U20038 (N_20038,N_19081,N_18615);
xor U20039 (N_20039,N_18173,N_18007);
nand U20040 (N_20040,N_19422,N_18160);
or U20041 (N_20041,N_19986,N_18726);
and U20042 (N_20042,N_19590,N_18958);
nand U20043 (N_20043,N_19782,N_19897);
nor U20044 (N_20044,N_18873,N_19371);
or U20045 (N_20045,N_19163,N_19728);
xnor U20046 (N_20046,N_19366,N_18901);
nor U20047 (N_20047,N_18911,N_19830);
or U20048 (N_20048,N_18593,N_19637);
nand U20049 (N_20049,N_18573,N_19653);
nor U20050 (N_20050,N_19367,N_18930);
or U20051 (N_20051,N_18364,N_19041);
nor U20052 (N_20052,N_19940,N_19707);
or U20053 (N_20053,N_18074,N_18326);
nand U20054 (N_20054,N_19103,N_18788);
xnor U20055 (N_20055,N_19177,N_18659);
or U20056 (N_20056,N_18616,N_19253);
or U20057 (N_20057,N_19072,N_19526);
nand U20058 (N_20058,N_18482,N_18775);
nor U20059 (N_20059,N_18921,N_19896);
xnor U20060 (N_20060,N_19669,N_19233);
nor U20061 (N_20061,N_18696,N_19443);
nor U20062 (N_20062,N_19374,N_18767);
or U20063 (N_20063,N_18916,N_18571);
and U20064 (N_20064,N_19819,N_18466);
or U20065 (N_20065,N_19414,N_19842);
and U20066 (N_20066,N_18744,N_19710);
or U20067 (N_20067,N_18974,N_18932);
xor U20068 (N_20068,N_18042,N_18650);
or U20069 (N_20069,N_18760,N_18931);
nor U20070 (N_20070,N_18026,N_18212);
and U20071 (N_20071,N_18349,N_18802);
and U20072 (N_20072,N_18344,N_19703);
nand U20073 (N_20073,N_19716,N_18555);
nand U20074 (N_20074,N_19416,N_18134);
xor U20075 (N_20075,N_19584,N_18486);
or U20076 (N_20076,N_19816,N_19425);
and U20077 (N_20077,N_19507,N_19126);
and U20078 (N_20078,N_18305,N_19377);
xnor U20079 (N_20079,N_19941,N_18537);
nor U20080 (N_20080,N_19219,N_18651);
nor U20081 (N_20081,N_19133,N_18610);
and U20082 (N_20082,N_18645,N_19238);
xnor U20083 (N_20083,N_19195,N_19724);
nand U20084 (N_20084,N_18097,N_19666);
and U20085 (N_20085,N_19596,N_19031);
nor U20086 (N_20086,N_19234,N_19158);
or U20087 (N_20087,N_19850,N_19739);
nand U20088 (N_20088,N_19650,N_18463);
xnor U20089 (N_20089,N_19586,N_18128);
or U20090 (N_20090,N_19457,N_19933);
and U20091 (N_20091,N_18941,N_18275);
xnor U20092 (N_20092,N_19828,N_19384);
nand U20093 (N_20093,N_19495,N_18303);
nand U20094 (N_20094,N_19589,N_18678);
nor U20095 (N_20095,N_18588,N_18842);
nor U20096 (N_20096,N_18478,N_18233);
nor U20097 (N_20097,N_19468,N_19761);
or U20098 (N_20098,N_19925,N_18604);
xor U20099 (N_20099,N_18693,N_18483);
or U20100 (N_20100,N_19752,N_19632);
or U20101 (N_20101,N_19309,N_18838);
nor U20102 (N_20102,N_18515,N_19286);
nand U20103 (N_20103,N_18957,N_19390);
nand U20104 (N_20104,N_19389,N_18589);
or U20105 (N_20105,N_18269,N_19517);
xnor U20106 (N_20106,N_19448,N_18152);
or U20107 (N_20107,N_19198,N_18291);
and U20108 (N_20108,N_18677,N_19591);
nor U20109 (N_20109,N_19854,N_18540);
and U20110 (N_20110,N_19415,N_18521);
xor U20111 (N_20111,N_18465,N_18689);
and U20112 (N_20112,N_18993,N_18113);
nor U20113 (N_20113,N_18129,N_19034);
or U20114 (N_20114,N_18220,N_19354);
and U20115 (N_20115,N_18820,N_18665);
nor U20116 (N_20116,N_18594,N_18239);
nand U20117 (N_20117,N_19581,N_19654);
and U20118 (N_20118,N_18982,N_19464);
nand U20119 (N_20119,N_18015,N_19644);
nand U20120 (N_20120,N_18263,N_18080);
xnor U20121 (N_20121,N_18554,N_19527);
nand U20122 (N_20122,N_19778,N_19529);
nor U20123 (N_20123,N_19076,N_18402);
nor U20124 (N_20124,N_19889,N_18886);
or U20125 (N_20125,N_19063,N_19958);
xor U20126 (N_20126,N_18582,N_18513);
xor U20127 (N_20127,N_18016,N_19070);
or U20128 (N_20128,N_18829,N_19292);
xor U20129 (N_20129,N_18411,N_18781);
xnor U20130 (N_20130,N_18968,N_18570);
nor U20131 (N_20131,N_19851,N_18193);
and U20132 (N_20132,N_18188,N_19593);
and U20133 (N_20133,N_18737,N_19797);
xnor U20134 (N_20134,N_19664,N_19601);
xor U20135 (N_20135,N_18860,N_19531);
xor U20136 (N_20136,N_19643,N_19683);
nand U20137 (N_20137,N_19411,N_18599);
nand U20138 (N_20138,N_18070,N_19395);
or U20139 (N_20139,N_19722,N_18255);
nor U20140 (N_20140,N_18048,N_18003);
nand U20141 (N_20141,N_18452,N_19540);
or U20142 (N_20142,N_18260,N_19522);
nor U20143 (N_20143,N_19614,N_18218);
nand U20144 (N_20144,N_19511,N_18613);
or U20145 (N_20145,N_18966,N_19821);
or U20146 (N_20146,N_18222,N_18306);
or U20147 (N_20147,N_19434,N_18713);
nor U20148 (N_20148,N_19200,N_19353);
nand U20149 (N_20149,N_19447,N_18531);
and U20150 (N_20150,N_18825,N_18283);
or U20151 (N_20151,N_19675,N_18964);
or U20152 (N_20152,N_18064,N_19329);
nand U20153 (N_20153,N_18102,N_18824);
nand U20154 (N_20154,N_18424,N_19969);
and U20155 (N_20155,N_19916,N_19843);
or U20156 (N_20156,N_18155,N_18747);
or U20157 (N_20157,N_18034,N_19698);
xor U20158 (N_20158,N_19680,N_19505);
nand U20159 (N_20159,N_18362,N_19067);
xor U20160 (N_20160,N_18150,N_18435);
nor U20161 (N_20161,N_19811,N_19695);
nand U20162 (N_20162,N_19004,N_18365);
and U20163 (N_20163,N_18598,N_19544);
or U20164 (N_20164,N_19311,N_19334);
or U20165 (N_20165,N_18679,N_19357);
nor U20166 (N_20166,N_19069,N_19386);
nor U20167 (N_20167,N_18994,N_18965);
or U20168 (N_20168,N_18211,N_18700);
nor U20169 (N_20169,N_19839,N_19024);
and U20170 (N_20170,N_18041,N_18823);
nand U20171 (N_20171,N_18244,N_18237);
nor U20172 (N_20172,N_19146,N_19406);
nand U20173 (N_20173,N_18487,N_19473);
nor U20174 (N_20174,N_18637,N_18423);
and U20175 (N_20175,N_18175,N_19691);
nand U20176 (N_20176,N_19770,N_19835);
nand U20177 (N_20177,N_19831,N_19116);
and U20178 (N_20178,N_19502,N_18415);
xor U20179 (N_20179,N_19316,N_19278);
and U20180 (N_20180,N_19400,N_18628);
or U20181 (N_20181,N_18116,N_18373);
xnor U20182 (N_20182,N_19912,N_19834);
or U20183 (N_20183,N_19700,N_19139);
nor U20184 (N_20184,N_18197,N_19143);
xnor U20185 (N_20185,N_19803,N_19676);
and U20186 (N_20186,N_19165,N_19350);
nor U20187 (N_20187,N_19312,N_19885);
xnor U20188 (N_20188,N_19972,N_19884);
nand U20189 (N_20189,N_19276,N_18101);
nor U20190 (N_20190,N_18107,N_19382);
nand U20191 (N_20191,N_19314,N_18387);
nor U20192 (N_20192,N_18315,N_19571);
and U20193 (N_20193,N_19627,N_18514);
or U20194 (N_20194,N_19167,N_18833);
or U20195 (N_20195,N_19240,N_19623);
and U20196 (N_20196,N_19156,N_18765);
nor U20197 (N_20197,N_18984,N_18380);
nand U20198 (N_20198,N_18472,N_19114);
and U20199 (N_20199,N_19423,N_19304);
nand U20200 (N_20200,N_18319,N_19483);
nor U20201 (N_20201,N_18928,N_18078);
nand U20202 (N_20202,N_19642,N_19258);
nand U20203 (N_20203,N_19702,N_19224);
or U20204 (N_20204,N_19943,N_19061);
nand U20205 (N_20205,N_18158,N_18271);
and U20206 (N_20206,N_19302,N_18115);
xnor U20207 (N_20207,N_19799,N_18835);
or U20208 (N_20208,N_18250,N_19837);
or U20209 (N_20209,N_18910,N_18159);
nand U20210 (N_20210,N_19921,N_18494);
nand U20211 (N_20211,N_19236,N_19757);
nand U20212 (N_20212,N_19725,N_18285);
or U20213 (N_20213,N_18827,N_19610);
nand U20214 (N_20214,N_19106,N_19300);
or U20215 (N_20215,N_19608,N_19585);
nor U20216 (N_20216,N_19364,N_18177);
or U20217 (N_20217,N_18161,N_18528);
and U20218 (N_20218,N_19111,N_19536);
xor U20219 (N_20219,N_19313,N_19478);
and U20220 (N_20220,N_18817,N_18664);
and U20221 (N_20221,N_18249,N_19399);
nor U20222 (N_20222,N_19569,N_19658);
nand U20223 (N_20223,N_18333,N_18338);
and U20224 (N_20224,N_18623,N_18058);
xnor U20225 (N_20225,N_19056,N_18277);
xor U20226 (N_20226,N_19849,N_19494);
nor U20227 (N_20227,N_18018,N_18273);
nor U20228 (N_20228,N_19318,N_18471);
and U20229 (N_20229,N_19065,N_19773);
xnor U20230 (N_20230,N_19170,N_19732);
nand U20231 (N_20231,N_19563,N_18795);
nor U20232 (N_20232,N_18684,N_19904);
xnor U20233 (N_20233,N_19039,N_19442);
nor U20234 (N_20234,N_18209,N_18290);
xnor U20235 (N_20235,N_19814,N_19089);
nor U20236 (N_20236,N_19005,N_19567);
nor U20237 (N_20237,N_18844,N_19613);
or U20238 (N_20238,N_19221,N_18138);
nand U20239 (N_20239,N_18025,N_19470);
xor U20240 (N_20240,N_19144,N_19462);
or U20241 (N_20241,N_18140,N_19346);
and U20242 (N_20242,N_18316,N_19518);
and U20243 (N_20243,N_18776,N_18027);
and U20244 (N_20244,N_18996,N_18722);
nand U20245 (N_20245,N_19378,N_18118);
and U20246 (N_20246,N_18766,N_18578);
nor U20247 (N_20247,N_18580,N_18553);
nor U20248 (N_20248,N_18717,N_18826);
nand U20249 (N_20249,N_19458,N_19127);
nand U20250 (N_20250,N_18350,N_19947);
xor U20251 (N_20251,N_18754,N_19772);
or U20252 (N_20252,N_18506,N_19417);
and U20253 (N_20253,N_18029,N_18718);
and U20254 (N_20254,N_18866,N_19264);
and U20255 (N_20255,N_19841,N_18146);
nand U20256 (N_20256,N_18060,N_18327);
nor U20257 (N_20257,N_19191,N_19135);
and U20258 (N_20258,N_19243,N_19784);
xnor U20259 (N_20259,N_18992,N_18205);
and U20260 (N_20260,N_18377,N_18192);
or U20261 (N_20261,N_18607,N_19351);
nor U20262 (N_20262,N_19895,N_18281);
nand U20263 (N_20263,N_19343,N_18559);
nor U20264 (N_20264,N_19731,N_19994);
nor U20265 (N_20265,N_18156,N_19844);
and U20266 (N_20266,N_19222,N_19398);
xnor U20267 (N_20267,N_19679,N_18575);
nand U20268 (N_20268,N_19790,N_18300);
xor U20269 (N_20269,N_19392,N_19881);
nand U20270 (N_20270,N_18227,N_19019);
nand U20271 (N_20271,N_19760,N_18800);
and U20272 (N_20272,N_19159,N_18467);
and U20273 (N_20273,N_19936,N_19101);
or U20274 (N_20274,N_18937,N_18938);
or U20275 (N_20275,N_19781,N_18654);
or U20276 (N_20276,N_18404,N_18927);
nor U20277 (N_20277,N_19751,N_19147);
xnor U20278 (N_20278,N_19391,N_19869);
xor U20279 (N_20279,N_19338,N_18977);
nor U20280 (N_20280,N_18186,N_18240);
xor U20281 (N_20281,N_19570,N_19882);
and U20282 (N_20282,N_18929,N_19682);
and U20283 (N_20283,N_19893,N_18956);
or U20284 (N_20284,N_18566,N_18169);
xor U20285 (N_20285,N_18307,N_18023);
nand U20286 (N_20286,N_18774,N_18301);
or U20287 (N_20287,N_19244,N_19847);
nor U20288 (N_20288,N_19694,N_18495);
xor U20289 (N_20289,N_18092,N_19934);
xnor U20290 (N_20290,N_18353,N_19520);
and U20291 (N_20291,N_18321,N_18550);
xor U20292 (N_20292,N_19331,N_19226);
nor U20293 (N_20293,N_18213,N_19824);
nand U20294 (N_20294,N_19651,N_18636);
and U20295 (N_20295,N_18071,N_19293);
and U20296 (N_20296,N_18065,N_19546);
xor U20297 (N_20297,N_18735,N_18000);
nor U20298 (N_20298,N_18953,N_19987);
or U20299 (N_20299,N_18224,N_19991);
xnor U20300 (N_20300,N_19574,N_18697);
xor U20301 (N_20301,N_18777,N_19192);
nor U20302 (N_20302,N_18661,N_19430);
or U20303 (N_20303,N_18125,N_19631);
or U20304 (N_20304,N_18312,N_19418);
xor U20305 (N_20305,N_19588,N_18597);
xnor U20306 (N_20306,N_19132,N_19685);
nor U20307 (N_20307,N_18475,N_19568);
nor U20308 (N_20308,N_19961,N_19503);
or U20309 (N_20309,N_18234,N_18818);
xnor U20310 (N_20310,N_18539,N_18302);
nor U20311 (N_20311,N_19104,N_18756);
nor U20312 (N_20312,N_18856,N_19310);
nand U20313 (N_20313,N_19216,N_18687);
nor U20314 (N_20314,N_18807,N_18520);
xnor U20315 (N_20315,N_18455,N_19467);
nand U20316 (N_20316,N_19917,N_19485);
nand U20317 (N_20317,N_18538,N_19469);
or U20318 (N_20318,N_19487,N_19022);
nor U20319 (N_20319,N_18581,N_19635);
nor U20320 (N_20320,N_19930,N_18769);
nor U20321 (N_20321,N_18715,N_18657);
xnor U20322 (N_20322,N_18725,N_18668);
xor U20323 (N_20323,N_19051,N_19050);
nor U20324 (N_20324,N_19124,N_18347);
or U20325 (N_20325,N_18527,N_19767);
or U20326 (N_20326,N_18081,N_19856);
xor U20327 (N_20327,N_18961,N_19184);
nand U20328 (N_20328,N_19628,N_19187);
or U20329 (N_20329,N_19361,N_19335);
or U20330 (N_20330,N_18088,N_18317);
nor U20331 (N_20331,N_19855,N_18858);
and U20332 (N_20332,N_19951,N_19538);
xnor U20333 (N_20333,N_19306,N_19681);
nor U20334 (N_20334,N_18459,N_18208);
and U20335 (N_20335,N_18557,N_19826);
xnor U20336 (N_20336,N_19575,N_19204);
nand U20337 (N_20337,N_19813,N_18453);
and U20338 (N_20338,N_18428,N_19677);
xnor U20339 (N_20339,N_19360,N_18682);
and U20340 (N_20340,N_18848,N_18174);
or U20341 (N_20341,N_19029,N_19603);
nand U20342 (N_20342,N_19848,N_18897);
nand U20343 (N_20343,N_19237,N_19129);
or U20344 (N_20344,N_19594,N_18840);
nand U20345 (N_20345,N_19136,N_19624);
nor U20346 (N_20346,N_19209,N_19214);
nand U20347 (N_20347,N_19937,N_18079);
or U20348 (N_20348,N_18987,N_19708);
nand U20349 (N_20349,N_19554,N_19138);
or U20350 (N_20350,N_18536,N_18278);
nor U20351 (N_20351,N_19213,N_18356);
nor U20352 (N_20352,N_19786,N_18367);
nand U20353 (N_20353,N_18199,N_19871);
and U20354 (N_20354,N_19674,N_18914);
or U20355 (N_20355,N_19924,N_18167);
and U20356 (N_20356,N_19976,N_18630);
xor U20357 (N_20357,N_18653,N_19975);
or U20358 (N_20358,N_18462,N_19862);
or U20359 (N_20359,N_18811,N_19965);
and U20360 (N_20360,N_19421,N_19564);
xnor U20361 (N_20361,N_18634,N_18625);
or U20362 (N_20362,N_19197,N_18279);
or U20363 (N_20363,N_19647,N_19110);
and U20364 (N_20364,N_19324,N_18343);
and U20365 (N_20365,N_18567,N_19438);
xor U20366 (N_20366,N_19973,N_18759);
nor U20367 (N_20367,N_18510,N_19966);
or U20368 (N_20368,N_19688,N_18892);
nand U20369 (N_20369,N_19606,N_18267);
xor U20370 (N_20370,N_19962,N_18389);
nand U20371 (N_20371,N_18099,N_18778);
and U20372 (N_20372,N_19307,N_18642);
nand U20373 (N_20373,N_19745,N_18532);
and U20374 (N_20374,N_18086,N_18813);
xor U20375 (N_20375,N_19530,N_18488);
and U20376 (N_20376,N_19193,N_19892);
nand U20377 (N_20377,N_18298,N_19189);
and U20378 (N_20378,N_18728,N_18590);
and U20379 (N_20379,N_19794,N_19274);
xnor U20380 (N_20380,N_18114,N_19995);
nor U20381 (N_20381,N_18900,N_19149);
nand U20382 (N_20382,N_19883,N_18434);
nand U20383 (N_20383,N_19979,N_18545);
or U20384 (N_20384,N_18410,N_18414);
nor U20385 (N_20385,N_18969,N_18256);
and U20386 (N_20386,N_18711,N_18368);
nor U20387 (N_20387,N_18806,N_19727);
xor U20388 (N_20388,N_18738,N_19742);
and U20389 (N_20389,N_18087,N_18028);
nor U20390 (N_20390,N_19454,N_19370);
and U20391 (N_20391,N_18342,N_19718);
and U20392 (N_20392,N_19074,N_19087);
and U20393 (N_20393,N_19678,N_18591);
nand U20394 (N_20394,N_19164,N_18336);
and U20395 (N_20395,N_18988,N_18006);
nand U20396 (N_20396,N_19989,N_19748);
nand U20397 (N_20397,N_19119,N_18874);
or U20398 (N_20398,N_18461,N_19036);
xnor U20399 (N_20399,N_19689,N_18878);
nor U20400 (N_20400,N_19394,N_19319);
and U20401 (N_20401,N_18460,N_19481);
or U20402 (N_20402,N_18194,N_19577);
xor U20403 (N_20403,N_19446,N_18324);
and U20404 (N_20404,N_18153,N_19121);
or U20405 (N_20405,N_18135,N_18764);
nand U20406 (N_20406,N_18309,N_19935);
nor U20407 (N_20407,N_18214,N_19915);
nand U20408 (N_20408,N_19117,N_18951);
nor U20409 (N_20409,N_19879,N_19931);
nor U20410 (N_20410,N_19403,N_19393);
and U20411 (N_20411,N_19141,N_19342);
nand U20412 (N_20412,N_18899,N_19058);
nand U20413 (N_20413,N_19323,N_18100);
nor U20414 (N_20414,N_18225,N_19380);
xnor U20415 (N_20415,N_18068,N_19426);
and U20416 (N_20416,N_18004,N_18119);
xor U20417 (N_20417,N_18917,N_18808);
nand U20418 (N_20418,N_18076,N_18740);
nor U20419 (N_20419,N_19515,N_18108);
or U20420 (N_20420,N_18762,N_18959);
nand U20421 (N_20421,N_19920,N_18656);
nand U20422 (N_20422,N_19479,N_19097);
nor U20423 (N_20423,N_19059,N_19376);
and U20424 (N_20424,N_19471,N_18403);
xor U20425 (N_20425,N_19489,N_19296);
or U20426 (N_20426,N_18758,N_18484);
nand U20427 (N_20427,N_18187,N_19550);
and U20428 (N_20428,N_18259,N_18323);
nor U20429 (N_20429,N_18091,N_18360);
xor U20430 (N_20430,N_19858,N_18676);
nand U20431 (N_20431,N_18832,N_18274);
nor U20432 (N_20432,N_18310,N_19512);
and U20433 (N_20433,N_19449,N_19809);
nand U20434 (N_20434,N_19611,N_19450);
and U20435 (N_20435,N_18647,N_18383);
nand U20436 (N_20436,N_18564,N_18147);
xnor U20437 (N_20437,N_18955,N_19043);
or U20438 (N_20438,N_19086,N_18366);
and U20439 (N_20439,N_18902,N_18096);
xor U20440 (N_20440,N_18293,N_18329);
xnor U20441 (N_20441,N_19295,N_18721);
nor U20442 (N_20442,N_18995,N_18978);
or U20443 (N_20443,N_18390,N_18533);
and U20444 (N_20444,N_18082,N_19134);
xnor U20445 (N_20445,N_18970,N_19118);
nand U20446 (N_20446,N_19340,N_19317);
nand U20447 (N_20447,N_19131,N_18952);
and U20448 (N_20448,N_19217,N_18215);
nand U20449 (N_20449,N_19257,N_18406);
nor U20450 (N_20450,N_19155,N_18526);
xor U20451 (N_20451,N_19665,N_18393);
nor U20452 (N_20452,N_19075,N_18809);
nor U20453 (N_20453,N_18816,N_18544);
xor U20454 (N_20454,N_18062,N_19952);
nand U20455 (N_20455,N_18083,N_18541);
and U20456 (N_20456,N_19833,N_18031);
nor U20457 (N_20457,N_18672,N_18865);
xnor U20458 (N_20458,N_18755,N_18106);
and U20459 (N_20459,N_18556,N_18529);
xor U20460 (N_20460,N_19763,N_19579);
or U20461 (N_20461,N_18891,N_18543);
and U20462 (N_20462,N_19369,N_19609);
and U20463 (N_20463,N_19359,N_19080);
or U20464 (N_20464,N_19115,N_19419);
nor U20465 (N_20465,N_19154,N_18392);
xnor U20466 (N_20466,N_18056,N_19804);
or U20467 (N_20467,N_18012,N_18370);
xnor U20468 (N_20468,N_19152,N_19789);
nor U20469 (N_20469,N_18960,N_19181);
and U20470 (N_20470,N_19242,N_18592);
or U20471 (N_20471,N_18375,N_19720);
or U20472 (N_20472,N_18221,N_18635);
nand U20473 (N_20473,N_19476,N_18669);
and U20474 (N_20474,N_19123,N_18439);
and U20475 (N_20475,N_18330,N_18855);
nor U20476 (N_20476,N_18986,N_18204);
or U20477 (N_20477,N_19301,N_18354);
xnor U20478 (N_20478,N_19053,N_19533);
nor U20479 (N_20479,N_18066,N_18525);
or U20480 (N_20480,N_19525,N_19451);
xnor U20481 (N_20481,N_18162,N_19771);
nor U20482 (N_20482,N_19501,N_19905);
or U20483 (N_20483,N_19160,N_18785);
nand U20484 (N_20484,N_19212,N_18803);
or U20485 (N_20485,N_18121,N_19641);
or U20486 (N_20486,N_18662,N_18334);
nand U20487 (N_20487,N_19829,N_19040);
xor U20488 (N_20488,N_18698,N_19970);
xor U20489 (N_20489,N_18145,N_18201);
and U20490 (N_20490,N_18178,N_19755);
or U20491 (N_20491,N_19218,N_18622);
and U20492 (N_20492,N_18862,N_19003);
nor U20493 (N_20493,N_18110,N_19545);
and U20494 (N_20494,N_19007,N_18845);
and U20495 (N_20495,N_18286,N_18949);
nor U20496 (N_20496,N_19713,N_18846);
nand U20497 (N_20497,N_18508,N_18761);
and U20498 (N_20498,N_18733,N_19145);
xor U20499 (N_20499,N_19140,N_19356);
nor U20500 (N_20500,N_19753,N_19281);
xor U20501 (N_20501,N_19348,N_19112);
nor U20502 (N_20502,N_18524,N_18417);
xnor U20503 (N_20503,N_18502,N_18339);
or U20504 (N_20504,N_19870,N_18479);
or U20505 (N_20505,N_19011,N_19514);
or U20506 (N_20506,N_19992,N_18745);
nor U20507 (N_20507,N_19998,N_18692);
or U20508 (N_20508,N_19322,N_18511);
nor U20509 (N_20509,N_19396,N_19865);
xor U20510 (N_20510,N_18388,N_19336);
or U20511 (N_20511,N_18702,N_19280);
or U20512 (N_20512,N_18111,N_19832);
nand U20513 (N_20513,N_18709,N_19743);
or U20514 (N_20514,N_18729,N_18743);
nor U20515 (N_20515,N_18516,N_19805);
nand U20516 (N_20516,N_18010,N_18923);
nor U20517 (N_20517,N_19566,N_19977);
nand U20518 (N_20518,N_18433,N_18105);
nand U20519 (N_20519,N_19899,N_19983);
or U20520 (N_20520,N_19779,N_18021);
nand U20521 (N_20521,N_19622,N_19345);
or U20522 (N_20522,N_19161,N_18407);
xnor U20523 (N_20523,N_19232,N_18624);
nand U20524 (N_20524,N_19246,N_18489);
and U20525 (N_20525,N_19082,N_19453);
xnor U20526 (N_20526,N_19981,N_19235);
and U20527 (N_20527,N_18126,N_18936);
nand U20528 (N_20528,N_19793,N_19482);
and U20529 (N_20529,N_19347,N_18967);
nand U20530 (N_20530,N_18699,N_18841);
and U20531 (N_20531,N_19723,N_19633);
or U20532 (N_20532,N_19352,N_18401);
and U20533 (N_20533,N_18207,N_18763);
nand U20534 (N_20534,N_18551,N_19048);
xnor U20535 (N_20535,N_19562,N_18837);
and U20536 (N_20536,N_18646,N_18067);
or U20537 (N_20537,N_19827,N_19898);
nor U20538 (N_20538,N_18605,N_19878);
or U20539 (N_20539,N_19409,N_19629);
or U20540 (N_20540,N_18094,N_19291);
nand U20541 (N_20541,N_19553,N_18024);
xor U20542 (N_20542,N_18331,N_18182);
nand U20543 (N_20543,N_19277,N_18660);
or U20544 (N_20544,N_18893,N_19052);
xor U20545 (N_20545,N_19012,N_18132);
and U20546 (N_20546,N_18050,N_18451);
xnor U20547 (N_20547,N_18355,N_19985);
nor U20548 (N_20548,N_18640,N_19496);
or U20549 (N_20549,N_18798,N_18834);
or U20550 (N_20550,N_19499,N_19079);
nand U20551 (N_20551,N_19867,N_19137);
xor U20552 (N_20552,N_18480,N_19735);
or U20553 (N_20553,N_18836,N_18266);
and U20554 (N_20554,N_18889,N_18202);
or U20555 (N_20555,N_19432,N_18688);
nand U20556 (N_20556,N_19903,N_19617);
nand U20557 (N_20557,N_19785,N_19288);
and U20558 (N_20558,N_19211,N_18680);
and U20559 (N_20559,N_19539,N_19460);
xnor U20560 (N_20560,N_18584,N_18382);
nor U20561 (N_20561,N_19194,N_18276);
nand U20562 (N_20562,N_19948,N_19874);
or U20563 (N_20563,N_19999,N_19166);
nor U20564 (N_20564,N_19696,N_19027);
nor U20565 (N_20565,N_18621,N_19456);
or U20566 (N_20566,N_19178,N_18629);
and U20567 (N_20567,N_19510,N_18627);
or U20568 (N_20568,N_18265,N_19017);
nor U20569 (N_20569,N_18036,N_19332);
or U20570 (N_20570,N_19180,N_18171);
nand U20571 (N_20571,N_18704,N_18141);
or U20572 (N_20572,N_19227,N_18247);
xor U20573 (N_20573,N_18179,N_19157);
and U20574 (N_20574,N_19521,N_18304);
xor U20575 (N_20575,N_18268,N_19488);
xnor U20576 (N_20576,N_19625,N_18548);
nand U20577 (N_20577,N_19592,N_18491);
nand U20578 (N_20578,N_19028,N_19887);
and U20579 (N_20579,N_18449,N_19297);
nor U20580 (N_20580,N_18719,N_19455);
nand U20581 (N_20581,N_19190,N_18013);
and U20582 (N_20582,N_19706,N_19960);
nor U20583 (N_20583,N_19894,N_19289);
or U20584 (N_20584,N_19825,N_19020);
or U20585 (N_20585,N_19648,N_19206);
nor U20586 (N_20586,N_19339,N_18231);
nor U20587 (N_20587,N_18493,N_18361);
nand U20588 (N_20588,N_18973,N_19565);
and U20589 (N_20589,N_18098,N_19910);
xnor U20590 (N_20590,N_18731,N_19498);
or U20591 (N_20591,N_18707,N_18020);
nand U20592 (N_20592,N_18985,N_19441);
and U20593 (N_20593,N_19699,N_18601);
xor U20594 (N_20594,N_19284,N_18444);
nor U20595 (N_20595,N_18440,N_19402);
xnor U20596 (N_20596,N_19477,N_18412);
nor U20597 (N_20597,N_18904,N_19740);
or U20598 (N_20598,N_19810,N_19255);
and U20599 (N_20599,N_19328,N_19045);
xor U20600 (N_20600,N_18261,N_18857);
and U20601 (N_20601,N_19967,N_19968);
nor U20602 (N_20602,N_19267,N_18876);
xor U20603 (N_20603,N_18503,N_18828);
nand U20604 (N_20604,N_19108,N_19942);
xnor U20605 (N_20605,N_18093,N_19093);
nand U20606 (N_20606,N_18882,N_19815);
or U20607 (N_20607,N_19955,N_19128);
nand U20608 (N_20608,N_18568,N_19791);
nand U20609 (N_20609,N_19618,N_19372);
nand U20610 (N_20610,N_18675,N_18340);
nor U20611 (N_20611,N_18796,N_18395);
nor U20612 (N_20612,N_18925,N_19737);
and U20613 (N_20613,N_19800,N_18819);
and U20614 (N_20614,N_18405,N_19573);
and U20615 (N_20615,N_18991,N_18445);
xnor U20616 (N_20616,N_18980,N_18504);
or U20617 (N_20617,N_19984,N_18191);
or U20618 (N_20618,N_18185,N_19262);
and U20619 (N_20619,N_19171,N_19057);
and U20620 (N_20620,N_18035,N_19580);
and U20621 (N_20621,N_18821,N_18345);
and U20622 (N_20622,N_18703,N_19668);
and U20623 (N_20623,N_19709,N_18009);
or U20624 (N_20624,N_18072,N_18228);
nand U20625 (N_20625,N_19555,N_19866);
or U20626 (N_20626,N_18369,N_19174);
nand U20627 (N_20627,N_19275,N_18501);
nor U20628 (N_20628,N_19251,N_18772);
xor U20629 (N_20629,N_18374,N_19500);
and U20630 (N_20630,N_18325,N_19271);
nand U20631 (N_20631,N_18574,N_19497);
nor U20632 (N_20632,N_19765,N_18385);
xor U20633 (N_20633,N_19549,N_19775);
xnor U20634 (N_20634,N_18934,N_18998);
nand U20635 (N_20635,N_19429,N_18014);
nor U20636 (N_20636,N_19294,N_19938);
nor U20637 (N_20637,N_18246,N_18311);
xnor U20638 (N_20638,N_19705,N_18418);
nor U20639 (N_20639,N_19558,N_18632);
nor U20640 (N_20640,N_18252,N_18341);
and U20641 (N_20641,N_18579,N_18909);
and U20642 (N_20642,N_19880,N_19210);
or U20643 (N_20643,N_19231,N_19646);
or U20644 (N_20644,N_18308,N_18413);
nor U20645 (N_20645,N_18288,N_18561);
xnor U20646 (N_20646,N_18398,N_19344);
or U20647 (N_20647,N_18716,N_18485);
nor U20648 (N_20648,N_18608,N_19465);
or U20649 (N_20649,N_19759,N_18861);
nor U20650 (N_20650,N_19408,N_19358);
or U20651 (N_20651,N_18168,N_19142);
or U20652 (N_20652,N_19777,N_19375);
and U20653 (N_20653,N_19466,N_18144);
xnor U20654 (N_20654,N_19600,N_18783);
nor U20655 (N_20655,N_19203,N_19185);
or U20656 (N_20656,N_19547,N_19762);
nor U20657 (N_20657,N_18045,N_18905);
and U20658 (N_20658,N_18674,N_18400);
or U20659 (N_20659,N_18940,N_19122);
xnor U20660 (N_20660,N_18104,N_18206);
and U20661 (N_20661,N_19774,N_19697);
nor U20662 (N_20662,N_19572,N_18872);
and U20663 (N_20663,N_18602,N_19605);
nor U20664 (N_20664,N_18854,N_18183);
xor U20665 (N_20665,N_18257,N_18791);
nor U20666 (N_20666,N_18648,N_18926);
and U20667 (N_20667,N_19037,N_18606);
or U20668 (N_20668,N_18127,N_19362);
or U20669 (N_20669,N_18061,N_18908);
and U20670 (N_20670,N_18875,N_18915);
or U20671 (N_20671,N_18251,N_18643);
xor U20672 (N_20672,N_19928,N_18163);
nor U20673 (N_20673,N_18457,N_18051);
and U20674 (N_20674,N_18572,N_18881);
and U20675 (N_20675,N_18396,N_19254);
or U20676 (N_20676,N_18438,N_18736);
nand U20677 (N_20677,N_19919,N_19172);
and U20678 (N_20678,N_19750,N_18500);
and U20679 (N_20679,N_19062,N_18033);
and U20680 (N_20680,N_19241,N_18569);
and U20681 (N_20681,N_18073,N_18454);
and U20682 (N_20682,N_18560,N_18948);
nor U20683 (N_20683,N_18999,N_19272);
xor U20684 (N_20684,N_19795,N_19188);
or U20685 (N_20685,N_18784,N_19741);
nor U20686 (N_20686,N_18850,N_19095);
nand U20687 (N_20687,N_18397,N_19754);
xor U20688 (N_20688,N_18851,N_18530);
xnor U20689 (N_20689,N_19717,N_18990);
nand U20690 (N_20690,N_18649,N_18890);
nand U20691 (N_20691,N_19186,N_18620);
or U20692 (N_20692,N_19864,N_19582);
nor U20693 (N_20693,N_19490,N_19877);
nor U20694 (N_20694,N_18372,N_18576);
and U20695 (N_20695,N_19412,N_18535);
nor U20696 (N_20696,N_18906,N_19693);
and U20697 (N_20697,N_18864,N_19151);
nor U20698 (N_20698,N_18830,N_18558);
and U20699 (N_20699,N_19634,N_19712);
xor U20700 (N_20700,N_19838,N_18464);
or U20701 (N_20701,N_18523,N_19265);
nand U20702 (N_20702,N_18469,N_18534);
xnor U20703 (N_20703,N_19630,N_19130);
nand U20704 (N_20704,N_18896,N_19913);
nor U20705 (N_20705,N_18658,N_19404);
nor U20706 (N_20706,N_18351,N_18335);
and U20707 (N_20707,N_19099,N_18443);
nand U20708 (N_20708,N_18295,N_19109);
and U20709 (N_20709,N_18328,N_18695);
or U20710 (N_20710,N_19537,N_18730);
and U20711 (N_20711,N_18706,N_18595);
xnor U20712 (N_20712,N_19173,N_18432);
nor U20713 (N_20713,N_18843,N_18235);
or U20714 (N_20714,N_19248,N_18612);
or U20715 (N_20715,N_19845,N_18853);
and U20716 (N_20716,N_18399,N_18032);
or U20717 (N_20717,N_19846,N_19015);
and U20718 (N_20718,N_19548,N_18712);
nand U20719 (N_20719,N_18148,N_19639);
and U20720 (N_20720,N_19888,N_18954);
xnor U20721 (N_20721,N_19379,N_19990);
xor U20722 (N_20722,N_19945,N_18371);
nand U20723 (N_20723,N_18723,N_19326);
or U20724 (N_20724,N_18496,N_18505);
xnor U20725 (N_20725,N_18922,N_19107);
xor U20726 (N_20726,N_19484,N_19162);
xor U20727 (N_20727,N_19261,N_18498);
xor U20728 (N_20728,N_19552,N_18195);
nand U20729 (N_20729,N_19472,N_18546);
nand U20730 (N_20730,N_18877,N_19452);
or U20731 (N_20731,N_19315,N_18318);
and U20732 (N_20732,N_19504,N_19259);
and U20733 (N_20733,N_19949,N_19268);
or U20734 (N_20734,N_18154,N_19780);
and U20735 (N_20735,N_19046,N_19385);
or U20736 (N_20736,N_19486,N_18732);
and U20737 (N_20737,N_18714,N_19776);
nor U20738 (N_20738,N_19808,N_19094);
nor U20739 (N_20739,N_18450,N_19125);
nand U20740 (N_20740,N_18431,N_19532);
nor U20741 (N_20741,N_19621,N_19652);
xnor U20742 (N_20742,N_19974,N_18549);
and U20743 (N_20743,N_18945,N_18357);
and U20744 (N_20744,N_19337,N_18289);
or U20745 (N_20745,N_18859,N_19493);
nand U20746 (N_20746,N_19239,N_18741);
or U20747 (N_20747,N_19749,N_18363);
nor U20748 (N_20748,N_18903,N_19055);
nand U20749 (N_20749,N_18779,N_18075);
and U20750 (N_20750,N_19341,N_18425);
and U20751 (N_20751,N_19439,N_19474);
xor U20752 (N_20752,N_18673,N_18379);
nand U20753 (N_20753,N_18200,N_18059);
and U20754 (N_20754,N_18789,N_19249);
or U20755 (N_20755,N_18436,N_18492);
xnor U20756 (N_20756,N_18084,N_19096);
or U20757 (N_20757,N_18519,N_19207);
nand U20758 (N_20758,N_19801,N_18198);
and U20759 (N_20759,N_18477,N_19982);
and U20760 (N_20760,N_18427,N_19308);
nor U20761 (N_20761,N_18196,N_18810);
nand U20762 (N_20762,N_18394,N_18039);
xnor U20763 (N_20763,N_18189,N_18771);
or U20764 (N_20764,N_19215,N_18609);
xnor U20765 (N_20765,N_19959,N_18942);
or U20766 (N_20766,N_18420,N_18044);
xnor U20767 (N_20767,N_19886,N_18946);
or U20768 (N_20768,N_19320,N_19299);
nand U20769 (N_20769,N_18751,N_19035);
and U20770 (N_20770,N_19325,N_18447);
nand U20771 (N_20771,N_18768,N_18069);
or U20772 (N_20772,N_18426,N_18793);
or U20773 (N_20773,N_18935,N_19953);
and U20774 (N_20774,N_19923,N_18691);
xor U20775 (N_20775,N_19085,N_18297);
xor U20776 (N_20776,N_18476,N_19516);
and U20777 (N_20777,N_18022,N_19672);
nand U20778 (N_20778,N_18143,N_19769);
or U20779 (N_20779,N_19491,N_19042);
nor U20780 (N_20780,N_18157,N_19661);
xor U20781 (N_20781,N_19298,N_19383);
xor U20782 (N_20782,N_19387,N_19875);
and U20783 (N_20783,N_18057,N_19671);
nor U20784 (N_20784,N_18490,N_18797);
xor U20785 (N_20785,N_18314,N_18253);
nand U20786 (N_20786,N_18381,N_18805);
nor U20787 (N_20787,N_18139,N_19000);
and U20788 (N_20788,N_18563,N_19807);
nand U20789 (N_20789,N_18884,N_18870);
nand U20790 (N_20790,N_18358,N_19247);
nand U20791 (N_20791,N_19655,N_18137);
nor U20792 (N_20792,N_19604,N_19806);
nand U20793 (N_20793,N_19440,N_19542);
xor U20794 (N_20794,N_18667,N_19078);
and U20795 (N_20795,N_18294,N_19863);
nand U20796 (N_20796,N_18280,N_18885);
nor U20797 (N_20797,N_18750,N_18619);
nor U20798 (N_20798,N_18391,N_18773);
or U20799 (N_20799,N_18710,N_19704);
nor U20800 (N_20800,N_18681,N_19583);
nand U20801 (N_20801,N_18077,N_18586);
xnor U20802 (N_20802,N_19636,N_18149);
nand U20803 (N_20803,N_18090,N_19701);
nor U20804 (N_20804,N_19543,N_19054);
xnor U20805 (N_20805,N_18831,N_19508);
nand U20806 (N_20806,N_18164,N_19026);
nand U20807 (N_20807,N_19169,N_19798);
nand U20808 (N_20808,N_18264,N_19822);
nand U20809 (N_20809,N_18046,N_18120);
nand U20810 (N_20810,N_18742,N_19327);
and U20811 (N_20811,N_18282,N_18522);
nor U20812 (N_20812,N_19002,N_18040);
nand U20813 (N_20813,N_18898,N_18008);
and U20814 (N_20814,N_18165,N_19016);
or U20815 (N_20815,N_19900,N_19657);
or U20816 (N_20816,N_18565,N_19175);
nor U20817 (N_20817,N_19023,N_19263);
nand U20818 (N_20818,N_19993,N_18230);
nor U20819 (N_20819,N_19183,N_19598);
xnor U20820 (N_20820,N_18441,N_18918);
nor U20821 (N_20821,N_18944,N_19321);
and U20822 (N_20822,N_18947,N_18652);
nand U20823 (N_20823,N_19964,N_19068);
xor U20824 (N_20824,N_18618,N_18421);
nor U20825 (N_20825,N_18962,N_19736);
or U20826 (N_20826,N_19220,N_19153);
xnor U20827 (N_20827,N_18663,N_18416);
nor U20828 (N_20828,N_18408,N_18517);
nand U20829 (N_20829,N_19475,N_19766);
or U20830 (N_20830,N_19616,N_18907);
or U20831 (N_20831,N_19073,N_19038);
and U20832 (N_20832,N_19876,N_18770);
or U20833 (N_20833,N_19506,N_18547);
nor U20834 (N_20834,N_19201,N_18641);
xor U20835 (N_20835,N_18151,N_19424);
xnor U20836 (N_20836,N_18815,N_18912);
and U20837 (N_20837,N_18284,N_19436);
or U20838 (N_20838,N_19640,N_18894);
and U20839 (N_20839,N_19252,N_18055);
xor U20840 (N_20840,N_18190,N_19980);
and U20841 (N_20841,N_19597,N_19349);
or U20842 (N_20842,N_19013,N_19872);
nand U20843 (N_20843,N_19908,N_19305);
nand U20844 (N_20844,N_18804,N_18971);
and U20845 (N_20845,N_19033,N_18448);
nor U20846 (N_20846,N_18880,N_19230);
and U20847 (N_20847,N_18801,N_18232);
nor U20848 (N_20848,N_19738,N_18983);
and U20849 (N_20849,N_18030,N_19363);
and U20850 (N_20850,N_18724,N_19519);
and U20851 (N_20851,N_19783,N_19927);
or U20852 (N_20852,N_19001,N_19578);
xor U20853 (N_20853,N_19150,N_19030);
nand U20854 (N_20854,N_18142,N_19279);
nor U20855 (N_20855,N_19857,N_19397);
or U20856 (N_20856,N_18631,N_19817);
xnor U20857 (N_20857,N_18429,N_19615);
xnor U20858 (N_20858,N_19256,N_18670);
nor U20859 (N_20859,N_18499,N_19853);
and U20860 (N_20860,N_19599,N_19787);
or U20861 (N_20861,N_18708,N_19551);
nor U20862 (N_20862,N_18655,N_19730);
and U20863 (N_20863,N_19330,N_19954);
nand U20864 (N_20864,N_19523,N_18509);
or U20865 (N_20865,N_18683,N_19859);
or U20866 (N_20866,N_19733,N_18600);
nand U20867 (N_20867,N_19090,N_19670);
nor U20868 (N_20868,N_18001,N_18133);
or U20869 (N_20869,N_18170,N_19978);
nor U20870 (N_20870,N_19018,N_18052);
or U20871 (N_20871,N_18292,N_18812);
xnor U20872 (N_20872,N_19638,N_19223);
or U20873 (N_20873,N_18320,N_18322);
nand U20874 (N_20874,N_19368,N_19902);
and U20875 (N_20875,N_19747,N_19196);
xor U20876 (N_20876,N_18124,N_18686);
nand U20877 (N_20877,N_18863,N_19405);
or U20878 (N_20878,N_19032,N_18346);
nor U20879 (N_20879,N_19064,N_19355);
nand U20880 (N_20880,N_18799,N_18869);
nor U20881 (N_20881,N_18112,N_19168);
nand U20882 (N_20882,N_19620,N_18603);
and U20883 (N_20883,N_18063,N_19245);
xor U20884 (N_20884,N_18920,N_19060);
xnor U20885 (N_20885,N_19270,N_18131);
or U20886 (N_20886,N_19287,N_18210);
nand U20887 (N_20887,N_19528,N_18752);
or U20888 (N_20888,N_18437,N_18749);
and U20889 (N_20889,N_19950,N_18248);
xnor U20890 (N_20890,N_18705,N_18241);
and U20891 (N_20891,N_19607,N_18296);
nand U20892 (N_20892,N_19282,N_19303);
nand U20893 (N_20893,N_18243,N_19071);
and U20894 (N_20894,N_18671,N_19649);
and U20895 (N_20895,N_19283,N_18270);
or U20896 (N_20896,N_18786,N_19105);
xnor U20897 (N_20897,N_19726,N_19612);
and U20898 (N_20898,N_18939,N_19660);
xnor U20899 (N_20899,N_19796,N_18887);
or U20900 (N_20900,N_18753,N_18223);
xor U20901 (N_20901,N_19818,N_18997);
nand U20902 (N_20902,N_18011,N_19077);
xor U20903 (N_20903,N_19714,N_19225);
xnor U20904 (N_20904,N_19176,N_19021);
xor U20905 (N_20905,N_18701,N_19102);
xnor U20906 (N_20906,N_18512,N_19205);
and U20907 (N_20907,N_19208,N_18313);
nor U20908 (N_20908,N_19929,N_18181);
nand U20909 (N_20909,N_18348,N_18109);
xor U20910 (N_20910,N_18611,N_19541);
and U20911 (N_20911,N_18203,N_19957);
and U20912 (N_20912,N_18242,N_18430);
nand U20913 (N_20913,N_19901,N_18386);
xnor U20914 (N_20914,N_18913,N_19823);
or U20915 (N_20915,N_19626,N_18219);
nor U20916 (N_20916,N_19561,N_19290);
nand U20917 (N_20917,N_18272,N_18054);
xor U20918 (N_20918,N_18888,N_18038);
xnor U20919 (N_20919,N_19891,N_18299);
and U20920 (N_20920,N_18497,N_18924);
nand U20921 (N_20921,N_19721,N_18644);
or U20922 (N_20922,N_19088,N_18748);
nor U20923 (N_20923,N_19645,N_18166);
and U20924 (N_20924,N_19008,N_18757);
nor U20925 (N_20925,N_18626,N_19595);
xor U20926 (N_20926,N_18456,N_18814);
nor U20927 (N_20927,N_19939,N_19049);
and U20928 (N_20928,N_18596,N_19266);
and U20929 (N_20929,N_19556,N_19719);
nand U20930 (N_20930,N_19840,N_18943);
or U20931 (N_20931,N_19534,N_18867);
and U20932 (N_20932,N_18790,N_18975);
xor U20933 (N_20933,N_18043,N_18245);
nand U20934 (N_20934,N_19480,N_18666);
xnor U20935 (N_20935,N_18473,N_18458);
nor U20936 (N_20936,N_19909,N_19711);
and U20937 (N_20937,N_19148,N_19768);
or U20938 (N_20938,N_19890,N_18089);
nor U20939 (N_20939,N_19734,N_19229);
nand U20940 (N_20940,N_18981,N_19025);
or U20941 (N_20941,N_19922,N_19861);
or U20942 (N_20942,N_19083,N_18258);
or U20943 (N_20943,N_19673,N_19868);
nor U20944 (N_20944,N_18049,N_18095);
xnor U20945 (N_20945,N_18002,N_18409);
nand U20946 (N_20946,N_18734,N_18419);
and U20947 (N_20947,N_19269,N_19010);
or U20948 (N_20948,N_19006,N_18871);
nor U20949 (N_20949,N_19946,N_19014);
nand U20950 (N_20950,N_19684,N_19963);
nor U20951 (N_20951,N_19557,N_19988);
nor U20952 (N_20952,N_19463,N_19365);
nand U20953 (N_20953,N_19996,N_18005);
nand U20954 (N_20954,N_18136,N_19758);
nor U20955 (N_20955,N_18468,N_19066);
nand U20956 (N_20956,N_19906,N_19535);
or U20957 (N_20957,N_19513,N_19509);
xor U20958 (N_20958,N_19182,N_18470);
nand U20959 (N_20959,N_18739,N_19373);
nor U20960 (N_20960,N_18950,N_18442);
xor U20961 (N_20961,N_18117,N_19179);
nor U20962 (N_20962,N_18507,N_18919);
nor U20963 (N_20963,N_18614,N_18446);
nor U20964 (N_20964,N_19914,N_18176);
and U20965 (N_20965,N_18852,N_19044);
nor U20966 (N_20966,N_18122,N_18792);
or U20967 (N_20967,N_19100,N_19729);
nor U20968 (N_20968,N_18216,N_18562);
nand U20969 (N_20969,N_19461,N_18587);
nand U20970 (N_20970,N_19576,N_19492);
nor U20971 (N_20971,N_18583,N_18577);
and U20972 (N_20972,N_19333,N_19662);
or U20973 (N_20973,N_18103,N_19410);
xnor U20974 (N_20974,N_18963,N_19459);
or U20975 (N_20975,N_19686,N_19009);
and U20976 (N_20976,N_19285,N_18287);
and U20977 (N_20977,N_19587,N_18542);
nor U20978 (N_20978,N_19690,N_19560);
xor U20979 (N_20979,N_18849,N_19091);
nor U20980 (N_20980,N_19437,N_19428);
or U20981 (N_20981,N_19120,N_19687);
nor U20982 (N_20982,N_18481,N_19764);
and U20983 (N_20983,N_18847,N_18518);
xnor U20984 (N_20984,N_18727,N_18172);
xnor U20985 (N_20985,N_19836,N_18585);
and U20986 (N_20986,N_19260,N_18895);
nand U20987 (N_20987,N_18883,N_18337);
nor U20988 (N_20988,N_19663,N_19113);
or U20989 (N_20989,N_19667,N_18184);
nor U20990 (N_20990,N_18238,N_18085);
nor U20991 (N_20991,N_18933,N_19413);
nand U20992 (N_20992,N_18053,N_18822);
xnor U20993 (N_20993,N_19559,N_18720);
xor U20994 (N_20994,N_19427,N_18989);
or U20995 (N_20995,N_18746,N_19250);
xor U20996 (N_20996,N_18639,N_19228);
and U20997 (N_20997,N_19852,N_19659);
and U20998 (N_20998,N_19911,N_19971);
nor U20999 (N_20999,N_19926,N_18617);
or U21000 (N_21000,N_19031,N_18146);
xor U21001 (N_21001,N_19946,N_19885);
nor U21002 (N_21002,N_18026,N_19225);
xor U21003 (N_21003,N_19547,N_18018);
and U21004 (N_21004,N_18146,N_18862);
xnor U21005 (N_21005,N_18334,N_19548);
nand U21006 (N_21006,N_18090,N_19363);
nand U21007 (N_21007,N_18138,N_19077);
nand U21008 (N_21008,N_18901,N_18048);
nor U21009 (N_21009,N_18878,N_19777);
or U21010 (N_21010,N_19459,N_19642);
nand U21011 (N_21011,N_18984,N_19073);
or U21012 (N_21012,N_19002,N_19761);
nand U21013 (N_21013,N_19817,N_19640);
xnor U21014 (N_21014,N_19038,N_19706);
nor U21015 (N_21015,N_18602,N_19456);
nand U21016 (N_21016,N_19354,N_19763);
or U21017 (N_21017,N_18709,N_18992);
nand U21018 (N_21018,N_19753,N_18888);
or U21019 (N_21019,N_19578,N_18487);
nor U21020 (N_21020,N_19001,N_18142);
nor U21021 (N_21021,N_18146,N_19620);
nand U21022 (N_21022,N_19376,N_18254);
or U21023 (N_21023,N_18336,N_18803);
or U21024 (N_21024,N_18805,N_18720);
nor U21025 (N_21025,N_18394,N_18649);
nor U21026 (N_21026,N_18135,N_18566);
nor U21027 (N_21027,N_18626,N_18983);
nand U21028 (N_21028,N_19939,N_18795);
nor U21029 (N_21029,N_19128,N_19809);
and U21030 (N_21030,N_18279,N_19018);
nor U21031 (N_21031,N_18261,N_19084);
nand U21032 (N_21032,N_18470,N_18034);
xor U21033 (N_21033,N_18760,N_18396);
xnor U21034 (N_21034,N_19778,N_19463);
or U21035 (N_21035,N_19179,N_18996);
nand U21036 (N_21036,N_19499,N_19588);
nand U21037 (N_21037,N_18711,N_18522);
nand U21038 (N_21038,N_19498,N_19914);
or U21039 (N_21039,N_19176,N_18257);
nor U21040 (N_21040,N_19355,N_19886);
and U21041 (N_21041,N_19334,N_19861);
and U21042 (N_21042,N_18498,N_18336);
xnor U21043 (N_21043,N_19504,N_19127);
and U21044 (N_21044,N_18760,N_18022);
and U21045 (N_21045,N_18338,N_18957);
nand U21046 (N_21046,N_18222,N_19302);
nand U21047 (N_21047,N_18497,N_19012);
nor U21048 (N_21048,N_18237,N_19770);
or U21049 (N_21049,N_18463,N_18950);
or U21050 (N_21050,N_18900,N_19476);
nor U21051 (N_21051,N_19787,N_18362);
nand U21052 (N_21052,N_19524,N_19839);
nor U21053 (N_21053,N_19169,N_18366);
or U21054 (N_21054,N_18193,N_19829);
xnor U21055 (N_21055,N_18109,N_18392);
nand U21056 (N_21056,N_18447,N_18846);
or U21057 (N_21057,N_19832,N_19205);
and U21058 (N_21058,N_18601,N_19152);
or U21059 (N_21059,N_19722,N_18130);
and U21060 (N_21060,N_18010,N_18714);
nor U21061 (N_21061,N_19484,N_19034);
nand U21062 (N_21062,N_19010,N_19654);
xnor U21063 (N_21063,N_18282,N_18737);
and U21064 (N_21064,N_18005,N_19008);
or U21065 (N_21065,N_18571,N_19899);
nand U21066 (N_21066,N_19362,N_18650);
xnor U21067 (N_21067,N_19954,N_19590);
or U21068 (N_21068,N_18440,N_18365);
and U21069 (N_21069,N_19257,N_19370);
nand U21070 (N_21070,N_19727,N_18232);
nor U21071 (N_21071,N_19305,N_19171);
or U21072 (N_21072,N_18935,N_19832);
nand U21073 (N_21073,N_18935,N_19215);
and U21074 (N_21074,N_19393,N_19364);
nor U21075 (N_21075,N_19390,N_19653);
nand U21076 (N_21076,N_19025,N_18785);
and U21077 (N_21077,N_19216,N_19219);
nor U21078 (N_21078,N_19537,N_19320);
and U21079 (N_21079,N_18022,N_18604);
xor U21080 (N_21080,N_19695,N_18733);
nand U21081 (N_21081,N_18949,N_19610);
nand U21082 (N_21082,N_19472,N_18415);
and U21083 (N_21083,N_18178,N_19476);
and U21084 (N_21084,N_19085,N_18394);
xnor U21085 (N_21085,N_19879,N_19088);
or U21086 (N_21086,N_19606,N_18608);
xor U21087 (N_21087,N_18646,N_18458);
nor U21088 (N_21088,N_18323,N_19553);
nand U21089 (N_21089,N_18403,N_19309);
nor U21090 (N_21090,N_19895,N_19678);
or U21091 (N_21091,N_19854,N_19578);
nor U21092 (N_21092,N_19102,N_19159);
nor U21093 (N_21093,N_18427,N_19714);
nor U21094 (N_21094,N_19197,N_18068);
and U21095 (N_21095,N_19935,N_19132);
nand U21096 (N_21096,N_18870,N_18335);
xnor U21097 (N_21097,N_19639,N_19446);
nand U21098 (N_21098,N_18025,N_19998);
and U21099 (N_21099,N_18846,N_18940);
nand U21100 (N_21100,N_19689,N_18711);
nor U21101 (N_21101,N_19969,N_19866);
and U21102 (N_21102,N_19658,N_19145);
and U21103 (N_21103,N_19278,N_19404);
or U21104 (N_21104,N_18954,N_19297);
and U21105 (N_21105,N_18418,N_19501);
or U21106 (N_21106,N_19616,N_19173);
nor U21107 (N_21107,N_19549,N_19332);
and U21108 (N_21108,N_19780,N_18014);
or U21109 (N_21109,N_18347,N_18508);
and U21110 (N_21110,N_18433,N_19451);
and U21111 (N_21111,N_18096,N_19851);
or U21112 (N_21112,N_18058,N_19788);
and U21113 (N_21113,N_19173,N_18293);
and U21114 (N_21114,N_18868,N_19927);
nor U21115 (N_21115,N_18257,N_18623);
nand U21116 (N_21116,N_18326,N_18300);
nor U21117 (N_21117,N_18283,N_18512);
nand U21118 (N_21118,N_19767,N_18835);
and U21119 (N_21119,N_19030,N_19533);
nand U21120 (N_21120,N_19979,N_18769);
and U21121 (N_21121,N_19901,N_18669);
and U21122 (N_21122,N_18238,N_18526);
xnor U21123 (N_21123,N_19861,N_19548);
nand U21124 (N_21124,N_19118,N_19198);
or U21125 (N_21125,N_19208,N_18718);
nor U21126 (N_21126,N_18793,N_19164);
xnor U21127 (N_21127,N_18806,N_18013);
nand U21128 (N_21128,N_19935,N_19790);
and U21129 (N_21129,N_19615,N_18530);
nor U21130 (N_21130,N_18056,N_18370);
nand U21131 (N_21131,N_18099,N_19970);
xnor U21132 (N_21132,N_19778,N_19276);
xnor U21133 (N_21133,N_19662,N_18218);
nand U21134 (N_21134,N_19075,N_19632);
or U21135 (N_21135,N_19986,N_18799);
or U21136 (N_21136,N_19087,N_18436);
nand U21137 (N_21137,N_18524,N_18431);
nand U21138 (N_21138,N_18546,N_18426);
nand U21139 (N_21139,N_19065,N_19398);
nor U21140 (N_21140,N_18956,N_19415);
or U21141 (N_21141,N_18043,N_19056);
xnor U21142 (N_21142,N_18146,N_19114);
and U21143 (N_21143,N_18374,N_19361);
or U21144 (N_21144,N_19039,N_18733);
nand U21145 (N_21145,N_19711,N_18617);
and U21146 (N_21146,N_18357,N_18806);
xnor U21147 (N_21147,N_19770,N_18638);
or U21148 (N_21148,N_18356,N_19028);
nand U21149 (N_21149,N_18263,N_18180);
or U21150 (N_21150,N_19235,N_19892);
nand U21151 (N_21151,N_19551,N_19370);
xor U21152 (N_21152,N_18563,N_18305);
and U21153 (N_21153,N_19442,N_19493);
or U21154 (N_21154,N_19112,N_19517);
nor U21155 (N_21155,N_18860,N_18145);
nor U21156 (N_21156,N_19747,N_18655);
nor U21157 (N_21157,N_18124,N_19101);
and U21158 (N_21158,N_19688,N_18798);
nor U21159 (N_21159,N_18440,N_18893);
xnor U21160 (N_21160,N_18374,N_18089);
nand U21161 (N_21161,N_19181,N_18735);
nor U21162 (N_21162,N_19618,N_19690);
nor U21163 (N_21163,N_18601,N_18485);
nand U21164 (N_21164,N_18459,N_19348);
xnor U21165 (N_21165,N_18722,N_18685);
nor U21166 (N_21166,N_19684,N_18039);
or U21167 (N_21167,N_19887,N_19746);
nand U21168 (N_21168,N_19674,N_19532);
nand U21169 (N_21169,N_18653,N_18119);
nor U21170 (N_21170,N_18446,N_18134);
nor U21171 (N_21171,N_18999,N_18318);
and U21172 (N_21172,N_18460,N_18820);
nand U21173 (N_21173,N_18396,N_19068);
and U21174 (N_21174,N_18338,N_18312);
nor U21175 (N_21175,N_18081,N_18685);
or U21176 (N_21176,N_19589,N_18887);
or U21177 (N_21177,N_19397,N_18258);
and U21178 (N_21178,N_18455,N_18139);
nand U21179 (N_21179,N_18437,N_19434);
xnor U21180 (N_21180,N_19342,N_18667);
and U21181 (N_21181,N_19554,N_18610);
nand U21182 (N_21182,N_19470,N_18991);
and U21183 (N_21183,N_18404,N_18488);
nand U21184 (N_21184,N_18231,N_19285);
nor U21185 (N_21185,N_18898,N_19581);
nand U21186 (N_21186,N_19766,N_18446);
and U21187 (N_21187,N_18334,N_19091);
or U21188 (N_21188,N_19261,N_19631);
nor U21189 (N_21189,N_19428,N_19367);
xnor U21190 (N_21190,N_19177,N_19595);
xor U21191 (N_21191,N_18424,N_19595);
nand U21192 (N_21192,N_18799,N_19434);
xnor U21193 (N_21193,N_18920,N_19676);
xnor U21194 (N_21194,N_19984,N_19760);
and U21195 (N_21195,N_18646,N_19531);
xnor U21196 (N_21196,N_18290,N_18543);
and U21197 (N_21197,N_19442,N_18618);
nand U21198 (N_21198,N_19470,N_19854);
and U21199 (N_21199,N_18283,N_19168);
or U21200 (N_21200,N_18691,N_18560);
and U21201 (N_21201,N_19906,N_18300);
and U21202 (N_21202,N_19577,N_19695);
or U21203 (N_21203,N_18237,N_19622);
nand U21204 (N_21204,N_18777,N_18203);
nor U21205 (N_21205,N_18291,N_18104);
xor U21206 (N_21206,N_18164,N_19873);
or U21207 (N_21207,N_18315,N_18402);
nor U21208 (N_21208,N_18395,N_19468);
nand U21209 (N_21209,N_19886,N_19032);
nor U21210 (N_21210,N_19884,N_18406);
xnor U21211 (N_21211,N_19779,N_18777);
nand U21212 (N_21212,N_18787,N_18677);
nor U21213 (N_21213,N_18944,N_19595);
and U21214 (N_21214,N_19912,N_19832);
and U21215 (N_21215,N_19856,N_18231);
xnor U21216 (N_21216,N_19753,N_19674);
or U21217 (N_21217,N_19213,N_18713);
or U21218 (N_21218,N_18046,N_18443);
nor U21219 (N_21219,N_18763,N_18419);
nand U21220 (N_21220,N_19336,N_18377);
nor U21221 (N_21221,N_19156,N_18602);
nor U21222 (N_21222,N_18142,N_18579);
nor U21223 (N_21223,N_19724,N_19198);
xor U21224 (N_21224,N_19451,N_19598);
nand U21225 (N_21225,N_18393,N_19043);
nor U21226 (N_21226,N_18864,N_19283);
xnor U21227 (N_21227,N_19819,N_18196);
xnor U21228 (N_21228,N_19912,N_19774);
and U21229 (N_21229,N_19411,N_18133);
and U21230 (N_21230,N_19494,N_19484);
or U21231 (N_21231,N_18821,N_18458);
nand U21232 (N_21232,N_18532,N_19787);
and U21233 (N_21233,N_19821,N_19454);
and U21234 (N_21234,N_18660,N_19992);
and U21235 (N_21235,N_18305,N_19308);
nor U21236 (N_21236,N_18004,N_19141);
and U21237 (N_21237,N_18280,N_19086);
nor U21238 (N_21238,N_18411,N_19303);
nor U21239 (N_21239,N_18780,N_18974);
nand U21240 (N_21240,N_18949,N_18704);
and U21241 (N_21241,N_19183,N_18948);
or U21242 (N_21242,N_18897,N_19144);
and U21243 (N_21243,N_19844,N_19371);
and U21244 (N_21244,N_19772,N_18681);
nor U21245 (N_21245,N_18561,N_18488);
xor U21246 (N_21246,N_19041,N_18547);
nor U21247 (N_21247,N_18684,N_19486);
nor U21248 (N_21248,N_19774,N_18802);
nand U21249 (N_21249,N_18691,N_18930);
and U21250 (N_21250,N_18501,N_18289);
and U21251 (N_21251,N_18743,N_19038);
or U21252 (N_21252,N_18287,N_18000);
nor U21253 (N_21253,N_18158,N_18880);
xnor U21254 (N_21254,N_18064,N_18555);
and U21255 (N_21255,N_18762,N_18346);
and U21256 (N_21256,N_18871,N_18362);
nor U21257 (N_21257,N_18342,N_18496);
or U21258 (N_21258,N_18829,N_18213);
xnor U21259 (N_21259,N_19550,N_18545);
and U21260 (N_21260,N_18623,N_19433);
or U21261 (N_21261,N_19338,N_18091);
and U21262 (N_21262,N_19411,N_19661);
or U21263 (N_21263,N_18489,N_19840);
and U21264 (N_21264,N_19800,N_19178);
nor U21265 (N_21265,N_18525,N_18284);
nor U21266 (N_21266,N_19088,N_19241);
nor U21267 (N_21267,N_18690,N_19115);
nand U21268 (N_21268,N_18088,N_18369);
nor U21269 (N_21269,N_18926,N_19626);
and U21270 (N_21270,N_18978,N_18272);
or U21271 (N_21271,N_18125,N_19621);
nor U21272 (N_21272,N_19743,N_18147);
nor U21273 (N_21273,N_19246,N_18725);
and U21274 (N_21274,N_18072,N_18815);
and U21275 (N_21275,N_19363,N_19625);
xor U21276 (N_21276,N_19359,N_18829);
xnor U21277 (N_21277,N_18664,N_19296);
xor U21278 (N_21278,N_19090,N_19216);
nand U21279 (N_21279,N_19722,N_18496);
and U21280 (N_21280,N_18448,N_19491);
or U21281 (N_21281,N_19639,N_19538);
nor U21282 (N_21282,N_18012,N_19235);
nand U21283 (N_21283,N_18747,N_19864);
or U21284 (N_21284,N_19794,N_19494);
nand U21285 (N_21285,N_19772,N_18413);
nor U21286 (N_21286,N_18892,N_18201);
nand U21287 (N_21287,N_18121,N_19192);
or U21288 (N_21288,N_18628,N_19633);
xor U21289 (N_21289,N_18560,N_18261);
xor U21290 (N_21290,N_19881,N_19139);
or U21291 (N_21291,N_19841,N_19221);
xor U21292 (N_21292,N_19050,N_18591);
or U21293 (N_21293,N_18699,N_18092);
xor U21294 (N_21294,N_18948,N_19411);
nor U21295 (N_21295,N_19710,N_19454);
nand U21296 (N_21296,N_19768,N_19708);
and U21297 (N_21297,N_18529,N_19437);
nand U21298 (N_21298,N_18409,N_18550);
xnor U21299 (N_21299,N_18290,N_19379);
or U21300 (N_21300,N_18248,N_18285);
nor U21301 (N_21301,N_18145,N_19735);
and U21302 (N_21302,N_19395,N_19322);
nand U21303 (N_21303,N_19997,N_19097);
nand U21304 (N_21304,N_18608,N_19875);
nand U21305 (N_21305,N_19814,N_19187);
nor U21306 (N_21306,N_19845,N_19470);
nor U21307 (N_21307,N_19658,N_19407);
xnor U21308 (N_21308,N_19930,N_18099);
xor U21309 (N_21309,N_18420,N_19608);
nand U21310 (N_21310,N_18714,N_18891);
or U21311 (N_21311,N_19096,N_18425);
xor U21312 (N_21312,N_18845,N_19035);
and U21313 (N_21313,N_18698,N_18225);
and U21314 (N_21314,N_19231,N_19423);
and U21315 (N_21315,N_19268,N_18090);
and U21316 (N_21316,N_19131,N_18975);
nand U21317 (N_21317,N_18392,N_18063);
xor U21318 (N_21318,N_18650,N_19944);
or U21319 (N_21319,N_18832,N_19837);
nand U21320 (N_21320,N_19526,N_19320);
or U21321 (N_21321,N_18846,N_19820);
or U21322 (N_21322,N_18277,N_19708);
xor U21323 (N_21323,N_19625,N_18070);
xor U21324 (N_21324,N_19848,N_19181);
nand U21325 (N_21325,N_18944,N_19469);
xnor U21326 (N_21326,N_18156,N_18898);
xor U21327 (N_21327,N_18747,N_18464);
xor U21328 (N_21328,N_18708,N_19931);
nand U21329 (N_21329,N_19084,N_18656);
and U21330 (N_21330,N_18748,N_19000);
or U21331 (N_21331,N_19389,N_18787);
or U21332 (N_21332,N_19794,N_18086);
and U21333 (N_21333,N_18437,N_19582);
and U21334 (N_21334,N_19489,N_19726);
nand U21335 (N_21335,N_19644,N_19393);
or U21336 (N_21336,N_19378,N_19171);
xor U21337 (N_21337,N_18645,N_19604);
nand U21338 (N_21338,N_18791,N_18370);
xnor U21339 (N_21339,N_18324,N_18095);
or U21340 (N_21340,N_19632,N_18300);
nand U21341 (N_21341,N_19919,N_19260);
or U21342 (N_21342,N_18173,N_18700);
nor U21343 (N_21343,N_18091,N_18329);
or U21344 (N_21344,N_19635,N_18727);
and U21345 (N_21345,N_19231,N_19116);
xor U21346 (N_21346,N_19802,N_18557);
and U21347 (N_21347,N_18430,N_18311);
or U21348 (N_21348,N_19982,N_19077);
nand U21349 (N_21349,N_18435,N_18941);
or U21350 (N_21350,N_18754,N_19809);
and U21351 (N_21351,N_19283,N_19183);
or U21352 (N_21352,N_19401,N_19744);
or U21353 (N_21353,N_19810,N_19100);
and U21354 (N_21354,N_18296,N_18563);
nand U21355 (N_21355,N_19797,N_19796);
nand U21356 (N_21356,N_19236,N_19589);
nor U21357 (N_21357,N_19714,N_18288);
nor U21358 (N_21358,N_18732,N_19495);
nand U21359 (N_21359,N_19517,N_19878);
nand U21360 (N_21360,N_19593,N_19654);
nand U21361 (N_21361,N_18398,N_19285);
and U21362 (N_21362,N_18807,N_18936);
or U21363 (N_21363,N_18929,N_19155);
nand U21364 (N_21364,N_19875,N_18430);
nand U21365 (N_21365,N_19123,N_19124);
xnor U21366 (N_21366,N_18905,N_19657);
nand U21367 (N_21367,N_19704,N_19989);
nor U21368 (N_21368,N_19575,N_18226);
xnor U21369 (N_21369,N_19002,N_19751);
nand U21370 (N_21370,N_19783,N_19470);
nand U21371 (N_21371,N_19791,N_19194);
and U21372 (N_21372,N_18155,N_18390);
nand U21373 (N_21373,N_19818,N_18042);
and U21374 (N_21374,N_19628,N_19780);
xnor U21375 (N_21375,N_19863,N_19713);
xor U21376 (N_21376,N_18184,N_18354);
nor U21377 (N_21377,N_18314,N_19923);
nand U21378 (N_21378,N_19294,N_18482);
nand U21379 (N_21379,N_18558,N_19839);
or U21380 (N_21380,N_18281,N_19561);
and U21381 (N_21381,N_18389,N_18276);
and U21382 (N_21382,N_18425,N_18290);
xor U21383 (N_21383,N_19360,N_19263);
nand U21384 (N_21384,N_19280,N_18482);
xor U21385 (N_21385,N_18550,N_19484);
nor U21386 (N_21386,N_19760,N_19061);
and U21387 (N_21387,N_18238,N_18914);
or U21388 (N_21388,N_19234,N_18329);
xnor U21389 (N_21389,N_18483,N_19125);
nand U21390 (N_21390,N_18302,N_19601);
xor U21391 (N_21391,N_18062,N_19765);
and U21392 (N_21392,N_18907,N_18722);
nand U21393 (N_21393,N_19458,N_18692);
xor U21394 (N_21394,N_18028,N_19043);
xnor U21395 (N_21395,N_19485,N_19393);
and U21396 (N_21396,N_18876,N_19740);
and U21397 (N_21397,N_19974,N_18779);
nand U21398 (N_21398,N_18749,N_18149);
nor U21399 (N_21399,N_19387,N_19539);
xnor U21400 (N_21400,N_18341,N_18321);
xor U21401 (N_21401,N_18276,N_18698);
nor U21402 (N_21402,N_19927,N_18609);
and U21403 (N_21403,N_19525,N_18338);
nor U21404 (N_21404,N_19752,N_18008);
nor U21405 (N_21405,N_18045,N_19031);
and U21406 (N_21406,N_18997,N_19505);
nor U21407 (N_21407,N_18432,N_19204);
or U21408 (N_21408,N_19427,N_19522);
or U21409 (N_21409,N_18774,N_19217);
xor U21410 (N_21410,N_19059,N_19463);
nor U21411 (N_21411,N_18976,N_18947);
or U21412 (N_21412,N_18616,N_19893);
xnor U21413 (N_21413,N_19818,N_18551);
or U21414 (N_21414,N_19198,N_18434);
and U21415 (N_21415,N_19431,N_18224);
nand U21416 (N_21416,N_18269,N_18065);
and U21417 (N_21417,N_19737,N_18154);
xor U21418 (N_21418,N_19184,N_19561);
or U21419 (N_21419,N_19532,N_19797);
xor U21420 (N_21420,N_18012,N_18580);
nand U21421 (N_21421,N_18784,N_18609);
nand U21422 (N_21422,N_18061,N_19072);
xor U21423 (N_21423,N_18041,N_18806);
xor U21424 (N_21424,N_18585,N_19762);
or U21425 (N_21425,N_18015,N_19717);
xor U21426 (N_21426,N_18405,N_18732);
xor U21427 (N_21427,N_18721,N_19596);
or U21428 (N_21428,N_19581,N_19019);
nor U21429 (N_21429,N_18237,N_18913);
xnor U21430 (N_21430,N_18886,N_18422);
nor U21431 (N_21431,N_18090,N_19606);
or U21432 (N_21432,N_19502,N_18914);
or U21433 (N_21433,N_18855,N_18150);
nor U21434 (N_21434,N_18813,N_18773);
nand U21435 (N_21435,N_19982,N_19576);
xor U21436 (N_21436,N_19427,N_19252);
nand U21437 (N_21437,N_19252,N_19491);
xor U21438 (N_21438,N_18914,N_18428);
nand U21439 (N_21439,N_19808,N_19564);
or U21440 (N_21440,N_18919,N_18694);
nand U21441 (N_21441,N_19808,N_18520);
xnor U21442 (N_21442,N_19770,N_18482);
xor U21443 (N_21443,N_19812,N_19213);
and U21444 (N_21444,N_18804,N_18280);
nand U21445 (N_21445,N_18377,N_19026);
or U21446 (N_21446,N_18851,N_19045);
nor U21447 (N_21447,N_18949,N_19000);
nand U21448 (N_21448,N_18099,N_18036);
nor U21449 (N_21449,N_19192,N_19536);
xnor U21450 (N_21450,N_18397,N_18590);
or U21451 (N_21451,N_18289,N_18164);
and U21452 (N_21452,N_19284,N_19511);
xnor U21453 (N_21453,N_19616,N_18364);
xor U21454 (N_21454,N_19848,N_19617);
and U21455 (N_21455,N_19765,N_18487);
nor U21456 (N_21456,N_19790,N_18284);
nor U21457 (N_21457,N_18745,N_19853);
nand U21458 (N_21458,N_18017,N_18196);
and U21459 (N_21459,N_19275,N_19151);
xor U21460 (N_21460,N_19678,N_19882);
xor U21461 (N_21461,N_18725,N_18987);
xor U21462 (N_21462,N_19347,N_19488);
and U21463 (N_21463,N_19047,N_18017);
xnor U21464 (N_21464,N_19047,N_19450);
nand U21465 (N_21465,N_19032,N_18664);
nor U21466 (N_21466,N_18790,N_18902);
or U21467 (N_21467,N_18136,N_19809);
nand U21468 (N_21468,N_19002,N_19631);
xor U21469 (N_21469,N_18554,N_19525);
and U21470 (N_21470,N_18284,N_18721);
nand U21471 (N_21471,N_18434,N_19043);
or U21472 (N_21472,N_18196,N_19040);
xnor U21473 (N_21473,N_18236,N_19050);
nand U21474 (N_21474,N_18349,N_18401);
nand U21475 (N_21475,N_18015,N_18300);
xnor U21476 (N_21476,N_18389,N_19118);
nor U21477 (N_21477,N_18310,N_18885);
nor U21478 (N_21478,N_18192,N_18025);
and U21479 (N_21479,N_18679,N_18454);
and U21480 (N_21480,N_18391,N_18251);
or U21481 (N_21481,N_19364,N_18582);
and U21482 (N_21482,N_19551,N_18025);
nor U21483 (N_21483,N_19842,N_19010);
nor U21484 (N_21484,N_19185,N_19580);
nor U21485 (N_21485,N_19156,N_18271);
nand U21486 (N_21486,N_18948,N_18474);
xnor U21487 (N_21487,N_18032,N_19895);
nor U21488 (N_21488,N_19267,N_18827);
xor U21489 (N_21489,N_18587,N_18623);
and U21490 (N_21490,N_18029,N_18888);
nor U21491 (N_21491,N_19669,N_18634);
or U21492 (N_21492,N_19676,N_19411);
nand U21493 (N_21493,N_19048,N_18762);
nand U21494 (N_21494,N_18945,N_18603);
or U21495 (N_21495,N_19297,N_19855);
or U21496 (N_21496,N_18671,N_19371);
nand U21497 (N_21497,N_19743,N_18655);
nand U21498 (N_21498,N_18005,N_19349);
nand U21499 (N_21499,N_18267,N_19602);
nor U21500 (N_21500,N_18122,N_18805);
nor U21501 (N_21501,N_18589,N_19427);
and U21502 (N_21502,N_18117,N_19087);
and U21503 (N_21503,N_18561,N_18821);
nand U21504 (N_21504,N_19327,N_19103);
nand U21505 (N_21505,N_19141,N_18369);
xor U21506 (N_21506,N_18115,N_18070);
nor U21507 (N_21507,N_18875,N_18690);
or U21508 (N_21508,N_18963,N_19537);
nor U21509 (N_21509,N_18692,N_18420);
xor U21510 (N_21510,N_19111,N_18494);
and U21511 (N_21511,N_19081,N_18231);
nand U21512 (N_21512,N_19343,N_19050);
nor U21513 (N_21513,N_18098,N_18608);
nand U21514 (N_21514,N_19407,N_18508);
nor U21515 (N_21515,N_19315,N_19017);
xor U21516 (N_21516,N_18850,N_19569);
nand U21517 (N_21517,N_18955,N_18378);
and U21518 (N_21518,N_18458,N_19862);
or U21519 (N_21519,N_18228,N_19732);
or U21520 (N_21520,N_18260,N_19997);
and U21521 (N_21521,N_18864,N_19006);
xnor U21522 (N_21522,N_18893,N_19012);
and U21523 (N_21523,N_18096,N_19780);
or U21524 (N_21524,N_19162,N_19834);
and U21525 (N_21525,N_18053,N_18103);
and U21526 (N_21526,N_18340,N_19336);
xor U21527 (N_21527,N_18390,N_18128);
and U21528 (N_21528,N_19066,N_18340);
or U21529 (N_21529,N_18390,N_18410);
or U21530 (N_21530,N_18313,N_18215);
xnor U21531 (N_21531,N_19389,N_19056);
or U21532 (N_21532,N_18555,N_19267);
or U21533 (N_21533,N_19463,N_18622);
and U21534 (N_21534,N_19843,N_19708);
xor U21535 (N_21535,N_18072,N_19056);
or U21536 (N_21536,N_19859,N_19913);
or U21537 (N_21537,N_18691,N_19121);
or U21538 (N_21538,N_18543,N_19765);
nand U21539 (N_21539,N_18243,N_18589);
nor U21540 (N_21540,N_19246,N_19031);
nand U21541 (N_21541,N_19751,N_18317);
and U21542 (N_21542,N_18580,N_19368);
and U21543 (N_21543,N_18373,N_19707);
nor U21544 (N_21544,N_18337,N_19376);
xor U21545 (N_21545,N_18019,N_19617);
nor U21546 (N_21546,N_18813,N_19615);
nand U21547 (N_21547,N_18120,N_19468);
nand U21548 (N_21548,N_18179,N_19115);
xor U21549 (N_21549,N_18325,N_19174);
or U21550 (N_21550,N_18855,N_18585);
nor U21551 (N_21551,N_19706,N_19890);
and U21552 (N_21552,N_18415,N_19122);
nor U21553 (N_21553,N_19344,N_19607);
nand U21554 (N_21554,N_18996,N_19707);
and U21555 (N_21555,N_18968,N_18629);
nor U21556 (N_21556,N_19640,N_18475);
xnor U21557 (N_21557,N_19805,N_19893);
xor U21558 (N_21558,N_19362,N_19798);
xnor U21559 (N_21559,N_18881,N_19459);
nand U21560 (N_21560,N_18413,N_19403);
and U21561 (N_21561,N_18445,N_19401);
nand U21562 (N_21562,N_19809,N_19919);
nand U21563 (N_21563,N_19486,N_19119);
xnor U21564 (N_21564,N_18974,N_19008);
and U21565 (N_21565,N_19076,N_19376);
and U21566 (N_21566,N_19905,N_18485);
nor U21567 (N_21567,N_19937,N_19008);
or U21568 (N_21568,N_19338,N_19496);
nand U21569 (N_21569,N_18973,N_18451);
or U21570 (N_21570,N_18042,N_18201);
or U21571 (N_21571,N_18153,N_18291);
xnor U21572 (N_21572,N_18484,N_19922);
xor U21573 (N_21573,N_18446,N_18380);
and U21574 (N_21574,N_18312,N_19730);
or U21575 (N_21575,N_18232,N_19828);
or U21576 (N_21576,N_19656,N_19491);
or U21577 (N_21577,N_19458,N_18972);
nor U21578 (N_21578,N_19753,N_18772);
nor U21579 (N_21579,N_19477,N_18353);
or U21580 (N_21580,N_18868,N_18831);
xnor U21581 (N_21581,N_18838,N_18361);
nand U21582 (N_21582,N_18019,N_19795);
and U21583 (N_21583,N_19615,N_18733);
or U21584 (N_21584,N_19406,N_18424);
and U21585 (N_21585,N_18711,N_18214);
and U21586 (N_21586,N_18174,N_18601);
nor U21587 (N_21587,N_18584,N_18695);
nand U21588 (N_21588,N_18749,N_18191);
and U21589 (N_21589,N_19383,N_19604);
or U21590 (N_21590,N_19030,N_19138);
nand U21591 (N_21591,N_19483,N_18869);
or U21592 (N_21592,N_18735,N_18953);
and U21593 (N_21593,N_18646,N_19227);
and U21594 (N_21594,N_18078,N_18363);
or U21595 (N_21595,N_18895,N_18530);
nand U21596 (N_21596,N_18607,N_19156);
xnor U21597 (N_21597,N_19000,N_18784);
and U21598 (N_21598,N_18252,N_18989);
nor U21599 (N_21599,N_18920,N_19554);
or U21600 (N_21600,N_18373,N_18568);
nand U21601 (N_21601,N_19658,N_18691);
xor U21602 (N_21602,N_18272,N_18220);
and U21603 (N_21603,N_18488,N_18703);
nand U21604 (N_21604,N_19937,N_19506);
nand U21605 (N_21605,N_18262,N_18348);
xnor U21606 (N_21606,N_18423,N_19581);
nand U21607 (N_21607,N_18298,N_19314);
nand U21608 (N_21608,N_18676,N_18191);
or U21609 (N_21609,N_18112,N_19425);
nand U21610 (N_21610,N_18376,N_18238);
xor U21611 (N_21611,N_18523,N_19668);
nand U21612 (N_21612,N_18582,N_19450);
and U21613 (N_21613,N_18595,N_19681);
xnor U21614 (N_21614,N_18698,N_18586);
and U21615 (N_21615,N_19392,N_18989);
nand U21616 (N_21616,N_18487,N_19650);
and U21617 (N_21617,N_18951,N_19122);
nand U21618 (N_21618,N_19366,N_19675);
nor U21619 (N_21619,N_19851,N_18540);
or U21620 (N_21620,N_18952,N_18338);
xor U21621 (N_21621,N_19991,N_18030);
nand U21622 (N_21622,N_19062,N_18332);
xnor U21623 (N_21623,N_18222,N_18641);
nor U21624 (N_21624,N_18104,N_18856);
nor U21625 (N_21625,N_18513,N_18452);
xor U21626 (N_21626,N_19363,N_19901);
xnor U21627 (N_21627,N_19586,N_19726);
nand U21628 (N_21628,N_19490,N_18514);
nor U21629 (N_21629,N_18557,N_18460);
nand U21630 (N_21630,N_18184,N_19723);
and U21631 (N_21631,N_19730,N_18856);
nand U21632 (N_21632,N_18332,N_19178);
or U21633 (N_21633,N_19277,N_18893);
and U21634 (N_21634,N_18524,N_19866);
nand U21635 (N_21635,N_19643,N_19868);
and U21636 (N_21636,N_19543,N_18868);
and U21637 (N_21637,N_19913,N_18072);
and U21638 (N_21638,N_18689,N_18384);
nor U21639 (N_21639,N_19838,N_18766);
xnor U21640 (N_21640,N_19954,N_18786);
nor U21641 (N_21641,N_19909,N_18788);
and U21642 (N_21642,N_19747,N_19708);
and U21643 (N_21643,N_19685,N_19414);
nand U21644 (N_21644,N_19002,N_19278);
nor U21645 (N_21645,N_18394,N_18515);
nand U21646 (N_21646,N_18500,N_18079);
and U21647 (N_21647,N_19557,N_19953);
nand U21648 (N_21648,N_19845,N_18308);
nor U21649 (N_21649,N_19877,N_18654);
nand U21650 (N_21650,N_19540,N_19624);
and U21651 (N_21651,N_18932,N_19993);
or U21652 (N_21652,N_18037,N_18381);
xnor U21653 (N_21653,N_18576,N_18470);
or U21654 (N_21654,N_19612,N_19762);
and U21655 (N_21655,N_19600,N_19476);
or U21656 (N_21656,N_19305,N_19856);
nand U21657 (N_21657,N_18710,N_19781);
and U21658 (N_21658,N_19141,N_19269);
and U21659 (N_21659,N_19673,N_19506);
or U21660 (N_21660,N_18518,N_18472);
nand U21661 (N_21661,N_18718,N_19259);
nand U21662 (N_21662,N_18131,N_18433);
nand U21663 (N_21663,N_18023,N_18714);
nand U21664 (N_21664,N_19762,N_18571);
nor U21665 (N_21665,N_18318,N_18416);
nor U21666 (N_21666,N_18559,N_18767);
nor U21667 (N_21667,N_19898,N_18249);
nand U21668 (N_21668,N_18383,N_19439);
xor U21669 (N_21669,N_18867,N_19552);
or U21670 (N_21670,N_19997,N_18575);
nand U21671 (N_21671,N_18218,N_19449);
or U21672 (N_21672,N_19421,N_19335);
and U21673 (N_21673,N_19504,N_18553);
and U21674 (N_21674,N_18325,N_19039);
nand U21675 (N_21675,N_19097,N_18841);
or U21676 (N_21676,N_19746,N_18499);
xnor U21677 (N_21677,N_18210,N_19467);
or U21678 (N_21678,N_18321,N_19364);
nor U21679 (N_21679,N_19979,N_18158);
xor U21680 (N_21680,N_18423,N_19153);
nand U21681 (N_21681,N_18127,N_18811);
nand U21682 (N_21682,N_18080,N_19779);
xor U21683 (N_21683,N_18715,N_19856);
xor U21684 (N_21684,N_18215,N_19359);
nand U21685 (N_21685,N_18848,N_19770);
and U21686 (N_21686,N_19205,N_18743);
and U21687 (N_21687,N_19742,N_19288);
nor U21688 (N_21688,N_19185,N_18171);
nor U21689 (N_21689,N_18338,N_19234);
xor U21690 (N_21690,N_19010,N_19671);
xor U21691 (N_21691,N_19816,N_18603);
xnor U21692 (N_21692,N_19805,N_19132);
nor U21693 (N_21693,N_19437,N_19858);
nor U21694 (N_21694,N_18554,N_18474);
and U21695 (N_21695,N_18394,N_19549);
nor U21696 (N_21696,N_18155,N_19807);
nand U21697 (N_21697,N_18064,N_18877);
nor U21698 (N_21698,N_19784,N_19627);
or U21699 (N_21699,N_18146,N_18227);
nand U21700 (N_21700,N_19930,N_18703);
or U21701 (N_21701,N_18472,N_18502);
and U21702 (N_21702,N_18797,N_18248);
nand U21703 (N_21703,N_19965,N_18949);
and U21704 (N_21704,N_18279,N_19069);
nand U21705 (N_21705,N_19460,N_18715);
xor U21706 (N_21706,N_19489,N_19786);
xor U21707 (N_21707,N_19636,N_19997);
or U21708 (N_21708,N_18831,N_18267);
or U21709 (N_21709,N_18097,N_19235);
nor U21710 (N_21710,N_19503,N_18668);
and U21711 (N_21711,N_18014,N_18591);
nand U21712 (N_21712,N_19464,N_19170);
nor U21713 (N_21713,N_18269,N_19120);
and U21714 (N_21714,N_19158,N_18109);
xnor U21715 (N_21715,N_19215,N_18971);
xnor U21716 (N_21716,N_19923,N_18688);
and U21717 (N_21717,N_18866,N_19771);
nor U21718 (N_21718,N_18763,N_18075);
nor U21719 (N_21719,N_19106,N_19921);
and U21720 (N_21720,N_19399,N_18052);
nand U21721 (N_21721,N_18447,N_18287);
xnor U21722 (N_21722,N_19170,N_18485);
xor U21723 (N_21723,N_19672,N_19466);
nand U21724 (N_21724,N_19370,N_19533);
or U21725 (N_21725,N_19096,N_19773);
xnor U21726 (N_21726,N_19979,N_19459);
nand U21727 (N_21727,N_18706,N_18389);
nand U21728 (N_21728,N_18469,N_18136);
nor U21729 (N_21729,N_18457,N_19540);
nand U21730 (N_21730,N_18099,N_18921);
nand U21731 (N_21731,N_19589,N_19122);
nand U21732 (N_21732,N_18149,N_18360);
and U21733 (N_21733,N_18362,N_18727);
xor U21734 (N_21734,N_19869,N_19281);
nand U21735 (N_21735,N_19557,N_19146);
or U21736 (N_21736,N_19498,N_18652);
nand U21737 (N_21737,N_19550,N_18673);
or U21738 (N_21738,N_19690,N_18712);
xnor U21739 (N_21739,N_19504,N_19926);
nor U21740 (N_21740,N_19035,N_19525);
xnor U21741 (N_21741,N_19508,N_18606);
nand U21742 (N_21742,N_18626,N_18938);
nand U21743 (N_21743,N_19310,N_19385);
nand U21744 (N_21744,N_19066,N_18732);
xor U21745 (N_21745,N_18819,N_19413);
nor U21746 (N_21746,N_19017,N_19772);
xor U21747 (N_21747,N_19142,N_18936);
nor U21748 (N_21748,N_19001,N_19822);
or U21749 (N_21749,N_18438,N_18731);
nor U21750 (N_21750,N_18519,N_18203);
nor U21751 (N_21751,N_18827,N_18575);
xor U21752 (N_21752,N_19705,N_18980);
or U21753 (N_21753,N_19171,N_18190);
and U21754 (N_21754,N_19658,N_18542);
xor U21755 (N_21755,N_19025,N_19188);
xnor U21756 (N_21756,N_19766,N_19920);
and U21757 (N_21757,N_19374,N_18453);
nand U21758 (N_21758,N_18925,N_18395);
or U21759 (N_21759,N_19832,N_18140);
xor U21760 (N_21760,N_19842,N_19724);
or U21761 (N_21761,N_18279,N_18524);
xnor U21762 (N_21762,N_18474,N_18294);
xor U21763 (N_21763,N_19260,N_18491);
or U21764 (N_21764,N_19011,N_19414);
xnor U21765 (N_21765,N_18326,N_18899);
and U21766 (N_21766,N_18951,N_18671);
xnor U21767 (N_21767,N_18409,N_19916);
or U21768 (N_21768,N_19101,N_18878);
or U21769 (N_21769,N_19399,N_19143);
xor U21770 (N_21770,N_18511,N_19791);
xor U21771 (N_21771,N_18339,N_18050);
nand U21772 (N_21772,N_18485,N_18955);
or U21773 (N_21773,N_19008,N_19501);
or U21774 (N_21774,N_19238,N_19089);
xor U21775 (N_21775,N_18575,N_18963);
nor U21776 (N_21776,N_18963,N_18705);
and U21777 (N_21777,N_19005,N_18995);
nand U21778 (N_21778,N_18402,N_19602);
xnor U21779 (N_21779,N_18410,N_18927);
and U21780 (N_21780,N_19851,N_19757);
nor U21781 (N_21781,N_19127,N_19762);
nand U21782 (N_21782,N_18163,N_19256);
xnor U21783 (N_21783,N_18577,N_19197);
xnor U21784 (N_21784,N_18958,N_18240);
nand U21785 (N_21785,N_19157,N_19662);
nor U21786 (N_21786,N_19187,N_19258);
and U21787 (N_21787,N_18499,N_19932);
nand U21788 (N_21788,N_19741,N_19275);
nand U21789 (N_21789,N_18164,N_19834);
or U21790 (N_21790,N_19935,N_19187);
nand U21791 (N_21791,N_19141,N_18623);
nor U21792 (N_21792,N_19593,N_18199);
xnor U21793 (N_21793,N_19321,N_19913);
or U21794 (N_21794,N_18135,N_18371);
and U21795 (N_21795,N_19549,N_19325);
and U21796 (N_21796,N_18133,N_18457);
nand U21797 (N_21797,N_19595,N_19795);
and U21798 (N_21798,N_18222,N_18055);
xnor U21799 (N_21799,N_18493,N_18448);
nand U21800 (N_21800,N_19004,N_19068);
xor U21801 (N_21801,N_18397,N_18557);
xnor U21802 (N_21802,N_18798,N_19107);
nand U21803 (N_21803,N_19372,N_18254);
xor U21804 (N_21804,N_19670,N_18393);
and U21805 (N_21805,N_19357,N_18300);
nor U21806 (N_21806,N_18603,N_19796);
xor U21807 (N_21807,N_18859,N_18682);
nor U21808 (N_21808,N_19487,N_18345);
or U21809 (N_21809,N_18115,N_18608);
or U21810 (N_21810,N_19482,N_18125);
nand U21811 (N_21811,N_19845,N_18253);
nand U21812 (N_21812,N_19638,N_18928);
and U21813 (N_21813,N_18299,N_19085);
nand U21814 (N_21814,N_19057,N_18489);
nand U21815 (N_21815,N_18388,N_19598);
nor U21816 (N_21816,N_19894,N_19409);
or U21817 (N_21817,N_18540,N_19638);
nor U21818 (N_21818,N_18831,N_19595);
nand U21819 (N_21819,N_18959,N_19792);
nand U21820 (N_21820,N_18319,N_19479);
or U21821 (N_21821,N_18808,N_18168);
xnor U21822 (N_21822,N_19282,N_19117);
nor U21823 (N_21823,N_19215,N_18149);
and U21824 (N_21824,N_19385,N_19550);
xnor U21825 (N_21825,N_19415,N_19429);
and U21826 (N_21826,N_18187,N_18945);
nand U21827 (N_21827,N_19415,N_18822);
and U21828 (N_21828,N_19766,N_18844);
or U21829 (N_21829,N_18693,N_18998);
xnor U21830 (N_21830,N_19924,N_19735);
or U21831 (N_21831,N_18596,N_18405);
nor U21832 (N_21832,N_19831,N_18412);
or U21833 (N_21833,N_18927,N_18630);
or U21834 (N_21834,N_18558,N_19271);
or U21835 (N_21835,N_18295,N_18590);
nand U21836 (N_21836,N_18057,N_18098);
nand U21837 (N_21837,N_18349,N_19523);
nand U21838 (N_21838,N_18356,N_18353);
xnor U21839 (N_21839,N_18026,N_18957);
or U21840 (N_21840,N_18554,N_19576);
and U21841 (N_21841,N_19566,N_19895);
xnor U21842 (N_21842,N_18659,N_19368);
and U21843 (N_21843,N_19905,N_19044);
and U21844 (N_21844,N_19963,N_19676);
or U21845 (N_21845,N_18917,N_18961);
or U21846 (N_21846,N_18728,N_19383);
and U21847 (N_21847,N_18941,N_19864);
and U21848 (N_21848,N_18319,N_18761);
and U21849 (N_21849,N_18934,N_18201);
nand U21850 (N_21850,N_18472,N_18482);
or U21851 (N_21851,N_18183,N_18955);
nand U21852 (N_21852,N_19716,N_19472);
and U21853 (N_21853,N_19702,N_18358);
and U21854 (N_21854,N_19890,N_19782);
nand U21855 (N_21855,N_19870,N_19536);
nand U21856 (N_21856,N_18334,N_18730);
nand U21857 (N_21857,N_18881,N_18818);
nand U21858 (N_21858,N_18280,N_18633);
xor U21859 (N_21859,N_19230,N_19195);
and U21860 (N_21860,N_19744,N_18064);
xnor U21861 (N_21861,N_18652,N_18856);
and U21862 (N_21862,N_18932,N_18086);
and U21863 (N_21863,N_19808,N_18855);
nand U21864 (N_21864,N_19900,N_19147);
and U21865 (N_21865,N_19038,N_18437);
xor U21866 (N_21866,N_19799,N_19996);
or U21867 (N_21867,N_18719,N_19575);
nand U21868 (N_21868,N_18199,N_19795);
nor U21869 (N_21869,N_19288,N_19646);
and U21870 (N_21870,N_18887,N_18804);
xnor U21871 (N_21871,N_18185,N_18593);
or U21872 (N_21872,N_18402,N_19001);
and U21873 (N_21873,N_19501,N_19480);
and U21874 (N_21874,N_18422,N_19602);
nand U21875 (N_21875,N_18561,N_18918);
xnor U21876 (N_21876,N_18262,N_18841);
xor U21877 (N_21877,N_19638,N_19030);
or U21878 (N_21878,N_18905,N_19075);
or U21879 (N_21879,N_18671,N_19872);
nor U21880 (N_21880,N_18872,N_19624);
nand U21881 (N_21881,N_19221,N_18634);
or U21882 (N_21882,N_18219,N_19307);
and U21883 (N_21883,N_18888,N_18453);
or U21884 (N_21884,N_18989,N_19496);
nor U21885 (N_21885,N_19138,N_19969);
or U21886 (N_21886,N_18377,N_18970);
xor U21887 (N_21887,N_19791,N_18412);
nor U21888 (N_21888,N_18256,N_18562);
or U21889 (N_21889,N_19853,N_19314);
xnor U21890 (N_21890,N_18796,N_18054);
or U21891 (N_21891,N_19297,N_19971);
nor U21892 (N_21892,N_18974,N_19356);
xnor U21893 (N_21893,N_18969,N_18809);
xnor U21894 (N_21894,N_19399,N_18890);
xor U21895 (N_21895,N_18654,N_19873);
or U21896 (N_21896,N_18188,N_19569);
nand U21897 (N_21897,N_19389,N_18358);
and U21898 (N_21898,N_18259,N_18742);
nand U21899 (N_21899,N_18834,N_19686);
xnor U21900 (N_21900,N_18192,N_18055);
or U21901 (N_21901,N_18204,N_19650);
nor U21902 (N_21902,N_19940,N_18165);
and U21903 (N_21903,N_18882,N_19403);
or U21904 (N_21904,N_19081,N_19255);
and U21905 (N_21905,N_19129,N_18199);
or U21906 (N_21906,N_19480,N_19985);
xnor U21907 (N_21907,N_19731,N_19872);
nand U21908 (N_21908,N_18834,N_19674);
and U21909 (N_21909,N_18082,N_19581);
xnor U21910 (N_21910,N_18960,N_19948);
nand U21911 (N_21911,N_19584,N_18161);
nand U21912 (N_21912,N_18164,N_19433);
and U21913 (N_21913,N_18842,N_18841);
and U21914 (N_21914,N_18686,N_18412);
and U21915 (N_21915,N_19449,N_19163);
xor U21916 (N_21916,N_18244,N_19587);
nor U21917 (N_21917,N_18101,N_18798);
nor U21918 (N_21918,N_18221,N_19606);
xor U21919 (N_21919,N_18422,N_19157);
xnor U21920 (N_21920,N_18723,N_19903);
nand U21921 (N_21921,N_18628,N_18881);
nand U21922 (N_21922,N_18414,N_18063);
or U21923 (N_21923,N_18130,N_19884);
nand U21924 (N_21924,N_19639,N_18739);
xnor U21925 (N_21925,N_19541,N_19854);
and U21926 (N_21926,N_19743,N_19323);
or U21927 (N_21927,N_19268,N_19265);
and U21928 (N_21928,N_19216,N_18791);
and U21929 (N_21929,N_19615,N_19218);
xor U21930 (N_21930,N_18852,N_19541);
and U21931 (N_21931,N_19712,N_18824);
nor U21932 (N_21932,N_19346,N_18744);
xor U21933 (N_21933,N_18544,N_19297);
xnor U21934 (N_21934,N_18205,N_19189);
xnor U21935 (N_21935,N_18017,N_19654);
xor U21936 (N_21936,N_18163,N_18076);
or U21937 (N_21937,N_19709,N_19052);
or U21938 (N_21938,N_19954,N_19355);
nor U21939 (N_21939,N_19743,N_19485);
and U21940 (N_21940,N_18851,N_19182);
xor U21941 (N_21941,N_19655,N_19689);
or U21942 (N_21942,N_18896,N_19669);
or U21943 (N_21943,N_18968,N_18948);
and U21944 (N_21944,N_18806,N_19224);
nor U21945 (N_21945,N_18713,N_19130);
xnor U21946 (N_21946,N_18799,N_19095);
and U21947 (N_21947,N_19558,N_18353);
nand U21948 (N_21948,N_18881,N_19200);
nand U21949 (N_21949,N_18506,N_19766);
nor U21950 (N_21950,N_19883,N_18563);
nor U21951 (N_21951,N_19548,N_18843);
or U21952 (N_21952,N_19461,N_18152);
or U21953 (N_21953,N_18403,N_19356);
or U21954 (N_21954,N_19029,N_19516);
xnor U21955 (N_21955,N_18383,N_18743);
xnor U21956 (N_21956,N_18016,N_18449);
nand U21957 (N_21957,N_19389,N_19643);
or U21958 (N_21958,N_18135,N_19524);
nor U21959 (N_21959,N_19056,N_19453);
nor U21960 (N_21960,N_19957,N_18957);
nand U21961 (N_21961,N_19351,N_18035);
or U21962 (N_21962,N_18414,N_18307);
or U21963 (N_21963,N_18442,N_19505);
nor U21964 (N_21964,N_19400,N_19320);
xnor U21965 (N_21965,N_18992,N_18954);
and U21966 (N_21966,N_19459,N_18247);
nand U21967 (N_21967,N_19070,N_18190);
xnor U21968 (N_21968,N_19400,N_18547);
and U21969 (N_21969,N_18386,N_19014);
nand U21970 (N_21970,N_18023,N_18286);
or U21971 (N_21971,N_19550,N_19048);
and U21972 (N_21972,N_19364,N_19536);
nand U21973 (N_21973,N_19361,N_18229);
or U21974 (N_21974,N_19100,N_18834);
nor U21975 (N_21975,N_18140,N_19200);
and U21976 (N_21976,N_18407,N_19409);
nand U21977 (N_21977,N_18768,N_19463);
xnor U21978 (N_21978,N_19850,N_18564);
xnor U21979 (N_21979,N_18024,N_19376);
or U21980 (N_21980,N_19410,N_19493);
nor U21981 (N_21981,N_18896,N_19274);
xor U21982 (N_21982,N_19965,N_19132);
or U21983 (N_21983,N_19288,N_19003);
nor U21984 (N_21984,N_18061,N_19278);
nor U21985 (N_21985,N_19953,N_19769);
and U21986 (N_21986,N_18428,N_18910);
or U21987 (N_21987,N_19742,N_19749);
or U21988 (N_21988,N_19177,N_19628);
nor U21989 (N_21989,N_19046,N_19438);
nor U21990 (N_21990,N_19260,N_18680);
xnor U21991 (N_21991,N_18211,N_19183);
or U21992 (N_21992,N_18177,N_18120);
nand U21993 (N_21993,N_19540,N_18717);
xor U21994 (N_21994,N_19778,N_19288);
nand U21995 (N_21995,N_18989,N_19498);
and U21996 (N_21996,N_18527,N_18477);
nor U21997 (N_21997,N_19451,N_19844);
nand U21998 (N_21998,N_18724,N_19653);
xor U21999 (N_21999,N_18453,N_18382);
or U22000 (N_22000,N_20188,N_20433);
and U22001 (N_22001,N_20034,N_20693);
xor U22002 (N_22002,N_21814,N_20618);
or U22003 (N_22003,N_21466,N_21597);
or U22004 (N_22004,N_21264,N_21228);
and U22005 (N_22005,N_21955,N_21988);
nand U22006 (N_22006,N_20157,N_21653);
nor U22007 (N_22007,N_21746,N_20089);
xnor U22008 (N_22008,N_21144,N_20612);
and U22009 (N_22009,N_20992,N_20844);
or U22010 (N_22010,N_20470,N_21017);
nand U22011 (N_22011,N_21733,N_20398);
nand U22012 (N_22012,N_20629,N_20885);
nand U22013 (N_22013,N_21420,N_21461);
nand U22014 (N_22014,N_20778,N_21661);
and U22015 (N_22015,N_20904,N_20045);
nor U22016 (N_22016,N_20742,N_20663);
xnor U22017 (N_22017,N_20113,N_20447);
nor U22018 (N_22018,N_21566,N_20633);
or U22019 (N_22019,N_20847,N_20175);
nand U22020 (N_22020,N_21359,N_20869);
and U22021 (N_22021,N_20653,N_21012);
or U22022 (N_22022,N_20625,N_21090);
xnor U22023 (N_22023,N_21647,N_20554);
and U22024 (N_22024,N_21612,N_21030);
nand U22025 (N_22025,N_20342,N_21022);
or U22026 (N_22026,N_21762,N_21790);
nor U22027 (N_22027,N_20003,N_21415);
and U22028 (N_22028,N_21188,N_21819);
nor U22029 (N_22029,N_21172,N_21037);
and U22030 (N_22030,N_20371,N_21718);
and U22031 (N_22031,N_21217,N_20775);
nand U22032 (N_22032,N_20086,N_20913);
and U22033 (N_22033,N_21399,N_21565);
xnor U22034 (N_22034,N_20182,N_21195);
or U22035 (N_22035,N_20132,N_20329);
nor U22036 (N_22036,N_21582,N_21501);
nor U22037 (N_22037,N_21044,N_21869);
nand U22038 (N_22038,N_21395,N_21673);
nor U22039 (N_22039,N_20899,N_21362);
and U22040 (N_22040,N_21475,N_21447);
nor U22041 (N_22041,N_20244,N_21478);
or U22042 (N_22042,N_21434,N_20834);
or U22043 (N_22043,N_21802,N_21868);
nand U22044 (N_22044,N_20199,N_20396);
nand U22045 (N_22045,N_20503,N_20088);
or U22046 (N_22046,N_20388,N_21282);
nand U22047 (N_22047,N_21943,N_21643);
or U22048 (N_22048,N_20627,N_20100);
nor U22049 (N_22049,N_20513,N_20831);
and U22050 (N_22050,N_20337,N_20134);
nand U22051 (N_22051,N_20631,N_20131);
nor U22052 (N_22052,N_20499,N_21816);
xor U22053 (N_22053,N_20839,N_20526);
or U22054 (N_22054,N_21484,N_20636);
or U22055 (N_22055,N_20039,N_21191);
and U22056 (N_22056,N_20278,N_21702);
nor U22057 (N_22057,N_20151,N_21440);
and U22058 (N_22058,N_21865,N_20280);
nor U22059 (N_22059,N_20282,N_21438);
or U22060 (N_22060,N_20428,N_20906);
and U22061 (N_22061,N_21644,N_21689);
nor U22062 (N_22062,N_20174,N_21700);
nand U22063 (N_22063,N_20385,N_20430);
and U22064 (N_22064,N_21716,N_21105);
or U22065 (N_22065,N_20827,N_20912);
and U22066 (N_22066,N_20845,N_21035);
nor U22067 (N_22067,N_20386,N_20475);
nor U22068 (N_22068,N_21132,N_21754);
xor U22069 (N_22069,N_21493,N_20208);
xor U22070 (N_22070,N_21633,N_20318);
and U22071 (N_22071,N_21637,N_20659);
or U22072 (N_22072,N_21927,N_20062);
or U22073 (N_22073,N_21098,N_21967);
nor U22074 (N_22074,N_21562,N_21801);
or U22075 (N_22075,N_21208,N_21928);
or U22076 (N_22076,N_20426,N_20190);
nor U22077 (N_22077,N_21518,N_20009);
nand U22078 (N_22078,N_20108,N_20984);
and U22079 (N_22079,N_21891,N_21249);
and U22080 (N_22080,N_21243,N_21036);
and U22081 (N_22081,N_21765,N_21898);
nand U22082 (N_22082,N_20795,N_21250);
nand U22083 (N_22083,N_21893,N_21956);
xor U22084 (N_22084,N_21608,N_21779);
nor U22085 (N_22085,N_20032,N_21656);
nand U22086 (N_22086,N_20158,N_21154);
nand U22087 (N_22087,N_20534,N_21987);
or U22088 (N_22088,N_20564,N_20734);
xnor U22089 (N_22089,N_21141,N_20766);
or U22090 (N_22090,N_20423,N_20583);
xor U22091 (N_22091,N_21999,N_21841);
nand U22092 (N_22092,N_21958,N_21425);
and U22093 (N_22093,N_20299,N_21525);
nor U22094 (N_22094,N_21023,N_21435);
or U22095 (N_22095,N_21680,N_21963);
xnor U22096 (N_22096,N_21005,N_21617);
or U22097 (N_22097,N_20105,N_20682);
xor U22098 (N_22098,N_20921,N_21285);
nand U22099 (N_22099,N_21140,N_20576);
xor U22100 (N_22100,N_21419,N_20012);
nor U22101 (N_22101,N_20245,N_21717);
or U22102 (N_22102,N_21166,N_21960);
xnor U22103 (N_22103,N_21632,N_20677);
nor U22104 (N_22104,N_21839,N_21010);
nand U22105 (N_22105,N_20973,N_20226);
and U22106 (N_22106,N_21374,N_21054);
nor U22107 (N_22107,N_20768,N_21863);
or U22108 (N_22108,N_20035,N_20991);
nand U22109 (N_22109,N_21183,N_20938);
nor U22110 (N_22110,N_20002,N_20943);
nand U22111 (N_22111,N_20241,N_20529);
nor U22112 (N_22112,N_20689,N_21629);
and U22113 (N_22113,N_20710,N_21185);
nand U22114 (N_22114,N_21248,N_20983);
xnor U22115 (N_22115,N_21757,N_21062);
or U22116 (N_22116,N_21735,N_21329);
nor U22117 (N_22117,N_21254,N_20044);
nor U22118 (N_22118,N_20261,N_21400);
and U22119 (N_22119,N_20441,N_20805);
and U22120 (N_22120,N_21178,N_20422);
xnor U22121 (N_22121,N_21111,N_21946);
and U22122 (N_22122,N_21009,N_21690);
nor U22123 (N_22123,N_20574,N_20535);
or U22124 (N_22124,N_20929,N_21535);
or U22125 (N_22125,N_20001,N_20007);
and U22126 (N_22126,N_20191,N_20286);
or U22127 (N_22127,N_20905,N_21021);
nor U22128 (N_22128,N_20995,N_21499);
xor U22129 (N_22129,N_20964,N_20661);
or U22130 (N_22130,N_21337,N_20866);
nor U22131 (N_22131,N_20019,N_21094);
nand U22132 (N_22132,N_20341,N_20977);
nor U22133 (N_22133,N_21711,N_21325);
nor U22134 (N_22134,N_20809,N_20058);
nand U22135 (N_22135,N_21338,N_21993);
or U22136 (N_22136,N_20066,N_20799);
nand U22137 (N_22137,N_21526,N_21991);
xor U22138 (N_22138,N_21843,N_21688);
or U22139 (N_22139,N_21571,N_20738);
nand U22140 (N_22140,N_21766,N_20613);
xnor U22141 (N_22141,N_20331,N_21628);
xnor U22142 (N_22142,N_21068,N_20023);
xnor U22143 (N_22143,N_20248,N_21724);
or U22144 (N_22144,N_21979,N_21184);
nand U22145 (N_22145,N_20882,N_20634);
nand U22146 (N_22146,N_21932,N_21907);
xor U22147 (N_22147,N_21970,N_20258);
or U22148 (N_22148,N_20487,N_20122);
and U22149 (N_22149,N_20265,N_21866);
and U22150 (N_22150,N_20184,N_20602);
nand U22151 (N_22151,N_20889,N_21524);
and U22152 (N_22152,N_20391,N_20203);
xor U22153 (N_22153,N_20681,N_21150);
or U22154 (N_22154,N_21623,N_20300);
nor U22155 (N_22155,N_20082,N_20963);
nor U22156 (N_22156,N_21830,N_21398);
and U22157 (N_22157,N_21048,N_20369);
xnor U22158 (N_22158,N_21821,N_21108);
and U22159 (N_22159,N_21778,N_20699);
and U22160 (N_22160,N_21749,N_20015);
or U22161 (N_22161,N_21468,N_20584);
xnor U22162 (N_22162,N_21215,N_20797);
nand U22163 (N_22163,N_20790,N_20745);
nand U22164 (N_22164,N_20668,N_21106);
and U22165 (N_22165,N_20085,N_20676);
and U22166 (N_22166,N_20011,N_21417);
or U22167 (N_22167,N_20059,N_20152);
or U22168 (N_22168,N_20419,N_20787);
and U22169 (N_22169,N_20617,N_20462);
nand U22170 (N_22170,N_20752,N_20107);
nor U22171 (N_22171,N_20941,N_21940);
and U22172 (N_22172,N_20662,N_21063);
nand U22173 (N_22173,N_21086,N_21600);
nand U22174 (N_22174,N_20459,N_21885);
or U22175 (N_22175,N_20514,N_21538);
and U22176 (N_22176,N_20140,N_20372);
or U22177 (N_22177,N_21649,N_20317);
nand U22178 (N_22178,N_20546,N_21840);
and U22179 (N_22179,N_20740,N_20970);
xnor U22180 (N_22180,N_21224,N_20200);
nor U22181 (N_22181,N_21070,N_20181);
nor U22182 (N_22182,N_20493,N_21259);
nand U22183 (N_22183,N_20565,N_21202);
nand U22184 (N_22184,N_20022,N_20148);
nor U22185 (N_22185,N_20497,N_20890);
or U22186 (N_22186,N_21505,N_21809);
or U22187 (N_22187,N_21810,N_20665);
xor U22188 (N_22188,N_21255,N_21409);
nand U22189 (N_22189,N_20109,N_21218);
nor U22190 (N_22190,N_21121,N_21096);
nor U22191 (N_22191,N_20166,N_21038);
nor U22192 (N_22192,N_21517,N_21130);
and U22193 (N_22193,N_20932,N_21805);
xnor U22194 (N_22194,N_20310,N_21658);
and U22195 (N_22195,N_20707,N_20269);
nand U22196 (N_22196,N_21823,N_21358);
nand U22197 (N_22197,N_20801,N_21675);
nor U22198 (N_22198,N_21996,N_20806);
xnor U22199 (N_22199,N_20373,N_20367);
or U22200 (N_22200,N_21167,N_21160);
xnor U22201 (N_22201,N_21482,N_20115);
nand U22202 (N_22202,N_20635,N_21732);
xnor U22203 (N_22203,N_21621,N_20581);
nand U22204 (N_22204,N_21206,N_21326);
xor U22205 (N_22205,N_21529,N_21334);
nor U22206 (N_22206,N_21448,N_20753);
nand U22207 (N_22207,N_21992,N_20524);
xnor U22208 (N_22208,N_21473,N_21857);
and U22209 (N_22209,N_20701,N_20956);
xnor U22210 (N_22210,N_20654,N_20256);
nor U22211 (N_22211,N_20561,N_20446);
nor U22212 (N_22212,N_20219,N_21910);
or U22213 (N_22213,N_21457,N_21464);
and U22214 (N_22214,N_21075,N_20875);
xor U22215 (N_22215,N_21222,N_20068);
xnor U22216 (N_22216,N_20480,N_21423);
or U22217 (N_22217,N_20348,N_21320);
and U22218 (N_22218,N_21053,N_21427);
nor U22219 (N_22219,N_21834,N_21936);
and U22220 (N_22220,N_21186,N_21568);
xor U22221 (N_22221,N_21546,N_21510);
or U22222 (N_22222,N_21290,N_21678);
or U22223 (N_22223,N_21583,N_20026);
nand U22224 (N_22224,N_21142,N_21383);
nand U22225 (N_22225,N_20533,N_21858);
and U22226 (N_22226,N_20380,N_20819);
or U22227 (N_22227,N_21470,N_20186);
xnor U22228 (N_22228,N_21231,N_21817);
nor U22229 (N_22229,N_20624,N_21407);
and U22230 (N_22230,N_20800,N_20918);
xor U22231 (N_22231,N_21961,N_21056);
nor U22232 (N_22232,N_21570,N_20767);
and U22233 (N_22233,N_21620,N_20358);
xor U22234 (N_22234,N_20072,N_20671);
nand U22235 (N_22235,N_20588,N_21990);
nor U22236 (N_22236,N_21860,N_21236);
or U22237 (N_22237,N_20409,N_20347);
nand U22238 (N_22238,N_21848,N_20814);
nor U22239 (N_22239,N_20050,N_20376);
xor U22240 (N_22240,N_20159,N_21997);
nand U22241 (N_22241,N_20461,N_20368);
nor U22242 (N_22242,N_20714,N_21755);
nand U22243 (N_22243,N_20339,N_20292);
and U22244 (N_22244,N_20065,N_21741);
nor U22245 (N_22245,N_21602,N_20336);
or U22246 (N_22246,N_21560,N_20512);
xnor U22247 (N_22247,N_20886,N_21567);
or U22248 (N_22248,N_20363,N_20868);
or U22249 (N_22249,N_21984,N_21607);
nor U22250 (N_22250,N_20284,N_21052);
nor U22251 (N_22251,N_20163,N_21281);
or U22252 (N_22252,N_21935,N_21625);
or U22253 (N_22253,N_20083,N_21346);
nand U22254 (N_22254,N_21684,N_20732);
nand U22255 (N_22255,N_21553,N_20123);
nor U22256 (N_22256,N_21704,N_20769);
or U22257 (N_22257,N_20403,N_21363);
nor U22258 (N_22258,N_20547,N_21115);
nand U22259 (N_22259,N_21837,N_21674);
nand U22260 (N_22260,N_21304,N_21698);
xnor U22261 (N_22261,N_20017,N_21751);
nor U22262 (N_22262,N_20669,N_20173);
xnor U22263 (N_22263,N_20975,N_20763);
nor U22264 (N_22264,N_21177,N_20674);
and U22265 (N_22265,N_21402,N_21155);
nand U22266 (N_22266,N_20104,N_21677);
and U22267 (N_22267,N_20686,N_21767);
and U22268 (N_22268,N_20794,N_20112);
nor U22269 (N_22269,N_20183,N_20733);
nand U22270 (N_22270,N_21951,N_21850);
or U22271 (N_22271,N_21827,N_20389);
or U22272 (N_22272,N_21060,N_21947);
nor U22273 (N_22273,N_21455,N_21855);
xor U22274 (N_22274,N_21345,N_20000);
xnor U22275 (N_22275,N_20703,N_20042);
or U22276 (N_22276,N_20047,N_21256);
nor U22277 (N_22277,N_20087,N_21066);
or U22278 (N_22278,N_20962,N_21340);
or U22279 (N_22279,N_20813,N_20415);
or U22280 (N_22280,N_20260,N_21199);
nor U22281 (N_22281,N_20364,N_20247);
nor U22282 (N_22282,N_21513,N_20855);
and U22283 (N_22283,N_21636,N_21011);
xnor U22284 (N_22284,N_20508,N_20860);
xor U22285 (N_22285,N_20754,N_21554);
nand U22286 (N_22286,N_21605,N_21648);
xor U22287 (N_22287,N_21116,N_20593);
xnor U22288 (N_22288,N_21710,N_20596);
or U22289 (N_22289,N_21983,N_20078);
and U22290 (N_22290,N_20755,N_21258);
or U22291 (N_22291,N_21950,N_21574);
nor U22292 (N_22292,N_20201,N_20563);
or U22293 (N_22293,N_20177,N_20037);
nor U22294 (N_22294,N_21503,N_21773);
nand U22295 (N_22295,N_21077,N_21219);
or U22296 (N_22296,N_21534,N_20725);
xor U22297 (N_22297,N_20252,N_21938);
nand U22298 (N_22298,N_20444,N_20916);
and U22299 (N_22299,N_21045,N_21693);
xor U22300 (N_22300,N_21786,N_20051);
and U22301 (N_22301,N_20021,N_21701);
nor U22302 (N_22302,N_21360,N_20859);
xnor U22303 (N_22303,N_21204,N_20440);
nor U22304 (N_22304,N_21692,N_21187);
and U22305 (N_22305,N_20379,N_20481);
xnor U22306 (N_22306,N_20285,N_20935);
nand U22307 (N_22307,N_20154,N_21251);
nand U22308 (N_22308,N_21995,N_20333);
nand U22309 (N_22309,N_20129,N_20987);
nand U22310 (N_22310,N_20053,N_21284);
or U22311 (N_22311,N_21739,N_20180);
nand U22312 (N_22312,N_21467,N_21135);
or U22313 (N_22313,N_20209,N_20095);
nand U22314 (N_22314,N_20116,N_20812);
nor U22315 (N_22315,N_21303,N_21306);
or U22316 (N_22316,N_20153,N_20067);
nor U22317 (N_22317,N_20578,N_20128);
nand U22318 (N_22318,N_20254,N_21169);
nor U22319 (N_22319,N_20908,N_20080);
nor U22320 (N_22320,N_21915,N_20678);
and U22321 (N_22321,N_21182,N_21978);
nor U22322 (N_22322,N_21107,N_21263);
and U22323 (N_22323,N_20909,N_20967);
nor U22324 (N_22324,N_21049,N_21158);
nand U22325 (N_22325,N_20298,N_21776);
nor U22326 (N_22326,N_20959,N_21028);
nor U22327 (N_22327,N_20783,N_20871);
or U22328 (N_22328,N_21432,N_21162);
and U22329 (N_22329,N_21799,N_21143);
or U22330 (N_22330,N_20509,N_20949);
nor U22331 (N_22331,N_20572,N_21181);
xnor U22332 (N_22332,N_20325,N_21120);
xnor U22333 (N_22333,N_21667,N_21452);
or U22334 (N_22334,N_20395,N_21272);
nor U22335 (N_22335,N_20084,N_21497);
nand U22336 (N_22336,N_21742,N_21516);
xnor U22337 (N_22337,N_20709,N_20867);
nand U22338 (N_22338,N_21373,N_20225);
and U22339 (N_22339,N_20472,N_20335);
xor U22340 (N_22340,N_20384,N_21532);
or U22341 (N_22341,N_20684,N_21171);
xor U22342 (N_22342,N_21521,N_21033);
or U22343 (N_22343,N_21424,N_21849);
and U22344 (N_22344,N_20735,N_21889);
nand U22345 (N_22345,N_21490,N_21515);
nor U22346 (N_22346,N_21727,N_21919);
or U22347 (N_22347,N_20429,N_20246);
nor U22348 (N_22348,N_21969,N_20155);
and U22349 (N_22349,N_21835,N_21787);
nand U22350 (N_22350,N_21933,N_21454);
nand U22351 (N_22351,N_20771,N_20272);
nand U22352 (N_22352,N_20532,N_21509);
or U22353 (N_22353,N_21707,N_20375);
and U22354 (N_22354,N_21543,N_20436);
or U22355 (N_22355,N_21234,N_20465);
nand U22356 (N_22356,N_20527,N_20505);
or U22357 (N_22357,N_20382,N_20450);
or U22358 (N_22358,N_20274,N_20397);
or U22359 (N_22359,N_20057,N_20837);
or U22360 (N_22360,N_20972,N_21292);
or U22361 (N_22361,N_20228,N_20550);
and U22362 (N_22362,N_20537,N_20897);
and U22363 (N_22363,N_20664,N_21634);
or U22364 (N_22364,N_21283,N_21469);
nor U22365 (N_22365,N_20762,N_20340);
nor U22366 (N_22366,N_20553,N_21074);
nor U22367 (N_22367,N_20273,N_21232);
nor U22368 (N_22368,N_21831,N_20729);
xnor U22369 (N_22369,N_20944,N_21924);
xnor U22370 (N_22370,N_20630,N_21065);
nor U22371 (N_22371,N_20434,N_20716);
xor U22372 (N_22372,N_20774,N_20070);
and U22373 (N_22373,N_21729,N_20796);
and U22374 (N_22374,N_20833,N_20570);
and U22375 (N_22375,N_21737,N_20607);
and U22376 (N_22376,N_21657,N_21370);
and U22377 (N_22377,N_21507,N_21721);
nor U22378 (N_22378,N_20823,N_21547);
nor U22379 (N_22379,N_21880,N_20777);
xnor U22380 (N_22380,N_21592,N_21088);
xnor U22381 (N_22381,N_21456,N_20931);
and U22382 (N_22382,N_20330,N_20840);
nand U22383 (N_22383,N_20585,N_21235);
xnor U22384 (N_22384,N_21609,N_21291);
xor U22385 (N_22385,N_21100,N_20071);
and U22386 (N_22386,N_20552,N_20748);
and U22387 (N_22387,N_21654,N_21382);
nand U22388 (N_22388,N_21321,N_21472);
nor U22389 (N_22389,N_21916,N_20915);
nor U22390 (N_22390,N_21085,N_20880);
and U22391 (N_22391,N_20571,N_20632);
nand U22392 (N_22392,N_21477,N_21895);
or U22393 (N_22393,N_20597,N_21890);
nor U22394 (N_22394,N_21930,N_21428);
nor U22395 (N_22395,N_20178,N_20390);
nand U22396 (N_22396,N_21528,N_20672);
or U22397 (N_22397,N_21311,N_20592);
and U22398 (N_22398,N_20160,N_20736);
nor U22399 (N_22399,N_21149,N_20016);
or U22400 (N_22400,N_20971,N_21929);
nor U22401 (N_22401,N_20704,N_20230);
xnor U22402 (N_22402,N_20054,N_21679);
nand U22403 (N_22403,N_20930,N_20721);
or U22404 (N_22404,N_20093,N_21000);
nand U22405 (N_22405,N_20515,N_20887);
nor U22406 (N_22406,N_21453,N_21945);
and U22407 (N_22407,N_20214,N_20639);
xnor U22408 (N_22408,N_21781,N_20655);
or U22409 (N_22409,N_20474,N_21165);
or U22410 (N_22410,N_21813,N_20642);
xnor U22411 (N_22411,N_20718,N_21591);
nor U22412 (N_22412,N_20960,N_20060);
xor U22413 (N_22413,N_20179,N_21811);
and U22414 (N_22414,N_21189,N_20722);
xor U22415 (N_22415,N_21844,N_21122);
nor U22416 (N_22416,N_20785,N_20197);
nor U22417 (N_22417,N_21125,N_21376);
xor U22418 (N_22418,N_21391,N_20234);
nor U22419 (N_22419,N_20792,N_20473);
and U22420 (N_22420,N_21297,N_21114);
xor U22421 (N_22421,N_20305,N_21163);
nor U22422 (N_22422,N_21216,N_20947);
nor U22423 (N_22423,N_20412,N_20951);
and U22424 (N_22424,N_21622,N_20892);
and U22425 (N_22425,N_20268,N_20328);
and U22426 (N_22426,N_20271,N_20857);
or U22427 (N_22427,N_21078,N_20969);
nand U22428 (N_22428,N_20287,N_20657);
or U22429 (N_22429,N_21223,N_21449);
and U22430 (N_22430,N_20435,N_21593);
nand U22431 (N_22431,N_20791,N_20135);
or U22432 (N_22432,N_20599,N_21709);
or U22433 (N_22433,N_20507,N_20646);
and U22434 (N_22434,N_20130,N_21064);
nand U22435 (N_22435,N_20124,N_20401);
or U22436 (N_22436,N_20934,N_21533);
nand U22437 (N_22437,N_20400,N_20548);
and U22438 (N_22438,N_21388,N_21371);
nor U22439 (N_22439,N_20843,N_20525);
and U22440 (N_22440,N_21743,N_21820);
or U22441 (N_22441,N_21315,N_21073);
and U22442 (N_22442,N_21211,N_20611);
and U22443 (N_22443,N_20118,N_21318);
xor U22444 (N_22444,N_20750,N_21877);
nor U22445 (N_22445,N_21829,N_20551);
or U22446 (N_22446,N_21879,N_20877);
or U22447 (N_22447,N_20405,N_21788);
xor U22448 (N_22448,N_20018,N_20764);
nor U22449 (N_22449,N_21007,N_20216);
or U22450 (N_22450,N_21462,N_21494);
or U22451 (N_22451,N_20049,N_20356);
xor U22452 (N_22452,N_21986,N_20222);
or U22453 (N_22453,N_20442,N_20293);
or U22454 (N_22454,N_20312,N_20950);
and U22455 (N_22455,N_20233,N_20720);
or U22456 (N_22456,N_20708,N_21752);
nor U22457 (N_22457,N_21894,N_20589);
nor U22458 (N_22458,N_20999,N_21753);
nor U22459 (N_22459,N_20120,N_20914);
xor U22460 (N_22460,N_20279,N_21557);
and U22461 (N_22461,N_21824,N_20321);
and U22462 (N_22462,N_21071,N_21495);
nand U22463 (N_22463,N_21659,N_21148);
or U22464 (N_22464,N_20189,N_21795);
xor U22465 (N_22465,N_20603,N_20161);
nor U22466 (N_22466,N_21587,N_20301);
or U22467 (N_22467,N_20788,N_20510);
or U22468 (N_22468,N_20531,N_21422);
xnor U22469 (N_22469,N_21396,N_20878);
nor U22470 (N_22470,N_20498,N_20986);
nand U22471 (N_22471,N_21798,N_20366);
xnor U22472 (N_22472,N_20454,N_20484);
nor U22473 (N_22473,N_20466,N_20776);
and U22474 (N_22474,N_21061,N_21353);
xor U22475 (N_22475,N_21595,N_21024);
nor U22476 (N_22476,N_20458,N_21414);
nor U22477 (N_22477,N_20779,N_21931);
or U22478 (N_22478,N_21578,N_20820);
nand U22479 (N_22479,N_21349,N_20598);
or U22480 (N_22480,N_21123,N_21134);
and U22481 (N_22481,N_21351,N_20683);
xor U22482 (N_22482,N_21463,N_20451);
xor U22483 (N_22483,N_20127,N_20647);
nor U22484 (N_22484,N_21964,N_21314);
or U22485 (N_22485,N_20239,N_21572);
xnor U22486 (N_22486,N_21926,N_20311);
xor U22487 (N_22487,N_20038,N_20147);
or U22488 (N_22488,N_21084,N_21888);
or U22489 (N_22489,N_20540,N_20096);
or U22490 (N_22490,N_21164,N_21792);
or U22491 (N_22491,N_20027,N_20036);
nor U22492 (N_22492,N_21278,N_20706);
nor U22493 (N_22493,N_21418,N_21020);
xnor U22494 (N_22494,N_20167,N_20888);
and U22495 (N_22495,N_21508,N_21335);
nand U22496 (N_22496,N_21613,N_21682);
nand U22497 (N_22497,N_21397,N_21856);
or U22498 (N_22498,N_20804,N_21246);
xnor U22499 (N_22499,N_20901,N_20211);
nand U22500 (N_22500,N_21873,N_20056);
or U22501 (N_22501,N_21341,N_21016);
or U22502 (N_22502,N_20357,N_21957);
nand U22503 (N_22503,N_20691,N_21635);
and U22504 (N_22504,N_21225,N_20715);
and U22505 (N_22505,N_20815,N_20680);
or U22506 (N_22506,N_20138,N_20437);
nand U22507 (N_22507,N_21270,N_20119);
and U22508 (N_22508,N_20575,N_21540);
nor U22509 (N_22509,N_20621,N_20121);
nand U22510 (N_22510,N_21610,N_21774);
xor U22511 (N_22511,N_21271,N_21378);
nor U22512 (N_22512,N_20232,N_20658);
nor U22513 (N_22513,N_21715,N_20431);
xnor U22514 (N_22514,N_21959,N_21796);
nor U22515 (N_22515,N_21145,N_21128);
xor U22516 (N_22516,N_21312,N_20852);
and U22517 (N_22517,N_20169,N_20488);
nor U22518 (N_22518,N_21082,N_21920);
nor U22519 (N_22519,N_21437,N_20610);
or U22520 (N_22520,N_21973,N_21156);
nand U22521 (N_22521,N_21392,N_21580);
nor U22522 (N_22522,N_20851,N_20922);
xor U22523 (N_22523,N_21934,N_20443);
xor U22524 (N_22524,N_21026,N_21734);
nand U22525 (N_22525,N_20378,N_20928);
nor U22526 (N_22526,N_20782,N_21443);
nor U22527 (N_22527,N_21584,N_21968);
nor U22528 (N_22528,N_20267,N_20711);
and U22529 (N_22529,N_21536,N_20902);
nand U22530 (N_22530,N_21459,N_21669);
nand U22531 (N_22531,N_20549,N_20925);
and U22532 (N_22532,N_20125,N_20206);
nor U22533 (N_22533,N_20591,N_21539);
and U22534 (N_22534,N_20468,N_21645);
or U22535 (N_22535,N_21559,N_21299);
or U22536 (N_22536,N_20452,N_21372);
and U22537 (N_22537,N_20025,N_20276);
xor U22538 (N_22538,N_20029,N_21265);
nor U22539 (N_22539,N_21589,N_20413);
xor U22540 (N_22540,N_21551,N_20545);
nand U22541 (N_22541,N_21047,N_20424);
or U22542 (N_22542,N_21705,N_20536);
nand U22543 (N_22543,N_21660,N_21298);
nor U22544 (N_22544,N_20308,N_21110);
nor U22545 (N_22545,N_21076,N_20319);
nand U22546 (N_22546,N_21377,N_21451);
nand U22547 (N_22547,N_21460,N_21646);
nand U22548 (N_22548,N_21029,N_20737);
or U22549 (N_22549,N_20486,N_20235);
nor U22550 (N_22550,N_20004,N_20694);
or U22551 (N_22551,N_20176,N_20353);
and U22552 (N_22552,N_21180,N_20538);
nand U22553 (N_22553,N_21596,N_20974);
nor U22554 (N_22554,N_20220,N_20789);
nor U22555 (N_22555,N_21681,N_20099);
nand U22556 (N_22556,N_21413,N_21379);
or U22557 (N_22557,N_20957,N_20041);
xor U22558 (N_22558,N_20221,N_21203);
and U22559 (N_22559,N_21624,N_21027);
nor U22560 (N_22560,N_21385,N_20609);
nor U22561 (N_22561,N_21952,N_20863);
nor U22562 (N_22562,N_20187,N_21683);
nor U22563 (N_22563,N_20165,N_20145);
xnor U22564 (N_22564,N_20238,N_20236);
nand U22565 (N_22565,N_21286,N_21722);
or U22566 (N_22566,N_20608,N_21925);
nor U22567 (N_22567,N_20289,N_20103);
or U22568 (N_22568,N_21498,N_21333);
and U22569 (N_22569,N_21836,N_21367);
nand U22570 (N_22570,N_21332,N_21579);
nor U22571 (N_22571,N_21577,N_21366);
xnor U22572 (N_22572,N_21685,N_20619);
and U22573 (N_22573,N_21833,N_21871);
nand U22574 (N_22574,N_21504,N_21319);
nand U22575 (N_22575,N_21205,N_21003);
xnor U22576 (N_22576,N_21238,N_20579);
nor U22577 (N_22577,N_20894,N_20828);
xor U22578 (N_22578,N_20420,N_21226);
xor U22579 (N_22579,N_21381,N_20670);
nor U22580 (N_22580,N_21761,N_21812);
xor U22581 (N_22581,N_20501,N_20489);
xor U22582 (N_22582,N_21826,N_20600);
xnor U22583 (N_22583,N_20985,N_20911);
xnor U22584 (N_22584,N_21760,N_20696);
or U22585 (N_22585,N_21867,N_20690);
or U22586 (N_22586,N_20557,N_20528);
or U22587 (N_22587,N_20924,N_21072);
xnor U22588 (N_22588,N_21853,N_20393);
xnor U22589 (N_22589,N_21793,N_21586);
nor U22590 (N_22590,N_21273,N_21471);
xor U22591 (N_22591,N_21387,N_20879);
and U22592 (N_22592,N_20688,N_20637);
xor U22593 (N_22593,N_21389,N_21213);
or U22594 (N_22594,N_20982,N_20993);
xnor U22595 (N_22595,N_20817,N_20781);
and U22596 (N_22596,N_20641,N_21117);
or U22597 (N_22597,N_20891,N_20978);
or U22598 (N_22598,N_20043,N_21146);
nor U22599 (N_22599,N_20604,N_21977);
xnor U22600 (N_22600,N_21791,N_21364);
or U22601 (N_22601,N_21652,N_20476);
nor U22602 (N_22602,N_21763,N_21046);
nand U22603 (N_22603,N_20544,N_21881);
nand U22604 (N_22604,N_21542,N_20907);
xor U22605 (N_22605,N_21687,N_20495);
nor U22606 (N_22606,N_20406,N_20543);
nand U22607 (N_22607,N_20351,N_20081);
nor U22608 (N_22608,N_21458,N_20832);
or U22609 (N_22609,N_20802,N_21882);
xor U22610 (N_22610,N_21386,N_20730);
nand U22611 (N_22611,N_21708,N_21887);
and U22612 (N_22612,N_20377,N_21118);
and U22613 (N_22613,N_21723,N_20990);
or U22614 (N_22614,N_21253,N_20302);
or U22615 (N_22615,N_21302,N_21832);
and U22616 (N_22616,N_20332,N_20826);
and U22617 (N_22617,N_20541,N_20309);
and U22618 (N_22618,N_21909,N_20283);
nand U22619 (N_22619,N_20077,N_21197);
and U22620 (N_22620,N_21361,N_21055);
nand U22621 (N_22621,N_21137,N_21903);
nand U22622 (N_22622,N_21745,N_21514);
nor U22623 (N_22623,N_20521,N_21606);
xnor U22624 (N_22624,N_21067,N_20784);
or U22625 (N_22625,N_20061,N_21998);
xnor U22626 (N_22626,N_21772,N_20580);
xnor U22627 (N_22627,N_20240,N_20387);
or U22628 (N_22628,N_21446,N_21244);
nor U22629 (N_22629,N_20595,N_21119);
and U22630 (N_22630,N_20024,N_20558);
nor U22631 (N_22631,N_20040,N_21851);
and U22632 (N_22632,N_20288,N_20212);
or U22633 (N_22633,N_21269,N_20030);
xnor U22634 (N_22634,N_21058,N_20940);
nand U22635 (N_22635,N_20196,N_21405);
xnor U22636 (N_22636,N_20213,N_21558);
xnor U22637 (N_22637,N_21083,N_20482);
nand U22638 (N_22638,N_20360,N_20836);
nand U22639 (N_22639,N_21069,N_21354);
nor U22640 (N_22640,N_20076,N_20411);
xnor U22641 (N_22641,N_21564,N_21295);
nand U22642 (N_22642,N_21001,N_21344);
xor U22643 (N_22643,N_21436,N_21902);
xnor U22644 (N_22644,N_21174,N_21093);
nor U22645 (N_22645,N_20614,N_20048);
and U22646 (N_22646,N_20757,N_21619);
or U22647 (N_22647,N_20231,N_20644);
and U22648 (N_22648,N_21489,N_20438);
or U22649 (N_22649,N_21981,N_20349);
and U22650 (N_22650,N_20052,N_21962);
and U22651 (N_22651,N_21097,N_21322);
and U22652 (N_22652,N_20955,N_21590);
nor U22653 (N_22653,N_21380,N_21274);
nand U22654 (N_22654,N_20760,N_21905);
xor U22655 (N_22655,N_21368,N_21252);
or U22656 (N_22656,N_20848,N_20075);
nand U22657 (N_22657,N_20793,N_21352);
or U22658 (N_22658,N_20858,N_21229);
and U22659 (N_22659,N_20953,N_20810);
and U22660 (N_22660,N_21237,N_21982);
and U22661 (N_22661,N_21267,N_20679);
nor U22662 (N_22662,N_20046,N_21728);
or U22663 (N_22663,N_20573,N_21937);
xor U22664 (N_22664,N_20477,N_20013);
and U22665 (N_22665,N_21697,N_21198);
nand U22666 (N_22666,N_21481,N_20751);
or U22667 (N_22667,N_20994,N_21492);
or U22668 (N_22668,N_21112,N_21091);
nor U22669 (N_22669,N_20110,N_21900);
or U22670 (N_22670,N_21550,N_20623);
xor U22671 (N_22671,N_20304,N_21691);
xnor U22672 (N_22672,N_21627,N_20303);
or U22673 (N_22673,N_21488,N_21347);
nor U22674 (N_22674,N_21942,N_21266);
nor U22675 (N_22675,N_21357,N_20150);
or U22676 (N_22676,N_20650,N_21276);
nand U22677 (N_22677,N_21331,N_21914);
and U22678 (N_22678,N_20900,N_20648);
and U22679 (N_22679,N_20846,N_21031);
nand U22680 (N_22680,N_20517,N_20761);
xnor U22681 (N_22681,N_20698,N_20242);
nor U22682 (N_22682,N_21300,N_20031);
nand U22683 (N_22683,N_21638,N_20893);
or U22684 (N_22684,N_21442,N_20896);
xor U22685 (N_22685,N_20590,N_21476);
or U22686 (N_22686,N_20417,N_20862);
and U22687 (N_22687,N_21555,N_21330);
or U22688 (N_22688,N_20825,N_20569);
or U22689 (N_22689,N_21941,N_20418);
nand U22690 (N_22690,N_21573,N_20937);
nor U22691 (N_22691,N_21151,N_20404);
xor U22692 (N_22692,N_21480,N_21519);
xnor U22693 (N_22693,N_20383,N_20917);
nor U22694 (N_22694,N_21113,N_20695);
nor U22695 (N_22695,N_21013,N_20359);
nand U22696 (N_22696,N_21756,N_20063);
or U22697 (N_22697,N_21859,N_21531);
or U22698 (N_22698,N_20731,N_20511);
nor U22699 (N_22699,N_20520,N_21642);
or U22700 (N_22700,N_21548,N_20811);
xnor U22701 (N_22701,N_20895,N_21549);
or U22702 (N_22702,N_21485,N_21838);
nand U22703 (N_22703,N_21109,N_21616);
nand U22704 (N_22704,N_21207,N_20006);
xor U22705 (N_22705,N_21736,N_20270);
nand U22706 (N_22706,N_20394,N_21416);
and U22707 (N_22707,N_20014,N_20346);
nor U22708 (N_22708,N_21444,N_21780);
xnor U22709 (N_22709,N_21327,N_20739);
nor U22710 (N_22710,N_20494,N_21971);
or U22711 (N_22711,N_21730,N_21944);
and U22712 (N_22712,N_20136,N_21870);
nor U22713 (N_22713,N_21129,N_21261);
and U22714 (N_22714,N_21923,N_20028);
nor U22715 (N_22715,N_20542,N_20218);
and U22716 (N_22716,N_21103,N_20881);
and U22717 (N_22717,N_21672,N_21209);
or U22718 (N_22718,N_20210,N_20568);
nor U22719 (N_22719,N_20747,N_20491);
nor U22720 (N_22720,N_21102,N_20483);
and U22721 (N_22721,N_21280,N_21014);
nor U22722 (N_22722,N_20719,N_20005);
nor U22723 (N_22723,N_21670,N_20455);
xnor U22724 (N_22724,N_21631,N_21355);
or U22725 (N_22725,N_20414,N_21974);
and U22726 (N_22726,N_20094,N_20249);
and U22727 (N_22727,N_21441,N_21601);
nor U22728 (N_22728,N_20724,N_20968);
nand U22729 (N_22729,N_21041,N_21313);
xor U22730 (N_22730,N_20323,N_21861);
or U22731 (N_22731,N_20560,N_20687);
and U22732 (N_22732,N_20432,N_21913);
xnor U22733 (N_22733,N_20374,N_21948);
nor U22734 (N_22734,N_20723,N_21401);
xor U22735 (N_22735,N_21544,N_20923);
and U22736 (N_22736,N_20702,N_20936);
xor U22737 (N_22737,N_21803,N_20864);
and U22738 (N_22738,N_21630,N_20133);
or U22739 (N_22739,N_20506,N_20622);
and U22740 (N_22740,N_21530,N_21139);
and U22741 (N_22741,N_20185,N_21748);
and U22742 (N_22742,N_21972,N_21176);
nor U22743 (N_22743,N_20496,N_20744);
nand U22744 (N_22744,N_21159,N_21569);
nor U22745 (N_22745,N_20324,N_20257);
nand U22746 (N_22746,N_21288,N_21153);
or U22747 (N_22747,N_20192,N_20898);
or U22748 (N_22748,N_20156,N_20996);
or U22749 (N_22749,N_21439,N_20079);
and U22750 (N_22750,N_21307,N_21651);
xor U22751 (N_22751,N_20416,N_21764);
and U22752 (N_22752,N_21512,N_21339);
or U22753 (N_22753,N_21500,N_20816);
nand U22754 (N_22754,N_20139,N_21002);
and U22755 (N_22755,N_21712,N_21575);
or U22756 (N_22756,N_20295,N_21663);
nand U22757 (N_22757,N_21664,N_21043);
nor U22758 (N_22758,N_21854,N_20074);
or U22759 (N_22759,N_21604,N_21845);
nand U22760 (N_22760,N_21874,N_20146);
and U22761 (N_22761,N_21328,N_21740);
xnor U22762 (N_22762,N_21878,N_21917);
nor U22763 (N_22763,N_21720,N_21912);
xor U22764 (N_22764,N_20945,N_20979);
and U22765 (N_22765,N_20586,N_20628);
nand U22766 (N_22766,N_20502,N_21147);
and U22767 (N_22767,N_20504,N_20098);
nand U22768 (N_22768,N_20556,N_20976);
nand U22769 (N_22769,N_20207,N_20361);
nor U22770 (N_22770,N_21896,N_21901);
nand U22771 (N_22771,N_21758,N_21210);
and U22772 (N_22772,N_20838,N_21157);
nor U22773 (N_22773,N_20835,N_21408);
xor U22774 (N_22774,N_21713,N_21662);
nor U22775 (N_22775,N_20297,N_20427);
or U22776 (N_22776,N_20277,N_21411);
and U22777 (N_22777,N_21561,N_20522);
xnor U22778 (N_22778,N_20263,N_20849);
xnor U22779 (N_22779,N_21316,N_20606);
xor U22780 (N_22780,N_21042,N_20856);
nand U22781 (N_22781,N_21911,N_21563);
or U22782 (N_22782,N_21846,N_21039);
and U22783 (N_22783,N_20876,N_21594);
and U22784 (N_22784,N_20281,N_21585);
and U22785 (N_22785,N_21431,N_20830);
nor U22786 (N_22786,N_21966,N_20010);
nand U22787 (N_22787,N_20202,N_20692);
and U22788 (N_22788,N_20673,N_20577);
nor U22789 (N_22789,N_21694,N_20168);
nor U22790 (N_22790,N_21980,N_21759);
nor U22791 (N_22791,N_20251,N_20728);
xor U22792 (N_22792,N_20854,N_21976);
nor U22793 (N_22793,N_21899,N_21350);
xnor U22794 (N_22794,N_20467,N_20861);
nor U22795 (N_22795,N_20954,N_21985);
or U22796 (N_22796,N_20195,N_21170);
nand U22797 (N_22797,N_21884,N_20587);
and U22798 (N_22798,N_20291,N_20652);
or U22799 (N_22799,N_20456,N_20601);
or U22800 (N_22800,N_21552,N_20343);
nor U22801 (N_22801,N_21864,N_20518);
xnor U22802 (N_22802,N_21598,N_20927);
xnor U22803 (N_22803,N_20989,N_21807);
and U22804 (N_22804,N_21275,N_21309);
xor U22805 (N_22805,N_21626,N_21875);
xnor U22806 (N_22806,N_20727,N_20966);
xor U22807 (N_22807,N_20117,N_20362);
nor U22808 (N_22808,N_21025,N_20469);
or U22809 (N_22809,N_20266,N_20243);
nand U22810 (N_22810,N_20322,N_21305);
xor U22811 (N_22811,N_21404,N_21406);
xor U22812 (N_22812,N_21375,N_21196);
nand U22813 (N_22813,N_20803,N_20645);
and U22814 (N_22814,N_21965,N_20355);
or U22815 (N_22815,N_21161,N_21131);
xor U22816 (N_22816,N_20217,N_21815);
and U22817 (N_22817,N_20262,N_21522);
xnor U22818 (N_22818,N_21393,N_20092);
and U22819 (N_22819,N_21650,N_21738);
nor U22820 (N_22820,N_21034,N_20798);
nand U22821 (N_22821,N_20069,N_21641);
nor U22822 (N_22822,N_21695,N_20408);
nor U22823 (N_22823,N_20345,N_20320);
nor U22824 (N_22824,N_21800,N_20910);
and U22825 (N_22825,N_20824,N_20765);
nand U22826 (N_22826,N_21192,N_20939);
xor U22827 (N_22827,N_21050,N_21581);
xor U22828 (N_22828,N_21260,N_20656);
xor U22829 (N_22829,N_21872,N_20478);
and U22830 (N_22830,N_21545,N_20566);
nand U22831 (N_22831,N_20758,N_21491);
nor U22832 (N_22832,N_20294,N_20114);
and U22833 (N_22833,N_21079,N_20275);
or U22834 (N_22834,N_20350,N_20853);
nand U22835 (N_22835,N_21092,N_20250);
xor U22836 (N_22836,N_20874,N_21918);
nor U22837 (N_22837,N_21921,N_20421);
xnor U22838 (N_22838,N_21296,N_21175);
or U22839 (N_22839,N_21032,N_20933);
or U22840 (N_22840,N_20594,N_20770);
xor U22841 (N_22841,N_21059,N_21725);
or U22842 (N_22842,N_21496,N_21770);
and U22843 (N_22843,N_20884,N_21523);
or U22844 (N_22844,N_21212,N_21671);
xor U22845 (N_22845,N_21057,N_21040);
or U22846 (N_22846,N_20883,N_20449);
and U22847 (N_22847,N_21429,N_21777);
or U22848 (N_22848,N_21747,N_21706);
xnor U22849 (N_22849,N_20582,N_20741);
or U22850 (N_22850,N_21804,N_21483);
nor U22851 (N_22851,N_21676,N_20988);
nor U22852 (N_22852,N_20425,N_20253);
nand U22853 (N_22853,N_20354,N_20313);
nand U22854 (N_22854,N_20713,N_21138);
xnor U22855 (N_22855,N_21336,N_20726);
and U22856 (N_22856,N_21989,N_21906);
and U22857 (N_22857,N_21101,N_21639);
and U22858 (N_22858,N_21287,N_20143);
nor U22859 (N_22859,N_20948,N_20850);
xor U22860 (N_22860,N_20170,N_20772);
or U22861 (N_22861,N_21949,N_21240);
or U22862 (N_22862,N_20020,N_20567);
xor U22863 (N_22863,N_21133,N_20643);
nor U22864 (N_22864,N_21245,N_21087);
or U22865 (N_22865,N_20326,N_21862);
xnor U22866 (N_22866,N_20842,N_20492);
and U22867 (N_22867,N_21686,N_20485);
nand U22868 (N_22868,N_21247,N_21775);
nand U22869 (N_22869,N_20162,N_21301);
xnor U22870 (N_22870,N_21310,N_20448);
and U22871 (N_22871,N_21655,N_21015);
xor U22872 (N_22872,N_21403,N_20743);
xnor U22873 (N_22873,N_21474,N_20090);
xor U22874 (N_22874,N_21487,N_21479);
nor U22875 (N_22875,N_21324,N_20149);
or U22876 (N_22876,N_20205,N_20101);
xor U22877 (N_22877,N_20198,N_20457);
and U22878 (N_22878,N_20224,N_21828);
xnor U22879 (N_22879,N_20370,N_21099);
nor U22880 (N_22880,N_21018,N_20407);
nor U22881 (N_22881,N_20164,N_21703);
nor U22882 (N_22882,N_21179,N_20344);
nor U22883 (N_22883,N_20998,N_20142);
nor U22884 (N_22884,N_21343,N_20903);
nor U22885 (N_22885,N_20471,N_21994);
xnor U22886 (N_22886,N_21421,N_20626);
nor U22887 (N_22887,N_20870,N_21719);
and U22888 (N_22888,N_20381,N_21227);
xnor U22889 (N_22889,N_20667,N_21369);
and U22890 (N_22890,N_20490,N_20193);
nor U22891 (N_22891,N_20296,N_21004);
or U22892 (N_22892,N_21214,N_20464);
or U22893 (N_22893,N_21168,N_21852);
and U22894 (N_22894,N_20555,N_21527);
nor U22895 (N_22895,N_20958,N_20872);
or U22896 (N_22896,N_21537,N_21239);
or U22897 (N_22897,N_21784,N_21445);
xnor U22898 (N_22898,N_21126,N_21666);
and U22899 (N_22899,N_21136,N_21611);
xnor U22900 (N_22900,N_21293,N_21886);
and U22901 (N_22901,N_20829,N_21588);
nand U22902 (N_22902,N_20649,N_20640);
nand U22903 (N_22903,N_20102,N_21789);
and U22904 (N_22904,N_21939,N_21257);
nand U22905 (N_22905,N_21426,N_21394);
nor U22906 (N_22906,N_20818,N_21412);
and U22907 (N_22907,N_20290,N_20314);
xor U22908 (N_22908,N_20091,N_21430);
nand U22909 (N_22909,N_20651,N_21410);
and U22910 (N_22910,N_21731,N_21576);
and U22911 (N_22911,N_20500,N_20997);
xnor U22912 (N_22912,N_21769,N_21904);
xnor U22913 (N_22913,N_21242,N_21744);
or U22914 (N_22914,N_20559,N_21782);
nor U22915 (N_22915,N_20255,N_20519);
nor U22916 (N_22916,N_21556,N_21750);
and U22917 (N_22917,N_20946,N_21806);
and U22918 (N_22918,N_20215,N_21954);
nor U22919 (N_22919,N_20980,N_21294);
or U22920 (N_22920,N_21317,N_21390);
xnor U22921 (N_22921,N_20172,N_21089);
or U22922 (N_22922,N_21384,N_20786);
nor U22923 (N_22923,N_20821,N_21173);
and U22924 (N_22924,N_21520,N_21908);
and U22925 (N_22925,N_20237,N_21808);
or U22926 (N_22926,N_21465,N_20402);
or U22927 (N_22927,N_21818,N_21618);
xnor U22928 (N_22928,N_20865,N_21541);
nand U22929 (N_22929,N_21897,N_21794);
and U22930 (N_22930,N_20952,N_20620);
or U22931 (N_22931,N_21506,N_20306);
xor U22932 (N_22932,N_20942,N_20338);
nor U22933 (N_22933,N_20638,N_21825);
and U22934 (N_22934,N_20264,N_21323);
xor U22935 (N_22935,N_21194,N_20097);
nor U22936 (N_22936,N_21127,N_21614);
and U22937 (N_22937,N_21220,N_20807);
nor U22938 (N_22938,N_21008,N_20073);
or U22939 (N_22939,N_21768,N_20756);
xnor U22940 (N_22940,N_21348,N_21640);
nor U22941 (N_22941,N_20259,N_21599);
xor U22942 (N_22942,N_20920,N_20697);
nor U22943 (N_22943,N_21502,N_20064);
and U22944 (N_22944,N_20712,N_20717);
xor U22945 (N_22945,N_20808,N_20315);
nand U22946 (N_22946,N_20307,N_20229);
nand U22947 (N_22947,N_21221,N_21668);
nor U22948 (N_22948,N_20410,N_20523);
nand U22949 (N_22949,N_21511,N_21277);
nand U22950 (N_22950,N_20144,N_20841);
xor U22951 (N_22951,N_20227,N_20965);
nand U22952 (N_22952,N_21365,N_20616);
nand U22953 (N_22953,N_21892,N_20055);
and U22954 (N_22954,N_21847,N_20961);
xor U22955 (N_22955,N_20615,N_21842);
nor U22956 (N_22956,N_21233,N_20516);
nor U22957 (N_22957,N_20126,N_20539);
or U22958 (N_22958,N_21006,N_21797);
and U22959 (N_22959,N_20460,N_20445);
nor U22960 (N_22960,N_21230,N_21289);
nor U22961 (N_22961,N_21356,N_20399);
and U22962 (N_22962,N_20822,N_20453);
xor U22963 (N_22963,N_21124,N_20773);
or U22964 (N_22964,N_21922,N_20685);
or U22965 (N_22965,N_20746,N_20749);
nor U22966 (N_22966,N_20141,N_20873);
nor U22967 (N_22967,N_21975,N_21152);
nand U22968 (N_22968,N_20137,N_21699);
xor U22969 (N_22969,N_21486,N_20780);
xnor U22970 (N_22970,N_21433,N_21200);
xnor U22971 (N_22971,N_20327,N_20605);
nand U22972 (N_22972,N_21450,N_20479);
and U22973 (N_22973,N_20666,N_20204);
nor U22974 (N_22974,N_20562,N_21726);
or U22975 (N_22975,N_20352,N_20223);
or U22976 (N_22976,N_20700,N_21051);
and U22977 (N_22977,N_21241,N_20171);
xor U22978 (N_22978,N_21308,N_21342);
nor U22979 (N_22979,N_21696,N_21201);
and U22980 (N_22980,N_21783,N_21771);
and U22981 (N_22981,N_20392,N_21019);
nor U22982 (N_22982,N_20365,N_21665);
or U22983 (N_22983,N_21104,N_21279);
or U22984 (N_22984,N_21080,N_20194);
and U22985 (N_22985,N_21822,N_20033);
nor U22986 (N_22986,N_20660,N_20705);
xnor U22987 (N_22987,N_21714,N_20759);
nor U22988 (N_22988,N_21190,N_21883);
or U22989 (N_22989,N_20334,N_21268);
nor U22990 (N_22990,N_20316,N_20439);
xnor U22991 (N_22991,N_21081,N_21193);
nand U22992 (N_22992,N_20530,N_20111);
or U22993 (N_22993,N_20675,N_21603);
nor U22994 (N_22994,N_20919,N_21953);
xnor U22995 (N_22995,N_21615,N_20926);
xnor U22996 (N_22996,N_21262,N_20463);
nor U22997 (N_22997,N_20106,N_21876);
or U22998 (N_22998,N_21785,N_20008);
xnor U22999 (N_22999,N_20981,N_21095);
and U23000 (N_23000,N_20444,N_21818);
and U23001 (N_23001,N_21139,N_21083);
nor U23002 (N_23002,N_21299,N_20526);
xor U23003 (N_23003,N_20304,N_21388);
or U23004 (N_23004,N_21180,N_20373);
or U23005 (N_23005,N_21135,N_21266);
xnor U23006 (N_23006,N_20192,N_20571);
nor U23007 (N_23007,N_21228,N_20940);
and U23008 (N_23008,N_21590,N_21230);
xor U23009 (N_23009,N_20464,N_21900);
xor U23010 (N_23010,N_21152,N_20976);
and U23011 (N_23011,N_20952,N_20035);
or U23012 (N_23012,N_20818,N_21004);
and U23013 (N_23013,N_20556,N_21700);
xnor U23014 (N_23014,N_20968,N_21130);
nand U23015 (N_23015,N_21765,N_20065);
and U23016 (N_23016,N_21681,N_20768);
nand U23017 (N_23017,N_21571,N_20408);
or U23018 (N_23018,N_20819,N_21517);
nor U23019 (N_23019,N_21548,N_21994);
xnor U23020 (N_23020,N_20539,N_21388);
or U23021 (N_23021,N_20959,N_20055);
or U23022 (N_23022,N_21469,N_20283);
nor U23023 (N_23023,N_20902,N_20141);
xnor U23024 (N_23024,N_21665,N_20253);
nor U23025 (N_23025,N_20507,N_21175);
or U23026 (N_23026,N_20158,N_20823);
nor U23027 (N_23027,N_20647,N_21170);
nand U23028 (N_23028,N_21819,N_20848);
xnor U23029 (N_23029,N_20653,N_21905);
or U23030 (N_23030,N_21070,N_21177);
nor U23031 (N_23031,N_21519,N_20842);
and U23032 (N_23032,N_21398,N_20226);
xnor U23033 (N_23033,N_21410,N_20768);
nand U23034 (N_23034,N_21154,N_21459);
or U23035 (N_23035,N_20923,N_20577);
and U23036 (N_23036,N_21181,N_20867);
or U23037 (N_23037,N_20368,N_21870);
or U23038 (N_23038,N_20490,N_21261);
nand U23039 (N_23039,N_21554,N_20010);
xnor U23040 (N_23040,N_20213,N_21643);
and U23041 (N_23041,N_20564,N_20042);
nand U23042 (N_23042,N_21934,N_20288);
nor U23043 (N_23043,N_20496,N_20862);
nand U23044 (N_23044,N_21497,N_20551);
and U23045 (N_23045,N_21274,N_21490);
nand U23046 (N_23046,N_21206,N_20804);
xor U23047 (N_23047,N_21373,N_20223);
and U23048 (N_23048,N_20524,N_20428);
nand U23049 (N_23049,N_20308,N_21246);
and U23050 (N_23050,N_21533,N_21750);
or U23051 (N_23051,N_20745,N_20486);
or U23052 (N_23052,N_21472,N_20649);
and U23053 (N_23053,N_20647,N_21957);
xnor U23054 (N_23054,N_20826,N_21874);
nor U23055 (N_23055,N_21349,N_21528);
nor U23056 (N_23056,N_20005,N_21955);
and U23057 (N_23057,N_20632,N_21581);
nand U23058 (N_23058,N_21151,N_20149);
and U23059 (N_23059,N_21181,N_21272);
nor U23060 (N_23060,N_20219,N_20216);
and U23061 (N_23061,N_20017,N_21231);
nand U23062 (N_23062,N_20551,N_21157);
xnor U23063 (N_23063,N_21383,N_20565);
nor U23064 (N_23064,N_21800,N_21555);
nor U23065 (N_23065,N_20488,N_20574);
and U23066 (N_23066,N_20703,N_20277);
nand U23067 (N_23067,N_21133,N_20360);
nand U23068 (N_23068,N_20408,N_20097);
nand U23069 (N_23069,N_21853,N_21457);
nor U23070 (N_23070,N_20812,N_21564);
xnor U23071 (N_23071,N_20659,N_20975);
nand U23072 (N_23072,N_20461,N_21204);
or U23073 (N_23073,N_21927,N_20934);
nand U23074 (N_23074,N_21135,N_21593);
or U23075 (N_23075,N_20966,N_20620);
nand U23076 (N_23076,N_21253,N_20189);
nand U23077 (N_23077,N_20802,N_20196);
nand U23078 (N_23078,N_21671,N_21757);
or U23079 (N_23079,N_20637,N_21252);
nor U23080 (N_23080,N_20504,N_21437);
nor U23081 (N_23081,N_21679,N_20958);
nand U23082 (N_23082,N_21140,N_21986);
or U23083 (N_23083,N_20294,N_20264);
and U23084 (N_23084,N_20845,N_20513);
and U23085 (N_23085,N_20045,N_20410);
or U23086 (N_23086,N_21677,N_20761);
or U23087 (N_23087,N_21338,N_20504);
nor U23088 (N_23088,N_20709,N_20635);
or U23089 (N_23089,N_21530,N_20149);
xnor U23090 (N_23090,N_20723,N_20470);
xor U23091 (N_23091,N_21199,N_21460);
and U23092 (N_23092,N_20508,N_21526);
and U23093 (N_23093,N_20120,N_20166);
xor U23094 (N_23094,N_21235,N_20680);
xor U23095 (N_23095,N_21307,N_20901);
and U23096 (N_23096,N_20621,N_20452);
and U23097 (N_23097,N_21859,N_21239);
or U23098 (N_23098,N_20204,N_20109);
and U23099 (N_23099,N_21098,N_21836);
xnor U23100 (N_23100,N_20318,N_20809);
and U23101 (N_23101,N_20918,N_20103);
nor U23102 (N_23102,N_20556,N_20613);
or U23103 (N_23103,N_21875,N_21624);
or U23104 (N_23104,N_21012,N_21596);
xor U23105 (N_23105,N_20363,N_20940);
xor U23106 (N_23106,N_21919,N_20800);
xor U23107 (N_23107,N_21322,N_20412);
and U23108 (N_23108,N_21106,N_20615);
or U23109 (N_23109,N_20411,N_21072);
and U23110 (N_23110,N_20972,N_20789);
nor U23111 (N_23111,N_20577,N_20419);
or U23112 (N_23112,N_20617,N_21329);
or U23113 (N_23113,N_20759,N_21776);
nand U23114 (N_23114,N_20746,N_21952);
or U23115 (N_23115,N_20007,N_20945);
or U23116 (N_23116,N_21447,N_21997);
nor U23117 (N_23117,N_20781,N_21954);
and U23118 (N_23118,N_20441,N_21831);
nand U23119 (N_23119,N_21867,N_21427);
xor U23120 (N_23120,N_21210,N_20840);
xor U23121 (N_23121,N_20861,N_20192);
xnor U23122 (N_23122,N_21409,N_21486);
xor U23123 (N_23123,N_21613,N_20614);
and U23124 (N_23124,N_20315,N_20652);
nor U23125 (N_23125,N_21902,N_21189);
and U23126 (N_23126,N_20679,N_21668);
nand U23127 (N_23127,N_21006,N_21874);
nand U23128 (N_23128,N_21243,N_21961);
nand U23129 (N_23129,N_20767,N_21695);
or U23130 (N_23130,N_21505,N_20078);
xor U23131 (N_23131,N_21914,N_21209);
xor U23132 (N_23132,N_20108,N_21594);
or U23133 (N_23133,N_21969,N_21757);
or U23134 (N_23134,N_20072,N_20177);
or U23135 (N_23135,N_20348,N_21691);
and U23136 (N_23136,N_20533,N_20457);
nand U23137 (N_23137,N_21078,N_20422);
nand U23138 (N_23138,N_21868,N_21384);
xor U23139 (N_23139,N_20354,N_21839);
nor U23140 (N_23140,N_20156,N_20213);
or U23141 (N_23141,N_21452,N_21111);
or U23142 (N_23142,N_21274,N_21046);
nand U23143 (N_23143,N_20394,N_20014);
and U23144 (N_23144,N_20739,N_20625);
and U23145 (N_23145,N_20253,N_20777);
xnor U23146 (N_23146,N_20715,N_21745);
and U23147 (N_23147,N_21061,N_20767);
and U23148 (N_23148,N_21851,N_20603);
and U23149 (N_23149,N_21635,N_21020);
or U23150 (N_23150,N_21727,N_21801);
and U23151 (N_23151,N_21431,N_21389);
and U23152 (N_23152,N_20101,N_21087);
xor U23153 (N_23153,N_21093,N_20877);
and U23154 (N_23154,N_21707,N_20417);
or U23155 (N_23155,N_21212,N_21907);
or U23156 (N_23156,N_21317,N_21607);
xor U23157 (N_23157,N_21861,N_21589);
or U23158 (N_23158,N_21216,N_20931);
or U23159 (N_23159,N_20450,N_21016);
and U23160 (N_23160,N_21078,N_20387);
or U23161 (N_23161,N_20564,N_21906);
and U23162 (N_23162,N_21970,N_20868);
nand U23163 (N_23163,N_21615,N_21217);
or U23164 (N_23164,N_20084,N_20666);
or U23165 (N_23165,N_20024,N_20054);
and U23166 (N_23166,N_20844,N_21227);
nor U23167 (N_23167,N_20699,N_20051);
nor U23168 (N_23168,N_20032,N_21509);
and U23169 (N_23169,N_20149,N_20653);
or U23170 (N_23170,N_20521,N_21800);
nand U23171 (N_23171,N_20959,N_20787);
or U23172 (N_23172,N_20655,N_21010);
and U23173 (N_23173,N_21112,N_20883);
nor U23174 (N_23174,N_21943,N_21064);
nor U23175 (N_23175,N_21194,N_20052);
nand U23176 (N_23176,N_20344,N_21160);
nand U23177 (N_23177,N_21153,N_21233);
nor U23178 (N_23178,N_20928,N_20080);
nor U23179 (N_23179,N_21193,N_20665);
xnor U23180 (N_23180,N_21241,N_21577);
and U23181 (N_23181,N_21711,N_21199);
nand U23182 (N_23182,N_20108,N_20826);
or U23183 (N_23183,N_20165,N_20881);
and U23184 (N_23184,N_20544,N_21596);
xnor U23185 (N_23185,N_21806,N_20930);
or U23186 (N_23186,N_20107,N_20052);
or U23187 (N_23187,N_20876,N_20273);
and U23188 (N_23188,N_21234,N_21181);
nor U23189 (N_23189,N_20307,N_21408);
nand U23190 (N_23190,N_21640,N_20246);
or U23191 (N_23191,N_21756,N_20978);
nand U23192 (N_23192,N_20310,N_20750);
nor U23193 (N_23193,N_20056,N_21838);
and U23194 (N_23194,N_21357,N_20832);
xnor U23195 (N_23195,N_20875,N_20175);
or U23196 (N_23196,N_20030,N_21316);
nor U23197 (N_23197,N_21216,N_21463);
and U23198 (N_23198,N_20296,N_20181);
or U23199 (N_23199,N_20665,N_20151);
nand U23200 (N_23200,N_20843,N_20923);
nand U23201 (N_23201,N_21405,N_21820);
or U23202 (N_23202,N_21079,N_20497);
nand U23203 (N_23203,N_21961,N_21975);
nor U23204 (N_23204,N_21779,N_20602);
nor U23205 (N_23205,N_21372,N_20405);
xnor U23206 (N_23206,N_21533,N_20667);
nor U23207 (N_23207,N_21868,N_20911);
xnor U23208 (N_23208,N_20995,N_21477);
or U23209 (N_23209,N_21722,N_20673);
xor U23210 (N_23210,N_21053,N_21020);
nand U23211 (N_23211,N_20092,N_21013);
and U23212 (N_23212,N_21369,N_20378);
xnor U23213 (N_23213,N_21638,N_20550);
xor U23214 (N_23214,N_21421,N_21048);
nor U23215 (N_23215,N_21062,N_20332);
xnor U23216 (N_23216,N_21871,N_21722);
and U23217 (N_23217,N_21460,N_20968);
nand U23218 (N_23218,N_20561,N_21159);
or U23219 (N_23219,N_21595,N_21713);
and U23220 (N_23220,N_21226,N_20953);
or U23221 (N_23221,N_20161,N_21107);
nor U23222 (N_23222,N_21083,N_20583);
xnor U23223 (N_23223,N_21246,N_20095);
xnor U23224 (N_23224,N_21673,N_20280);
nor U23225 (N_23225,N_20619,N_20268);
xor U23226 (N_23226,N_20170,N_20516);
or U23227 (N_23227,N_20511,N_20068);
xnor U23228 (N_23228,N_20082,N_20116);
or U23229 (N_23229,N_21780,N_21946);
and U23230 (N_23230,N_20399,N_21659);
xnor U23231 (N_23231,N_20269,N_21231);
xnor U23232 (N_23232,N_20377,N_20553);
nor U23233 (N_23233,N_20674,N_20865);
xor U23234 (N_23234,N_21144,N_20424);
nand U23235 (N_23235,N_20701,N_20135);
nor U23236 (N_23236,N_21933,N_21320);
nand U23237 (N_23237,N_20739,N_21364);
or U23238 (N_23238,N_21497,N_21616);
or U23239 (N_23239,N_20930,N_20399);
xor U23240 (N_23240,N_21133,N_21063);
nor U23241 (N_23241,N_20450,N_20457);
xor U23242 (N_23242,N_21404,N_20025);
or U23243 (N_23243,N_20988,N_20081);
or U23244 (N_23244,N_20571,N_21485);
nor U23245 (N_23245,N_21739,N_20026);
or U23246 (N_23246,N_20297,N_20007);
xor U23247 (N_23247,N_21545,N_21503);
or U23248 (N_23248,N_20627,N_21804);
nand U23249 (N_23249,N_20622,N_20705);
and U23250 (N_23250,N_21272,N_21961);
or U23251 (N_23251,N_20736,N_20621);
nor U23252 (N_23252,N_20164,N_21885);
nand U23253 (N_23253,N_21391,N_21144);
and U23254 (N_23254,N_21271,N_21141);
and U23255 (N_23255,N_20205,N_20068);
nand U23256 (N_23256,N_21940,N_20334);
and U23257 (N_23257,N_21201,N_20026);
nand U23258 (N_23258,N_21176,N_20351);
nor U23259 (N_23259,N_20566,N_20879);
or U23260 (N_23260,N_20453,N_21079);
xor U23261 (N_23261,N_21939,N_20293);
and U23262 (N_23262,N_21590,N_21066);
nor U23263 (N_23263,N_20482,N_20475);
and U23264 (N_23264,N_21209,N_21799);
xor U23265 (N_23265,N_21308,N_20044);
or U23266 (N_23266,N_20343,N_21572);
or U23267 (N_23267,N_21009,N_20712);
or U23268 (N_23268,N_20587,N_21883);
xnor U23269 (N_23269,N_21759,N_21646);
nor U23270 (N_23270,N_20258,N_21305);
nor U23271 (N_23271,N_20580,N_21975);
nor U23272 (N_23272,N_21692,N_20316);
and U23273 (N_23273,N_21052,N_20252);
nand U23274 (N_23274,N_21986,N_21908);
nor U23275 (N_23275,N_21036,N_20927);
nand U23276 (N_23276,N_20228,N_21306);
nand U23277 (N_23277,N_20445,N_21096);
nand U23278 (N_23278,N_20580,N_20081);
and U23279 (N_23279,N_21971,N_20098);
xor U23280 (N_23280,N_20752,N_20048);
and U23281 (N_23281,N_20146,N_21109);
nand U23282 (N_23282,N_20785,N_21632);
nand U23283 (N_23283,N_21789,N_21986);
xnor U23284 (N_23284,N_20665,N_20278);
xnor U23285 (N_23285,N_20956,N_21256);
nand U23286 (N_23286,N_20364,N_20607);
and U23287 (N_23287,N_21631,N_21296);
xor U23288 (N_23288,N_21241,N_21380);
or U23289 (N_23289,N_21456,N_21467);
or U23290 (N_23290,N_20560,N_20302);
xor U23291 (N_23291,N_20183,N_20439);
and U23292 (N_23292,N_21779,N_20834);
nor U23293 (N_23293,N_20551,N_20993);
nor U23294 (N_23294,N_20105,N_21702);
or U23295 (N_23295,N_20533,N_20681);
and U23296 (N_23296,N_21156,N_21984);
nand U23297 (N_23297,N_20566,N_20590);
nand U23298 (N_23298,N_20623,N_21038);
xnor U23299 (N_23299,N_21657,N_21091);
and U23300 (N_23300,N_20951,N_21689);
and U23301 (N_23301,N_20247,N_20790);
nand U23302 (N_23302,N_20031,N_20332);
xor U23303 (N_23303,N_21835,N_21967);
or U23304 (N_23304,N_21051,N_21407);
or U23305 (N_23305,N_21395,N_20903);
xor U23306 (N_23306,N_21143,N_21064);
and U23307 (N_23307,N_21857,N_21649);
and U23308 (N_23308,N_21929,N_21508);
and U23309 (N_23309,N_21292,N_21792);
nand U23310 (N_23310,N_20150,N_20631);
or U23311 (N_23311,N_21873,N_20262);
xnor U23312 (N_23312,N_20160,N_20373);
nor U23313 (N_23313,N_21941,N_20265);
and U23314 (N_23314,N_21449,N_21650);
nand U23315 (N_23315,N_20767,N_21025);
or U23316 (N_23316,N_20200,N_21930);
and U23317 (N_23317,N_21007,N_20855);
xor U23318 (N_23318,N_20520,N_21976);
xor U23319 (N_23319,N_21254,N_20824);
nor U23320 (N_23320,N_20373,N_20593);
and U23321 (N_23321,N_21737,N_21988);
and U23322 (N_23322,N_20422,N_21024);
nand U23323 (N_23323,N_21569,N_20467);
xnor U23324 (N_23324,N_20726,N_20223);
xnor U23325 (N_23325,N_21582,N_20359);
xor U23326 (N_23326,N_21688,N_21112);
xor U23327 (N_23327,N_21137,N_21673);
and U23328 (N_23328,N_21782,N_21619);
or U23329 (N_23329,N_20103,N_20826);
and U23330 (N_23330,N_21064,N_20089);
or U23331 (N_23331,N_21747,N_20150);
nand U23332 (N_23332,N_20551,N_21015);
nor U23333 (N_23333,N_21581,N_21268);
and U23334 (N_23334,N_21359,N_20607);
nor U23335 (N_23335,N_21973,N_20662);
nor U23336 (N_23336,N_20422,N_21218);
nand U23337 (N_23337,N_20210,N_21944);
xor U23338 (N_23338,N_20716,N_20407);
and U23339 (N_23339,N_20232,N_21964);
nand U23340 (N_23340,N_20878,N_21483);
nand U23341 (N_23341,N_20910,N_21920);
nand U23342 (N_23342,N_20721,N_21141);
or U23343 (N_23343,N_21475,N_21664);
or U23344 (N_23344,N_21935,N_20518);
xnor U23345 (N_23345,N_21472,N_20004);
and U23346 (N_23346,N_21689,N_20236);
or U23347 (N_23347,N_21139,N_21771);
or U23348 (N_23348,N_20267,N_21756);
nand U23349 (N_23349,N_20833,N_21071);
nand U23350 (N_23350,N_21238,N_20903);
xnor U23351 (N_23351,N_20951,N_21836);
nor U23352 (N_23352,N_21426,N_20105);
xor U23353 (N_23353,N_20892,N_21691);
nand U23354 (N_23354,N_20576,N_21303);
xor U23355 (N_23355,N_20512,N_21834);
xor U23356 (N_23356,N_20550,N_20053);
nand U23357 (N_23357,N_20331,N_20059);
xnor U23358 (N_23358,N_20004,N_20106);
and U23359 (N_23359,N_20604,N_21398);
xor U23360 (N_23360,N_20017,N_20167);
nand U23361 (N_23361,N_21117,N_20986);
or U23362 (N_23362,N_20294,N_20578);
or U23363 (N_23363,N_20504,N_20158);
or U23364 (N_23364,N_20727,N_20138);
and U23365 (N_23365,N_21079,N_21986);
xor U23366 (N_23366,N_20374,N_20306);
and U23367 (N_23367,N_20088,N_20876);
or U23368 (N_23368,N_20227,N_21666);
and U23369 (N_23369,N_21442,N_20257);
nand U23370 (N_23370,N_20471,N_21301);
nor U23371 (N_23371,N_21448,N_20590);
nor U23372 (N_23372,N_21514,N_21969);
xnor U23373 (N_23373,N_20451,N_21516);
or U23374 (N_23374,N_21287,N_20567);
nand U23375 (N_23375,N_21180,N_21480);
xor U23376 (N_23376,N_21698,N_20549);
nor U23377 (N_23377,N_20479,N_20078);
xor U23378 (N_23378,N_21816,N_20248);
and U23379 (N_23379,N_21482,N_20435);
xor U23380 (N_23380,N_20878,N_21077);
nor U23381 (N_23381,N_20771,N_20172);
and U23382 (N_23382,N_21920,N_21443);
and U23383 (N_23383,N_20700,N_20822);
nor U23384 (N_23384,N_21705,N_20269);
xor U23385 (N_23385,N_20251,N_20129);
nor U23386 (N_23386,N_21166,N_21249);
nor U23387 (N_23387,N_20132,N_21155);
nand U23388 (N_23388,N_21949,N_20840);
and U23389 (N_23389,N_20577,N_21826);
nor U23390 (N_23390,N_20086,N_21119);
nor U23391 (N_23391,N_21030,N_20794);
xor U23392 (N_23392,N_21071,N_20367);
nand U23393 (N_23393,N_21535,N_20800);
xnor U23394 (N_23394,N_21379,N_20801);
xor U23395 (N_23395,N_20321,N_20156);
nor U23396 (N_23396,N_20658,N_20488);
nor U23397 (N_23397,N_21479,N_21209);
xor U23398 (N_23398,N_21417,N_21702);
and U23399 (N_23399,N_20706,N_21348);
nand U23400 (N_23400,N_20048,N_20795);
xnor U23401 (N_23401,N_21088,N_20480);
nor U23402 (N_23402,N_20764,N_21358);
xor U23403 (N_23403,N_20150,N_20680);
and U23404 (N_23404,N_21382,N_21093);
nor U23405 (N_23405,N_21141,N_20300);
and U23406 (N_23406,N_20508,N_21827);
nand U23407 (N_23407,N_21607,N_21285);
nand U23408 (N_23408,N_20166,N_21358);
and U23409 (N_23409,N_20160,N_21081);
or U23410 (N_23410,N_20278,N_21971);
or U23411 (N_23411,N_20102,N_20931);
nor U23412 (N_23412,N_20966,N_21947);
or U23413 (N_23413,N_21728,N_20192);
nor U23414 (N_23414,N_21390,N_21845);
xnor U23415 (N_23415,N_21790,N_20098);
or U23416 (N_23416,N_21925,N_20184);
or U23417 (N_23417,N_20728,N_20118);
xor U23418 (N_23418,N_20858,N_21911);
or U23419 (N_23419,N_21754,N_20149);
or U23420 (N_23420,N_20240,N_20909);
nor U23421 (N_23421,N_20193,N_21053);
nor U23422 (N_23422,N_21144,N_21717);
xnor U23423 (N_23423,N_21319,N_21251);
xor U23424 (N_23424,N_21016,N_21340);
and U23425 (N_23425,N_21722,N_20981);
nand U23426 (N_23426,N_21665,N_20039);
nor U23427 (N_23427,N_20936,N_21411);
nand U23428 (N_23428,N_21625,N_20350);
nand U23429 (N_23429,N_21452,N_21355);
and U23430 (N_23430,N_21841,N_20714);
or U23431 (N_23431,N_21117,N_21631);
xor U23432 (N_23432,N_20215,N_20035);
and U23433 (N_23433,N_21371,N_20116);
and U23434 (N_23434,N_20881,N_20164);
or U23435 (N_23435,N_20644,N_20307);
nor U23436 (N_23436,N_21213,N_20171);
nand U23437 (N_23437,N_20442,N_21626);
and U23438 (N_23438,N_20399,N_20188);
or U23439 (N_23439,N_20807,N_20529);
nand U23440 (N_23440,N_20499,N_21796);
xnor U23441 (N_23441,N_20063,N_20278);
and U23442 (N_23442,N_21330,N_21412);
and U23443 (N_23443,N_20737,N_21800);
nand U23444 (N_23444,N_21539,N_20457);
nand U23445 (N_23445,N_20415,N_20059);
nor U23446 (N_23446,N_20250,N_21055);
xnor U23447 (N_23447,N_20977,N_20476);
xnor U23448 (N_23448,N_20744,N_20537);
and U23449 (N_23449,N_21903,N_20260);
xor U23450 (N_23450,N_20249,N_21041);
and U23451 (N_23451,N_20884,N_20575);
xnor U23452 (N_23452,N_20870,N_21441);
xnor U23453 (N_23453,N_21048,N_20012);
or U23454 (N_23454,N_20020,N_21508);
or U23455 (N_23455,N_20258,N_21762);
xor U23456 (N_23456,N_20190,N_21596);
and U23457 (N_23457,N_20444,N_21380);
nand U23458 (N_23458,N_21647,N_20536);
or U23459 (N_23459,N_20640,N_21544);
xor U23460 (N_23460,N_20213,N_21797);
nor U23461 (N_23461,N_20899,N_21149);
or U23462 (N_23462,N_21811,N_20797);
nor U23463 (N_23463,N_20373,N_21118);
nor U23464 (N_23464,N_20204,N_20927);
nand U23465 (N_23465,N_20150,N_20051);
nand U23466 (N_23466,N_21935,N_20924);
nand U23467 (N_23467,N_21311,N_21871);
and U23468 (N_23468,N_21192,N_20037);
xnor U23469 (N_23469,N_21619,N_20649);
nor U23470 (N_23470,N_20285,N_21366);
xor U23471 (N_23471,N_21350,N_21039);
nor U23472 (N_23472,N_21420,N_20124);
xor U23473 (N_23473,N_21423,N_20460);
nor U23474 (N_23474,N_20648,N_21182);
xor U23475 (N_23475,N_20915,N_21394);
xnor U23476 (N_23476,N_20754,N_20719);
nand U23477 (N_23477,N_21081,N_21195);
or U23478 (N_23478,N_21592,N_20748);
xnor U23479 (N_23479,N_21483,N_20957);
and U23480 (N_23480,N_20769,N_21795);
or U23481 (N_23481,N_20422,N_21947);
or U23482 (N_23482,N_20335,N_20705);
nor U23483 (N_23483,N_20778,N_21523);
xor U23484 (N_23484,N_20136,N_21595);
nor U23485 (N_23485,N_20215,N_21617);
and U23486 (N_23486,N_21401,N_20958);
and U23487 (N_23487,N_21911,N_20985);
nor U23488 (N_23488,N_20362,N_20131);
nor U23489 (N_23489,N_21971,N_20908);
xor U23490 (N_23490,N_20577,N_20744);
xnor U23491 (N_23491,N_21237,N_21618);
and U23492 (N_23492,N_21399,N_21470);
nor U23493 (N_23493,N_21508,N_20900);
or U23494 (N_23494,N_20149,N_21654);
or U23495 (N_23495,N_20277,N_21511);
and U23496 (N_23496,N_20065,N_20175);
xor U23497 (N_23497,N_20655,N_21935);
nand U23498 (N_23498,N_21226,N_20708);
nor U23499 (N_23499,N_20735,N_20953);
and U23500 (N_23500,N_21245,N_20034);
xnor U23501 (N_23501,N_21470,N_20278);
nor U23502 (N_23502,N_21886,N_20767);
xnor U23503 (N_23503,N_21994,N_20407);
or U23504 (N_23504,N_20238,N_21179);
xnor U23505 (N_23505,N_21008,N_21313);
nand U23506 (N_23506,N_20952,N_21085);
nand U23507 (N_23507,N_20043,N_20147);
xor U23508 (N_23508,N_20211,N_20609);
and U23509 (N_23509,N_21395,N_20720);
xor U23510 (N_23510,N_20665,N_20171);
nor U23511 (N_23511,N_21180,N_21593);
nand U23512 (N_23512,N_20466,N_20707);
and U23513 (N_23513,N_20775,N_20804);
and U23514 (N_23514,N_21772,N_21913);
nor U23515 (N_23515,N_20164,N_20321);
and U23516 (N_23516,N_21257,N_21960);
nand U23517 (N_23517,N_21019,N_21074);
nand U23518 (N_23518,N_21356,N_21705);
and U23519 (N_23519,N_20490,N_21281);
nand U23520 (N_23520,N_21319,N_20359);
xnor U23521 (N_23521,N_21337,N_21950);
nor U23522 (N_23522,N_20247,N_20464);
or U23523 (N_23523,N_20223,N_20146);
and U23524 (N_23524,N_21666,N_21438);
and U23525 (N_23525,N_20503,N_20750);
or U23526 (N_23526,N_20338,N_20855);
or U23527 (N_23527,N_21371,N_21851);
nand U23528 (N_23528,N_20835,N_20088);
nor U23529 (N_23529,N_20224,N_21992);
nand U23530 (N_23530,N_21458,N_21152);
nand U23531 (N_23531,N_20463,N_21052);
or U23532 (N_23532,N_21898,N_21719);
nand U23533 (N_23533,N_20068,N_20679);
and U23534 (N_23534,N_21528,N_20796);
nor U23535 (N_23535,N_20646,N_20355);
nand U23536 (N_23536,N_21025,N_21551);
or U23537 (N_23537,N_21854,N_20150);
and U23538 (N_23538,N_20879,N_21457);
nand U23539 (N_23539,N_20668,N_21750);
and U23540 (N_23540,N_20649,N_20624);
nor U23541 (N_23541,N_21553,N_20261);
and U23542 (N_23542,N_21421,N_21986);
or U23543 (N_23543,N_20324,N_20568);
nand U23544 (N_23544,N_20055,N_20358);
or U23545 (N_23545,N_21825,N_20792);
and U23546 (N_23546,N_21756,N_20100);
and U23547 (N_23547,N_21149,N_20487);
or U23548 (N_23548,N_20101,N_21480);
nand U23549 (N_23549,N_21526,N_21353);
nor U23550 (N_23550,N_20985,N_20010);
xnor U23551 (N_23551,N_20096,N_21342);
xor U23552 (N_23552,N_20221,N_21128);
or U23553 (N_23553,N_21248,N_21497);
and U23554 (N_23554,N_21143,N_21532);
nand U23555 (N_23555,N_21683,N_20513);
and U23556 (N_23556,N_20211,N_20500);
nand U23557 (N_23557,N_20794,N_20843);
and U23558 (N_23558,N_21020,N_21750);
xnor U23559 (N_23559,N_20642,N_20987);
nor U23560 (N_23560,N_20317,N_20586);
xnor U23561 (N_23561,N_20479,N_21260);
xnor U23562 (N_23562,N_21816,N_20244);
nand U23563 (N_23563,N_20049,N_20821);
nand U23564 (N_23564,N_21847,N_21815);
nor U23565 (N_23565,N_21379,N_21622);
and U23566 (N_23566,N_21692,N_20625);
and U23567 (N_23567,N_20192,N_21246);
nor U23568 (N_23568,N_21839,N_20672);
xor U23569 (N_23569,N_20539,N_21308);
xnor U23570 (N_23570,N_21696,N_20647);
or U23571 (N_23571,N_21957,N_20301);
nand U23572 (N_23572,N_21386,N_20622);
and U23573 (N_23573,N_21644,N_21542);
xor U23574 (N_23574,N_20480,N_20080);
nor U23575 (N_23575,N_21554,N_21323);
xnor U23576 (N_23576,N_21687,N_20239);
xor U23577 (N_23577,N_20428,N_21527);
nand U23578 (N_23578,N_21015,N_20571);
or U23579 (N_23579,N_20681,N_20592);
nor U23580 (N_23580,N_20961,N_21948);
or U23581 (N_23581,N_21864,N_21121);
nand U23582 (N_23582,N_20755,N_21084);
xnor U23583 (N_23583,N_21540,N_21796);
nor U23584 (N_23584,N_20457,N_21329);
nand U23585 (N_23585,N_20183,N_20578);
and U23586 (N_23586,N_21638,N_21936);
and U23587 (N_23587,N_20286,N_20838);
and U23588 (N_23588,N_21844,N_20022);
xnor U23589 (N_23589,N_21303,N_20264);
and U23590 (N_23590,N_21368,N_20695);
nor U23591 (N_23591,N_20071,N_20363);
xor U23592 (N_23592,N_21512,N_21394);
xnor U23593 (N_23593,N_20341,N_20122);
nand U23594 (N_23594,N_21268,N_21629);
and U23595 (N_23595,N_20048,N_21337);
nor U23596 (N_23596,N_20607,N_21745);
nor U23597 (N_23597,N_21338,N_20590);
and U23598 (N_23598,N_21127,N_20287);
xnor U23599 (N_23599,N_20328,N_20019);
nor U23600 (N_23600,N_20372,N_21436);
xnor U23601 (N_23601,N_20285,N_21106);
and U23602 (N_23602,N_20890,N_21440);
xnor U23603 (N_23603,N_20930,N_20672);
nor U23604 (N_23604,N_20406,N_20504);
or U23605 (N_23605,N_20886,N_20228);
nor U23606 (N_23606,N_20348,N_21901);
nand U23607 (N_23607,N_21683,N_21243);
and U23608 (N_23608,N_21302,N_20378);
or U23609 (N_23609,N_20493,N_20950);
xnor U23610 (N_23610,N_20668,N_20106);
xnor U23611 (N_23611,N_20319,N_21500);
or U23612 (N_23612,N_20159,N_20967);
nor U23613 (N_23613,N_21173,N_20226);
nand U23614 (N_23614,N_20253,N_20957);
nor U23615 (N_23615,N_21384,N_20409);
nor U23616 (N_23616,N_20064,N_20914);
or U23617 (N_23617,N_20926,N_20884);
and U23618 (N_23618,N_21910,N_20964);
xnor U23619 (N_23619,N_20971,N_21996);
xor U23620 (N_23620,N_21198,N_20951);
xnor U23621 (N_23621,N_21659,N_21664);
or U23622 (N_23622,N_21397,N_20334);
nand U23623 (N_23623,N_20118,N_21086);
nor U23624 (N_23624,N_20450,N_21635);
xor U23625 (N_23625,N_21841,N_20333);
nand U23626 (N_23626,N_20563,N_20396);
nor U23627 (N_23627,N_21856,N_20760);
and U23628 (N_23628,N_20884,N_21573);
nor U23629 (N_23629,N_21019,N_20928);
or U23630 (N_23630,N_20226,N_20891);
and U23631 (N_23631,N_21918,N_21887);
and U23632 (N_23632,N_21905,N_20936);
xnor U23633 (N_23633,N_20279,N_21225);
or U23634 (N_23634,N_20987,N_21009);
xnor U23635 (N_23635,N_20646,N_20104);
nand U23636 (N_23636,N_21705,N_21547);
and U23637 (N_23637,N_20004,N_20478);
and U23638 (N_23638,N_20454,N_20621);
and U23639 (N_23639,N_20501,N_21079);
and U23640 (N_23640,N_21107,N_21332);
or U23641 (N_23641,N_20031,N_20555);
nor U23642 (N_23642,N_20463,N_20229);
nor U23643 (N_23643,N_21715,N_20814);
or U23644 (N_23644,N_21661,N_20609);
and U23645 (N_23645,N_20429,N_20768);
or U23646 (N_23646,N_21196,N_20962);
nand U23647 (N_23647,N_20533,N_21418);
nor U23648 (N_23648,N_21820,N_21233);
xor U23649 (N_23649,N_20439,N_21454);
and U23650 (N_23650,N_21295,N_20293);
nand U23651 (N_23651,N_21829,N_21851);
and U23652 (N_23652,N_20934,N_20832);
and U23653 (N_23653,N_20587,N_21419);
xnor U23654 (N_23654,N_21399,N_20998);
nand U23655 (N_23655,N_20297,N_20829);
nor U23656 (N_23656,N_20182,N_20083);
xnor U23657 (N_23657,N_20997,N_20706);
xnor U23658 (N_23658,N_21945,N_21726);
and U23659 (N_23659,N_20197,N_21956);
and U23660 (N_23660,N_20092,N_20442);
and U23661 (N_23661,N_20891,N_21257);
nor U23662 (N_23662,N_21955,N_21267);
and U23663 (N_23663,N_20581,N_20041);
and U23664 (N_23664,N_21827,N_20597);
and U23665 (N_23665,N_21037,N_20226);
and U23666 (N_23666,N_21444,N_21323);
nand U23667 (N_23667,N_20974,N_21624);
or U23668 (N_23668,N_21473,N_21113);
nor U23669 (N_23669,N_20406,N_20976);
or U23670 (N_23670,N_21130,N_21390);
and U23671 (N_23671,N_21039,N_20895);
or U23672 (N_23672,N_20512,N_21512);
nand U23673 (N_23673,N_21095,N_21175);
nand U23674 (N_23674,N_21159,N_20431);
and U23675 (N_23675,N_20507,N_21600);
or U23676 (N_23676,N_21733,N_20998);
and U23677 (N_23677,N_21681,N_20667);
nor U23678 (N_23678,N_20989,N_21114);
and U23679 (N_23679,N_21920,N_21056);
nor U23680 (N_23680,N_20658,N_21499);
and U23681 (N_23681,N_21257,N_20421);
nor U23682 (N_23682,N_21657,N_20121);
nand U23683 (N_23683,N_20801,N_20932);
nand U23684 (N_23684,N_21322,N_20700);
nand U23685 (N_23685,N_21152,N_20670);
nand U23686 (N_23686,N_20393,N_20725);
and U23687 (N_23687,N_20541,N_21983);
or U23688 (N_23688,N_21238,N_21621);
nand U23689 (N_23689,N_21559,N_21576);
or U23690 (N_23690,N_21384,N_21326);
and U23691 (N_23691,N_20761,N_21406);
nand U23692 (N_23692,N_21122,N_21693);
and U23693 (N_23693,N_20523,N_20662);
nand U23694 (N_23694,N_21781,N_20783);
and U23695 (N_23695,N_21941,N_21198);
and U23696 (N_23696,N_20441,N_20238);
and U23697 (N_23697,N_20655,N_21404);
and U23698 (N_23698,N_21382,N_21429);
or U23699 (N_23699,N_21624,N_21818);
or U23700 (N_23700,N_21287,N_20294);
xor U23701 (N_23701,N_20104,N_20507);
nor U23702 (N_23702,N_20209,N_21736);
nand U23703 (N_23703,N_20344,N_20606);
xor U23704 (N_23704,N_21015,N_20101);
and U23705 (N_23705,N_20713,N_21264);
and U23706 (N_23706,N_21564,N_21031);
nand U23707 (N_23707,N_21378,N_20979);
nand U23708 (N_23708,N_20867,N_20950);
nand U23709 (N_23709,N_21827,N_20519);
xor U23710 (N_23710,N_21054,N_21056);
xor U23711 (N_23711,N_21042,N_20478);
nand U23712 (N_23712,N_21906,N_20105);
nor U23713 (N_23713,N_20640,N_20525);
and U23714 (N_23714,N_20683,N_20442);
xor U23715 (N_23715,N_21303,N_20488);
nand U23716 (N_23716,N_21691,N_21702);
and U23717 (N_23717,N_20569,N_20163);
and U23718 (N_23718,N_20129,N_20278);
nor U23719 (N_23719,N_20159,N_20202);
nor U23720 (N_23720,N_21883,N_21026);
nand U23721 (N_23721,N_20019,N_20867);
and U23722 (N_23722,N_21071,N_20033);
nor U23723 (N_23723,N_20887,N_20648);
and U23724 (N_23724,N_21978,N_20582);
or U23725 (N_23725,N_20583,N_20572);
nor U23726 (N_23726,N_21317,N_20221);
xnor U23727 (N_23727,N_21787,N_20290);
and U23728 (N_23728,N_20853,N_20230);
or U23729 (N_23729,N_20653,N_21115);
nor U23730 (N_23730,N_20617,N_21864);
nand U23731 (N_23731,N_21936,N_20655);
nand U23732 (N_23732,N_20744,N_20920);
nand U23733 (N_23733,N_21516,N_21757);
nor U23734 (N_23734,N_20559,N_20634);
nor U23735 (N_23735,N_21639,N_21258);
nor U23736 (N_23736,N_20826,N_20542);
nor U23737 (N_23737,N_20415,N_21385);
nor U23738 (N_23738,N_21417,N_20219);
or U23739 (N_23739,N_21972,N_20083);
and U23740 (N_23740,N_20497,N_20740);
xor U23741 (N_23741,N_21335,N_20593);
or U23742 (N_23742,N_21079,N_21803);
xor U23743 (N_23743,N_21291,N_21722);
nor U23744 (N_23744,N_20996,N_20894);
or U23745 (N_23745,N_21117,N_20348);
xor U23746 (N_23746,N_20437,N_20299);
xnor U23747 (N_23747,N_21850,N_21673);
and U23748 (N_23748,N_21248,N_21988);
nand U23749 (N_23749,N_20237,N_20343);
and U23750 (N_23750,N_20142,N_21123);
nor U23751 (N_23751,N_20888,N_21505);
or U23752 (N_23752,N_21012,N_21414);
or U23753 (N_23753,N_21084,N_21318);
xor U23754 (N_23754,N_21736,N_20331);
xnor U23755 (N_23755,N_21852,N_21014);
xor U23756 (N_23756,N_21919,N_21432);
nor U23757 (N_23757,N_20419,N_20180);
nand U23758 (N_23758,N_21466,N_20141);
xnor U23759 (N_23759,N_20887,N_21251);
or U23760 (N_23760,N_21799,N_21843);
and U23761 (N_23761,N_20829,N_21820);
or U23762 (N_23762,N_21745,N_20006);
or U23763 (N_23763,N_20647,N_20479);
xnor U23764 (N_23764,N_20775,N_20747);
or U23765 (N_23765,N_21137,N_21198);
or U23766 (N_23766,N_21715,N_20977);
or U23767 (N_23767,N_21414,N_21988);
or U23768 (N_23768,N_21669,N_20231);
or U23769 (N_23769,N_21812,N_20417);
or U23770 (N_23770,N_20768,N_21482);
nand U23771 (N_23771,N_20390,N_21433);
nor U23772 (N_23772,N_20620,N_20282);
and U23773 (N_23773,N_21964,N_20685);
or U23774 (N_23774,N_21076,N_20879);
nand U23775 (N_23775,N_20336,N_20940);
xor U23776 (N_23776,N_20101,N_20345);
and U23777 (N_23777,N_20932,N_21366);
or U23778 (N_23778,N_20763,N_21307);
or U23779 (N_23779,N_20981,N_20787);
nand U23780 (N_23780,N_20119,N_20409);
and U23781 (N_23781,N_20737,N_21449);
or U23782 (N_23782,N_20399,N_21913);
nor U23783 (N_23783,N_20537,N_21842);
or U23784 (N_23784,N_20090,N_21238);
nor U23785 (N_23785,N_20093,N_20724);
nand U23786 (N_23786,N_21341,N_21223);
or U23787 (N_23787,N_20180,N_20964);
xnor U23788 (N_23788,N_20819,N_20304);
xnor U23789 (N_23789,N_20572,N_21370);
nor U23790 (N_23790,N_21700,N_20620);
nor U23791 (N_23791,N_20725,N_21306);
nor U23792 (N_23792,N_20329,N_21635);
and U23793 (N_23793,N_20936,N_21564);
and U23794 (N_23794,N_20793,N_21219);
nand U23795 (N_23795,N_21271,N_21548);
nand U23796 (N_23796,N_21540,N_21937);
xnor U23797 (N_23797,N_21596,N_21739);
nor U23798 (N_23798,N_20489,N_21605);
or U23799 (N_23799,N_20628,N_20538);
nor U23800 (N_23800,N_21947,N_20914);
and U23801 (N_23801,N_20568,N_20565);
nor U23802 (N_23802,N_21751,N_20903);
and U23803 (N_23803,N_21862,N_20396);
nor U23804 (N_23804,N_21661,N_20058);
and U23805 (N_23805,N_21114,N_21820);
nand U23806 (N_23806,N_21244,N_20450);
nand U23807 (N_23807,N_20109,N_21337);
and U23808 (N_23808,N_20688,N_21280);
nor U23809 (N_23809,N_21474,N_20618);
nor U23810 (N_23810,N_20142,N_20818);
nor U23811 (N_23811,N_20593,N_20422);
nand U23812 (N_23812,N_21285,N_21976);
xor U23813 (N_23813,N_20881,N_20212);
nor U23814 (N_23814,N_21598,N_21232);
or U23815 (N_23815,N_21871,N_20825);
nand U23816 (N_23816,N_21526,N_20115);
and U23817 (N_23817,N_20186,N_20835);
nand U23818 (N_23818,N_20566,N_20108);
and U23819 (N_23819,N_21586,N_21295);
nand U23820 (N_23820,N_20341,N_21176);
xnor U23821 (N_23821,N_20385,N_20832);
xor U23822 (N_23822,N_21433,N_21745);
nor U23823 (N_23823,N_20626,N_20525);
or U23824 (N_23824,N_21311,N_21802);
nand U23825 (N_23825,N_20654,N_20283);
and U23826 (N_23826,N_21728,N_21291);
and U23827 (N_23827,N_21282,N_20248);
or U23828 (N_23828,N_21714,N_21421);
nand U23829 (N_23829,N_20251,N_20855);
nand U23830 (N_23830,N_20478,N_21346);
nand U23831 (N_23831,N_21306,N_21395);
and U23832 (N_23832,N_21841,N_20136);
xor U23833 (N_23833,N_21384,N_20987);
or U23834 (N_23834,N_21355,N_20437);
or U23835 (N_23835,N_20582,N_21399);
or U23836 (N_23836,N_21595,N_20338);
nor U23837 (N_23837,N_21251,N_20400);
or U23838 (N_23838,N_20892,N_20798);
and U23839 (N_23839,N_20037,N_20794);
xor U23840 (N_23840,N_20188,N_21206);
nor U23841 (N_23841,N_20319,N_20124);
nor U23842 (N_23842,N_21748,N_20621);
or U23843 (N_23843,N_20984,N_21158);
xor U23844 (N_23844,N_21550,N_21547);
nor U23845 (N_23845,N_21652,N_21089);
and U23846 (N_23846,N_21402,N_20131);
nand U23847 (N_23847,N_21451,N_21224);
or U23848 (N_23848,N_21234,N_20346);
or U23849 (N_23849,N_20349,N_21790);
xor U23850 (N_23850,N_21020,N_20493);
xnor U23851 (N_23851,N_21192,N_21721);
nand U23852 (N_23852,N_20414,N_20884);
and U23853 (N_23853,N_21727,N_21015);
nor U23854 (N_23854,N_21110,N_21689);
xor U23855 (N_23855,N_21257,N_21923);
and U23856 (N_23856,N_20309,N_21413);
and U23857 (N_23857,N_20232,N_21711);
nor U23858 (N_23858,N_21031,N_20634);
nand U23859 (N_23859,N_20715,N_20841);
and U23860 (N_23860,N_21437,N_21064);
and U23861 (N_23861,N_20087,N_20005);
xor U23862 (N_23862,N_21210,N_20281);
nor U23863 (N_23863,N_21943,N_21656);
nand U23864 (N_23864,N_20859,N_21723);
xor U23865 (N_23865,N_21449,N_21866);
nand U23866 (N_23866,N_21438,N_20491);
nand U23867 (N_23867,N_21020,N_21328);
or U23868 (N_23868,N_20454,N_21501);
xor U23869 (N_23869,N_21865,N_21235);
nand U23870 (N_23870,N_20837,N_21149);
nand U23871 (N_23871,N_20774,N_21715);
nor U23872 (N_23872,N_20231,N_21418);
or U23873 (N_23873,N_20202,N_21714);
nor U23874 (N_23874,N_20992,N_21555);
xnor U23875 (N_23875,N_20034,N_20223);
and U23876 (N_23876,N_21125,N_21021);
nand U23877 (N_23877,N_21356,N_20567);
nand U23878 (N_23878,N_21764,N_20325);
nor U23879 (N_23879,N_21910,N_21961);
and U23880 (N_23880,N_21948,N_21449);
nand U23881 (N_23881,N_21832,N_20053);
and U23882 (N_23882,N_20978,N_20452);
and U23883 (N_23883,N_21122,N_20957);
nor U23884 (N_23884,N_20497,N_21209);
nor U23885 (N_23885,N_21997,N_20518);
nor U23886 (N_23886,N_21435,N_20272);
nand U23887 (N_23887,N_20788,N_21859);
nand U23888 (N_23888,N_21624,N_20025);
nand U23889 (N_23889,N_20475,N_21927);
and U23890 (N_23890,N_20765,N_20209);
nand U23891 (N_23891,N_20621,N_21931);
nand U23892 (N_23892,N_20436,N_21495);
and U23893 (N_23893,N_20168,N_20026);
nand U23894 (N_23894,N_21556,N_21331);
nand U23895 (N_23895,N_20149,N_21275);
nand U23896 (N_23896,N_20264,N_21497);
or U23897 (N_23897,N_21589,N_21939);
xor U23898 (N_23898,N_21962,N_20786);
nand U23899 (N_23899,N_20031,N_20718);
or U23900 (N_23900,N_21657,N_20961);
and U23901 (N_23901,N_21943,N_21285);
nand U23902 (N_23902,N_21158,N_20387);
nand U23903 (N_23903,N_20135,N_20681);
and U23904 (N_23904,N_20540,N_21507);
nor U23905 (N_23905,N_21295,N_21691);
and U23906 (N_23906,N_21165,N_20530);
nand U23907 (N_23907,N_21311,N_21818);
nand U23908 (N_23908,N_20884,N_20542);
nor U23909 (N_23909,N_20332,N_20999);
or U23910 (N_23910,N_21768,N_20374);
nand U23911 (N_23911,N_21939,N_20306);
and U23912 (N_23912,N_21003,N_20012);
xnor U23913 (N_23913,N_20769,N_20549);
and U23914 (N_23914,N_20258,N_20954);
and U23915 (N_23915,N_21540,N_21464);
and U23916 (N_23916,N_20866,N_21619);
nand U23917 (N_23917,N_21741,N_21370);
and U23918 (N_23918,N_20433,N_20653);
nor U23919 (N_23919,N_20536,N_20456);
nor U23920 (N_23920,N_21834,N_21415);
nand U23921 (N_23921,N_21451,N_21824);
nand U23922 (N_23922,N_21287,N_20753);
or U23923 (N_23923,N_21818,N_21673);
xnor U23924 (N_23924,N_20987,N_20527);
nor U23925 (N_23925,N_21786,N_21851);
nand U23926 (N_23926,N_21029,N_20068);
nor U23927 (N_23927,N_21422,N_20242);
and U23928 (N_23928,N_20773,N_21549);
and U23929 (N_23929,N_20767,N_20574);
nor U23930 (N_23930,N_21672,N_21804);
nor U23931 (N_23931,N_20160,N_21550);
or U23932 (N_23932,N_21442,N_21743);
nor U23933 (N_23933,N_20621,N_21137);
nand U23934 (N_23934,N_21974,N_20941);
nand U23935 (N_23935,N_21896,N_21007);
or U23936 (N_23936,N_20059,N_20199);
and U23937 (N_23937,N_21190,N_20461);
or U23938 (N_23938,N_21106,N_20580);
or U23939 (N_23939,N_21041,N_20129);
and U23940 (N_23940,N_21560,N_21261);
nand U23941 (N_23941,N_21053,N_20760);
or U23942 (N_23942,N_20059,N_21121);
nor U23943 (N_23943,N_20560,N_20151);
xor U23944 (N_23944,N_20332,N_20022);
nand U23945 (N_23945,N_20586,N_21291);
nand U23946 (N_23946,N_20844,N_21129);
nor U23947 (N_23947,N_21622,N_20360);
nor U23948 (N_23948,N_20845,N_20351);
and U23949 (N_23949,N_21414,N_21350);
or U23950 (N_23950,N_21029,N_20872);
and U23951 (N_23951,N_20484,N_21464);
and U23952 (N_23952,N_20046,N_20871);
and U23953 (N_23953,N_20057,N_20655);
and U23954 (N_23954,N_21752,N_21400);
nand U23955 (N_23955,N_20349,N_20637);
xor U23956 (N_23956,N_20375,N_21486);
xor U23957 (N_23957,N_21587,N_20388);
xor U23958 (N_23958,N_21861,N_20981);
xor U23959 (N_23959,N_21642,N_20281);
nand U23960 (N_23960,N_21260,N_21629);
nor U23961 (N_23961,N_21536,N_20585);
nor U23962 (N_23962,N_21687,N_20366);
xor U23963 (N_23963,N_20544,N_20812);
xnor U23964 (N_23964,N_20792,N_20381);
nand U23965 (N_23965,N_20300,N_20108);
nand U23966 (N_23966,N_20187,N_20989);
nand U23967 (N_23967,N_20906,N_20050);
nand U23968 (N_23968,N_20387,N_21049);
xnor U23969 (N_23969,N_21294,N_21279);
nand U23970 (N_23970,N_20651,N_21414);
and U23971 (N_23971,N_20268,N_20701);
and U23972 (N_23972,N_20844,N_21880);
nor U23973 (N_23973,N_21438,N_20000);
or U23974 (N_23974,N_21418,N_20822);
or U23975 (N_23975,N_21112,N_20617);
xnor U23976 (N_23976,N_21168,N_20687);
or U23977 (N_23977,N_20423,N_20212);
or U23978 (N_23978,N_20833,N_21465);
and U23979 (N_23979,N_20821,N_20797);
or U23980 (N_23980,N_20292,N_21639);
or U23981 (N_23981,N_20441,N_21648);
nor U23982 (N_23982,N_20893,N_21934);
nand U23983 (N_23983,N_20912,N_21060);
nand U23984 (N_23984,N_20829,N_20934);
or U23985 (N_23985,N_20411,N_20394);
nand U23986 (N_23986,N_21764,N_20378);
and U23987 (N_23987,N_20073,N_21936);
nand U23988 (N_23988,N_20195,N_21132);
nor U23989 (N_23989,N_21705,N_21747);
xor U23990 (N_23990,N_21244,N_20674);
and U23991 (N_23991,N_20467,N_21643);
nor U23992 (N_23992,N_20810,N_20331);
xnor U23993 (N_23993,N_20137,N_21347);
xnor U23994 (N_23994,N_21444,N_20923);
and U23995 (N_23995,N_21631,N_21814);
nand U23996 (N_23996,N_21719,N_20510);
and U23997 (N_23997,N_20589,N_21595);
or U23998 (N_23998,N_21440,N_20329);
and U23999 (N_23999,N_21761,N_21236);
and U24000 (N_24000,N_22175,N_23801);
or U24001 (N_24001,N_22209,N_23366);
and U24002 (N_24002,N_23594,N_22020);
xnor U24003 (N_24003,N_22512,N_23315);
and U24004 (N_24004,N_23168,N_23376);
xor U24005 (N_24005,N_23737,N_23600);
nor U24006 (N_24006,N_23441,N_22719);
and U24007 (N_24007,N_23920,N_22038);
and U24008 (N_24008,N_23443,N_22960);
or U24009 (N_24009,N_22758,N_22154);
nand U24010 (N_24010,N_22176,N_23005);
or U24011 (N_24011,N_23375,N_23985);
or U24012 (N_24012,N_23291,N_22032);
nand U24013 (N_24013,N_22065,N_22316);
nand U24014 (N_24014,N_22818,N_23653);
xor U24015 (N_24015,N_22448,N_22507);
or U24016 (N_24016,N_22616,N_23983);
and U24017 (N_24017,N_23553,N_22618);
or U24018 (N_24018,N_23473,N_23405);
xnor U24019 (N_24019,N_23141,N_22643);
and U24020 (N_24020,N_23064,N_23084);
nand U24021 (N_24021,N_23794,N_22264);
nand U24022 (N_24022,N_23911,N_22619);
nor U24023 (N_24023,N_22040,N_22509);
xor U24024 (N_24024,N_22735,N_23847);
and U24025 (N_24025,N_22183,N_23127);
nor U24026 (N_24026,N_23555,N_22345);
nor U24027 (N_24027,N_23055,N_22901);
nor U24028 (N_24028,N_23446,N_22674);
nand U24029 (N_24029,N_23837,N_22562);
nand U24030 (N_24030,N_23433,N_23564);
or U24031 (N_24031,N_23213,N_23595);
and U24032 (N_24032,N_22381,N_23276);
and U24033 (N_24033,N_23768,N_23569);
nand U24034 (N_24034,N_23043,N_23807);
nand U24035 (N_24035,N_23943,N_23512);
xnor U24036 (N_24036,N_22339,N_23390);
xnor U24037 (N_24037,N_22829,N_23821);
or U24038 (N_24038,N_23026,N_22320);
xnor U24039 (N_24039,N_22426,N_23840);
nand U24040 (N_24040,N_22514,N_23571);
nor U24041 (N_24041,N_23203,N_23301);
and U24042 (N_24042,N_22579,N_23058);
and U24043 (N_24043,N_23435,N_23293);
or U24044 (N_24044,N_22539,N_23228);
xnor U24045 (N_24045,N_23237,N_22041);
nor U24046 (N_24046,N_22469,N_23897);
and U24047 (N_24047,N_23535,N_22855);
nand U24048 (N_24048,N_22178,N_22170);
and U24049 (N_24049,N_23580,N_22651);
nand U24050 (N_24050,N_22993,N_22105);
or U24051 (N_24051,N_23965,N_23490);
nand U24052 (N_24052,N_23025,N_22498);
nor U24053 (N_24053,N_22683,N_23835);
nor U24054 (N_24054,N_22204,N_22408);
xor U24055 (N_24055,N_22113,N_22473);
or U24056 (N_24056,N_23744,N_22784);
or U24057 (N_24057,N_23368,N_22091);
or U24058 (N_24058,N_23697,N_22368);
nand U24059 (N_24059,N_23392,N_23621);
and U24060 (N_24060,N_22648,N_22018);
and U24061 (N_24061,N_23789,N_23513);
nand U24062 (N_24062,N_22827,N_22314);
nor U24063 (N_24063,N_22751,N_22394);
xnor U24064 (N_24064,N_23129,N_23545);
xor U24065 (N_24065,N_23982,N_22110);
xnor U24066 (N_24066,N_22047,N_23485);
or U24067 (N_24067,N_23028,N_22013);
or U24068 (N_24068,N_23489,N_22627);
xnor U24069 (N_24069,N_23936,N_22897);
nand U24070 (N_24070,N_22021,N_23908);
nand U24071 (N_24071,N_22807,N_22131);
xor U24072 (N_24072,N_22198,N_23461);
and U24073 (N_24073,N_23664,N_23302);
and U24074 (N_24074,N_22816,N_22395);
or U24075 (N_24075,N_23748,N_23822);
or U24076 (N_24076,N_22919,N_23811);
nand U24077 (N_24077,N_23330,N_23316);
xnor U24078 (N_24078,N_23514,N_22104);
nor U24079 (N_24079,N_22242,N_23635);
xnor U24080 (N_24080,N_23468,N_23479);
nand U24081 (N_24081,N_22798,N_23460);
nor U24082 (N_24082,N_23373,N_22281);
or U24083 (N_24083,N_23296,N_23264);
xnor U24084 (N_24084,N_23171,N_23824);
and U24085 (N_24085,N_23627,N_23029);
nand U24086 (N_24086,N_23888,N_22039);
xor U24087 (N_24087,N_23367,N_23357);
and U24088 (N_24088,N_22321,N_22950);
or U24089 (N_24089,N_22666,N_22903);
nor U24090 (N_24090,N_23363,N_22348);
nand U24091 (N_24091,N_22747,N_23284);
nand U24092 (N_24092,N_22467,N_22443);
nor U24093 (N_24093,N_23123,N_23205);
xnor U24094 (N_24094,N_22911,N_22981);
nor U24095 (N_24095,N_23458,N_22384);
nor U24096 (N_24096,N_22416,N_23322);
nand U24097 (N_24097,N_23387,N_23371);
nand U24098 (N_24098,N_22315,N_22307);
and U24099 (N_24099,N_22774,N_22062);
and U24100 (N_24100,N_23360,N_22262);
or U24101 (N_24101,N_23786,N_23834);
and U24102 (N_24102,N_22725,N_23260);
nand U24103 (N_24103,N_23364,N_22077);
xnor U24104 (N_24104,N_23581,N_23465);
xnor U24105 (N_24105,N_22708,N_22332);
and U24106 (N_24106,N_22777,N_22780);
or U24107 (N_24107,N_22924,N_23544);
nor U24108 (N_24108,N_22210,N_23082);
or U24109 (N_24109,N_22859,N_23754);
or U24110 (N_24110,N_22485,N_23727);
nor U24111 (N_24111,N_23157,N_23286);
nand U24112 (N_24112,N_22613,N_23212);
or U24113 (N_24113,N_23350,N_23527);
nor U24114 (N_24114,N_22603,N_23843);
xor U24115 (N_24115,N_22707,N_22456);
or U24116 (N_24116,N_22940,N_22205);
nor U24117 (N_24117,N_23399,N_22119);
nor U24118 (N_24118,N_23955,N_22896);
nor U24119 (N_24119,N_23742,N_22145);
nor U24120 (N_24120,N_22904,N_22334);
or U24121 (N_24121,N_23230,N_23942);
and U24122 (N_24122,N_22082,N_22474);
or U24123 (N_24123,N_23875,N_22789);
xnor U24124 (N_24124,N_23802,N_22785);
xor U24125 (N_24125,N_22948,N_22906);
and U24126 (N_24126,N_22809,N_23677);
xnor U24127 (N_24127,N_22609,N_22560);
and U24128 (N_24128,N_22865,N_23803);
and U24129 (N_24129,N_22084,N_22050);
or U24130 (N_24130,N_23753,N_22826);
or U24131 (N_24131,N_23013,N_23074);
nand U24132 (N_24132,N_23238,N_23975);
nor U24133 (N_24133,N_22893,N_23844);
or U24134 (N_24134,N_22515,N_22757);
and U24135 (N_24135,N_22773,N_23019);
nor U24136 (N_24136,N_22994,N_22716);
and U24137 (N_24137,N_23703,N_22420);
or U24138 (N_24138,N_22094,N_22941);
nand U24139 (N_24139,N_23234,N_23765);
or U24140 (N_24140,N_22524,N_23928);
or U24141 (N_24141,N_22186,N_23109);
xnor U24142 (N_24142,N_23216,N_22962);
and U24143 (N_24143,N_23472,N_22997);
or U24144 (N_24144,N_22857,N_22260);
or U24145 (N_24145,N_23440,N_22202);
nor U24146 (N_24146,N_23892,N_23944);
or U24147 (N_24147,N_22935,N_22810);
nand U24148 (N_24148,N_22429,N_22023);
xor U24149 (N_24149,N_22567,N_23693);
xor U24150 (N_24150,N_22814,N_23099);
xnor U24151 (N_24151,N_23759,N_23780);
nor U24152 (N_24152,N_22561,N_22090);
or U24153 (N_24153,N_22134,N_22410);
nor U24154 (N_24154,N_23561,N_22949);
or U24155 (N_24155,N_22190,N_22532);
nand U24156 (N_24156,N_23201,N_22102);
nor U24157 (N_24157,N_23529,N_23917);
nand U24158 (N_24158,N_23377,N_23143);
xor U24159 (N_24159,N_23991,N_22054);
xor U24160 (N_24160,N_23404,N_22852);
xor U24161 (N_24161,N_22885,N_22843);
nand U24162 (N_24162,N_22379,N_22750);
nand U24163 (N_24163,N_23935,N_23263);
or U24164 (N_24164,N_22057,N_23140);
nor U24165 (N_24165,N_23723,N_22215);
and U24166 (N_24166,N_22024,N_22098);
or U24167 (N_24167,N_23117,N_23102);
nor U24168 (N_24168,N_22166,N_22076);
nor U24169 (N_24169,N_22414,N_22171);
nor U24170 (N_24170,N_22046,N_23321);
or U24171 (N_24171,N_22733,N_22646);
xnor U24172 (N_24172,N_23610,N_22053);
nand U24173 (N_24173,N_23093,N_23503);
nand U24174 (N_24174,N_23732,N_22351);
nor U24175 (N_24175,N_22069,N_23617);
nand U24176 (N_24176,N_23320,N_23439);
or U24177 (N_24177,N_22159,N_22302);
nand U24178 (N_24178,N_23338,N_23968);
xnor U24179 (N_24179,N_22397,N_23332);
nand U24180 (N_24180,N_22476,N_22608);
nor U24181 (N_24181,N_22718,N_22662);
xor U24182 (N_24182,N_23724,N_22804);
and U24183 (N_24183,N_22959,N_23671);
nor U24184 (N_24184,N_23730,N_22311);
xnor U24185 (N_24185,N_22723,N_22991);
nor U24186 (N_24186,N_22915,N_23656);
nor U24187 (N_24187,N_23112,N_23662);
nor U24188 (N_24188,N_22495,N_23182);
or U24189 (N_24189,N_23583,N_22724);
xor U24190 (N_24190,N_22889,N_22005);
xnor U24191 (N_24191,N_23997,N_22520);
nand U24192 (N_24192,N_22530,N_23506);
nor U24193 (N_24193,N_23156,N_22235);
nand U24194 (N_24194,N_23006,N_23938);
or U24195 (N_24195,N_22390,N_22582);
and U24196 (N_24196,N_23590,N_22160);
xnor U24197 (N_24197,N_22033,N_23962);
nor U24198 (N_24198,N_22820,N_23195);
xor U24199 (N_24199,N_23577,N_22398);
nand U24200 (N_24200,N_22667,N_22905);
or U24201 (N_24201,N_22064,N_23179);
or U24202 (N_24202,N_22161,N_23176);
xor U24203 (N_24203,N_22966,N_23777);
nand U24204 (N_24204,N_23136,N_23873);
nand U24205 (N_24205,N_22342,N_22846);
nand U24206 (N_24206,N_22551,N_22872);
nor U24207 (N_24207,N_23563,N_23045);
and U24208 (N_24208,N_22549,N_22523);
nor U24209 (N_24209,N_23694,N_23153);
xor U24210 (N_24210,N_23356,N_22477);
and U24211 (N_24211,N_23898,N_22411);
nand U24212 (N_24212,N_22006,N_23189);
nand U24213 (N_24213,N_23731,N_23313);
or U24214 (N_24214,N_23670,N_22769);
or U24215 (N_24215,N_22251,N_22120);
and U24216 (N_24216,N_22987,N_22317);
nor U24217 (N_24217,N_23023,N_23741);
nor U24218 (N_24218,N_22830,N_23954);
and U24219 (N_24219,N_23809,N_23776);
nand U24220 (N_24220,N_23124,N_22799);
and U24221 (N_24221,N_23094,N_23036);
and U24222 (N_24222,N_22553,N_22241);
nor U24223 (N_24223,N_23134,N_23532);
nor U24224 (N_24224,N_22211,N_23980);
xnor U24225 (N_24225,N_22179,N_23781);
nand U24226 (N_24226,N_22552,N_22833);
nor U24227 (N_24227,N_22934,N_23509);
and U24228 (N_24228,N_22276,N_23862);
or U24229 (N_24229,N_22459,N_22151);
nor U24230 (N_24230,N_23174,N_23418);
and U24231 (N_24231,N_23582,N_23714);
nor U24232 (N_24232,N_22462,N_23804);
or U24233 (N_24233,N_22030,N_23778);
or U24234 (N_24234,N_22431,N_22932);
nor U24235 (N_24235,N_23300,N_22045);
nor U24236 (N_24236,N_23256,N_22984);
or U24237 (N_24237,N_23130,N_23218);
nand U24238 (N_24238,N_23848,N_23783);
xnor U24239 (N_24239,N_22741,N_23831);
xor U24240 (N_24240,N_22870,N_23388);
and U24241 (N_24241,N_23374,N_23918);
or U24242 (N_24242,N_22709,N_22936);
xnor U24243 (N_24243,N_23990,N_22008);
or U24244 (N_24244,N_23961,N_23312);
nand U24245 (N_24245,N_23568,N_23247);
and U24246 (N_24246,N_23257,N_22300);
xnor U24247 (N_24247,N_22093,N_22261);
and U24248 (N_24248,N_23262,N_22740);
xnor U24249 (N_24249,N_23103,N_23370);
xor U24250 (N_24250,N_23608,N_22029);
xor U24251 (N_24251,N_23163,N_22330);
nor U24252 (N_24252,N_23429,N_22336);
and U24253 (N_24253,N_23198,N_22765);
nand U24254 (N_24254,N_23210,N_23947);
xor U24255 (N_24255,N_23842,N_23530);
nor U24256 (N_24256,N_23447,N_22286);
and U24257 (N_24257,N_22571,N_22191);
nor U24258 (N_24258,N_22611,N_23869);
and U24259 (N_24259,N_23823,N_23927);
nor U24260 (N_24260,N_22668,N_22726);
and U24261 (N_24261,N_23814,N_22764);
and U24262 (N_24262,N_22458,N_22468);
nor U24263 (N_24263,N_22306,N_22989);
nor U24264 (N_24264,N_22886,N_22871);
xnor U24265 (N_24265,N_22631,N_22676);
nand U24266 (N_24266,N_23164,N_22890);
nor U24267 (N_24267,N_22192,N_23067);
or U24268 (N_24268,N_23646,N_22635);
nor U24269 (N_24269,N_22877,N_22388);
nor U24270 (N_24270,N_23243,N_22963);
nand U24271 (N_24271,N_23524,N_23734);
nand U24272 (N_24272,N_23402,N_23540);
nor U24273 (N_24273,N_22358,N_23434);
or U24274 (N_24274,N_22437,N_23861);
xnor U24275 (N_24275,N_22930,N_23069);
and U24276 (N_24276,N_23467,N_23596);
nand U24277 (N_24277,N_23208,N_22895);
or U24278 (N_24278,N_23283,N_22569);
or U24279 (N_24279,N_23348,N_22548);
and U24280 (N_24280,N_22768,N_22137);
and U24281 (N_24281,N_23755,N_23122);
nand U24282 (N_24282,N_23705,N_23516);
xor U24283 (N_24283,N_22664,N_22689);
and U24284 (N_24284,N_23624,N_22292);
or U24285 (N_24285,N_22815,N_23344);
nand U24286 (N_24286,N_23591,N_22428);
nand U24287 (N_24287,N_22386,N_23976);
nand U24288 (N_24288,N_23452,N_22898);
xnor U24289 (N_24289,N_22783,N_22844);
nor U24290 (N_24290,N_22506,N_22673);
and U24291 (N_24291,N_22834,N_23340);
or U24292 (N_24292,N_22913,N_23598);
or U24293 (N_24293,N_22229,N_23630);
xor U24294 (N_24294,N_23901,N_22187);
nand U24295 (N_24295,N_23265,N_22055);
nor U24296 (N_24296,N_23793,N_23269);
or U24297 (N_24297,N_23159,N_23343);
or U24298 (N_24298,N_23412,N_22189);
or U24299 (N_24299,N_22049,N_23702);
xor U24300 (N_24300,N_22801,N_23658);
nor U24301 (N_24301,N_22604,N_22883);
or U24302 (N_24302,N_23011,N_22167);
xor U24303 (N_24303,N_23915,N_23096);
xor U24304 (N_24304,N_23791,N_23144);
nand U24305 (N_24305,N_23424,N_23764);
and U24306 (N_24306,N_23682,N_23054);
nand U24307 (N_24307,N_23491,N_22923);
and U24308 (N_24308,N_22945,N_22858);
or U24309 (N_24309,N_22121,N_23053);
or U24310 (N_24310,N_23146,N_22944);
or U24311 (N_24311,N_23692,N_23119);
nor U24312 (N_24312,N_23634,N_23337);
xnor U24313 (N_24313,N_22142,N_22586);
xor U24314 (N_24314,N_22168,N_22968);
nand U24315 (N_24315,N_22628,N_22811);
or U24316 (N_24316,N_22231,N_23197);
xnor U24317 (N_24317,N_22266,N_22755);
nand U24318 (N_24318,N_23819,N_23139);
nand U24319 (N_24319,N_22412,N_22600);
and U24320 (N_24320,N_22624,N_22658);
nand U24321 (N_24321,N_23044,N_23346);
nor U24322 (N_24322,N_22869,N_22237);
nand U24323 (N_24323,N_22224,N_22117);
nor U24324 (N_24324,N_23014,N_23537);
and U24325 (N_24325,N_23267,N_22044);
nand U24326 (N_24326,N_23929,N_22744);
nor U24327 (N_24327,N_22291,N_22681);
nor U24328 (N_24328,N_22756,N_23871);
nor U24329 (N_24329,N_23609,N_23946);
and U24330 (N_24330,N_23355,N_23104);
and U24331 (N_24331,N_22988,N_23105);
or U24332 (N_24332,N_23413,N_23685);
and U24333 (N_24333,N_22075,N_23451);
nand U24334 (N_24334,N_23747,N_23017);
nor U24335 (N_24335,N_22123,N_22761);
nor U24336 (N_24336,N_22165,N_23684);
xnor U24337 (N_24337,N_23533,N_23718);
nand U24338 (N_24338,N_22876,N_23739);
xnor U24339 (N_24339,N_23242,N_22699);
or U24340 (N_24340,N_22639,N_22116);
and U24341 (N_24341,N_23538,N_23632);
nor U24342 (N_24342,N_23675,N_23852);
and U24343 (N_24343,N_23279,N_22650);
nand U24344 (N_24344,N_22684,N_23554);
or U24345 (N_24345,N_23957,N_22440);
nor U24346 (N_24346,N_23637,N_22956);
nand U24347 (N_24347,N_23978,N_23445);
xnor U24348 (N_24348,N_22982,N_22796);
nor U24349 (N_24349,N_22623,N_23361);
xnor U24350 (N_24350,N_23573,N_22554);
and U24351 (N_24351,N_23190,N_23880);
xor U24352 (N_24352,N_22418,N_22902);
nor U24353 (N_24353,N_23057,N_23650);
nand U24354 (N_24354,N_22433,N_23981);
xor U24355 (N_24355,N_23798,N_22965);
nor U24356 (N_24356,N_22655,N_23454);
xnor U24357 (N_24357,N_22369,N_22068);
or U24358 (N_24358,N_22775,N_23347);
or U24359 (N_24359,N_23743,N_23790);
xnor U24360 (N_24360,N_23108,N_23953);
or U24361 (N_24361,N_22878,N_23958);
nand U24362 (N_24362,N_23972,N_23241);
nand U24363 (N_24363,N_22017,N_22975);
and U24364 (N_24364,N_23261,N_22702);
and U24365 (N_24365,N_22337,N_22731);
xor U24366 (N_24366,N_22759,N_23235);
xnor U24367 (N_24367,N_23772,N_23004);
xor U24368 (N_24368,N_23504,N_23931);
nor U24369 (N_24369,N_23900,N_23073);
nand U24370 (N_24370,N_22971,N_22313);
xnor U24371 (N_24371,N_23948,N_23172);
or U24372 (N_24372,N_22977,N_23353);
or U24373 (N_24373,N_23906,N_22602);
and U24374 (N_24374,N_22239,N_22067);
xnor U24375 (N_24375,N_22483,N_22823);
xor U24376 (N_24376,N_22481,N_23185);
and U24377 (N_24377,N_22347,N_23184);
xor U24378 (N_24378,N_22464,N_22280);
nand U24379 (N_24379,N_22095,N_23706);
nor U24380 (N_24380,N_23863,N_22625);
and U24381 (N_24381,N_23531,N_22088);
nor U24382 (N_24382,N_22802,N_22103);
xor U24383 (N_24383,N_23226,N_22772);
and U24384 (N_24384,N_22853,N_22144);
and U24385 (N_24385,N_22370,N_23521);
nand U24386 (N_24386,N_23660,N_22972);
or U24387 (N_24387,N_22387,N_23922);
xor U24388 (N_24388,N_23052,N_23090);
or U24389 (N_24389,N_22907,N_22626);
xnor U24390 (N_24390,N_22063,N_23619);
nand U24391 (N_24391,N_23258,N_23274);
or U24392 (N_24392,N_22453,N_22455);
and U24393 (N_24393,N_23175,N_22705);
xor U24394 (N_24394,N_22174,N_22866);
nand U24395 (N_24395,N_22685,N_23562);
and U24396 (N_24396,N_22640,N_23956);
or U24397 (N_24397,N_22502,N_23034);
nor U24398 (N_24398,N_23173,N_23904);
or U24399 (N_24399,N_22503,N_22736);
nor U24400 (N_24400,N_22533,N_22487);
xnor U24401 (N_24401,N_23116,N_23252);
or U24402 (N_24402,N_23314,N_22158);
nor U24403 (N_24403,N_22457,N_22873);
nand U24404 (N_24404,N_22504,N_23622);
or U24405 (N_24405,N_22929,N_23643);
and U24406 (N_24406,N_23566,N_22636);
nor U24407 (N_24407,N_23391,N_22665);
and U24408 (N_24408,N_23215,N_23010);
or U24409 (N_24409,N_23066,N_23408);
nor U24410 (N_24410,N_23507,N_23950);
nand U24411 (N_24411,N_23576,N_22312);
nor U24412 (N_24412,N_23552,N_22610);
nand U24413 (N_24413,N_23268,N_22590);
nand U24414 (N_24414,N_23987,N_23921);
or U24415 (N_24415,N_23186,N_23690);
nor U24416 (N_24416,N_23385,N_23494);
or U24417 (N_24417,N_22450,N_23147);
xor U24418 (N_24418,N_23463,N_22223);
and U24419 (N_24419,N_23795,N_23395);
nand U24420 (N_24420,N_22288,N_23394);
nand U24421 (N_24421,N_23647,N_23855);
nor U24422 (N_24422,N_23416,N_22700);
and U24423 (N_24423,N_22701,N_23966);
nor U24424 (N_24424,N_22425,N_23015);
or U24425 (N_24425,N_23351,N_23120);
or U24426 (N_24426,N_23502,N_23128);
nor U24427 (N_24427,N_22212,N_22236);
xnor U24428 (N_24428,N_22779,N_23254);
nor U24429 (N_24429,N_23565,N_23180);
nor U24430 (N_24430,N_23497,N_22421);
nand U24431 (N_24431,N_23805,N_22607);
xnor U24432 (N_24432,N_22819,N_22193);
and U24433 (N_24433,N_23719,N_22333);
xnor U24434 (N_24434,N_22432,N_22822);
xor U24435 (N_24435,N_22715,N_22559);
nand U24436 (N_24436,N_22256,N_23003);
and U24437 (N_24437,N_22541,N_22014);
and U24438 (N_24438,N_22407,N_23113);
nand U24439 (N_24439,N_22615,N_22845);
xor U24440 (N_24440,N_22998,N_22854);
nor U24441 (N_24441,N_23035,N_22252);
xor U24442 (N_24442,N_22598,N_23221);
or U24443 (N_24443,N_23560,N_22697);
or U24444 (N_24444,N_22728,N_23278);
xor U24445 (N_24445,N_23415,N_23661);
xnor U24446 (N_24446,N_23750,N_22364);
and U24447 (N_24447,N_23895,N_23763);
or U24448 (N_24448,N_22670,N_23550);
xor U24449 (N_24449,N_22920,N_23098);
nand U24450 (N_24450,N_22856,N_22752);
or U24451 (N_24451,N_23559,N_23070);
or U24452 (N_24452,N_23160,N_22126);
and U24453 (N_24453,N_22279,N_23602);
or U24454 (N_24454,N_22806,N_23499);
xor U24455 (N_24455,N_23700,N_23841);
xor U24456 (N_24456,N_23192,N_22732);
xor U24457 (N_24457,N_22257,N_22568);
xnor U24458 (N_24458,N_22680,N_22888);
and U24459 (N_24459,N_23018,N_22226);
or U24460 (N_24460,N_23217,N_23579);
xor U24461 (N_24461,N_22423,N_23325);
nor U24462 (N_24462,N_23645,N_23785);
and U24463 (N_24463,N_23155,N_22200);
or U24464 (N_24464,N_22862,N_22596);
or U24465 (N_24465,N_22213,N_22344);
xor U24466 (N_24466,N_23501,N_22910);
xnor U24467 (N_24467,N_22588,N_23253);
xor U24468 (N_24468,N_22995,N_22155);
and U24469 (N_24469,N_22273,N_23308);
and U24470 (N_24470,N_23001,N_23649);
nand U24471 (N_24471,N_23607,N_22617);
nor U24472 (N_24472,N_23097,N_23792);
nor U24473 (N_24473,N_22353,N_22173);
nor U24474 (N_24474,N_23349,N_23816);
xor U24475 (N_24475,N_23683,N_23095);
or U24476 (N_24476,N_22136,N_23856);
nor U24477 (N_24477,N_23547,N_23085);
and U24478 (N_24478,N_23442,N_22690);
nor U24479 (N_24479,N_23305,N_23183);
nand U24480 (N_24480,N_23817,N_22400);
and U24481 (N_24481,N_22641,N_23362);
and U24482 (N_24482,N_23774,N_23167);
nor U24483 (N_24483,N_23339,N_23967);
and U24484 (N_24484,N_22363,N_22621);
and U24485 (N_24485,N_22274,N_22831);
and U24486 (N_24486,N_23652,N_23912);
xnor U24487 (N_24487,N_22392,N_23427);
and U24488 (N_24488,N_22882,N_23492);
and U24489 (N_24489,N_22565,N_22880);
nor U24490 (N_24490,N_23868,N_23797);
nor U24491 (N_24491,N_22794,N_23909);
or U24492 (N_24492,N_22422,N_22486);
and U24493 (N_24493,N_22947,N_22753);
nor U24494 (N_24494,N_23236,N_22647);
xnor U24495 (N_24495,N_22034,N_22074);
xnor U24496 (N_24496,N_22220,N_22955);
or U24497 (N_24497,N_23345,N_22682);
or U24498 (N_24498,N_22985,N_23735);
or U24499 (N_24499,N_23292,N_23916);
xnor U24500 (N_24500,N_22976,N_22534);
nand U24501 (N_24501,N_22821,N_23905);
xor U24502 (N_24502,N_22092,N_23914);
nor U24503 (N_24503,N_22505,N_23449);
or U24504 (N_24504,N_22837,N_22805);
nand U24505 (N_24505,N_23383,N_22232);
and U24506 (N_24506,N_22106,N_22513);
nor U24507 (N_24507,N_22185,N_23425);
nor U24508 (N_24508,N_22060,N_23818);
and U24509 (N_24509,N_23558,N_22323);
xor U24510 (N_24510,N_23101,N_23761);
xnor U24511 (N_24511,N_22986,N_22494);
nand U24512 (N_24512,N_22409,N_22148);
nor U24513 (N_24513,N_22557,N_23359);
or U24514 (N_24514,N_22214,N_23572);
nor U24515 (N_24515,N_23482,N_22704);
nand U24516 (N_24516,N_22580,N_23114);
xor U24517 (N_24517,N_22620,N_22424);
or U24518 (N_24518,N_22954,N_22442);
and U24519 (N_24519,N_23083,N_22112);
nor U24520 (N_24520,N_22864,N_22766);
xor U24521 (N_24521,N_23138,N_22938);
nor U24522 (N_24522,N_23773,N_22927);
and U24523 (N_24523,N_22227,N_23629);
xor U24524 (N_24524,N_23668,N_22206);
or U24525 (N_24525,N_23246,N_23769);
and U24526 (N_24526,N_22653,N_23845);
and U24527 (N_24527,N_23612,N_22025);
nor U24528 (N_24528,N_22999,N_22654);
or U24529 (N_24529,N_22415,N_23224);
xor U24530 (N_24530,N_23886,N_23992);
nand U24531 (N_24531,N_22367,N_23462);
xor U24532 (N_24532,N_23369,N_23169);
nand U24533 (N_24533,N_22016,N_22096);
xnor U24534 (N_24534,N_22478,N_22525);
xor U24535 (N_24535,N_23951,N_22380);
xnor U24536 (N_24536,N_23681,N_22385);
nor U24537 (N_24537,N_23358,N_22884);
xnor U24538 (N_24538,N_22727,N_23199);
nor U24539 (N_24539,N_23086,N_23523);
nor U24540 (N_24540,N_22656,N_22787);
and U24541 (N_24541,N_22659,N_23024);
nor U24542 (N_24542,N_22359,N_23567);
or U24543 (N_24543,N_23187,N_22441);
xnor U24544 (N_24544,N_23738,N_22737);
and U24545 (N_24545,N_22140,N_23341);
and U24546 (N_24546,N_22842,N_23384);
xor U24547 (N_24547,N_23932,N_23166);
nor U24548 (N_24548,N_22052,N_22484);
nor U24549 (N_24549,N_22851,N_22003);
and U24550 (N_24550,N_22078,N_22566);
and U24551 (N_24551,N_23455,N_23232);
or U24552 (N_24552,N_22713,N_23317);
nor U24553 (N_24553,N_23088,N_22308);
nor U24554 (N_24554,N_23994,N_22517);
and U24555 (N_24555,N_23575,N_23225);
or U24556 (N_24556,N_22634,N_22354);
xnor U24557 (N_24557,N_22153,N_22942);
xnor U24558 (N_24558,N_23698,N_22436);
or U24559 (N_24559,N_22199,N_22246);
xnor U24560 (N_24560,N_22742,N_23365);
or U24561 (N_24561,N_22734,N_23403);
and U24562 (N_24562,N_22921,N_23304);
nand U24563 (N_24563,N_23048,N_22538);
nand U24564 (N_24564,N_23059,N_23728);
and U24565 (N_24565,N_23973,N_23471);
nor U24566 (N_24566,N_22382,N_23860);
and U24567 (N_24567,N_22838,N_23611);
and U24568 (N_24568,N_23872,N_23409);
or U24569 (N_24569,N_22839,N_23679);
and U24570 (N_24570,N_23638,N_23328);
or U24571 (N_24571,N_23273,N_23851);
nor U24572 (N_24572,N_22863,N_22564);
and U24573 (N_24573,N_23636,N_23758);
and U24574 (N_24574,N_22022,N_23046);
nand U24575 (N_24575,N_23154,N_23644);
or U24576 (N_24576,N_23181,N_23335);
xnor U24577 (N_24577,N_23828,N_23704);
nor U24578 (N_24578,N_23628,N_22238);
and U24579 (N_24579,N_23420,N_22378);
nor U24580 (N_24580,N_23515,N_23089);
nand U24581 (N_24581,N_22341,N_22555);
and U24582 (N_24582,N_22472,N_23870);
xnor U24583 (N_24583,N_23775,N_22244);
nor U24584 (N_24584,N_23633,N_23270);
or U24585 (N_24585,N_22340,N_22230);
or U24586 (N_24586,N_22240,N_22601);
nand U24587 (N_24587,N_23266,N_22357);
or U24588 (N_24588,N_22973,N_23726);
nand U24589 (N_24589,N_22219,N_23526);
nand U24590 (N_24590,N_23436,N_23557);
and U24591 (N_24591,N_23307,N_23708);
or U24592 (N_24592,N_22763,N_23989);
nand U24593 (N_24593,N_22522,N_23641);
xor U24594 (N_24594,N_23924,N_23038);
nor U24595 (N_24595,N_23812,N_23717);
nor U24596 (N_24596,N_23756,N_22129);
or U24597 (N_24597,N_22338,N_22518);
and U24598 (N_24598,N_23838,N_22983);
and U24599 (N_24599,N_22585,N_23810);
nor U24600 (N_24600,N_22536,N_23481);
nor U24601 (N_24601,N_22632,N_22926);
and U24602 (N_24602,N_22143,N_23354);
nand U24603 (N_24603,N_23282,N_22194);
or U24604 (N_24604,N_23620,N_22669);
nor U24605 (N_24605,N_22275,N_23616);
nor U24606 (N_24606,N_23546,N_23229);
or U24607 (N_24607,N_22836,N_23760);
or U24608 (N_24608,N_23275,N_22754);
nand U24609 (N_24609,N_23655,N_22622);
and U24610 (N_24610,N_23200,N_22157);
and U24611 (N_24611,N_22004,N_23170);
nand U24612 (N_24612,N_22800,N_23907);
nor U24613 (N_24613,N_23280,N_23713);
nand U24614 (N_24614,N_22383,N_23517);
nand U24615 (N_24615,N_22449,N_23864);
nand U24616 (N_24616,N_22605,N_23574);
and U24617 (N_24617,N_22792,N_23222);
or U24618 (N_24618,N_23782,N_22491);
xor U24619 (N_24619,N_22346,N_23428);
xnor U24620 (N_24620,N_22061,N_22508);
or U24621 (N_24621,N_22245,N_23757);
nand U24622 (N_24622,N_23080,N_23642);
and U24623 (N_24623,N_23297,N_22482);
or U24624 (N_24624,N_22259,N_22048);
and U24625 (N_24625,N_22026,N_23289);
nand U24626 (N_24626,N_23854,N_22141);
nor U24627 (N_24627,N_23239,N_23827);
xnor U24628 (N_24628,N_23110,N_23423);
nand U24629 (N_24629,N_22526,N_22729);
or U24630 (N_24630,N_22961,N_23784);
or U24631 (N_24631,N_23988,N_23839);
and U24632 (N_24632,N_22748,N_22746);
or U24633 (N_24633,N_22909,N_22574);
or U24634 (N_24634,N_23826,N_22563);
nor U24635 (N_24635,N_23964,N_23993);
or U24636 (N_24636,N_22931,N_22297);
xnor U24637 (N_24637,N_22606,N_23890);
nor U24638 (N_24638,N_23771,N_23585);
nand U24639 (N_24639,N_23520,N_23716);
and U24640 (N_24640,N_22328,N_22164);
and U24641 (N_24641,N_22027,N_23220);
nand U24642 (N_24642,N_22133,N_23281);
nor U24643 (N_24643,N_22066,N_23830);
xor U24644 (N_24644,N_22460,N_23974);
xnor U24645 (N_24645,N_22100,N_23115);
nand U24646 (N_24646,N_22115,N_23543);
nor U24647 (N_24647,N_22511,N_23271);
nor U24648 (N_24648,N_23487,N_22510);
and U24649 (N_24649,N_22356,N_22760);
nor U24650 (N_24650,N_22591,N_23039);
or U24651 (N_24651,N_22036,N_23008);
and U24652 (N_24652,N_22277,N_22135);
xnor U24653 (N_24653,N_23519,N_23396);
and U24654 (N_24654,N_23865,N_23148);
xor U24655 (N_24655,N_23729,N_22162);
or U24656 (N_24656,N_23406,N_22499);
and U24657 (N_24657,N_23227,N_22545);
xnor U24658 (N_24658,N_23882,N_23250);
or U24659 (N_24659,N_23939,N_22743);
nand U24660 (N_24660,N_23587,N_23722);
and U24661 (N_24661,N_23709,N_23584);
and U24662 (N_24662,N_23245,N_22720);
nand U24663 (N_24663,N_22122,N_23631);
or U24664 (N_24664,N_23687,N_22043);
nor U24665 (N_24665,N_22083,N_23295);
xor U24666 (N_24666,N_22009,N_22916);
xor U24667 (N_24667,N_23032,N_23829);
or U24668 (N_24668,N_22813,N_23068);
or U24669 (N_24669,N_22918,N_23002);
nor U24670 (N_24670,N_22828,N_23959);
nand U24671 (N_24671,N_22225,N_23137);
xnor U24672 (N_24672,N_23240,N_23178);
xor U24673 (N_24673,N_22071,N_23615);
nor U24674 (N_24674,N_23979,N_23528);
xor U24675 (N_24675,N_22325,N_22577);
xnor U24676 (N_24676,N_23299,N_22492);
nand U24677 (N_24677,N_22452,N_23152);
xnor U24678 (N_24678,N_22782,N_23480);
nand U24679 (N_24679,N_23853,N_22221);
nand U24680 (N_24680,N_23298,N_22572);
nor U24681 (N_24681,N_22612,N_22156);
nand U24682 (N_24682,N_22138,N_22575);
and U24683 (N_24683,N_22216,N_23352);
xnor U24684 (N_24684,N_23720,N_22738);
and U24685 (N_24685,N_23626,N_22686);
xor U24686 (N_24686,N_22974,N_23334);
and U24687 (N_24687,N_22404,N_23259);
or U24688 (N_24688,N_23913,N_23779);
and U24689 (N_24689,N_22461,N_23495);
and U24690 (N_24690,N_22250,N_23211);
nor U24691 (N_24691,N_23733,N_23142);
nand U24692 (N_24692,N_23378,N_23255);
or U24693 (N_24693,N_23475,N_23131);
nor U24694 (N_24694,N_22891,N_23800);
nor U24695 (N_24695,N_23923,N_22406);
and U24696 (N_24696,N_22128,N_22967);
and U24697 (N_24697,N_23191,N_22645);
xor U24698 (N_24698,N_23977,N_22149);
nand U24699 (N_24699,N_22660,N_22980);
xnor U24700 (N_24700,N_22445,N_23331);
and U24701 (N_24701,N_23806,N_23878);
and U24702 (N_24702,N_22770,N_23091);
and U24703 (N_24703,N_23752,N_22578);
nor U24704 (N_24704,N_23711,N_22964);
xor U24705 (N_24705,N_22019,N_23715);
xnor U24706 (N_24706,N_23056,N_23407);
xor U24707 (N_24707,N_23121,N_23666);
xor U24708 (N_24708,N_23926,N_22305);
nor U24709 (N_24709,N_23770,N_22365);
and U24710 (N_24710,N_23721,N_22319);
or U24711 (N_24711,N_23382,N_23061);
nand U24712 (N_24712,N_22207,N_22299);
xnor U24713 (N_24713,N_23963,N_23593);
nand U24714 (N_24714,N_22583,N_22996);
nor U24715 (N_24715,N_22677,N_22150);
or U24716 (N_24716,N_22265,N_22085);
or U24717 (N_24717,N_22879,N_23075);
xnor U24718 (N_24718,N_22012,N_22335);
xnor U24719 (N_24719,N_22638,N_22489);
xor U24720 (N_24720,N_23027,N_22007);
nand U24721 (N_24721,N_23448,N_22470);
or U24722 (N_24722,N_23209,N_22446);
nand U24723 (N_24723,N_23466,N_22688);
and U24724 (N_24724,N_22454,N_23393);
and U24725 (N_24725,N_22290,N_22233);
or U24726 (N_24726,N_23815,N_22519);
and U24727 (N_24727,N_22722,N_23588);
or U24728 (N_24728,N_22778,N_23893);
or U24729 (N_24729,N_23751,N_23022);
xnor U24730 (N_24730,N_22349,N_22633);
xor U24731 (N_24731,N_23597,N_22573);
or U24732 (N_24732,N_22630,N_22272);
or U24733 (N_24733,N_23496,N_22413);
xor U24734 (N_24734,N_23903,N_23126);
xnor U24735 (N_24735,N_22745,N_22692);
nand U24736 (N_24736,N_23318,N_22584);
and U24737 (N_24737,N_22287,N_22255);
xor U24738 (N_24738,N_23876,N_23695);
nand U24739 (N_24739,N_22739,N_23431);
xor U24740 (N_24740,N_23421,N_23033);
and U24741 (N_24741,N_22592,N_22712);
and U24742 (N_24742,N_23767,N_22310);
xnor U24743 (N_24743,N_23505,N_23012);
and U24744 (N_24744,N_22301,N_23081);
xnor U24745 (N_24745,N_22825,N_23060);
nand U24746 (N_24746,N_23076,N_23899);
or U24747 (N_24747,N_23483,N_22217);
nor U24748 (N_24748,N_23919,N_23850);
xnor U24749 (N_24749,N_22637,N_22599);
and U24750 (N_24750,N_22848,N_22762);
and U24751 (N_24751,N_22696,N_23077);
and U24752 (N_24752,N_22547,N_23342);
xor U24753 (N_24753,N_23202,N_22374);
nand U24754 (N_24754,N_23410,N_23984);
and U24755 (N_24755,N_23372,N_22051);
xor U24756 (N_24756,N_23165,N_22389);
or U24757 (N_24757,N_23135,N_22979);
and U24758 (N_24758,N_23960,N_22841);
xnor U24759 (N_24759,N_23161,N_23050);
nand U24760 (N_24760,N_23016,N_22874);
nor U24761 (N_24761,N_22550,N_22928);
nor U24762 (N_24762,N_23578,N_23688);
or U24763 (N_24763,N_22694,N_22730);
or U24764 (N_24764,N_22480,N_23930);
nor U24765 (N_24765,N_22035,N_23614);
and U24766 (N_24766,N_23820,N_22111);
xnor U24767 (N_24767,N_23219,N_22322);
or U24768 (N_24768,N_23592,N_22263);
nand U24769 (N_24769,N_23288,N_22081);
nor U24770 (N_24770,N_22447,N_22419);
nand U24771 (N_24771,N_23400,N_22037);
or U24772 (N_24772,N_22405,N_22253);
nor U24773 (N_24773,N_22671,N_22527);
nor U24774 (N_24774,N_22840,N_22130);
and U24775 (N_24775,N_23319,N_23618);
nor U24776 (N_24776,N_23149,N_23078);
nand U24777 (N_24777,N_23042,N_22139);
nor U24778 (N_24778,N_23231,N_22516);
xor U24779 (N_24779,N_22894,N_22970);
nand U24780 (N_24780,N_22152,N_23836);
nor U24781 (N_24781,N_22109,N_23746);
nand U24782 (N_24782,N_22114,N_22969);
nand U24783 (N_24783,N_22254,N_23087);
nor U24784 (N_24784,N_22282,N_22399);
nand U24785 (N_24785,N_23889,N_22296);
and U24786 (N_24786,N_23411,N_22249);
nor U24787 (N_24787,N_22070,N_22781);
xnor U24788 (N_24788,N_23648,N_22146);
nand U24789 (N_24789,N_23925,N_23787);
xor U24790 (N_24790,N_22797,N_23303);
xnor U24791 (N_24791,N_22721,N_22900);
xor U24792 (N_24792,N_23877,N_23710);
nand U24793 (N_24793,N_23477,N_22698);
and U24794 (N_24794,N_23125,N_22500);
and U24795 (N_24795,N_23500,N_23518);
or U24796 (N_24796,N_23401,N_23952);
and U24797 (N_24797,N_23030,N_22195);
nand U24798 (N_24798,N_23937,N_22295);
nor U24799 (N_24799,N_23031,N_23707);
nor U24800 (N_24800,N_23333,N_22285);
nand U24801 (N_24801,N_23426,N_23676);
nand U24802 (N_24802,N_22269,N_23037);
and U24803 (N_24803,N_22393,N_22703);
nand U24804 (N_24804,N_22396,N_23745);
or U24805 (N_24805,N_23417,N_22177);
or U24806 (N_24806,N_23586,N_22375);
and U24807 (N_24807,N_23606,N_22011);
xor U24808 (N_24808,N_23162,N_23324);
xor U24809 (N_24809,N_23749,N_22172);
nor U24810 (N_24810,N_22917,N_22309);
nor U24811 (N_24811,N_23063,N_23858);
nor U24812 (N_24812,N_22371,N_23881);
nand U24813 (N_24813,N_23788,N_23311);
nor U24814 (N_24814,N_23398,N_23386);
or U24815 (N_24815,N_22479,N_23310);
or U24816 (N_24816,N_22329,N_23672);
or U24817 (N_24817,N_22391,N_22101);
or U24818 (N_24818,N_22644,N_23223);
nand U24819 (N_24819,N_22706,N_23945);
nand U24820 (N_24820,N_22203,N_23498);
or U24821 (N_24821,N_22933,N_23437);
and U24822 (N_24822,N_22908,N_22465);
xnor U24823 (N_24823,N_22939,N_23065);
nand U24824 (N_24824,N_23651,N_22593);
xor U24825 (N_24825,N_22471,N_23736);
nor U24826 (N_24826,N_23551,N_23486);
nor U24827 (N_24827,N_23397,N_22540);
or U24828 (N_24828,N_23680,N_23894);
or U24829 (N_24829,N_23457,N_22978);
or U24830 (N_24830,N_23450,N_22132);
xnor U24831 (N_24831,N_23092,N_22543);
or U24832 (N_24832,N_22362,N_22679);
or U24833 (N_24833,N_22318,N_22267);
xnor U24834 (N_24834,N_22293,N_22587);
and U24835 (N_24835,N_23522,N_23047);
or U24836 (N_24836,N_22268,N_23542);
or U24837 (N_24837,N_23474,N_23294);
xnor U24838 (N_24838,N_23640,N_23188);
or U24839 (N_24839,N_23476,N_23207);
nand U24840 (N_24840,N_22990,N_22952);
and U24841 (N_24841,N_23686,N_23290);
and U24842 (N_24842,N_23277,N_22401);
and U24843 (N_24843,N_22127,N_23469);
nand U24844 (N_24844,N_23493,N_22614);
xor U24845 (N_24845,N_23072,N_23986);
or U24846 (N_24846,N_22058,N_23874);
xor U24847 (N_24847,N_23456,N_22953);
xor U24848 (N_24848,N_22788,N_22373);
xor U24849 (N_24849,N_22808,N_23879);
and U24850 (N_24850,N_23251,N_22248);
and U24851 (N_24851,N_23766,N_23625);
nor U24852 (N_24852,N_23691,N_23657);
and U24853 (N_24853,N_22946,N_22000);
xnor U24854 (N_24854,N_23444,N_23678);
or U24855 (N_24855,N_23459,N_22294);
nor U24856 (N_24856,N_22595,N_22861);
nor U24857 (N_24857,N_22652,N_23740);
or U24858 (N_24858,N_22529,N_23430);
nor U24859 (N_24859,N_23151,N_22497);
xnor U24860 (N_24860,N_22010,N_23389);
nor U24861 (N_24861,N_23857,N_23453);
nand U24862 (N_24862,N_23589,N_23601);
nor U24863 (N_24863,N_22710,N_23825);
xnor U24864 (N_24864,N_22528,N_23995);
nand U24865 (N_24865,N_22793,N_22403);
and U24866 (N_24866,N_23419,N_23118);
or U24867 (N_24867,N_22695,N_22343);
or U24868 (N_24868,N_23177,N_22691);
nor U24869 (N_24869,N_22490,N_22451);
nand U24870 (N_24870,N_22892,N_22544);
and U24871 (N_24871,N_22570,N_23214);
xnor U24872 (N_24872,N_22776,N_22080);
and U24873 (N_24873,N_23323,N_22922);
nand U24874 (N_24874,N_22372,N_22169);
xor U24875 (N_24875,N_22496,N_22108);
nor U24876 (N_24876,N_23941,N_22958);
or U24877 (N_24877,N_22860,N_22711);
or U24878 (N_24878,N_22298,N_22849);
nand U24879 (N_24879,N_22531,N_23249);
xnor U24880 (N_24880,N_22749,N_23158);
nor U24881 (N_24881,N_23866,N_22957);
nand U24882 (N_24882,N_22832,N_22188);
nand U24883 (N_24883,N_23665,N_23808);
and U24884 (N_24884,N_23539,N_23883);
nor U24885 (N_24885,N_23106,N_23422);
or U24886 (N_24886,N_22824,N_22835);
nand U24887 (N_24887,N_23570,N_23604);
or U24888 (N_24888,N_23510,N_23891);
or U24889 (N_24889,N_22488,N_22283);
nand U24890 (N_24890,N_23762,N_23327);
nand U24891 (N_24891,N_23603,N_22887);
and U24892 (N_24892,N_22417,N_22672);
nor U24893 (N_24893,N_23204,N_22201);
and U24894 (N_24894,N_22182,N_23949);
nor U24895 (N_24895,N_23654,N_22402);
and U24896 (N_24896,N_22118,N_22326);
xnor U24897 (N_24897,N_22850,N_22271);
and U24898 (N_24898,N_22925,N_23832);
nand U24899 (N_24899,N_22795,N_22438);
or U24900 (N_24900,N_22228,N_23623);
and U24901 (N_24901,N_22002,N_22355);
nor U24902 (N_24902,N_22791,N_23381);
nor U24903 (N_24903,N_22868,N_22284);
nor U24904 (N_24904,N_22218,N_23910);
xor U24905 (N_24905,N_22817,N_22867);
and U24906 (N_24906,N_23071,N_22196);
or U24907 (N_24907,N_23100,N_22594);
nor U24908 (N_24908,N_23549,N_23062);
or U24909 (N_24909,N_23150,N_23934);
xnor U24910 (N_24910,N_22327,N_22943);
or U24911 (N_24911,N_22350,N_22501);
and U24912 (N_24912,N_22079,N_23536);
xnor U24913 (N_24913,N_23849,N_22444);
or U24914 (N_24914,N_23699,N_22767);
xnor U24915 (N_24915,N_23021,N_22087);
xnor U24916 (N_24916,N_22180,N_23111);
nor U24917 (N_24917,N_23673,N_23041);
nand U24918 (N_24918,N_22537,N_23133);
nor U24919 (N_24919,N_22558,N_22714);
xnor U24920 (N_24920,N_23244,N_22099);
nand U24921 (N_24921,N_23548,N_23488);
xor U24922 (N_24922,N_23508,N_22912);
nor U24923 (N_24923,N_23233,N_22521);
and U24924 (N_24924,N_23887,N_22001);
or U24925 (N_24925,N_22803,N_23525);
xnor U24926 (N_24926,N_22475,N_23000);
nand U24927 (N_24927,N_23272,N_23040);
nor U24928 (N_24928,N_22430,N_23884);
nor U24929 (N_24929,N_23833,N_22222);
xnor U24930 (N_24930,N_22197,N_22678);
xnor U24931 (N_24931,N_23145,N_23998);
nor U24932 (N_24932,N_23336,N_22303);
and U24933 (N_24933,N_23484,N_23613);
nand U24934 (N_24934,N_23438,N_23669);
xnor U24935 (N_24935,N_22717,N_22360);
nor U24936 (N_24936,N_22031,N_22576);
nor U24937 (N_24937,N_23464,N_22427);
or U24938 (N_24938,N_23940,N_23193);
or U24939 (N_24939,N_22687,N_22466);
and U24940 (N_24940,N_23079,N_22015);
xor U24941 (N_24941,N_23725,N_22028);
xnor U24942 (N_24942,N_23696,N_23196);
nor U24943 (N_24943,N_23326,N_22289);
and U24944 (N_24944,N_22097,N_23867);
nor U24945 (N_24945,N_23799,N_23689);
or U24946 (N_24946,N_23896,N_22258);
xor U24947 (N_24947,N_23051,N_22642);
nand U24948 (N_24948,N_23667,N_22147);
or U24949 (N_24949,N_22352,N_23206);
xnor U24950 (N_24950,N_22542,N_22181);
and U24951 (N_24951,N_23859,N_22086);
nand U24952 (N_24952,N_23287,N_23470);
or U24953 (N_24953,N_23379,N_23511);
and U24954 (N_24954,N_22125,N_23846);
nand U24955 (N_24955,N_23933,N_23248);
and U24956 (N_24956,N_22366,N_22331);
nor U24957 (N_24957,N_22073,N_22270);
xnor U24958 (N_24958,N_22493,N_22304);
and U24959 (N_24959,N_23885,N_22597);
nor U24960 (N_24960,N_22059,N_22649);
nand U24961 (N_24961,N_23701,N_22589);
and U24962 (N_24962,N_22324,N_23007);
nor U24963 (N_24963,N_22951,N_23478);
xnor U24964 (N_24964,N_22376,N_22629);
nor U24965 (N_24965,N_22899,N_22535);
or U24966 (N_24966,N_22937,N_22675);
or U24967 (N_24967,N_23969,N_23970);
xor U24968 (N_24968,N_23712,N_23813);
nor U24969 (N_24969,N_23285,N_23049);
or U24970 (N_24970,N_23309,N_22581);
or U24971 (N_24971,N_22435,N_23605);
xor U24972 (N_24972,N_23796,N_23194);
nand U24973 (N_24973,N_23599,N_22992);
or U24974 (N_24974,N_23639,N_22786);
and U24975 (N_24975,N_22089,N_22361);
or U24976 (N_24976,N_23132,N_23414);
nor U24977 (N_24977,N_23020,N_23674);
nand U24978 (N_24978,N_22463,N_22042);
xnor U24979 (N_24979,N_23009,N_22847);
or U24980 (N_24980,N_22377,N_23999);
and U24981 (N_24981,N_23541,N_22693);
nor U24982 (N_24982,N_22771,N_22243);
nand U24983 (N_24983,N_23996,N_22914);
xnor U24984 (N_24984,N_23107,N_22124);
xnor U24985 (N_24985,N_23902,N_22107);
nand U24986 (N_24986,N_22875,N_22556);
xnor U24987 (N_24987,N_23432,N_23663);
or U24988 (N_24988,N_22163,N_22657);
xor U24989 (N_24989,N_22234,N_22546);
nor U24990 (N_24990,N_23380,N_22812);
nand U24991 (N_24991,N_22056,N_22434);
and U24992 (N_24992,N_23556,N_22184);
nand U24993 (N_24993,N_23306,N_23971);
or U24994 (N_24994,N_22439,N_23659);
nand U24995 (N_24995,N_22072,N_22208);
nand U24996 (N_24996,N_22881,N_22663);
nor U24997 (N_24997,N_22278,N_22247);
and U24998 (N_24998,N_23329,N_23534);
and U24999 (N_24999,N_22790,N_22661);
nand U25000 (N_25000,N_22910,N_22309);
or U25001 (N_25001,N_22967,N_22030);
nor U25002 (N_25002,N_22444,N_23612);
or U25003 (N_25003,N_22190,N_22841);
and U25004 (N_25004,N_22650,N_22765);
nand U25005 (N_25005,N_23708,N_22566);
nand U25006 (N_25006,N_23396,N_22135);
and U25007 (N_25007,N_22038,N_23627);
nand U25008 (N_25008,N_23349,N_22297);
xor U25009 (N_25009,N_22556,N_22424);
or U25010 (N_25010,N_22300,N_22856);
nand U25011 (N_25011,N_23209,N_22447);
xnor U25012 (N_25012,N_23835,N_22532);
and U25013 (N_25013,N_22845,N_23270);
or U25014 (N_25014,N_22850,N_23392);
and U25015 (N_25015,N_22026,N_22293);
or U25016 (N_25016,N_23282,N_23001);
nor U25017 (N_25017,N_22700,N_22922);
nand U25018 (N_25018,N_22152,N_22224);
and U25019 (N_25019,N_22480,N_23718);
nor U25020 (N_25020,N_23940,N_23792);
xnor U25021 (N_25021,N_22552,N_23654);
and U25022 (N_25022,N_23543,N_22122);
or U25023 (N_25023,N_22865,N_22941);
xor U25024 (N_25024,N_23012,N_22258);
xnor U25025 (N_25025,N_22152,N_22426);
and U25026 (N_25026,N_22588,N_23143);
xnor U25027 (N_25027,N_22655,N_23136);
nor U25028 (N_25028,N_22437,N_23689);
nor U25029 (N_25029,N_22507,N_23145);
or U25030 (N_25030,N_22142,N_23236);
or U25031 (N_25031,N_22406,N_23408);
nor U25032 (N_25032,N_22298,N_23766);
xnor U25033 (N_25033,N_22924,N_22696);
nand U25034 (N_25034,N_22602,N_23779);
and U25035 (N_25035,N_22386,N_23810);
and U25036 (N_25036,N_22780,N_22679);
nor U25037 (N_25037,N_23956,N_23132);
nand U25038 (N_25038,N_22433,N_23988);
nor U25039 (N_25039,N_23968,N_22951);
nor U25040 (N_25040,N_23494,N_23540);
nand U25041 (N_25041,N_22642,N_22283);
nand U25042 (N_25042,N_23433,N_22465);
nor U25043 (N_25043,N_22646,N_22778);
and U25044 (N_25044,N_23013,N_22952);
nand U25045 (N_25045,N_22006,N_22081);
or U25046 (N_25046,N_22330,N_22141);
or U25047 (N_25047,N_23623,N_23936);
xnor U25048 (N_25048,N_23753,N_22610);
nand U25049 (N_25049,N_22299,N_23232);
xor U25050 (N_25050,N_23584,N_22248);
or U25051 (N_25051,N_22668,N_23376);
xor U25052 (N_25052,N_23516,N_23642);
xnor U25053 (N_25053,N_23258,N_22642);
nand U25054 (N_25054,N_22266,N_23830);
nand U25055 (N_25055,N_22183,N_22120);
or U25056 (N_25056,N_22191,N_23780);
and U25057 (N_25057,N_22210,N_22758);
xnor U25058 (N_25058,N_23784,N_22499);
xnor U25059 (N_25059,N_22787,N_22413);
or U25060 (N_25060,N_22070,N_23584);
nor U25061 (N_25061,N_23376,N_23503);
nand U25062 (N_25062,N_23337,N_23260);
nor U25063 (N_25063,N_23224,N_22791);
and U25064 (N_25064,N_23166,N_23752);
nor U25065 (N_25065,N_23780,N_22207);
xnor U25066 (N_25066,N_23744,N_22530);
or U25067 (N_25067,N_22197,N_23096);
nand U25068 (N_25068,N_22476,N_23322);
nand U25069 (N_25069,N_23852,N_22839);
nand U25070 (N_25070,N_22601,N_22763);
and U25071 (N_25071,N_22057,N_22606);
xnor U25072 (N_25072,N_22811,N_22032);
and U25073 (N_25073,N_22918,N_23873);
xnor U25074 (N_25074,N_23237,N_23936);
nor U25075 (N_25075,N_23051,N_23515);
nor U25076 (N_25076,N_22368,N_22256);
nor U25077 (N_25077,N_22127,N_23606);
nand U25078 (N_25078,N_22059,N_22013);
and U25079 (N_25079,N_22713,N_22414);
and U25080 (N_25080,N_22630,N_23923);
and U25081 (N_25081,N_22868,N_22573);
nand U25082 (N_25082,N_23173,N_22945);
nor U25083 (N_25083,N_22189,N_23802);
nor U25084 (N_25084,N_23978,N_23001);
nand U25085 (N_25085,N_22041,N_22126);
and U25086 (N_25086,N_22540,N_22853);
or U25087 (N_25087,N_23657,N_23441);
or U25088 (N_25088,N_22990,N_22911);
or U25089 (N_25089,N_23213,N_22129);
nand U25090 (N_25090,N_22783,N_22693);
nor U25091 (N_25091,N_22508,N_22932);
and U25092 (N_25092,N_22102,N_23459);
xor U25093 (N_25093,N_23326,N_23584);
nor U25094 (N_25094,N_22804,N_22244);
xor U25095 (N_25095,N_22977,N_23879);
nor U25096 (N_25096,N_22469,N_23267);
nand U25097 (N_25097,N_22338,N_22867);
nor U25098 (N_25098,N_22468,N_22492);
and U25099 (N_25099,N_23894,N_22488);
nor U25100 (N_25100,N_22977,N_22628);
nand U25101 (N_25101,N_23689,N_22375);
or U25102 (N_25102,N_23064,N_22775);
and U25103 (N_25103,N_22768,N_22414);
nor U25104 (N_25104,N_23601,N_23319);
or U25105 (N_25105,N_22819,N_22033);
and U25106 (N_25106,N_22320,N_23912);
xnor U25107 (N_25107,N_22203,N_22660);
nor U25108 (N_25108,N_22810,N_22372);
or U25109 (N_25109,N_22925,N_23119);
or U25110 (N_25110,N_22087,N_23515);
nor U25111 (N_25111,N_22279,N_22072);
nor U25112 (N_25112,N_22209,N_22751);
xnor U25113 (N_25113,N_22576,N_22450);
or U25114 (N_25114,N_22784,N_22264);
xor U25115 (N_25115,N_22446,N_23956);
or U25116 (N_25116,N_23851,N_23617);
xor U25117 (N_25117,N_22870,N_22979);
xor U25118 (N_25118,N_22510,N_23493);
nor U25119 (N_25119,N_23657,N_22296);
xnor U25120 (N_25120,N_22226,N_22506);
nand U25121 (N_25121,N_23185,N_22205);
nand U25122 (N_25122,N_23495,N_22797);
and U25123 (N_25123,N_23547,N_22070);
xnor U25124 (N_25124,N_23195,N_22365);
or U25125 (N_25125,N_22062,N_23024);
xor U25126 (N_25126,N_22873,N_22651);
nor U25127 (N_25127,N_23673,N_22402);
or U25128 (N_25128,N_22735,N_22359);
nand U25129 (N_25129,N_22210,N_23870);
and U25130 (N_25130,N_23118,N_22450);
or U25131 (N_25131,N_23766,N_23878);
xor U25132 (N_25132,N_22586,N_22013);
and U25133 (N_25133,N_22417,N_23063);
or U25134 (N_25134,N_23525,N_22047);
nand U25135 (N_25135,N_22551,N_23929);
and U25136 (N_25136,N_23805,N_23824);
or U25137 (N_25137,N_22491,N_22152);
nor U25138 (N_25138,N_22032,N_23132);
nand U25139 (N_25139,N_22962,N_22430);
nor U25140 (N_25140,N_23621,N_22579);
nor U25141 (N_25141,N_23637,N_22019);
and U25142 (N_25142,N_22985,N_22047);
or U25143 (N_25143,N_22859,N_22304);
nor U25144 (N_25144,N_22353,N_22748);
or U25145 (N_25145,N_22920,N_23570);
nor U25146 (N_25146,N_22747,N_22613);
nor U25147 (N_25147,N_22646,N_23459);
nand U25148 (N_25148,N_23937,N_22570);
xnor U25149 (N_25149,N_23101,N_23371);
or U25150 (N_25150,N_22744,N_22767);
and U25151 (N_25151,N_23107,N_23754);
nand U25152 (N_25152,N_22223,N_22014);
nand U25153 (N_25153,N_22066,N_22152);
nand U25154 (N_25154,N_23106,N_22243);
and U25155 (N_25155,N_23742,N_23089);
nor U25156 (N_25156,N_23674,N_22366);
or U25157 (N_25157,N_22809,N_22207);
or U25158 (N_25158,N_22030,N_22741);
nor U25159 (N_25159,N_22173,N_22150);
nand U25160 (N_25160,N_23101,N_22388);
or U25161 (N_25161,N_23595,N_22393);
nor U25162 (N_25162,N_22995,N_22687);
xnor U25163 (N_25163,N_22019,N_23278);
and U25164 (N_25164,N_22364,N_23223);
and U25165 (N_25165,N_23022,N_22044);
nand U25166 (N_25166,N_23243,N_22137);
or U25167 (N_25167,N_23961,N_23877);
and U25168 (N_25168,N_22708,N_22276);
xnor U25169 (N_25169,N_22488,N_22049);
or U25170 (N_25170,N_22997,N_23995);
and U25171 (N_25171,N_22484,N_23923);
nand U25172 (N_25172,N_23677,N_22402);
and U25173 (N_25173,N_22870,N_22690);
or U25174 (N_25174,N_22506,N_22663);
nand U25175 (N_25175,N_23555,N_22136);
or U25176 (N_25176,N_23460,N_22070);
xnor U25177 (N_25177,N_23265,N_22173);
nand U25178 (N_25178,N_22292,N_23504);
nor U25179 (N_25179,N_22626,N_23376);
or U25180 (N_25180,N_23544,N_22470);
or U25181 (N_25181,N_23405,N_23850);
and U25182 (N_25182,N_23999,N_23072);
and U25183 (N_25183,N_22839,N_22763);
nand U25184 (N_25184,N_22322,N_23269);
xor U25185 (N_25185,N_23367,N_22443);
or U25186 (N_25186,N_22744,N_22958);
xor U25187 (N_25187,N_22162,N_23519);
or U25188 (N_25188,N_22711,N_22843);
nor U25189 (N_25189,N_23330,N_22398);
nand U25190 (N_25190,N_22421,N_23073);
and U25191 (N_25191,N_23937,N_23179);
xor U25192 (N_25192,N_23288,N_23896);
and U25193 (N_25193,N_23024,N_23466);
nor U25194 (N_25194,N_22867,N_23008);
or U25195 (N_25195,N_22334,N_23474);
nand U25196 (N_25196,N_22977,N_22222);
xnor U25197 (N_25197,N_23192,N_23545);
and U25198 (N_25198,N_23300,N_22923);
or U25199 (N_25199,N_23796,N_23958);
and U25200 (N_25200,N_22607,N_23182);
nand U25201 (N_25201,N_23020,N_23043);
xnor U25202 (N_25202,N_23933,N_22220);
and U25203 (N_25203,N_23201,N_22425);
and U25204 (N_25204,N_23946,N_22694);
nor U25205 (N_25205,N_23172,N_23996);
xnor U25206 (N_25206,N_22868,N_22992);
xor U25207 (N_25207,N_22962,N_22076);
nand U25208 (N_25208,N_23590,N_23833);
xor U25209 (N_25209,N_22334,N_22879);
and U25210 (N_25210,N_22480,N_22096);
nand U25211 (N_25211,N_22459,N_23455);
and U25212 (N_25212,N_23293,N_23200);
nor U25213 (N_25213,N_22477,N_23694);
or U25214 (N_25214,N_23690,N_22818);
or U25215 (N_25215,N_22022,N_22285);
or U25216 (N_25216,N_23507,N_22256);
nor U25217 (N_25217,N_22721,N_23905);
or U25218 (N_25218,N_23955,N_22975);
and U25219 (N_25219,N_22578,N_22829);
xnor U25220 (N_25220,N_22099,N_23936);
and U25221 (N_25221,N_23488,N_23381);
and U25222 (N_25222,N_22229,N_23358);
xnor U25223 (N_25223,N_22119,N_23044);
xnor U25224 (N_25224,N_22389,N_23532);
or U25225 (N_25225,N_22566,N_23547);
and U25226 (N_25226,N_23173,N_22393);
xor U25227 (N_25227,N_22064,N_23892);
and U25228 (N_25228,N_22926,N_23809);
nor U25229 (N_25229,N_22701,N_23707);
xor U25230 (N_25230,N_23418,N_23709);
nor U25231 (N_25231,N_23686,N_23217);
xnor U25232 (N_25232,N_23058,N_22175);
nand U25233 (N_25233,N_23134,N_22952);
and U25234 (N_25234,N_23811,N_23034);
nor U25235 (N_25235,N_23769,N_22846);
and U25236 (N_25236,N_23562,N_23144);
nand U25237 (N_25237,N_22683,N_22551);
or U25238 (N_25238,N_22916,N_23747);
xnor U25239 (N_25239,N_22962,N_23525);
nand U25240 (N_25240,N_23750,N_23379);
nor U25241 (N_25241,N_22004,N_23671);
xnor U25242 (N_25242,N_22056,N_23348);
or U25243 (N_25243,N_23690,N_22195);
xnor U25244 (N_25244,N_22720,N_23874);
nand U25245 (N_25245,N_22796,N_23630);
nand U25246 (N_25246,N_22407,N_23553);
xnor U25247 (N_25247,N_23816,N_23231);
nor U25248 (N_25248,N_23212,N_23328);
nor U25249 (N_25249,N_22049,N_23785);
xor U25250 (N_25250,N_23691,N_22522);
nand U25251 (N_25251,N_23133,N_23325);
xor U25252 (N_25252,N_23479,N_23298);
xnor U25253 (N_25253,N_23007,N_23994);
and U25254 (N_25254,N_22692,N_23050);
nor U25255 (N_25255,N_23817,N_23783);
nor U25256 (N_25256,N_23468,N_23633);
or U25257 (N_25257,N_22415,N_22895);
or U25258 (N_25258,N_23860,N_22038);
or U25259 (N_25259,N_22604,N_23490);
or U25260 (N_25260,N_22590,N_22770);
and U25261 (N_25261,N_23854,N_23301);
or U25262 (N_25262,N_22965,N_23568);
nand U25263 (N_25263,N_23504,N_22738);
nor U25264 (N_25264,N_22369,N_23320);
nor U25265 (N_25265,N_23656,N_22784);
or U25266 (N_25266,N_22643,N_22792);
nand U25267 (N_25267,N_22598,N_23829);
nand U25268 (N_25268,N_22914,N_23292);
xor U25269 (N_25269,N_23623,N_22380);
or U25270 (N_25270,N_22308,N_23385);
xnor U25271 (N_25271,N_23124,N_23471);
or U25272 (N_25272,N_22148,N_23099);
xnor U25273 (N_25273,N_22777,N_23498);
or U25274 (N_25274,N_23346,N_23238);
nor U25275 (N_25275,N_23532,N_23351);
and U25276 (N_25276,N_23207,N_22989);
and U25277 (N_25277,N_23279,N_22611);
and U25278 (N_25278,N_23578,N_22296);
and U25279 (N_25279,N_23503,N_22246);
nand U25280 (N_25280,N_22113,N_22311);
nor U25281 (N_25281,N_22340,N_23684);
nand U25282 (N_25282,N_22873,N_23887);
and U25283 (N_25283,N_23836,N_23920);
xnor U25284 (N_25284,N_22897,N_23225);
and U25285 (N_25285,N_23483,N_23241);
xor U25286 (N_25286,N_23293,N_22678);
xor U25287 (N_25287,N_22968,N_23656);
or U25288 (N_25288,N_23843,N_22915);
nor U25289 (N_25289,N_22748,N_23483);
and U25290 (N_25290,N_23440,N_23349);
xor U25291 (N_25291,N_23856,N_22653);
xor U25292 (N_25292,N_22813,N_22790);
xnor U25293 (N_25293,N_22319,N_22605);
nor U25294 (N_25294,N_22997,N_22885);
and U25295 (N_25295,N_23502,N_22655);
or U25296 (N_25296,N_23555,N_23389);
xor U25297 (N_25297,N_22226,N_22160);
and U25298 (N_25298,N_23136,N_22762);
or U25299 (N_25299,N_23314,N_23262);
nor U25300 (N_25300,N_23576,N_22625);
nand U25301 (N_25301,N_22757,N_23990);
and U25302 (N_25302,N_22725,N_22813);
xor U25303 (N_25303,N_22115,N_22930);
nor U25304 (N_25304,N_22122,N_23628);
and U25305 (N_25305,N_22051,N_22504);
nand U25306 (N_25306,N_23775,N_23044);
or U25307 (N_25307,N_23643,N_22962);
xnor U25308 (N_25308,N_22957,N_23812);
xnor U25309 (N_25309,N_23789,N_22942);
xnor U25310 (N_25310,N_22716,N_23893);
xnor U25311 (N_25311,N_22212,N_23934);
nand U25312 (N_25312,N_23168,N_23017);
or U25313 (N_25313,N_22821,N_22282);
and U25314 (N_25314,N_23777,N_23367);
or U25315 (N_25315,N_23367,N_23171);
xor U25316 (N_25316,N_22699,N_22089);
and U25317 (N_25317,N_22867,N_23047);
nand U25318 (N_25318,N_22025,N_23128);
and U25319 (N_25319,N_22738,N_23764);
nand U25320 (N_25320,N_23580,N_22603);
nand U25321 (N_25321,N_23318,N_23862);
nand U25322 (N_25322,N_22498,N_23335);
and U25323 (N_25323,N_22947,N_22494);
xor U25324 (N_25324,N_23643,N_23522);
or U25325 (N_25325,N_23547,N_22195);
nor U25326 (N_25326,N_22483,N_22616);
nand U25327 (N_25327,N_22073,N_22094);
and U25328 (N_25328,N_22487,N_22232);
xor U25329 (N_25329,N_23549,N_22858);
nand U25330 (N_25330,N_23431,N_22566);
nor U25331 (N_25331,N_23272,N_23547);
nor U25332 (N_25332,N_22041,N_23354);
or U25333 (N_25333,N_23710,N_22368);
nor U25334 (N_25334,N_22063,N_22091);
nor U25335 (N_25335,N_22918,N_22692);
or U25336 (N_25336,N_23174,N_23908);
and U25337 (N_25337,N_23103,N_23770);
nand U25338 (N_25338,N_22736,N_23704);
xnor U25339 (N_25339,N_23605,N_23193);
or U25340 (N_25340,N_22297,N_22088);
xnor U25341 (N_25341,N_23207,N_22036);
nand U25342 (N_25342,N_23118,N_23088);
and U25343 (N_25343,N_22133,N_22053);
xnor U25344 (N_25344,N_23693,N_23422);
nor U25345 (N_25345,N_23535,N_22954);
nand U25346 (N_25346,N_23101,N_22639);
and U25347 (N_25347,N_23835,N_23923);
and U25348 (N_25348,N_23934,N_23158);
nand U25349 (N_25349,N_23805,N_23252);
xnor U25350 (N_25350,N_23756,N_23452);
nand U25351 (N_25351,N_22486,N_22662);
nand U25352 (N_25352,N_22318,N_23959);
nor U25353 (N_25353,N_23157,N_23096);
or U25354 (N_25354,N_23264,N_22550);
nand U25355 (N_25355,N_23929,N_23825);
xnor U25356 (N_25356,N_23457,N_22809);
nor U25357 (N_25357,N_23047,N_23350);
xnor U25358 (N_25358,N_23363,N_23253);
xnor U25359 (N_25359,N_23576,N_22955);
nor U25360 (N_25360,N_22768,N_23472);
or U25361 (N_25361,N_23347,N_23138);
nor U25362 (N_25362,N_22230,N_23575);
or U25363 (N_25363,N_23127,N_22126);
or U25364 (N_25364,N_23813,N_23941);
xnor U25365 (N_25365,N_23223,N_22983);
and U25366 (N_25366,N_23532,N_23380);
nor U25367 (N_25367,N_23094,N_22218);
and U25368 (N_25368,N_22749,N_22325);
nor U25369 (N_25369,N_22388,N_23672);
nor U25370 (N_25370,N_23212,N_23442);
xnor U25371 (N_25371,N_23922,N_23775);
xor U25372 (N_25372,N_23886,N_22186);
and U25373 (N_25373,N_22712,N_23906);
nor U25374 (N_25374,N_23212,N_23080);
nor U25375 (N_25375,N_22325,N_23874);
or U25376 (N_25376,N_22354,N_23024);
nor U25377 (N_25377,N_23010,N_22053);
or U25378 (N_25378,N_23848,N_22740);
and U25379 (N_25379,N_23919,N_23521);
or U25380 (N_25380,N_23572,N_22735);
or U25381 (N_25381,N_23614,N_23297);
nor U25382 (N_25382,N_23187,N_23051);
nor U25383 (N_25383,N_22527,N_22269);
xor U25384 (N_25384,N_22953,N_22719);
and U25385 (N_25385,N_23770,N_23790);
xor U25386 (N_25386,N_23378,N_23048);
nor U25387 (N_25387,N_22698,N_23679);
xor U25388 (N_25388,N_22005,N_22262);
and U25389 (N_25389,N_23427,N_22431);
nor U25390 (N_25390,N_22140,N_23835);
xnor U25391 (N_25391,N_22072,N_23356);
xor U25392 (N_25392,N_22805,N_23190);
or U25393 (N_25393,N_22463,N_23385);
and U25394 (N_25394,N_23669,N_22290);
nand U25395 (N_25395,N_22129,N_23975);
or U25396 (N_25396,N_22934,N_23471);
and U25397 (N_25397,N_22680,N_22574);
nor U25398 (N_25398,N_22626,N_22716);
or U25399 (N_25399,N_23321,N_22954);
nand U25400 (N_25400,N_23662,N_23342);
xor U25401 (N_25401,N_23461,N_22762);
nand U25402 (N_25402,N_22637,N_23582);
nor U25403 (N_25403,N_23910,N_22592);
or U25404 (N_25404,N_22646,N_23645);
or U25405 (N_25405,N_22716,N_23176);
or U25406 (N_25406,N_22553,N_22255);
nor U25407 (N_25407,N_23589,N_22886);
xor U25408 (N_25408,N_22170,N_22502);
and U25409 (N_25409,N_23846,N_22303);
nand U25410 (N_25410,N_23998,N_23902);
and U25411 (N_25411,N_23860,N_23499);
or U25412 (N_25412,N_22874,N_23042);
and U25413 (N_25413,N_23635,N_23867);
nand U25414 (N_25414,N_23715,N_22399);
xor U25415 (N_25415,N_22481,N_22052);
nor U25416 (N_25416,N_22607,N_23974);
nor U25417 (N_25417,N_23096,N_22976);
xnor U25418 (N_25418,N_23133,N_22546);
nand U25419 (N_25419,N_22971,N_22045);
or U25420 (N_25420,N_22353,N_23644);
or U25421 (N_25421,N_22453,N_23303);
xor U25422 (N_25422,N_22107,N_22417);
or U25423 (N_25423,N_23834,N_23581);
xor U25424 (N_25424,N_23326,N_22242);
and U25425 (N_25425,N_22699,N_23635);
or U25426 (N_25426,N_23479,N_23393);
and U25427 (N_25427,N_22577,N_23652);
nand U25428 (N_25428,N_23378,N_22258);
and U25429 (N_25429,N_22528,N_22905);
or U25430 (N_25430,N_22112,N_23674);
nand U25431 (N_25431,N_22272,N_22909);
nor U25432 (N_25432,N_22510,N_22176);
or U25433 (N_25433,N_22366,N_23501);
nor U25434 (N_25434,N_23231,N_22446);
nand U25435 (N_25435,N_23250,N_22983);
nand U25436 (N_25436,N_23118,N_23820);
or U25437 (N_25437,N_23879,N_22624);
xnor U25438 (N_25438,N_23364,N_22125);
or U25439 (N_25439,N_22606,N_22435);
and U25440 (N_25440,N_23263,N_22389);
nand U25441 (N_25441,N_23772,N_23914);
nand U25442 (N_25442,N_22371,N_22686);
nand U25443 (N_25443,N_23210,N_22194);
nand U25444 (N_25444,N_23997,N_23353);
and U25445 (N_25445,N_23104,N_23250);
or U25446 (N_25446,N_22980,N_22480);
xnor U25447 (N_25447,N_23729,N_23464);
nor U25448 (N_25448,N_22775,N_23938);
xnor U25449 (N_25449,N_22457,N_23377);
xnor U25450 (N_25450,N_22742,N_23766);
nand U25451 (N_25451,N_23532,N_23523);
xor U25452 (N_25452,N_22689,N_23390);
xor U25453 (N_25453,N_22629,N_22150);
xor U25454 (N_25454,N_22233,N_23245);
xnor U25455 (N_25455,N_22518,N_23094);
or U25456 (N_25456,N_22592,N_23471);
or U25457 (N_25457,N_23232,N_22983);
and U25458 (N_25458,N_23282,N_23173);
and U25459 (N_25459,N_22408,N_22577);
xor U25460 (N_25460,N_22497,N_22682);
and U25461 (N_25461,N_23787,N_23508);
nor U25462 (N_25462,N_22080,N_22886);
xor U25463 (N_25463,N_23578,N_22172);
or U25464 (N_25464,N_23856,N_23918);
and U25465 (N_25465,N_22930,N_22659);
xnor U25466 (N_25466,N_22591,N_22544);
nand U25467 (N_25467,N_23907,N_23256);
nor U25468 (N_25468,N_22635,N_23194);
nand U25469 (N_25469,N_23723,N_22819);
nand U25470 (N_25470,N_23718,N_22814);
xnor U25471 (N_25471,N_23378,N_23704);
nor U25472 (N_25472,N_22447,N_23099);
nor U25473 (N_25473,N_23247,N_22895);
nor U25474 (N_25474,N_23881,N_23344);
nor U25475 (N_25475,N_22373,N_22193);
nand U25476 (N_25476,N_23011,N_23623);
nor U25477 (N_25477,N_22561,N_23696);
nand U25478 (N_25478,N_23589,N_23319);
nor U25479 (N_25479,N_22941,N_22690);
nor U25480 (N_25480,N_23369,N_23898);
or U25481 (N_25481,N_22709,N_23182);
nand U25482 (N_25482,N_22007,N_22747);
or U25483 (N_25483,N_22687,N_22186);
nor U25484 (N_25484,N_23693,N_22929);
or U25485 (N_25485,N_23432,N_23066);
or U25486 (N_25486,N_23140,N_22181);
nor U25487 (N_25487,N_23799,N_22989);
and U25488 (N_25488,N_23984,N_22942);
xnor U25489 (N_25489,N_22287,N_22279);
or U25490 (N_25490,N_23959,N_22411);
and U25491 (N_25491,N_22528,N_22841);
and U25492 (N_25492,N_22461,N_23590);
and U25493 (N_25493,N_23087,N_23753);
and U25494 (N_25494,N_22547,N_22181);
or U25495 (N_25495,N_23857,N_22311);
or U25496 (N_25496,N_23083,N_22887);
or U25497 (N_25497,N_23198,N_23187);
nor U25498 (N_25498,N_22109,N_23790);
xnor U25499 (N_25499,N_22806,N_22860);
or U25500 (N_25500,N_22325,N_22206);
nand U25501 (N_25501,N_23314,N_23127);
nor U25502 (N_25502,N_23048,N_22478);
and U25503 (N_25503,N_22998,N_22016);
and U25504 (N_25504,N_22926,N_22879);
and U25505 (N_25505,N_23220,N_23439);
nand U25506 (N_25506,N_22671,N_22892);
nor U25507 (N_25507,N_23007,N_22877);
nand U25508 (N_25508,N_22577,N_22672);
or U25509 (N_25509,N_22690,N_22418);
nand U25510 (N_25510,N_23504,N_22815);
nand U25511 (N_25511,N_23739,N_23334);
xor U25512 (N_25512,N_22488,N_23552);
nand U25513 (N_25513,N_22503,N_23691);
nor U25514 (N_25514,N_22937,N_22441);
xor U25515 (N_25515,N_22814,N_23387);
and U25516 (N_25516,N_22469,N_22855);
or U25517 (N_25517,N_22430,N_23590);
or U25518 (N_25518,N_23235,N_22513);
and U25519 (N_25519,N_23666,N_22287);
xnor U25520 (N_25520,N_22025,N_22482);
nor U25521 (N_25521,N_23437,N_22352);
and U25522 (N_25522,N_23174,N_23613);
and U25523 (N_25523,N_22992,N_22796);
nand U25524 (N_25524,N_23839,N_22848);
and U25525 (N_25525,N_22857,N_23182);
or U25526 (N_25526,N_23577,N_22594);
nand U25527 (N_25527,N_22350,N_23672);
and U25528 (N_25528,N_23247,N_22765);
or U25529 (N_25529,N_22919,N_22297);
or U25530 (N_25530,N_23378,N_23748);
and U25531 (N_25531,N_22345,N_22463);
and U25532 (N_25532,N_22330,N_23459);
and U25533 (N_25533,N_23611,N_22747);
and U25534 (N_25534,N_22999,N_22389);
and U25535 (N_25535,N_22612,N_23688);
xnor U25536 (N_25536,N_22609,N_22960);
xor U25537 (N_25537,N_23244,N_22108);
xor U25538 (N_25538,N_22718,N_23483);
nand U25539 (N_25539,N_22244,N_22497);
nand U25540 (N_25540,N_23040,N_23695);
nor U25541 (N_25541,N_22442,N_23323);
nand U25542 (N_25542,N_22243,N_23936);
xnor U25543 (N_25543,N_22606,N_23666);
and U25544 (N_25544,N_22654,N_23510);
or U25545 (N_25545,N_22226,N_23694);
and U25546 (N_25546,N_23311,N_23259);
xnor U25547 (N_25547,N_23120,N_23348);
or U25548 (N_25548,N_23929,N_23049);
and U25549 (N_25549,N_22320,N_23975);
nor U25550 (N_25550,N_22956,N_22982);
nor U25551 (N_25551,N_22665,N_23789);
nor U25552 (N_25552,N_23786,N_23304);
nor U25553 (N_25553,N_22344,N_23366);
or U25554 (N_25554,N_23010,N_22593);
nor U25555 (N_25555,N_23469,N_23612);
and U25556 (N_25556,N_22100,N_23157);
nor U25557 (N_25557,N_23479,N_23456);
and U25558 (N_25558,N_22205,N_23148);
and U25559 (N_25559,N_23386,N_23212);
xor U25560 (N_25560,N_22107,N_22352);
xor U25561 (N_25561,N_23054,N_22173);
or U25562 (N_25562,N_23368,N_22805);
xnor U25563 (N_25563,N_23812,N_22486);
and U25564 (N_25564,N_22022,N_23257);
nor U25565 (N_25565,N_23262,N_23297);
nor U25566 (N_25566,N_22234,N_22286);
nand U25567 (N_25567,N_23590,N_22676);
or U25568 (N_25568,N_23292,N_22615);
xor U25569 (N_25569,N_22540,N_23333);
or U25570 (N_25570,N_23786,N_22188);
and U25571 (N_25571,N_23019,N_22342);
or U25572 (N_25572,N_22588,N_23022);
nor U25573 (N_25573,N_23361,N_23607);
nand U25574 (N_25574,N_23871,N_22429);
nand U25575 (N_25575,N_22295,N_22430);
or U25576 (N_25576,N_22285,N_22062);
nand U25577 (N_25577,N_23470,N_22691);
or U25578 (N_25578,N_22625,N_22480);
xor U25579 (N_25579,N_23707,N_22661);
nand U25580 (N_25580,N_22435,N_23145);
or U25581 (N_25581,N_22189,N_22192);
xnor U25582 (N_25582,N_22134,N_23115);
xnor U25583 (N_25583,N_23159,N_23740);
xnor U25584 (N_25584,N_22160,N_23045);
or U25585 (N_25585,N_23147,N_23386);
xnor U25586 (N_25586,N_23607,N_22293);
nor U25587 (N_25587,N_22409,N_23866);
and U25588 (N_25588,N_22609,N_23469);
nand U25589 (N_25589,N_22265,N_22302);
and U25590 (N_25590,N_23338,N_23580);
xor U25591 (N_25591,N_22997,N_22356);
nor U25592 (N_25592,N_22948,N_23754);
nor U25593 (N_25593,N_23795,N_23774);
nand U25594 (N_25594,N_22107,N_22683);
nor U25595 (N_25595,N_23896,N_23160);
or U25596 (N_25596,N_22986,N_23516);
or U25597 (N_25597,N_23609,N_22321);
xor U25598 (N_25598,N_22604,N_23731);
or U25599 (N_25599,N_23921,N_23982);
or U25600 (N_25600,N_23342,N_22817);
or U25601 (N_25601,N_23655,N_23106);
or U25602 (N_25602,N_22642,N_23174);
or U25603 (N_25603,N_23790,N_22978);
and U25604 (N_25604,N_23207,N_23353);
nor U25605 (N_25605,N_23192,N_22763);
xor U25606 (N_25606,N_23945,N_22619);
nor U25607 (N_25607,N_22060,N_23619);
and U25608 (N_25608,N_22450,N_23711);
nand U25609 (N_25609,N_23534,N_23947);
nor U25610 (N_25610,N_22955,N_22899);
nor U25611 (N_25611,N_23768,N_22019);
or U25612 (N_25612,N_22014,N_22725);
xnor U25613 (N_25613,N_23357,N_23084);
and U25614 (N_25614,N_23701,N_23329);
and U25615 (N_25615,N_23223,N_22536);
and U25616 (N_25616,N_23357,N_23667);
xnor U25617 (N_25617,N_22645,N_22714);
nand U25618 (N_25618,N_22821,N_23716);
nand U25619 (N_25619,N_23910,N_23196);
or U25620 (N_25620,N_23548,N_23421);
nor U25621 (N_25621,N_23963,N_23479);
nor U25622 (N_25622,N_23950,N_22854);
and U25623 (N_25623,N_22481,N_23328);
xnor U25624 (N_25624,N_23901,N_22213);
and U25625 (N_25625,N_22212,N_23289);
or U25626 (N_25626,N_23737,N_23901);
xor U25627 (N_25627,N_22210,N_23828);
nor U25628 (N_25628,N_23981,N_22192);
or U25629 (N_25629,N_22677,N_23494);
nand U25630 (N_25630,N_23672,N_23532);
nand U25631 (N_25631,N_23628,N_23824);
nand U25632 (N_25632,N_23895,N_22949);
nor U25633 (N_25633,N_23470,N_22735);
and U25634 (N_25634,N_22479,N_23308);
xor U25635 (N_25635,N_22442,N_22240);
nor U25636 (N_25636,N_23868,N_23363);
nor U25637 (N_25637,N_22091,N_23768);
and U25638 (N_25638,N_22730,N_22213);
xor U25639 (N_25639,N_22915,N_22522);
nor U25640 (N_25640,N_22146,N_23536);
nor U25641 (N_25641,N_22341,N_23416);
and U25642 (N_25642,N_22065,N_22769);
nor U25643 (N_25643,N_22957,N_23109);
and U25644 (N_25644,N_23933,N_23882);
xnor U25645 (N_25645,N_23606,N_23968);
or U25646 (N_25646,N_22257,N_22189);
nand U25647 (N_25647,N_22614,N_23621);
and U25648 (N_25648,N_23169,N_23726);
nor U25649 (N_25649,N_23537,N_22279);
or U25650 (N_25650,N_22303,N_23407);
nand U25651 (N_25651,N_22238,N_22435);
xor U25652 (N_25652,N_23085,N_23485);
nor U25653 (N_25653,N_22485,N_23187);
nor U25654 (N_25654,N_22922,N_23636);
nand U25655 (N_25655,N_23066,N_23526);
xnor U25656 (N_25656,N_23548,N_22541);
xor U25657 (N_25657,N_23646,N_23004);
nor U25658 (N_25658,N_23914,N_23385);
nor U25659 (N_25659,N_23895,N_22891);
or U25660 (N_25660,N_22551,N_23264);
or U25661 (N_25661,N_22662,N_23808);
nand U25662 (N_25662,N_22708,N_22812);
xnor U25663 (N_25663,N_23933,N_22722);
and U25664 (N_25664,N_23584,N_22531);
nor U25665 (N_25665,N_23225,N_22101);
xor U25666 (N_25666,N_23633,N_22476);
nor U25667 (N_25667,N_22951,N_22823);
nor U25668 (N_25668,N_22633,N_23070);
xnor U25669 (N_25669,N_23681,N_22376);
nor U25670 (N_25670,N_22786,N_23092);
or U25671 (N_25671,N_23825,N_22070);
xnor U25672 (N_25672,N_23476,N_22096);
and U25673 (N_25673,N_22943,N_23553);
and U25674 (N_25674,N_22281,N_22688);
nor U25675 (N_25675,N_22942,N_22055);
xnor U25676 (N_25676,N_23322,N_22712);
nand U25677 (N_25677,N_23830,N_22632);
xor U25678 (N_25678,N_22570,N_23136);
nand U25679 (N_25679,N_22105,N_23559);
nand U25680 (N_25680,N_23580,N_22066);
nand U25681 (N_25681,N_23844,N_23564);
or U25682 (N_25682,N_23158,N_22309);
or U25683 (N_25683,N_23942,N_22362);
and U25684 (N_25684,N_23457,N_22043);
nor U25685 (N_25685,N_22071,N_22558);
nor U25686 (N_25686,N_23934,N_22479);
nor U25687 (N_25687,N_23239,N_22074);
nand U25688 (N_25688,N_22318,N_23376);
nand U25689 (N_25689,N_23836,N_22742);
xor U25690 (N_25690,N_23534,N_23678);
nand U25691 (N_25691,N_22956,N_23200);
and U25692 (N_25692,N_22397,N_22656);
and U25693 (N_25693,N_22687,N_22263);
and U25694 (N_25694,N_23465,N_22890);
xor U25695 (N_25695,N_23098,N_22740);
and U25696 (N_25696,N_22474,N_22030);
and U25697 (N_25697,N_23152,N_22478);
or U25698 (N_25698,N_22276,N_22935);
or U25699 (N_25699,N_22312,N_22027);
nand U25700 (N_25700,N_23599,N_22484);
nand U25701 (N_25701,N_23455,N_22929);
or U25702 (N_25702,N_23358,N_23991);
and U25703 (N_25703,N_23893,N_23336);
xnor U25704 (N_25704,N_22266,N_22154);
nor U25705 (N_25705,N_22219,N_23432);
nor U25706 (N_25706,N_22623,N_23483);
or U25707 (N_25707,N_22733,N_23440);
xnor U25708 (N_25708,N_23435,N_22153);
or U25709 (N_25709,N_23217,N_23634);
or U25710 (N_25710,N_22727,N_22191);
nor U25711 (N_25711,N_22413,N_23190);
nand U25712 (N_25712,N_22800,N_23322);
nor U25713 (N_25713,N_22660,N_22749);
and U25714 (N_25714,N_22139,N_22485);
xnor U25715 (N_25715,N_22674,N_22128);
or U25716 (N_25716,N_23963,N_22224);
nand U25717 (N_25717,N_22440,N_23981);
nand U25718 (N_25718,N_23332,N_23828);
or U25719 (N_25719,N_23290,N_23426);
or U25720 (N_25720,N_22417,N_23085);
or U25721 (N_25721,N_23383,N_23658);
nand U25722 (N_25722,N_23146,N_22281);
xor U25723 (N_25723,N_22389,N_23349);
nand U25724 (N_25724,N_22697,N_23507);
nand U25725 (N_25725,N_23620,N_23693);
and U25726 (N_25726,N_22328,N_23775);
nand U25727 (N_25727,N_23370,N_22016);
nand U25728 (N_25728,N_22246,N_23657);
xor U25729 (N_25729,N_23891,N_23019);
or U25730 (N_25730,N_23425,N_22680);
nor U25731 (N_25731,N_22607,N_23510);
nand U25732 (N_25732,N_23159,N_23691);
xnor U25733 (N_25733,N_23886,N_23228);
nor U25734 (N_25734,N_22301,N_23726);
nand U25735 (N_25735,N_22919,N_22825);
nor U25736 (N_25736,N_22471,N_22398);
nand U25737 (N_25737,N_23314,N_23518);
and U25738 (N_25738,N_23943,N_22414);
and U25739 (N_25739,N_22499,N_23969);
and U25740 (N_25740,N_22599,N_22495);
and U25741 (N_25741,N_23144,N_22093);
and U25742 (N_25742,N_22725,N_22021);
and U25743 (N_25743,N_23721,N_23676);
or U25744 (N_25744,N_22870,N_22635);
nand U25745 (N_25745,N_22069,N_22990);
nand U25746 (N_25746,N_23437,N_22622);
nor U25747 (N_25747,N_23549,N_23995);
nor U25748 (N_25748,N_22788,N_22429);
and U25749 (N_25749,N_22318,N_22732);
and U25750 (N_25750,N_23641,N_22446);
nand U25751 (N_25751,N_22877,N_23351);
nor U25752 (N_25752,N_23690,N_22990);
and U25753 (N_25753,N_23995,N_23493);
or U25754 (N_25754,N_22922,N_22012);
or U25755 (N_25755,N_23439,N_22924);
nand U25756 (N_25756,N_22312,N_23958);
xnor U25757 (N_25757,N_22733,N_22105);
nand U25758 (N_25758,N_23506,N_23704);
or U25759 (N_25759,N_22631,N_22035);
xor U25760 (N_25760,N_22321,N_23308);
nor U25761 (N_25761,N_22350,N_23784);
xnor U25762 (N_25762,N_22798,N_23692);
nor U25763 (N_25763,N_22655,N_22261);
and U25764 (N_25764,N_22719,N_23782);
nand U25765 (N_25765,N_23817,N_22581);
nand U25766 (N_25766,N_23375,N_23020);
nor U25767 (N_25767,N_23265,N_23898);
xor U25768 (N_25768,N_23295,N_22035);
nor U25769 (N_25769,N_23053,N_23763);
or U25770 (N_25770,N_23376,N_22454);
xnor U25771 (N_25771,N_23529,N_23062);
nor U25772 (N_25772,N_22260,N_22337);
xnor U25773 (N_25773,N_22026,N_22249);
and U25774 (N_25774,N_23745,N_23143);
and U25775 (N_25775,N_23109,N_23507);
xor U25776 (N_25776,N_23760,N_22918);
and U25777 (N_25777,N_22400,N_22505);
xor U25778 (N_25778,N_23011,N_23084);
and U25779 (N_25779,N_23018,N_23877);
or U25780 (N_25780,N_23407,N_23278);
or U25781 (N_25781,N_23653,N_22275);
xor U25782 (N_25782,N_23173,N_22130);
nor U25783 (N_25783,N_22865,N_23817);
xor U25784 (N_25784,N_22353,N_22451);
or U25785 (N_25785,N_22885,N_23121);
xnor U25786 (N_25786,N_22638,N_22897);
and U25787 (N_25787,N_23718,N_22460);
xnor U25788 (N_25788,N_22309,N_23819);
nand U25789 (N_25789,N_22951,N_22601);
and U25790 (N_25790,N_22269,N_23615);
and U25791 (N_25791,N_22817,N_22354);
and U25792 (N_25792,N_23674,N_23113);
nor U25793 (N_25793,N_23418,N_22611);
or U25794 (N_25794,N_23395,N_22576);
or U25795 (N_25795,N_22055,N_22256);
nor U25796 (N_25796,N_23912,N_23496);
xnor U25797 (N_25797,N_22163,N_23331);
nand U25798 (N_25798,N_23962,N_22298);
or U25799 (N_25799,N_22705,N_22746);
and U25800 (N_25800,N_23033,N_22525);
nand U25801 (N_25801,N_23600,N_23174);
nor U25802 (N_25802,N_22723,N_23880);
xor U25803 (N_25803,N_23084,N_23235);
nor U25804 (N_25804,N_23660,N_22496);
nor U25805 (N_25805,N_22043,N_23029);
nor U25806 (N_25806,N_23806,N_22730);
and U25807 (N_25807,N_22554,N_23519);
nor U25808 (N_25808,N_22448,N_23579);
nor U25809 (N_25809,N_23947,N_23967);
or U25810 (N_25810,N_23172,N_23661);
nand U25811 (N_25811,N_23201,N_22546);
or U25812 (N_25812,N_23516,N_23648);
nand U25813 (N_25813,N_23767,N_22377);
xor U25814 (N_25814,N_23102,N_23013);
xnor U25815 (N_25815,N_23956,N_22775);
xnor U25816 (N_25816,N_22096,N_23068);
xnor U25817 (N_25817,N_22206,N_22273);
nand U25818 (N_25818,N_22331,N_22771);
nor U25819 (N_25819,N_23334,N_23674);
nor U25820 (N_25820,N_22639,N_23628);
nand U25821 (N_25821,N_22512,N_22346);
and U25822 (N_25822,N_23703,N_23528);
or U25823 (N_25823,N_23290,N_22400);
and U25824 (N_25824,N_22529,N_23968);
and U25825 (N_25825,N_22896,N_22933);
or U25826 (N_25826,N_23318,N_23795);
nand U25827 (N_25827,N_23935,N_22424);
xor U25828 (N_25828,N_22440,N_22312);
or U25829 (N_25829,N_23462,N_22779);
or U25830 (N_25830,N_22941,N_23846);
xnor U25831 (N_25831,N_23286,N_23916);
or U25832 (N_25832,N_22941,N_23750);
xnor U25833 (N_25833,N_22750,N_22252);
xnor U25834 (N_25834,N_22829,N_22096);
xor U25835 (N_25835,N_22298,N_22538);
nand U25836 (N_25836,N_22405,N_23738);
and U25837 (N_25837,N_23078,N_22669);
xor U25838 (N_25838,N_22950,N_22505);
and U25839 (N_25839,N_23446,N_23822);
or U25840 (N_25840,N_22401,N_23928);
nor U25841 (N_25841,N_22212,N_22444);
nand U25842 (N_25842,N_22436,N_23253);
nor U25843 (N_25843,N_23120,N_23171);
xnor U25844 (N_25844,N_22862,N_22414);
nor U25845 (N_25845,N_22000,N_22150);
nand U25846 (N_25846,N_23046,N_22217);
nand U25847 (N_25847,N_22645,N_23766);
xnor U25848 (N_25848,N_22950,N_23583);
nor U25849 (N_25849,N_22943,N_23999);
nand U25850 (N_25850,N_23490,N_23218);
or U25851 (N_25851,N_22411,N_23865);
or U25852 (N_25852,N_23782,N_23383);
nor U25853 (N_25853,N_22860,N_22151);
or U25854 (N_25854,N_22437,N_23663);
and U25855 (N_25855,N_23143,N_23505);
or U25856 (N_25856,N_22600,N_22569);
and U25857 (N_25857,N_22319,N_22517);
nor U25858 (N_25858,N_22485,N_23852);
xor U25859 (N_25859,N_23298,N_23404);
and U25860 (N_25860,N_23316,N_23188);
or U25861 (N_25861,N_22223,N_23028);
or U25862 (N_25862,N_22308,N_23634);
and U25863 (N_25863,N_23389,N_22225);
nor U25864 (N_25864,N_22619,N_22753);
or U25865 (N_25865,N_23430,N_22763);
xnor U25866 (N_25866,N_23638,N_22091);
nand U25867 (N_25867,N_23492,N_23556);
and U25868 (N_25868,N_22249,N_22253);
nand U25869 (N_25869,N_22111,N_22919);
nand U25870 (N_25870,N_22570,N_22318);
nand U25871 (N_25871,N_22277,N_23279);
xor U25872 (N_25872,N_23721,N_23375);
and U25873 (N_25873,N_23658,N_23951);
nand U25874 (N_25874,N_23902,N_23721);
nor U25875 (N_25875,N_23448,N_23010);
nand U25876 (N_25876,N_22610,N_23006);
and U25877 (N_25877,N_23064,N_22505);
nand U25878 (N_25878,N_22165,N_23871);
nand U25879 (N_25879,N_22303,N_22404);
nand U25880 (N_25880,N_22789,N_23879);
or U25881 (N_25881,N_23856,N_22916);
xnor U25882 (N_25882,N_22464,N_22051);
or U25883 (N_25883,N_23713,N_23978);
nor U25884 (N_25884,N_23811,N_22430);
nor U25885 (N_25885,N_23895,N_23314);
or U25886 (N_25886,N_23736,N_23299);
and U25887 (N_25887,N_23610,N_22385);
or U25888 (N_25888,N_22490,N_22064);
nand U25889 (N_25889,N_22612,N_22560);
xor U25890 (N_25890,N_22114,N_23889);
xnor U25891 (N_25891,N_23034,N_22885);
nor U25892 (N_25892,N_22226,N_23751);
and U25893 (N_25893,N_23430,N_22916);
nand U25894 (N_25894,N_22450,N_23771);
or U25895 (N_25895,N_23934,N_23608);
nand U25896 (N_25896,N_23203,N_23752);
or U25897 (N_25897,N_23267,N_23902);
nor U25898 (N_25898,N_22046,N_23874);
nand U25899 (N_25899,N_23765,N_23354);
and U25900 (N_25900,N_23212,N_23479);
nor U25901 (N_25901,N_22965,N_23670);
nand U25902 (N_25902,N_22998,N_23283);
or U25903 (N_25903,N_22949,N_23138);
xor U25904 (N_25904,N_23089,N_23389);
nor U25905 (N_25905,N_23348,N_23307);
and U25906 (N_25906,N_23710,N_23336);
and U25907 (N_25907,N_22795,N_22001);
or U25908 (N_25908,N_23166,N_23573);
xor U25909 (N_25909,N_22418,N_22133);
and U25910 (N_25910,N_23906,N_23860);
xnor U25911 (N_25911,N_22196,N_22427);
or U25912 (N_25912,N_23761,N_23608);
nand U25913 (N_25913,N_23214,N_22626);
nand U25914 (N_25914,N_22702,N_23154);
or U25915 (N_25915,N_22900,N_23008);
or U25916 (N_25916,N_22219,N_23799);
xnor U25917 (N_25917,N_23662,N_23976);
xnor U25918 (N_25918,N_23369,N_22827);
nand U25919 (N_25919,N_22469,N_22104);
and U25920 (N_25920,N_23988,N_23300);
nand U25921 (N_25921,N_22983,N_22600);
nor U25922 (N_25922,N_22866,N_23301);
xor U25923 (N_25923,N_23545,N_23343);
xnor U25924 (N_25924,N_22315,N_23572);
nand U25925 (N_25925,N_22228,N_23680);
or U25926 (N_25926,N_23997,N_23390);
nand U25927 (N_25927,N_23572,N_23767);
xor U25928 (N_25928,N_22400,N_23174);
nand U25929 (N_25929,N_22714,N_23048);
nand U25930 (N_25930,N_23618,N_22269);
nor U25931 (N_25931,N_22707,N_23456);
and U25932 (N_25932,N_22571,N_23752);
or U25933 (N_25933,N_22600,N_22230);
nor U25934 (N_25934,N_23796,N_23637);
nand U25935 (N_25935,N_23726,N_23932);
or U25936 (N_25936,N_23819,N_22884);
and U25937 (N_25937,N_22766,N_23216);
and U25938 (N_25938,N_22516,N_22889);
nand U25939 (N_25939,N_22895,N_22469);
and U25940 (N_25940,N_23722,N_23358);
or U25941 (N_25941,N_23407,N_22316);
and U25942 (N_25942,N_22441,N_22604);
and U25943 (N_25943,N_23082,N_23461);
or U25944 (N_25944,N_22736,N_23610);
xnor U25945 (N_25945,N_22130,N_22468);
nor U25946 (N_25946,N_22805,N_23703);
and U25947 (N_25947,N_22953,N_22878);
nand U25948 (N_25948,N_23371,N_22708);
nor U25949 (N_25949,N_23575,N_23434);
nand U25950 (N_25950,N_23047,N_23043);
or U25951 (N_25951,N_22112,N_23609);
xor U25952 (N_25952,N_23394,N_23049);
nand U25953 (N_25953,N_22869,N_22740);
xor U25954 (N_25954,N_23704,N_22436);
and U25955 (N_25955,N_23811,N_23569);
nand U25956 (N_25956,N_23842,N_22771);
or U25957 (N_25957,N_22232,N_22090);
nor U25958 (N_25958,N_23145,N_23420);
xnor U25959 (N_25959,N_22993,N_22759);
nand U25960 (N_25960,N_22386,N_22028);
nor U25961 (N_25961,N_23607,N_23036);
nand U25962 (N_25962,N_22248,N_22739);
and U25963 (N_25963,N_22475,N_23382);
nand U25964 (N_25964,N_23140,N_22635);
and U25965 (N_25965,N_22173,N_23236);
or U25966 (N_25966,N_23939,N_22447);
nor U25967 (N_25967,N_23924,N_23531);
nand U25968 (N_25968,N_23508,N_22443);
nand U25969 (N_25969,N_23353,N_22216);
xnor U25970 (N_25970,N_23046,N_23268);
nor U25971 (N_25971,N_22894,N_23769);
nor U25972 (N_25972,N_22116,N_23393);
xnor U25973 (N_25973,N_23320,N_22217);
and U25974 (N_25974,N_23890,N_22950);
nand U25975 (N_25975,N_23450,N_23784);
xnor U25976 (N_25976,N_22570,N_23892);
xnor U25977 (N_25977,N_23609,N_22723);
xor U25978 (N_25978,N_22684,N_23342);
and U25979 (N_25979,N_23275,N_23403);
and U25980 (N_25980,N_23959,N_23452);
and U25981 (N_25981,N_22944,N_23179);
and U25982 (N_25982,N_22165,N_23629);
xor U25983 (N_25983,N_22585,N_22727);
or U25984 (N_25984,N_23954,N_23112);
xor U25985 (N_25985,N_23901,N_23819);
nor U25986 (N_25986,N_23440,N_23619);
and U25987 (N_25987,N_23210,N_22852);
and U25988 (N_25988,N_22785,N_23645);
nand U25989 (N_25989,N_22573,N_23020);
nor U25990 (N_25990,N_22288,N_23277);
nand U25991 (N_25991,N_22487,N_23200);
and U25992 (N_25992,N_23649,N_22292);
nand U25993 (N_25993,N_22046,N_22977);
and U25994 (N_25994,N_23088,N_23486);
nor U25995 (N_25995,N_22764,N_23249);
and U25996 (N_25996,N_22236,N_23872);
xnor U25997 (N_25997,N_23549,N_23960);
or U25998 (N_25998,N_22736,N_22339);
and U25999 (N_25999,N_23086,N_23400);
or U26000 (N_26000,N_24978,N_25600);
xor U26001 (N_26001,N_25541,N_25474);
and U26002 (N_26002,N_25222,N_25763);
and U26003 (N_26003,N_24675,N_24210);
and U26004 (N_26004,N_24533,N_24437);
and U26005 (N_26005,N_24269,N_24400);
nand U26006 (N_26006,N_25574,N_25736);
xnor U26007 (N_26007,N_24149,N_25581);
or U26008 (N_26008,N_25213,N_24871);
nand U26009 (N_26009,N_25792,N_24282);
xnor U26010 (N_26010,N_25329,N_24514);
or U26011 (N_26011,N_24952,N_25592);
nor U26012 (N_26012,N_25523,N_25983);
and U26013 (N_26013,N_25793,N_25399);
nand U26014 (N_26014,N_24196,N_25454);
and U26015 (N_26015,N_25150,N_24671);
and U26016 (N_26016,N_24133,N_24470);
or U26017 (N_26017,N_24647,N_25760);
xnor U26018 (N_26018,N_24251,N_25543);
nor U26019 (N_26019,N_25400,N_24369);
xor U26020 (N_26020,N_24655,N_25841);
nor U26021 (N_26021,N_24834,N_24016);
or U26022 (N_26022,N_24773,N_24505);
nor U26023 (N_26023,N_24605,N_24979);
xnor U26024 (N_26024,N_24967,N_25549);
and U26025 (N_26025,N_24167,N_24005);
and U26026 (N_26026,N_24614,N_24752);
xor U26027 (N_26027,N_25065,N_24803);
xor U26028 (N_26028,N_25250,N_25082);
nand U26029 (N_26029,N_25708,N_24218);
nand U26030 (N_26030,N_24715,N_25071);
nand U26031 (N_26031,N_25243,N_24071);
xor U26032 (N_26032,N_25432,N_24636);
nor U26033 (N_26033,N_25401,N_24989);
nand U26034 (N_26034,N_24646,N_24777);
nor U26035 (N_26035,N_24556,N_24964);
nand U26036 (N_26036,N_25623,N_25709);
xnor U26037 (N_26037,N_25025,N_24613);
or U26038 (N_26038,N_25010,N_24105);
and U26039 (N_26039,N_25402,N_25536);
and U26040 (N_26040,N_24631,N_25113);
and U26041 (N_26041,N_25202,N_25964);
nand U26042 (N_26042,N_24254,N_25811);
or U26043 (N_26043,N_25864,N_25188);
nand U26044 (N_26044,N_24085,N_24199);
nand U26045 (N_26045,N_24447,N_25285);
nor U26046 (N_26046,N_24540,N_24585);
and U26047 (N_26047,N_25386,N_24442);
xor U26048 (N_26048,N_25049,N_24142);
xor U26049 (N_26049,N_25733,N_24281);
xor U26050 (N_26050,N_24096,N_25157);
nor U26051 (N_26051,N_25994,N_24541);
nor U26052 (N_26052,N_25815,N_24579);
nor U26053 (N_26053,N_25052,N_24279);
xor U26054 (N_26054,N_25293,N_24880);
or U26055 (N_26055,N_24306,N_24924);
nand U26056 (N_26056,N_25120,N_25347);
xnor U26057 (N_26057,N_24986,N_25012);
nor U26058 (N_26058,N_24980,N_25149);
xnor U26059 (N_26059,N_25894,N_25738);
nor U26060 (N_26060,N_25415,N_25699);
xnor U26061 (N_26061,N_25911,N_25999);
xnor U26062 (N_26062,N_25606,N_24366);
nand U26063 (N_26063,N_24238,N_24991);
and U26064 (N_26064,N_25365,N_24955);
nand U26065 (N_26065,N_24152,N_25987);
or U26066 (N_26066,N_25234,N_25859);
xor U26067 (N_26067,N_25725,N_25836);
nor U26068 (N_26068,N_24239,N_25018);
xor U26069 (N_26069,N_25308,N_24602);
nor U26070 (N_26070,N_25086,N_25253);
or U26071 (N_26071,N_24582,N_25033);
nor U26072 (N_26072,N_25895,N_25102);
nor U26073 (N_26073,N_25445,N_24345);
nor U26074 (N_26074,N_24274,N_25573);
or U26075 (N_26075,N_25115,N_24225);
and U26076 (N_26076,N_24235,N_24736);
or U26077 (N_26077,N_25818,N_24748);
nor U26078 (N_26078,N_24686,N_25050);
xor U26079 (N_26079,N_25156,N_24053);
nor U26080 (N_26080,N_24350,N_24531);
or U26081 (N_26081,N_24034,N_25603);
nand U26082 (N_26082,N_25460,N_25459);
or U26083 (N_26083,N_24909,N_25970);
and U26084 (N_26084,N_24323,N_25967);
and U26085 (N_26085,N_25788,N_24129);
nand U26086 (N_26086,N_24520,N_25302);
and U26087 (N_26087,N_25363,N_25048);
nor U26088 (N_26088,N_25391,N_24000);
and U26089 (N_26089,N_25502,N_25403);
nor U26090 (N_26090,N_24993,N_25320);
xnor U26091 (N_26091,N_24289,N_24185);
nor U26092 (N_26092,N_25147,N_24312);
and U26093 (N_26093,N_24676,N_24878);
nand U26094 (N_26094,N_25580,N_25439);
or U26095 (N_26095,N_25642,N_25548);
xor U26096 (N_26096,N_24396,N_24120);
xor U26097 (N_26097,N_24855,N_25241);
or U26098 (N_26098,N_25628,N_25865);
nor U26099 (N_26099,N_25912,N_25722);
or U26100 (N_26100,N_24528,N_24764);
and U26101 (N_26101,N_25977,N_24162);
xnor U26102 (N_26102,N_25526,N_24672);
nand U26103 (N_26103,N_25638,N_25996);
xor U26104 (N_26104,N_25923,N_25879);
nor U26105 (N_26105,N_24895,N_24427);
and U26106 (N_26106,N_25404,N_24551);
and U26107 (N_26107,N_25383,N_24190);
nand U26108 (N_26108,N_25267,N_25579);
and U26109 (N_26109,N_24692,N_24667);
and U26110 (N_26110,N_25101,N_25051);
nor U26111 (N_26111,N_24829,N_25944);
nor U26112 (N_26112,N_24694,N_25896);
or U26113 (N_26113,N_25099,N_25719);
and U26114 (N_26114,N_24604,N_24285);
nor U26115 (N_26115,N_25428,N_25007);
xnor U26116 (N_26116,N_25845,N_25910);
or U26117 (N_26117,N_25244,N_24429);
xnor U26118 (N_26118,N_25986,N_25494);
xor U26119 (N_26119,N_25472,N_24224);
or U26120 (N_26120,N_25332,N_24554);
xnor U26121 (N_26121,N_25956,N_25255);
or U26122 (N_26122,N_24450,N_24992);
and U26123 (N_26123,N_25905,N_25118);
nor U26124 (N_26124,N_24297,N_25351);
nor U26125 (N_26125,N_24590,N_24738);
and U26126 (N_26126,N_24789,N_25350);
xnor U26127 (N_26127,N_24823,N_24500);
xnor U26128 (N_26128,N_25930,N_25920);
nor U26129 (N_26129,N_24355,N_25798);
xnor U26130 (N_26130,N_25181,N_24147);
and U26131 (N_26131,N_24161,N_24349);
nor U26132 (N_26132,N_25254,N_25624);
and U26133 (N_26133,N_24184,N_25989);
nand U26134 (N_26134,N_25416,N_25500);
and U26135 (N_26135,N_25395,N_24697);
and U26136 (N_26136,N_24765,N_24290);
or U26137 (N_26137,N_24869,N_25616);
and U26138 (N_26138,N_24130,N_24191);
nand U26139 (N_26139,N_25665,N_24775);
xnor U26140 (N_26140,N_24673,N_25433);
or U26141 (N_26141,N_24173,N_25177);
or U26142 (N_26142,N_24507,N_24592);
and U26143 (N_26143,N_24017,N_25870);
and U26144 (N_26144,N_25852,N_24305);
xor U26145 (N_26145,N_25377,N_25611);
nand U26146 (N_26146,N_24918,N_24325);
and U26147 (N_26147,N_24719,N_24601);
and U26148 (N_26148,N_25278,N_25040);
nor U26149 (N_26149,N_25078,N_24808);
or U26150 (N_26150,N_24578,N_25368);
nand U26151 (N_26151,N_25069,N_25701);
xnor U26152 (N_26152,N_24916,N_25819);
xnor U26153 (N_26153,N_25483,N_24768);
xor U26154 (N_26154,N_24820,N_25307);
nand U26155 (N_26155,N_25371,N_25979);
xor U26156 (N_26156,N_25245,N_25199);
nand U26157 (N_26157,N_25675,N_25272);
and U26158 (N_26158,N_25676,N_24093);
and U26159 (N_26159,N_25785,N_24308);
xor U26160 (N_26160,N_25858,N_25876);
and U26161 (N_26161,N_24075,N_25723);
nor U26162 (N_26162,N_24669,N_24856);
nand U26163 (N_26163,N_25620,N_25715);
nor U26164 (N_26164,N_24351,N_24957);
nor U26165 (N_26165,N_24213,N_24063);
nor U26166 (N_26166,N_24230,N_25506);
nor U26167 (N_26167,N_24391,N_24243);
nor U26168 (N_26168,N_24004,N_25759);
and U26169 (N_26169,N_25200,N_25087);
or U26170 (N_26170,N_25303,N_25937);
and U26171 (N_26171,N_24203,N_24996);
nand U26172 (N_26172,N_25093,N_24890);
nand U26173 (N_26173,N_25651,N_25497);
nand U26174 (N_26174,N_24244,N_25140);
nand U26175 (N_26175,N_25597,N_24713);
or U26176 (N_26176,N_25995,N_25521);
nand U26177 (N_26177,N_25513,N_24958);
or U26178 (N_26178,N_24268,N_25569);
nor U26179 (N_26179,N_25297,N_25367);
xnor U26180 (N_26180,N_25074,N_25327);
nand U26181 (N_26181,N_25323,N_25027);
or U26182 (N_26182,N_25343,N_24641);
nand U26183 (N_26183,N_25288,N_24946);
nand U26184 (N_26184,N_24035,N_24570);
or U26185 (N_26185,N_25583,N_24402);
nor U26186 (N_26186,N_25957,N_24569);
or U26187 (N_26187,N_24644,N_24434);
or U26188 (N_26188,N_25528,N_24907);
nor U26189 (N_26189,N_25008,N_25850);
or U26190 (N_26190,N_24490,N_24705);
nor U26191 (N_26191,N_25560,N_24198);
or U26192 (N_26192,N_25516,N_25717);
xor U26193 (N_26193,N_25387,N_25290);
nor U26194 (N_26194,N_25389,N_24801);
nand U26195 (N_26195,N_24215,N_25262);
or U26196 (N_26196,N_24553,N_24538);
or U26197 (N_26197,N_25982,N_25265);
nand U26198 (N_26198,N_24475,N_25384);
nor U26199 (N_26199,N_24148,N_25457);
or U26200 (N_26200,N_24114,N_25807);
nor U26201 (N_26201,N_24441,N_25270);
and U26202 (N_26202,N_25268,N_24685);
and U26203 (N_26203,N_25927,N_24720);
nor U26204 (N_26204,N_24583,N_25015);
and U26205 (N_26205,N_25183,N_25503);
nand U26206 (N_26206,N_25796,N_24742);
or U26207 (N_26207,N_24248,N_25237);
and U26208 (N_26208,N_25598,N_24192);
nor U26209 (N_26209,N_25236,N_24492);
nand U26210 (N_26210,N_24885,N_24990);
or U26211 (N_26211,N_24087,N_24943);
or U26212 (N_26212,N_24621,N_25767);
nor U26213 (N_26213,N_25164,N_24517);
nand U26214 (N_26214,N_25451,N_24240);
and U26215 (N_26215,N_25517,N_25992);
and U26216 (N_26216,N_24187,N_25555);
and U26217 (N_26217,N_24280,N_24363);
nor U26218 (N_26218,N_25975,N_25107);
or U26219 (N_26219,N_25336,N_25248);
nand U26220 (N_26220,N_25810,N_25637);
xor U26221 (N_26221,N_24863,N_24693);
nand U26222 (N_26222,N_25197,N_25782);
nand U26223 (N_26223,N_25430,N_24197);
xor U26224 (N_26224,N_24416,N_25512);
nor U26225 (N_26225,N_25129,N_24638);
and U26226 (N_26226,N_25249,N_24409);
and U26227 (N_26227,N_24684,N_24832);
xnor U26228 (N_26228,N_24571,N_24296);
xnor U26229 (N_26229,N_25463,N_25641);
nand U26230 (N_26230,N_25470,N_24870);
and U26231 (N_26231,N_25418,N_25802);
and U26232 (N_26232,N_24221,N_24352);
and U26233 (N_26233,N_25116,N_25670);
or U26234 (N_26234,N_24932,N_24449);
or U26235 (N_26235,N_25754,N_25238);
or U26236 (N_26236,N_25411,N_24746);
and U26237 (N_26237,N_24668,N_24830);
nor U26238 (N_26238,N_24887,N_24371);
and U26239 (N_26239,N_24155,N_25703);
nor U26240 (N_26240,N_25885,N_25640);
nand U26241 (N_26241,N_24118,N_25607);
or U26242 (N_26242,N_25901,N_25198);
xor U26243 (N_26243,N_24506,N_24178);
nor U26244 (N_26244,N_24923,N_25914);
or U26245 (N_26245,N_25632,N_25458);
nand U26246 (N_26246,N_25872,N_25654);
nand U26247 (N_26247,N_24395,N_24902);
or U26248 (N_26248,N_25877,N_24353);
xnor U26249 (N_26249,N_25938,N_24458);
nor U26250 (N_26250,N_25867,N_24726);
nor U26251 (N_26251,N_24645,N_25275);
and U26252 (N_26252,N_25408,N_25161);
nor U26253 (N_26253,N_25821,N_25294);
and U26254 (N_26254,N_25731,N_24753);
xnor U26255 (N_26255,N_25419,N_24334);
or U26256 (N_26256,N_25761,N_25205);
nand U26257 (N_26257,N_25595,N_24354);
xnor U26258 (N_26258,N_25535,N_24117);
xor U26259 (N_26259,N_24080,N_24654);
xnor U26260 (N_26260,N_24626,N_24717);
xor U26261 (N_26261,N_24088,N_25452);
nor U26262 (N_26262,N_25013,N_25083);
xor U26263 (N_26263,N_25273,N_24700);
nor U26264 (N_26264,N_24205,N_24612);
nor U26265 (N_26265,N_24660,N_25287);
nand U26266 (N_26266,N_25662,N_25064);
or U26267 (N_26267,N_24013,N_25469);
xnor U26268 (N_26268,N_25909,N_25942);
or U26269 (N_26269,N_24260,N_24574);
nor U26270 (N_26270,N_24915,N_24301);
nand U26271 (N_26271,N_25413,N_25728);
or U26272 (N_26272,N_25047,N_25225);
nor U26273 (N_26273,N_25321,N_25732);
nand U26274 (N_26274,N_24875,N_25133);
or U26275 (N_26275,N_25724,N_24904);
or U26276 (N_26276,N_25322,N_25565);
nand U26277 (N_26277,N_24896,N_24273);
xor U26278 (N_26278,N_25768,N_24956);
xnor U26279 (N_26279,N_25130,N_25524);
xor U26280 (N_26280,N_24982,N_24357);
or U26281 (N_26281,N_25515,N_25185);
nor U26282 (N_26282,N_24844,N_24581);
or U26283 (N_26283,N_24639,N_25863);
and U26284 (N_26284,N_25137,N_24519);
xor U26285 (N_26285,N_24543,N_24104);
or U26286 (N_26286,N_24237,N_24023);
nand U26287 (N_26287,N_24478,N_24776);
nand U26288 (N_26288,N_25981,N_24236);
nand U26289 (N_26289,N_25550,N_25846);
nand U26290 (N_26290,N_24392,N_25174);
nand U26291 (N_26291,N_24365,N_24651);
xor U26292 (N_26292,N_24948,N_24284);
or U26293 (N_26293,N_24794,N_25786);
xor U26294 (N_26294,N_25939,N_24873);
or U26295 (N_26295,N_24689,N_24799);
xnor U26296 (N_26296,N_25769,N_25121);
or U26297 (N_26297,N_24589,N_24228);
and U26298 (N_26298,N_24787,N_25965);
or U26299 (N_26299,N_24398,N_24928);
nor U26300 (N_26300,N_24405,N_25209);
nor U26301 (N_26301,N_24984,N_24128);
xor U26302 (N_26302,N_25167,N_24960);
nor U26303 (N_26303,N_24143,N_24643);
and U26304 (N_26304,N_25274,N_24078);
and U26305 (N_26305,N_25593,N_25097);
nor U26306 (N_26306,N_25406,N_24866);
xor U26307 (N_26307,N_25698,N_25720);
and U26308 (N_26308,N_24183,N_25166);
nand U26309 (N_26309,N_24811,N_25379);
or U26310 (N_26310,N_24145,N_24411);
xnor U26311 (N_26311,N_24122,N_24326);
nor U26312 (N_26312,N_25073,N_25545);
xnor U26313 (N_26313,N_25695,N_24368);
xnor U26314 (N_26314,N_25639,N_25737);
and U26315 (N_26315,N_24337,N_25424);
nand U26316 (N_26316,N_25357,N_25284);
and U26317 (N_26317,N_25485,N_25465);
xnor U26318 (N_26318,N_25043,N_24101);
nor U26319 (N_26319,N_25189,N_24467);
nor U26320 (N_26320,N_25660,N_24482);
and U26321 (N_26321,N_24508,N_24015);
and U26322 (N_26322,N_24793,N_24327);
xor U26323 (N_26323,N_25081,N_25615);
xor U26324 (N_26324,N_24862,N_24730);
nand U26325 (N_26325,N_25563,N_24051);
nand U26326 (N_26326,N_25777,N_25498);
nor U26327 (N_26327,N_24919,N_24295);
nand U26328 (N_26328,N_24100,N_25770);
and U26329 (N_26329,N_25678,N_24359);
xor U26330 (N_26330,N_25435,N_25749);
nand U26331 (N_26331,N_25890,N_25330);
or U26332 (N_26332,N_24291,N_24318);
nor U26333 (N_26333,N_24833,N_25544);
and U26334 (N_26334,N_24997,N_25354);
nand U26335 (N_26335,N_25745,N_25918);
or U26336 (N_26336,N_24681,N_24930);
xor U26337 (N_26337,N_25940,N_24406);
or U26338 (N_26338,N_24032,N_25491);
nand U26339 (N_26339,N_24370,N_24941);
or U26340 (N_26340,N_24172,N_24790);
nor U26341 (N_26341,N_24330,N_24620);
nand U26342 (N_26342,N_25833,N_24180);
or U26343 (N_26343,N_24329,N_25172);
xor U26344 (N_26344,N_25562,N_24929);
and U26345 (N_26345,N_25571,N_25257);
or U26346 (N_26346,N_25029,N_25893);
nor U26347 (N_26347,N_25366,N_24688);
xnor U26348 (N_26348,N_25501,N_24358);
xor U26349 (N_26349,N_24175,N_25705);
or U26350 (N_26350,N_25570,N_24464);
and U26351 (N_26351,N_24632,N_24868);
xnor U26352 (N_26352,N_24486,N_24336);
nor U26353 (N_26353,N_24891,N_25903);
nor U26354 (N_26354,N_25056,N_25668);
xnor U26355 (N_26355,N_25828,N_24860);
and U26356 (N_26356,N_24033,N_24292);
nor U26357 (N_26357,N_25602,N_24189);
nand U26358 (N_26358,N_25809,N_25860);
or U26359 (N_26359,N_24293,N_25212);
nand U26360 (N_26360,N_24973,N_24496);
nor U26361 (N_26361,N_25577,N_25648);
and U26362 (N_26362,N_24373,N_25296);
nor U26363 (N_26363,N_24342,N_25829);
xnor U26364 (N_26364,N_25352,N_25479);
xnor U26365 (N_26365,N_25407,N_25163);
nor U26366 (N_26366,N_25612,N_25684);
nor U26367 (N_26367,N_25496,N_25936);
or U26368 (N_26368,N_25362,N_24022);
xnor U26369 (N_26369,N_24125,N_25666);
nor U26370 (N_26370,N_24403,N_24126);
or U26371 (N_26371,N_24159,N_25084);
or U26372 (N_26372,N_24419,N_25588);
nor U26373 (N_26373,N_24339,N_25036);
or U26374 (N_26374,N_25392,N_24098);
nor U26375 (N_26375,N_24261,N_24944);
xor U26376 (N_26376,N_24439,N_24749);
xor U26377 (N_26377,N_25929,N_24810);
or U26378 (N_26378,N_25683,N_25300);
nand U26379 (N_26379,N_24949,N_24822);
xor U26380 (N_26380,N_24750,N_24091);
or U26381 (N_26381,N_24488,N_25553);
nor U26382 (N_26382,N_25928,N_25063);
nand U26383 (N_26383,N_25947,N_25144);
nor U26384 (N_26384,N_24831,N_24287);
xnor U26385 (N_26385,N_24038,N_25280);
nand U26386 (N_26386,N_24060,N_24674);
nand U26387 (N_26387,N_25669,N_25539);
nand U26388 (N_26388,N_25264,N_25090);
xnor U26389 (N_26389,N_25978,N_24076);
or U26390 (N_26390,N_25486,N_24055);
nand U26391 (N_26391,N_24664,N_25168);
nand U26392 (N_26392,N_25045,N_24484);
nand U26393 (N_26393,N_24375,N_25904);
or U26394 (N_26394,N_24223,N_25286);
nor U26395 (N_26395,N_24382,N_25783);
nand U26396 (N_26396,N_24766,N_24445);
and U26397 (N_26397,N_25546,N_24255);
and U26398 (N_26398,N_24791,N_24277);
or U26399 (N_26399,N_24272,N_24857);
xor U26400 (N_26400,N_25726,N_25608);
nand U26401 (N_26401,N_24418,N_25659);
nor U26402 (N_26402,N_24608,N_24181);
or U26403 (N_26403,N_25943,N_25825);
and U26404 (N_26404,N_24968,N_24906);
nor U26405 (N_26405,N_24652,N_25138);
xnor U26406 (N_26406,N_24779,N_24425);
nor U26407 (N_26407,N_25889,N_24942);
or U26408 (N_26408,N_25751,N_25649);
xor U26409 (N_26409,N_24438,N_24430);
nor U26410 (N_26410,N_25437,N_25568);
nand U26411 (N_26411,N_25958,N_24317);
nand U26412 (N_26412,N_24547,N_24321);
or U26413 (N_26413,N_24850,N_25663);
nor U26414 (N_26414,N_25688,N_25369);
or U26415 (N_26415,N_24423,N_24135);
xor U26416 (N_26416,N_25128,N_25412);
or U26417 (N_26417,N_24931,N_25271);
nand U26418 (N_26418,N_24754,N_25488);
or U26419 (N_26419,N_25306,N_24657);
nor U26420 (N_26420,N_25446,N_24435);
nor U26421 (N_26421,N_24732,N_24288);
nand U26422 (N_26422,N_24920,N_25566);
nor U26423 (N_26423,N_25499,N_24962);
and U26424 (N_26424,N_25482,N_24650);
and U26425 (N_26425,N_25949,N_24884);
and U26426 (N_26426,N_25032,N_25653);
nand U26427 (N_26427,N_24842,N_25655);
or U26428 (N_26428,N_25921,N_24933);
nor U26429 (N_26429,N_25151,N_25233);
and U26430 (N_26430,N_24950,N_25256);
or U26431 (N_26431,N_25279,N_24247);
xnor U26432 (N_26432,N_25743,N_25826);
or U26433 (N_26433,N_24988,N_24839);
xnor U26434 (N_26434,N_24220,N_24275);
nand U26435 (N_26435,N_25532,N_24062);
or U26436 (N_26436,N_25298,N_25551);
nand U26437 (N_26437,N_25834,N_24227);
xnor U26438 (N_26438,N_25039,N_24745);
xor U26439 (N_26439,N_25299,N_24234);
or U26440 (N_26440,N_24335,N_24854);
xnor U26441 (N_26441,N_24537,N_25991);
or U26442 (N_26442,N_25016,N_25173);
xor U26443 (N_26443,N_24256,N_24026);
or U26444 (N_26444,N_24858,N_25376);
or U26445 (N_26445,N_24510,N_25861);
xor U26446 (N_26446,N_25755,N_25721);
or U26447 (N_26447,N_25421,N_25787);
nand U26448 (N_26448,N_25394,N_25552);
xnor U26449 (N_26449,N_25908,N_25434);
or U26450 (N_26450,N_25934,N_25667);
and U26451 (N_26451,N_24266,N_24985);
or U26452 (N_26452,N_24555,N_25110);
or U26453 (N_26453,N_24549,N_24042);
xnor U26454 (N_26454,N_25191,N_24231);
nand U26455 (N_26455,N_24061,N_24577);
xor U26456 (N_26456,N_24491,N_25337);
or U26457 (N_26457,N_25373,N_25781);
or U26458 (N_26458,N_24444,N_24047);
nor U26459 (N_26459,N_24969,N_24030);
xor U26460 (N_26460,N_24739,N_24797);
xor U26461 (N_26461,N_24807,N_24755);
or U26462 (N_26462,N_24154,N_25219);
nand U26463 (N_26463,N_25948,N_24961);
and U26464 (N_26464,N_25589,N_25390);
xnor U26465 (N_26465,N_24559,N_25672);
xnor U26466 (N_26466,N_24166,N_25812);
xnor U26467 (N_26467,N_25510,N_25710);
xnor U26468 (N_26468,N_25348,N_24136);
and U26469 (N_26469,N_24193,N_25311);
xnor U26470 (N_26470,N_24217,N_24113);
nand U26471 (N_26471,N_24509,N_25913);
nand U26472 (N_26472,N_24804,N_25338);
xor U26473 (N_26473,N_24138,N_24721);
nand U26474 (N_26474,N_25201,N_25801);
nand U26475 (N_26475,N_25734,N_25089);
nor U26476 (N_26476,N_25331,N_25175);
nand U26477 (N_26477,N_25832,N_24760);
xor U26478 (N_26478,N_24921,N_25554);
or U26479 (N_26479,N_25633,N_24412);
and U26480 (N_26480,N_24963,N_24007);
xnor U26481 (N_26481,N_25897,N_24846);
and U26482 (N_26482,N_24640,N_25134);
nand U26483 (N_26483,N_25924,N_25229);
nand U26484 (N_26484,N_24081,N_25873);
xnor U26485 (N_26485,N_25643,N_25974);
nor U26486 (N_26486,N_25690,N_25292);
xor U26487 (N_26487,N_24938,N_24625);
xor U26488 (N_26488,N_24324,N_24037);
and U26489 (N_26489,N_25746,N_24550);
xor U26490 (N_26490,N_24258,N_25650);
nand U26491 (N_26491,N_25953,N_25594);
nor U26492 (N_26492,N_24629,N_24882);
nor U26493 (N_26493,N_25310,N_24436);
nor U26494 (N_26494,N_25289,N_24202);
nand U26495 (N_26495,N_25883,N_24975);
xor U26496 (N_26496,N_24747,N_24170);
nor U26497 (N_26497,N_25169,N_24597);
nor U26498 (N_26498,N_24530,N_25467);
nand U26499 (N_26499,N_24343,N_25117);
and U26500 (N_26500,N_25537,N_24927);
and U26501 (N_26501,N_25687,N_24598);
and U26502 (N_26502,N_24708,N_25816);
and U26503 (N_26503,N_25077,N_25489);
xor U26504 (N_26504,N_24111,N_24270);
nand U26505 (N_26505,N_25207,N_24137);
nand U26506 (N_26506,N_24707,N_25022);
and U26507 (N_26507,N_24386,N_25963);
or U26508 (N_26508,N_24901,N_24498);
xnor U26509 (N_26509,N_25044,N_24724);
nand U26510 (N_26510,N_25410,N_24782);
nand U26511 (N_26511,N_24567,N_24910);
and U26512 (N_26512,N_24089,N_25037);
nor U26513 (N_26513,N_24821,N_24529);
nor U26514 (N_26514,N_25335,N_24966);
xor U26515 (N_26515,N_24798,N_24723);
or U26516 (N_26516,N_25533,N_25954);
nand U26517 (N_26517,N_25396,N_25441);
nor U26518 (N_26518,N_25747,N_25473);
nor U26519 (N_26519,N_24515,N_25774);
or U26520 (N_26520,N_25661,N_25578);
or U26521 (N_26521,N_25797,N_24788);
or U26522 (N_26522,N_25520,N_24840);
nand U26523 (N_26523,N_25853,N_25827);
xnor U26524 (N_26524,N_25131,N_24695);
and U26525 (N_26525,N_24083,N_24501);
nand U26526 (N_26526,N_24222,N_25538);
and U26527 (N_26527,N_24743,N_25193);
xnor U26528 (N_26528,N_24770,N_25182);
and U26529 (N_26529,N_24049,N_24678);
and U26530 (N_26530,N_25142,N_25773);
nand U26531 (N_26531,N_25179,N_24466);
xnor U26532 (N_26532,N_24828,N_24795);
nand U26533 (N_26533,N_25026,N_25076);
nand U26534 (N_26534,N_24360,N_24511);
nand U26535 (N_26535,N_24841,N_24474);
or U26536 (N_26536,N_25824,N_25360);
xnor U26537 (N_26537,N_25752,N_24622);
nor U26538 (N_26538,N_24572,N_25125);
or U26539 (N_26539,N_25180,N_24763);
or U26540 (N_26540,N_24711,N_25214);
nor U26541 (N_26541,N_25849,N_25034);
or U26542 (N_26542,N_24401,N_24397);
or U26543 (N_26543,N_25440,N_24319);
xor U26544 (N_26544,N_24112,N_24132);
nand U26545 (N_26545,N_24413,N_25941);
nor U26546 (N_26546,N_25375,N_24294);
and U26547 (N_26547,N_25425,N_24211);
and U26548 (N_26548,N_24157,N_25266);
nand U26549 (N_26549,N_25057,N_24552);
and U26550 (N_26550,N_25711,N_25933);
xnor U26551 (N_26551,N_25780,N_24428);
and U26552 (N_26552,N_24513,N_24340);
and U26553 (N_26553,N_24607,N_25971);
and U26554 (N_26554,N_24729,N_25626);
xor U26555 (N_26555,N_24024,N_25508);
xor U26556 (N_26556,N_25252,N_25339);
nand U26557 (N_26557,N_24393,N_24179);
xnor U26558 (N_26558,N_25126,N_25028);
nand U26559 (N_26559,N_24591,N_24769);
or U26560 (N_26560,N_25844,N_24311);
xnor U26561 (N_26561,N_24599,N_24865);
nand U26562 (N_26562,N_25997,N_25031);
xnor U26563 (N_26563,N_24476,N_24084);
or U26564 (N_26564,N_25609,N_24837);
nand U26565 (N_26565,N_25647,N_25744);
and U26566 (N_26566,N_25917,N_25382);
nand U26567 (N_26567,N_24903,N_25968);
or U26568 (N_26568,N_25658,N_24817);
xor U26569 (N_26569,N_24099,N_24587);
or U26570 (N_26570,N_25124,N_24463);
or U26571 (N_26571,N_24816,N_25464);
or U26572 (N_26572,N_25216,N_25511);
or U26573 (N_26573,N_25224,N_25223);
and U26574 (N_26574,N_24633,N_24036);
nor U26575 (N_26575,N_24440,N_25707);
nand U26576 (N_26576,N_24457,N_24586);
or U26577 (N_26577,N_25915,N_25240);
nand U26578 (N_26578,N_24704,N_24278);
and U26579 (N_26579,N_25575,N_24699);
xor U26580 (N_26580,N_24618,N_25492);
nand U26581 (N_26581,N_24610,N_24422);
and U26582 (N_26582,N_25631,N_24524);
nand U26583 (N_26583,N_25059,N_25247);
xnor U26584 (N_26584,N_24263,N_24523);
nand U26585 (N_26585,N_24709,N_24127);
and U26586 (N_26586,N_25961,N_25312);
and U26587 (N_26587,N_25477,N_25966);
nor U26588 (N_26588,N_25231,N_24826);
and U26589 (N_26589,N_24977,N_25696);
and U26590 (N_26590,N_25874,N_24558);
nand U26591 (N_26591,N_24257,N_25694);
and U26592 (N_26592,N_24905,N_24983);
or U26593 (N_26593,N_24451,N_25276);
nor U26594 (N_26594,N_25789,N_25053);
nor U26595 (N_26595,N_24054,N_25309);
nand U26596 (N_26596,N_25364,N_24594);
nor U26597 (N_26597,N_25493,N_25114);
nor U26598 (N_26598,N_24922,N_25319);
xnor U26599 (N_26599,N_25907,N_25599);
nand U26600 (N_26600,N_25304,N_24043);
or U26601 (N_26601,N_24648,N_24503);
or U26602 (N_26602,N_25261,N_24947);
and U26603 (N_26603,N_25251,N_24461);
nand U26604 (N_26604,N_24725,N_25353);
nand U26605 (N_26605,N_25344,N_24546);
xnor U26606 (N_26606,N_25067,N_24774);
nor U26607 (N_26607,N_25886,N_24315);
nor U26608 (N_26608,N_25091,N_25505);
or U26609 (N_26609,N_25945,N_25951);
and U26610 (N_26610,N_24972,N_24454);
nor U26611 (N_26611,N_25686,N_25345);
nand U26612 (N_26612,N_24443,N_24453);
nor U26613 (N_26613,N_24121,N_25652);
and U26614 (N_26614,N_24264,N_24852);
nand U26615 (N_26615,N_24344,N_25226);
and U26616 (N_26616,N_24316,N_25906);
xnor U26617 (N_26617,N_25629,N_24999);
nor U26618 (N_26618,N_24727,N_24381);
and U26619 (N_26619,N_24864,N_25080);
or U26620 (N_26620,N_24838,N_24532);
and U26621 (N_26621,N_25916,N_24265);
nor U26622 (N_26622,N_25227,N_25475);
or U26623 (N_26623,N_24242,N_24566);
or U26624 (N_26624,N_24011,N_25095);
or U26625 (N_26625,N_24981,N_25105);
and U26626 (N_26626,N_25657,N_25449);
xor U26627 (N_26627,N_24102,N_25625);
or U26628 (N_26628,N_24756,N_25840);
nor U26629 (N_26629,N_24542,N_24718);
nor U26630 (N_26630,N_25764,N_24092);
and U26631 (N_26631,N_24536,N_24388);
nor U26632 (N_26632,N_24843,N_25313);
nor U26633 (N_26633,N_24825,N_24954);
xor U26634 (N_26634,N_24204,N_24377);
xor U26635 (N_26635,N_25714,N_24346);
nand U26636 (N_26636,N_25507,N_24913);
xnor U26637 (N_26637,N_25269,N_24029);
or U26638 (N_26638,N_24883,N_24761);
or U26639 (N_26639,N_24462,N_24050);
or U26640 (N_26640,N_25153,N_25478);
xnor U26641 (N_26641,N_25618,N_25634);
or U26642 (N_26642,N_24703,N_25514);
nor U26643 (N_26643,N_25221,N_24103);
or U26644 (N_26644,N_25572,N_24331);
nor U26645 (N_26645,N_24452,N_25718);
and U26646 (N_26646,N_25619,N_24012);
and U26647 (N_26647,N_24086,N_25892);
nor U26648 (N_26648,N_25817,N_25122);
and U26649 (N_26649,N_25355,N_25692);
or U26650 (N_26650,N_24521,N_24731);
nand U26651 (N_26651,N_25341,N_25586);
or U26652 (N_26652,N_24073,N_25960);
xnor U26653 (N_26653,N_25232,N_24195);
nand U26654 (N_26654,N_25204,N_25729);
nor U26655 (N_26655,N_24469,N_24959);
or U26656 (N_26656,N_24151,N_25534);
nor U26657 (N_26657,N_25455,N_24259);
nor U26658 (N_26658,N_25871,N_25561);
xor U26659 (N_26659,N_24489,N_24888);
and U26660 (N_26660,N_24207,N_25127);
nor U26661 (N_26661,N_24848,N_24176);
and U26662 (N_26662,N_24045,N_24851);
or U26663 (N_26663,N_25108,N_24836);
or U26664 (N_26664,N_24814,N_25888);
and U26665 (N_26665,N_25556,N_24019);
nand U26666 (N_26666,N_24512,N_25291);
nor U26667 (N_26667,N_24067,N_25436);
nor U26668 (N_26668,N_24595,N_24642);
nand U26669 (N_26669,N_25487,N_25697);
or U26670 (N_26670,N_25504,N_24106);
nor U26671 (N_26671,N_24853,N_25471);
and U26672 (N_26672,N_24737,N_25019);
or U26673 (N_26673,N_24468,N_25146);
nand U26674 (N_26674,N_25935,N_25476);
xnor U26675 (N_26675,N_24534,N_24472);
nand U26676 (N_26676,N_24953,N_24995);
xor U26677 (N_26677,N_24653,N_24861);
and U26678 (N_26678,N_24562,N_24813);
or U26679 (N_26679,N_25590,N_24394);
or U26680 (N_26680,N_25931,N_25866);
xnor U26681 (N_26681,N_24876,N_24680);
and U26682 (N_26682,N_24611,N_24568);
or U26683 (N_26683,N_24328,N_24169);
nor U26684 (N_26684,N_24052,N_25187);
nor U26685 (N_26685,N_25359,N_24998);
xnor U26686 (N_26686,N_25211,N_25854);
or U26687 (N_26687,N_24072,N_25217);
xnor U26688 (N_26688,N_24399,N_24751);
nor U26689 (N_26689,N_24206,N_25856);
nand U26690 (N_26690,N_25741,N_25750);
or U26691 (N_26691,N_25984,N_25004);
or U26692 (N_26692,N_24214,N_24348);
nor U26693 (N_26693,N_25753,N_24003);
xor U26694 (N_26694,N_24070,N_24722);
nand U26695 (N_26695,N_25950,N_25862);
nor U26696 (N_26696,N_24314,N_25838);
and U26697 (N_26697,N_24874,N_25035);
and U26698 (N_26698,N_24208,N_25215);
and U26699 (N_26699,N_25259,N_25461);
nand U26700 (N_26700,N_25380,N_24710);
nor U26701 (N_26701,N_24580,N_25980);
nor U26702 (N_26702,N_24827,N_24588);
and U26703 (N_26703,N_24970,N_24188);
and U26704 (N_26704,N_24792,N_25447);
and U26705 (N_26705,N_24683,N_25195);
nand U26706 (N_26706,N_25431,N_24186);
and U26707 (N_26707,N_24174,N_24603);
or U26708 (N_26708,N_25154,N_24165);
and U26709 (N_26709,N_25072,N_24387);
and U26710 (N_26710,N_25260,N_24448);
or U26711 (N_26711,N_24735,N_25143);
nor U26712 (N_26712,N_25263,N_25689);
nand U26713 (N_26713,N_25239,N_24900);
or U26714 (N_26714,N_25756,N_24819);
or U26715 (N_26715,N_25993,N_24298);
nor U26716 (N_26716,N_25988,N_25576);
nand U26717 (N_26717,N_24200,N_25058);
xnor U26718 (N_26718,N_25900,N_24303);
or U26719 (N_26719,N_24241,N_24031);
or U26720 (N_26720,N_25795,N_25316);
xor U26721 (N_26721,N_24156,N_25055);
nand U26722 (N_26722,N_24628,N_25591);
nor U26723 (N_26723,N_25218,N_25884);
xnor U26724 (N_26724,N_25210,N_25645);
nand U26725 (N_26725,N_25691,N_25295);
xor U26726 (N_26726,N_25794,N_24417);
xnor U26727 (N_26727,N_24216,N_25448);
nor U26728 (N_26728,N_24624,N_24119);
nor U26729 (N_26729,N_24233,N_25682);
and U26730 (N_26730,N_25020,N_25716);
xor U26731 (N_26731,N_24935,N_24565);
nor U26732 (N_26732,N_25062,N_25617);
nand U26733 (N_26733,N_24596,N_24018);
or U26734 (N_26734,N_25962,N_25621);
or U26735 (N_26735,N_24160,N_25671);
and U26736 (N_26736,N_25094,N_24741);
nand U26737 (N_26737,N_25531,N_25054);
and U26738 (N_26738,N_24911,N_25830);
xor U26739 (N_26739,N_25808,N_25527);
nand U26740 (N_26740,N_25070,N_24131);
nor U26741 (N_26741,N_24925,N_24665);
and U26742 (N_26742,N_25822,N_24593);
or U26743 (N_26743,N_25601,N_25000);
and U26744 (N_26744,N_25973,N_25148);
nor U26745 (N_26745,N_25342,N_25203);
and U26746 (N_26746,N_24495,N_25162);
xor U26747 (N_26747,N_24634,N_25220);
nand U26748 (N_26748,N_24459,N_24473);
nand U26749 (N_26749,N_24229,N_24716);
or U26750 (N_26750,N_25326,N_24249);
xor U26751 (N_26751,N_24322,N_24649);
nand U26752 (N_26752,N_25042,N_24702);
nor U26753 (N_26753,N_24276,N_24663);
nand U26754 (N_26754,N_24041,N_24976);
or U26755 (N_26755,N_25735,N_25922);
or U26756 (N_26756,N_25522,N_25804);
nor U26757 (N_26757,N_25946,N_24300);
and U26758 (N_26758,N_24656,N_24039);
or U26759 (N_26759,N_24937,N_25899);
nand U26760 (N_26760,N_25727,N_24433);
xnor U26761 (N_26761,N_25145,N_25800);
nand U26762 (N_26762,N_25358,N_25881);
xor U26763 (N_26763,N_24177,N_25813);
xnor U26764 (N_26764,N_24805,N_25397);
nor U26765 (N_26765,N_24815,N_24494);
xnor U26766 (N_26766,N_25791,N_25420);
and U26767 (N_26767,N_24758,N_24897);
or U26768 (N_26768,N_24372,N_25775);
or U26769 (N_26769,N_25926,N_24090);
or U26770 (N_26770,N_24201,N_24912);
nand U26771 (N_26771,N_25700,N_25334);
and U26772 (N_26772,N_25160,N_24824);
nor U26773 (N_26773,N_24364,N_25835);
and U26774 (N_26774,N_25605,N_25887);
nor U26775 (N_26775,N_25820,N_24835);
xor U26776 (N_26776,N_25305,N_25192);
nor U26777 (N_26777,N_24194,N_24109);
xnor U26778 (N_26778,N_24144,N_24771);
nand U26779 (N_26779,N_24800,N_25159);
and U26780 (N_26780,N_24573,N_24246);
nand U26781 (N_26781,N_24849,N_24845);
xnor U26782 (N_26782,N_24304,N_25017);
nand U26783 (N_26783,N_24376,N_25880);
nor U26784 (N_26784,N_24518,N_24940);
and U26785 (N_26785,N_24410,N_24232);
or U26786 (N_26786,N_24107,N_25006);
and U26787 (N_26787,N_24347,N_24414);
nand U26788 (N_26788,N_25713,N_25636);
nor U26789 (N_26789,N_25875,N_25170);
nor U26790 (N_26790,N_25372,N_24994);
or U26791 (N_26791,N_24123,N_25847);
or U26792 (N_26792,N_24691,N_25990);
xnor U26793 (N_26793,N_24485,N_25060);
xnor U26794 (N_26794,N_24380,N_25361);
and U26795 (N_26795,N_24146,N_25656);
nand U26796 (N_26796,N_24516,N_24010);
or U26797 (N_26797,N_24390,N_24168);
and U26798 (N_26798,N_25096,N_24535);
nor U26799 (N_26799,N_24158,N_24781);
xnor U26800 (N_26800,N_24333,N_24630);
nor U26801 (N_26801,N_24690,N_24914);
nor U26802 (N_26802,N_24481,N_25075);
nand U26803 (N_26803,N_25061,N_24701);
or U26804 (N_26804,N_25426,N_24796);
nor U26805 (N_26805,N_24493,N_25068);
and U26806 (N_26806,N_24483,N_25814);
nor U26807 (N_26807,N_25283,N_24802);
nor U26808 (N_26808,N_24971,N_25171);
or U26809 (N_26809,N_24056,N_25635);
nand U26810 (N_26810,N_25427,N_24974);
nand U26811 (N_26811,N_25318,N_24431);
nand U26812 (N_26812,N_24021,N_24785);
or U26813 (N_26813,N_25730,N_25878);
nor U26814 (N_26814,N_24893,N_24733);
xor U26815 (N_26815,N_24762,N_25325);
or U26816 (N_26816,N_24313,N_25757);
xor U26817 (N_26817,N_25558,N_24548);
or U26818 (N_26818,N_25704,N_24666);
and U26819 (N_26819,N_24908,N_25136);
xor U26820 (N_26820,N_25340,N_25585);
nor U26821 (N_26821,N_25104,N_24385);
nand U26822 (N_26822,N_25564,N_25518);
xnor U26823 (N_26823,N_24499,N_25186);
nand U26824 (N_26824,N_25582,N_25141);
xor U26825 (N_26825,N_24002,N_24384);
xnor U26826 (N_26826,N_24812,N_25370);
nand U26827 (N_26827,N_25024,N_25281);
nor U26828 (N_26828,N_24623,N_24066);
or U26829 (N_26829,N_25443,N_25919);
or U26830 (N_26830,N_25196,N_24679);
xor U26831 (N_26831,N_24164,N_25484);
nand U26832 (N_26832,N_24082,N_24637);
nand U26833 (N_26833,N_24014,N_25778);
or U26834 (N_26834,N_24898,N_25627);
and U26835 (N_26835,N_25679,N_25855);
nand U26836 (N_26836,N_25103,N_25429);
xnor U26837 (N_26837,N_25258,N_24212);
nand U26838 (N_26838,N_24141,N_24847);
nand U26839 (N_26839,N_25001,N_24378);
nor U26840 (N_26840,N_25112,N_24374);
and U26841 (N_26841,N_24025,N_24759);
or U26842 (N_26842,N_24881,N_24057);
and U26843 (N_26843,N_25851,N_24698);
or U26844 (N_26844,N_24446,N_24527);
or U26845 (N_26845,N_25242,N_25976);
xnor U26846 (N_26846,N_25613,N_25674);
and U26847 (N_26847,N_25417,N_24163);
nor U26848 (N_26848,N_24600,N_24635);
nand U26849 (N_26849,N_24028,N_25739);
and U26850 (N_26850,N_24712,N_24757);
or U26851 (N_26851,N_25547,N_24252);
nand U26852 (N_26852,N_24818,N_24545);
xor U26853 (N_26853,N_25450,N_24065);
xor U26854 (N_26854,N_24046,N_24662);
or U26855 (N_26855,N_25374,N_25423);
nand U26856 (N_26856,N_25038,N_24404);
xor U26857 (N_26857,N_24945,N_24124);
or U26858 (N_26858,N_25784,N_25194);
nand U26859 (N_26859,N_24150,N_25481);
or U26860 (N_26860,N_25630,N_24479);
nor U26861 (N_26861,N_24714,N_24892);
xnor U26862 (N_26862,N_25857,N_25584);
and U26863 (N_26863,N_25014,N_25466);
nor U26864 (N_26864,N_25030,N_24987);
or U26865 (N_26865,N_24074,N_24728);
and U26866 (N_26866,N_24407,N_25955);
nor U26867 (N_26867,N_24783,N_25139);
xnor U26868 (N_26868,N_25100,N_24670);
or U26869 (N_26869,N_25023,N_25003);
xnor U26870 (N_26870,N_25530,N_25388);
nand U26871 (N_26871,N_24310,N_24471);
or U26872 (N_26872,N_24108,N_25646);
xnor U26873 (N_26873,N_25046,N_25559);
or U26874 (N_26874,N_24383,N_25005);
or U26875 (N_26875,N_24068,N_25409);
nor U26876 (N_26876,N_24778,N_25925);
nor U26877 (N_26877,N_25779,N_25414);
or U26878 (N_26878,N_24367,N_24153);
nand U26879 (N_26879,N_24139,N_24116);
nor U26880 (N_26880,N_24389,N_25444);
xor U26881 (N_26881,N_25456,N_25898);
nor U26882 (N_26882,N_24557,N_24886);
nand U26883 (N_26883,N_25843,N_24362);
or U26884 (N_26884,N_25333,N_25587);
xnor U26885 (N_26885,N_25677,N_24283);
and U26886 (N_26886,N_24609,N_24182);
nor U26887 (N_26887,N_24934,N_24661);
and U26888 (N_26888,N_25158,N_25098);
nand U26889 (N_26889,N_24575,N_24706);
nor U26890 (N_26890,N_24734,N_25969);
and U26891 (N_26891,N_24302,N_24867);
xor U26892 (N_26892,N_25282,N_25041);
xnor U26893 (N_26893,N_25184,N_24421);
xnor U26894 (N_26894,N_25385,N_24001);
nor U26895 (N_26895,N_25315,N_24806);
nor U26896 (N_26896,N_25480,N_25805);
or U26897 (N_26897,N_25381,N_24064);
or U26898 (N_26898,N_25109,N_25610);
nand U26899 (N_26899,N_25021,N_24040);
or U26900 (N_26900,N_25328,N_25693);
or U26901 (N_26901,N_25790,N_25766);
nand U26902 (N_26902,N_24487,N_25806);
and U26903 (N_26903,N_24286,N_24563);
xor U26904 (N_26904,N_24617,N_25540);
nand U26905 (N_26905,N_24426,N_24219);
nand U26906 (N_26906,N_24253,N_24379);
and U26907 (N_26907,N_25985,N_24338);
and U26908 (N_26908,N_25596,N_25823);
nand U26909 (N_26909,N_24460,N_24226);
nor U26910 (N_26910,N_24209,N_25178);
and U26911 (N_26911,N_24320,N_24740);
or U26912 (N_26912,N_25803,N_24951);
xnor U26913 (N_26913,N_24584,N_24767);
or U26914 (N_26914,N_25868,N_25119);
xor U26915 (N_26915,N_25132,N_24250);
or U26916 (N_26916,N_25664,N_24408);
and U26917 (N_26917,N_24522,N_24059);
nand U26918 (N_26918,N_24872,N_24008);
or U26919 (N_26919,N_25776,N_25176);
and U26920 (N_26920,N_24544,N_24307);
nand U26921 (N_26921,N_24616,N_24696);
or U26922 (N_26922,N_24659,N_25882);
nor U26923 (N_26923,N_25230,N_25206);
nor U26924 (N_26924,N_25301,N_24744);
and U26925 (N_26925,N_24627,N_24424);
and U26926 (N_26926,N_25356,N_24097);
nor U26927 (N_26927,N_25438,N_25740);
or U26928 (N_26928,N_24027,N_25509);
or U26929 (N_26929,N_25525,N_24786);
nor U26930 (N_26930,N_24455,N_25277);
nor U26931 (N_26931,N_24477,N_24965);
xnor U26932 (N_26932,N_24140,N_24095);
and U26933 (N_26933,N_25972,N_25622);
xor U26934 (N_26934,N_24110,N_25842);
and U26935 (N_26935,N_25208,N_25011);
nand U26936 (N_26936,N_25869,N_24415);
xor U26937 (N_26937,N_25762,N_24309);
or U26938 (N_26938,N_25085,N_25190);
nor U26939 (N_26939,N_25088,N_25228);
nor U26940 (N_26940,N_25495,N_25839);
nand U26941 (N_26941,N_25891,N_25771);
nor U26942 (N_26942,N_24936,N_25772);
nor U26943 (N_26943,N_24879,N_25314);
xor U26944 (N_26944,N_25468,N_24877);
nor U26945 (N_26945,N_24615,N_25346);
nor U26946 (N_26946,N_25837,N_25706);
nand U26947 (N_26947,N_24606,N_25712);
and U26948 (N_26948,N_25932,N_25758);
or U26949 (N_26949,N_24809,N_24079);
nor U26950 (N_26950,N_24171,N_24859);
or U26951 (N_26951,N_24564,N_24262);
xor U26952 (N_26952,N_24271,N_25959);
nand U26953 (N_26953,N_25848,N_24420);
and U26954 (N_26954,N_25106,N_25092);
nor U26955 (N_26955,N_25453,N_24077);
or U26956 (N_26956,N_24465,N_25604);
nand U26957 (N_26957,N_25685,N_25681);
nor U26958 (N_26958,N_24772,N_24504);
xor U26959 (N_26959,N_25155,N_24560);
nor U26960 (N_26960,N_24069,N_25235);
xnor U26961 (N_26961,N_24561,N_24480);
or U26962 (N_26962,N_25111,N_25519);
nand U26963 (N_26963,N_25748,N_24687);
xor U26964 (N_26964,N_25246,N_25123);
xor U26965 (N_26965,N_25066,N_24341);
nand U26966 (N_26966,N_25614,N_25673);
xnor U26967 (N_26967,N_25422,N_24894);
or U26968 (N_26968,N_24784,N_25135);
and U26969 (N_26969,N_24780,N_24456);
nand U26970 (N_26970,N_25009,N_24539);
nor U26971 (N_26971,N_24048,N_24889);
xor U26972 (N_26972,N_25152,N_25742);
nand U26973 (N_26973,N_25902,N_24134);
or U26974 (N_26974,N_24502,N_24299);
nand U26975 (N_26975,N_25542,N_25998);
nand U26976 (N_26976,N_25529,N_25349);
and U26977 (N_26977,N_25952,N_25462);
or U26978 (N_26978,N_25317,N_24926);
and U26979 (N_26979,N_24267,N_24939);
nand U26980 (N_26980,N_25799,N_24899);
nand U26981 (N_26981,N_25831,N_24094);
xor U26982 (N_26982,N_24058,N_24356);
and U26983 (N_26983,N_25398,N_24576);
or U26984 (N_26984,N_25765,N_25165);
and U26985 (N_26985,N_25324,N_25405);
nand U26986 (N_26986,N_24432,N_24009);
or U26987 (N_26987,N_24115,N_25002);
nand U26988 (N_26988,N_25490,N_24332);
nand U26989 (N_26989,N_24006,N_24658);
and U26990 (N_26990,N_24361,N_25702);
or U26991 (N_26991,N_24682,N_24525);
xnor U26992 (N_26992,N_25393,N_24020);
nand U26993 (N_26993,N_24677,N_25567);
xor U26994 (N_26994,N_24044,N_25079);
nand U26995 (N_26995,N_24619,N_25644);
or U26996 (N_26996,N_24497,N_25680);
nand U26997 (N_26997,N_25557,N_24526);
xnor U26998 (N_26998,N_24917,N_24245);
and U26999 (N_26999,N_25442,N_25378);
xnor U27000 (N_27000,N_25767,N_25070);
or U27001 (N_27001,N_24845,N_24119);
nand U27002 (N_27002,N_25319,N_25215);
and U27003 (N_27003,N_25457,N_24932);
xor U27004 (N_27004,N_25657,N_24220);
and U27005 (N_27005,N_24845,N_25051);
nor U27006 (N_27006,N_24641,N_25540);
and U27007 (N_27007,N_25703,N_24522);
nand U27008 (N_27008,N_25405,N_25422);
nand U27009 (N_27009,N_24164,N_24011);
nand U27010 (N_27010,N_25547,N_25991);
and U27011 (N_27011,N_24719,N_25869);
nand U27012 (N_27012,N_24394,N_24071);
or U27013 (N_27013,N_24708,N_24159);
xnor U27014 (N_27014,N_25769,N_25724);
and U27015 (N_27015,N_24102,N_24712);
xor U27016 (N_27016,N_24515,N_24909);
nor U27017 (N_27017,N_24059,N_25082);
or U27018 (N_27018,N_24371,N_25081);
or U27019 (N_27019,N_25454,N_24694);
nand U27020 (N_27020,N_25260,N_25749);
nand U27021 (N_27021,N_24439,N_25410);
or U27022 (N_27022,N_25640,N_25222);
nor U27023 (N_27023,N_25568,N_24832);
and U27024 (N_27024,N_25594,N_25150);
and U27025 (N_27025,N_24285,N_25646);
or U27026 (N_27026,N_24931,N_25357);
and U27027 (N_27027,N_25132,N_24806);
nor U27028 (N_27028,N_25290,N_25509);
nor U27029 (N_27029,N_24005,N_24565);
or U27030 (N_27030,N_24598,N_24091);
nor U27031 (N_27031,N_25253,N_25199);
xnor U27032 (N_27032,N_25869,N_25269);
xnor U27033 (N_27033,N_25322,N_25094);
xnor U27034 (N_27034,N_24081,N_24604);
nand U27035 (N_27035,N_24495,N_24833);
or U27036 (N_27036,N_25159,N_25230);
and U27037 (N_27037,N_25753,N_25363);
xnor U27038 (N_27038,N_25650,N_25543);
nand U27039 (N_27039,N_25770,N_25910);
and U27040 (N_27040,N_25974,N_25223);
nor U27041 (N_27041,N_25316,N_24424);
nand U27042 (N_27042,N_25646,N_25330);
xnor U27043 (N_27043,N_24872,N_24778);
xor U27044 (N_27044,N_25211,N_24838);
xor U27045 (N_27045,N_25443,N_24718);
or U27046 (N_27046,N_24832,N_24984);
nand U27047 (N_27047,N_25641,N_24361);
or U27048 (N_27048,N_25428,N_25938);
nand U27049 (N_27049,N_25646,N_25192);
or U27050 (N_27050,N_24617,N_24169);
and U27051 (N_27051,N_25863,N_24348);
and U27052 (N_27052,N_25101,N_24170);
and U27053 (N_27053,N_24140,N_24291);
and U27054 (N_27054,N_25283,N_24350);
nand U27055 (N_27055,N_24472,N_25785);
nand U27056 (N_27056,N_25901,N_25597);
and U27057 (N_27057,N_24362,N_25007);
nor U27058 (N_27058,N_25117,N_25952);
nor U27059 (N_27059,N_25710,N_25196);
and U27060 (N_27060,N_24350,N_24526);
nor U27061 (N_27061,N_25652,N_25119);
or U27062 (N_27062,N_24335,N_24328);
nor U27063 (N_27063,N_24608,N_25417);
or U27064 (N_27064,N_24441,N_25027);
and U27065 (N_27065,N_25192,N_24280);
xor U27066 (N_27066,N_25954,N_24591);
nor U27067 (N_27067,N_25686,N_24740);
xor U27068 (N_27068,N_25751,N_24989);
and U27069 (N_27069,N_24634,N_25805);
or U27070 (N_27070,N_25823,N_25972);
xor U27071 (N_27071,N_24142,N_24214);
xnor U27072 (N_27072,N_24655,N_24011);
xor U27073 (N_27073,N_24306,N_25422);
nand U27074 (N_27074,N_24004,N_25940);
and U27075 (N_27075,N_25910,N_25927);
nand U27076 (N_27076,N_25366,N_24832);
xnor U27077 (N_27077,N_24853,N_24322);
xnor U27078 (N_27078,N_25843,N_24020);
nor U27079 (N_27079,N_24638,N_25917);
and U27080 (N_27080,N_24643,N_25747);
and U27081 (N_27081,N_24698,N_25865);
xnor U27082 (N_27082,N_24253,N_24704);
and U27083 (N_27083,N_25260,N_24280);
or U27084 (N_27084,N_24889,N_25270);
or U27085 (N_27085,N_24333,N_24831);
nand U27086 (N_27086,N_25835,N_24962);
nor U27087 (N_27087,N_24572,N_25765);
nor U27088 (N_27088,N_25669,N_24754);
and U27089 (N_27089,N_24592,N_24634);
or U27090 (N_27090,N_25670,N_25891);
nor U27091 (N_27091,N_25645,N_24034);
nand U27092 (N_27092,N_24682,N_25342);
nor U27093 (N_27093,N_25751,N_25985);
nor U27094 (N_27094,N_24819,N_24912);
xor U27095 (N_27095,N_24911,N_25188);
or U27096 (N_27096,N_24410,N_25055);
nand U27097 (N_27097,N_25621,N_24168);
or U27098 (N_27098,N_24835,N_25161);
xnor U27099 (N_27099,N_24589,N_25424);
or U27100 (N_27100,N_24536,N_24610);
xnor U27101 (N_27101,N_24683,N_24370);
or U27102 (N_27102,N_24740,N_24748);
xor U27103 (N_27103,N_25480,N_24321);
or U27104 (N_27104,N_25979,N_24656);
nand U27105 (N_27105,N_24404,N_25984);
nor U27106 (N_27106,N_25234,N_25609);
nand U27107 (N_27107,N_25645,N_25109);
xor U27108 (N_27108,N_25435,N_25785);
xor U27109 (N_27109,N_25767,N_24412);
nor U27110 (N_27110,N_24064,N_25597);
nand U27111 (N_27111,N_24268,N_24006);
or U27112 (N_27112,N_25452,N_24968);
xor U27113 (N_27113,N_24386,N_24423);
xor U27114 (N_27114,N_24283,N_24883);
xnor U27115 (N_27115,N_25643,N_25892);
or U27116 (N_27116,N_24894,N_25140);
or U27117 (N_27117,N_25713,N_25321);
xor U27118 (N_27118,N_24895,N_24538);
nor U27119 (N_27119,N_24668,N_24175);
or U27120 (N_27120,N_25728,N_24177);
or U27121 (N_27121,N_25285,N_25958);
nand U27122 (N_27122,N_24243,N_25037);
and U27123 (N_27123,N_24727,N_25705);
or U27124 (N_27124,N_25657,N_24561);
and U27125 (N_27125,N_24168,N_24614);
nor U27126 (N_27126,N_25194,N_25287);
and U27127 (N_27127,N_24218,N_24997);
or U27128 (N_27128,N_24850,N_24982);
and U27129 (N_27129,N_24676,N_25573);
nand U27130 (N_27130,N_24783,N_25716);
or U27131 (N_27131,N_24450,N_24583);
nand U27132 (N_27132,N_25195,N_25292);
and U27133 (N_27133,N_25106,N_24853);
and U27134 (N_27134,N_24889,N_25313);
or U27135 (N_27135,N_24880,N_25527);
or U27136 (N_27136,N_24706,N_24169);
and U27137 (N_27137,N_24505,N_24916);
xor U27138 (N_27138,N_24361,N_25230);
nand U27139 (N_27139,N_25684,N_24192);
and U27140 (N_27140,N_24150,N_24439);
and U27141 (N_27141,N_24433,N_24057);
xnor U27142 (N_27142,N_25020,N_25744);
or U27143 (N_27143,N_24278,N_24171);
nand U27144 (N_27144,N_25547,N_25306);
and U27145 (N_27145,N_25655,N_25321);
xnor U27146 (N_27146,N_25447,N_24198);
nor U27147 (N_27147,N_25662,N_25777);
xnor U27148 (N_27148,N_24879,N_24258);
nor U27149 (N_27149,N_25106,N_25411);
and U27150 (N_27150,N_24299,N_25643);
or U27151 (N_27151,N_25360,N_24202);
nand U27152 (N_27152,N_24790,N_24660);
nor U27153 (N_27153,N_25321,N_25136);
or U27154 (N_27154,N_25975,N_24071);
nand U27155 (N_27155,N_24815,N_25218);
and U27156 (N_27156,N_24513,N_24510);
or U27157 (N_27157,N_24427,N_25289);
or U27158 (N_27158,N_25435,N_25896);
xnor U27159 (N_27159,N_25721,N_24851);
or U27160 (N_27160,N_24464,N_25483);
xor U27161 (N_27161,N_24912,N_25073);
nor U27162 (N_27162,N_25720,N_24367);
and U27163 (N_27163,N_24112,N_25163);
xor U27164 (N_27164,N_24428,N_24711);
nor U27165 (N_27165,N_25768,N_25386);
nor U27166 (N_27166,N_24666,N_24736);
xor U27167 (N_27167,N_24187,N_24317);
nor U27168 (N_27168,N_24176,N_24464);
and U27169 (N_27169,N_25576,N_24224);
nand U27170 (N_27170,N_25164,N_24180);
nor U27171 (N_27171,N_24139,N_25726);
nor U27172 (N_27172,N_24909,N_25338);
nand U27173 (N_27173,N_24543,N_24314);
or U27174 (N_27174,N_24200,N_25028);
nor U27175 (N_27175,N_25445,N_24420);
xnor U27176 (N_27176,N_25017,N_24864);
nor U27177 (N_27177,N_24183,N_24142);
nor U27178 (N_27178,N_25479,N_25096);
and U27179 (N_27179,N_25870,N_24675);
xor U27180 (N_27180,N_24976,N_25606);
xnor U27181 (N_27181,N_25004,N_24554);
xor U27182 (N_27182,N_25975,N_24080);
or U27183 (N_27183,N_24243,N_24532);
xnor U27184 (N_27184,N_25516,N_25172);
xor U27185 (N_27185,N_25833,N_24330);
nor U27186 (N_27186,N_25023,N_25684);
and U27187 (N_27187,N_25680,N_25235);
nand U27188 (N_27188,N_24206,N_24456);
nor U27189 (N_27189,N_24853,N_24417);
nand U27190 (N_27190,N_24569,N_25334);
nand U27191 (N_27191,N_25193,N_24806);
nor U27192 (N_27192,N_25662,N_24349);
nand U27193 (N_27193,N_24033,N_24008);
nor U27194 (N_27194,N_25491,N_24271);
or U27195 (N_27195,N_25683,N_24830);
nand U27196 (N_27196,N_24337,N_25610);
nand U27197 (N_27197,N_25772,N_24130);
nor U27198 (N_27198,N_25412,N_24097);
nor U27199 (N_27199,N_25431,N_25928);
nor U27200 (N_27200,N_24293,N_25050);
and U27201 (N_27201,N_24715,N_24732);
and U27202 (N_27202,N_25315,N_25740);
or U27203 (N_27203,N_25132,N_24398);
and U27204 (N_27204,N_25088,N_24144);
xor U27205 (N_27205,N_24909,N_24170);
and U27206 (N_27206,N_25396,N_24046);
and U27207 (N_27207,N_24471,N_25890);
xnor U27208 (N_27208,N_24174,N_24871);
nor U27209 (N_27209,N_24713,N_25234);
or U27210 (N_27210,N_24025,N_25714);
nor U27211 (N_27211,N_24600,N_25866);
or U27212 (N_27212,N_24925,N_25937);
nor U27213 (N_27213,N_24160,N_25072);
nor U27214 (N_27214,N_25634,N_24185);
xor U27215 (N_27215,N_24057,N_24292);
nand U27216 (N_27216,N_25161,N_24654);
nor U27217 (N_27217,N_24249,N_25022);
and U27218 (N_27218,N_24180,N_24071);
xor U27219 (N_27219,N_24597,N_25448);
nor U27220 (N_27220,N_25220,N_25019);
xor U27221 (N_27221,N_24494,N_25148);
nand U27222 (N_27222,N_25427,N_24136);
or U27223 (N_27223,N_24469,N_24832);
xnor U27224 (N_27224,N_25956,N_25369);
xor U27225 (N_27225,N_25671,N_25894);
and U27226 (N_27226,N_25361,N_24371);
nand U27227 (N_27227,N_24461,N_25658);
nor U27228 (N_27228,N_25662,N_25952);
nor U27229 (N_27229,N_25920,N_24207);
nor U27230 (N_27230,N_24228,N_24734);
nor U27231 (N_27231,N_24510,N_24669);
xnor U27232 (N_27232,N_24074,N_25732);
and U27233 (N_27233,N_25576,N_24594);
and U27234 (N_27234,N_25141,N_24113);
nor U27235 (N_27235,N_25232,N_24831);
or U27236 (N_27236,N_24503,N_24159);
or U27237 (N_27237,N_24723,N_24408);
or U27238 (N_27238,N_25781,N_25080);
or U27239 (N_27239,N_24096,N_25802);
or U27240 (N_27240,N_25416,N_24301);
or U27241 (N_27241,N_25182,N_25352);
nor U27242 (N_27242,N_25188,N_25129);
xnor U27243 (N_27243,N_24417,N_24321);
or U27244 (N_27244,N_24975,N_25948);
nand U27245 (N_27245,N_25961,N_24191);
nand U27246 (N_27246,N_24417,N_25342);
and U27247 (N_27247,N_25758,N_25602);
nand U27248 (N_27248,N_25804,N_24877);
xnor U27249 (N_27249,N_24971,N_25618);
and U27250 (N_27250,N_24604,N_24837);
nand U27251 (N_27251,N_24243,N_24868);
nand U27252 (N_27252,N_24200,N_25418);
nand U27253 (N_27253,N_25536,N_25377);
and U27254 (N_27254,N_24490,N_25262);
and U27255 (N_27255,N_24102,N_25498);
xor U27256 (N_27256,N_25294,N_24606);
nand U27257 (N_27257,N_25590,N_25065);
or U27258 (N_27258,N_24426,N_25216);
nand U27259 (N_27259,N_25269,N_25745);
xnor U27260 (N_27260,N_24253,N_24991);
nand U27261 (N_27261,N_25790,N_25133);
nor U27262 (N_27262,N_24834,N_25251);
and U27263 (N_27263,N_24515,N_24318);
and U27264 (N_27264,N_25821,N_25799);
and U27265 (N_27265,N_25768,N_25769);
or U27266 (N_27266,N_24072,N_24455);
or U27267 (N_27267,N_25662,N_24890);
and U27268 (N_27268,N_24811,N_25408);
and U27269 (N_27269,N_24686,N_25081);
nor U27270 (N_27270,N_25436,N_24622);
and U27271 (N_27271,N_24994,N_25380);
nor U27272 (N_27272,N_25682,N_25191);
and U27273 (N_27273,N_24627,N_24282);
or U27274 (N_27274,N_24026,N_24908);
nand U27275 (N_27275,N_24729,N_25037);
and U27276 (N_27276,N_24047,N_25589);
xor U27277 (N_27277,N_24417,N_25882);
nand U27278 (N_27278,N_25443,N_24837);
nor U27279 (N_27279,N_25479,N_25924);
nor U27280 (N_27280,N_25239,N_25584);
xor U27281 (N_27281,N_25248,N_24239);
nand U27282 (N_27282,N_25741,N_25593);
xnor U27283 (N_27283,N_24786,N_25468);
nand U27284 (N_27284,N_24229,N_25829);
or U27285 (N_27285,N_25636,N_25837);
and U27286 (N_27286,N_25690,N_25851);
xor U27287 (N_27287,N_25219,N_24562);
nand U27288 (N_27288,N_25898,N_24369);
nor U27289 (N_27289,N_25298,N_25804);
nor U27290 (N_27290,N_25265,N_24427);
nand U27291 (N_27291,N_25299,N_25415);
nor U27292 (N_27292,N_25800,N_24061);
xnor U27293 (N_27293,N_24570,N_24428);
nand U27294 (N_27294,N_24928,N_24421);
or U27295 (N_27295,N_24612,N_25147);
and U27296 (N_27296,N_24737,N_25094);
nor U27297 (N_27297,N_24208,N_24983);
and U27298 (N_27298,N_25974,N_25768);
nor U27299 (N_27299,N_25663,N_25907);
xnor U27300 (N_27300,N_25321,N_25139);
or U27301 (N_27301,N_24146,N_25122);
nand U27302 (N_27302,N_24223,N_24561);
and U27303 (N_27303,N_25643,N_24723);
xnor U27304 (N_27304,N_25355,N_24895);
xor U27305 (N_27305,N_24066,N_24604);
xor U27306 (N_27306,N_25679,N_25020);
xnor U27307 (N_27307,N_24855,N_24105);
nand U27308 (N_27308,N_24035,N_25904);
or U27309 (N_27309,N_25690,N_25827);
nand U27310 (N_27310,N_25957,N_24279);
nand U27311 (N_27311,N_24866,N_24466);
nand U27312 (N_27312,N_24997,N_24345);
nand U27313 (N_27313,N_25476,N_25132);
or U27314 (N_27314,N_24445,N_25954);
or U27315 (N_27315,N_25025,N_25039);
nand U27316 (N_27316,N_24804,N_25359);
or U27317 (N_27317,N_24069,N_25507);
nor U27318 (N_27318,N_24720,N_24455);
nand U27319 (N_27319,N_24028,N_24893);
xnor U27320 (N_27320,N_24618,N_24928);
nand U27321 (N_27321,N_24212,N_25767);
and U27322 (N_27322,N_25801,N_25665);
and U27323 (N_27323,N_24734,N_25143);
nand U27324 (N_27324,N_25393,N_25447);
and U27325 (N_27325,N_25419,N_24532);
nor U27326 (N_27326,N_25433,N_25146);
nand U27327 (N_27327,N_24489,N_24574);
nand U27328 (N_27328,N_25587,N_24597);
nand U27329 (N_27329,N_25255,N_24388);
nand U27330 (N_27330,N_24133,N_25139);
or U27331 (N_27331,N_24203,N_24858);
nor U27332 (N_27332,N_24760,N_25398);
nor U27333 (N_27333,N_25970,N_25175);
nor U27334 (N_27334,N_25656,N_24776);
or U27335 (N_27335,N_24820,N_24222);
or U27336 (N_27336,N_25810,N_25041);
nor U27337 (N_27337,N_24550,N_25465);
and U27338 (N_27338,N_24127,N_25615);
and U27339 (N_27339,N_24121,N_24553);
nand U27340 (N_27340,N_25896,N_25422);
and U27341 (N_27341,N_24267,N_25436);
nor U27342 (N_27342,N_25527,N_24840);
and U27343 (N_27343,N_24503,N_25020);
xor U27344 (N_27344,N_24474,N_25162);
and U27345 (N_27345,N_25587,N_25858);
xor U27346 (N_27346,N_24620,N_24169);
nand U27347 (N_27347,N_25526,N_25107);
and U27348 (N_27348,N_24585,N_24095);
nor U27349 (N_27349,N_25485,N_25428);
xor U27350 (N_27350,N_24617,N_25774);
nor U27351 (N_27351,N_25766,N_24776);
nor U27352 (N_27352,N_24123,N_24953);
nand U27353 (N_27353,N_25468,N_24596);
nor U27354 (N_27354,N_25622,N_24906);
xor U27355 (N_27355,N_25350,N_24634);
nor U27356 (N_27356,N_24315,N_24638);
xor U27357 (N_27357,N_24904,N_24935);
xnor U27358 (N_27358,N_25070,N_24403);
and U27359 (N_27359,N_24239,N_25471);
and U27360 (N_27360,N_25603,N_25730);
nor U27361 (N_27361,N_25311,N_25473);
nand U27362 (N_27362,N_24014,N_25254);
and U27363 (N_27363,N_25560,N_25840);
nand U27364 (N_27364,N_24382,N_25296);
nor U27365 (N_27365,N_24661,N_24995);
nor U27366 (N_27366,N_24773,N_25707);
nand U27367 (N_27367,N_24558,N_24035);
or U27368 (N_27368,N_24591,N_24114);
or U27369 (N_27369,N_25352,N_24660);
and U27370 (N_27370,N_25252,N_24597);
or U27371 (N_27371,N_24401,N_24502);
nor U27372 (N_27372,N_25212,N_25321);
nand U27373 (N_27373,N_24712,N_24310);
nand U27374 (N_27374,N_25122,N_24533);
and U27375 (N_27375,N_24702,N_25597);
or U27376 (N_27376,N_24399,N_25446);
nand U27377 (N_27377,N_25674,N_25065);
xnor U27378 (N_27378,N_25585,N_25056);
xor U27379 (N_27379,N_25701,N_25747);
nor U27380 (N_27380,N_25579,N_24915);
xnor U27381 (N_27381,N_25452,N_24286);
nor U27382 (N_27382,N_24385,N_25091);
or U27383 (N_27383,N_24709,N_25096);
nand U27384 (N_27384,N_24007,N_24070);
nand U27385 (N_27385,N_25121,N_24252);
xnor U27386 (N_27386,N_24256,N_24864);
and U27387 (N_27387,N_24869,N_24034);
and U27388 (N_27388,N_24979,N_25394);
xnor U27389 (N_27389,N_25345,N_25831);
or U27390 (N_27390,N_25405,N_24651);
and U27391 (N_27391,N_25182,N_25362);
nand U27392 (N_27392,N_25617,N_24897);
nand U27393 (N_27393,N_25047,N_24676);
or U27394 (N_27394,N_24915,N_25150);
xor U27395 (N_27395,N_25442,N_24416);
nor U27396 (N_27396,N_24327,N_25598);
or U27397 (N_27397,N_24002,N_24016);
nor U27398 (N_27398,N_24458,N_24687);
nand U27399 (N_27399,N_25506,N_25250);
nor U27400 (N_27400,N_24342,N_25400);
nand U27401 (N_27401,N_25560,N_24764);
nand U27402 (N_27402,N_25774,N_24028);
nand U27403 (N_27403,N_24429,N_25572);
xor U27404 (N_27404,N_24219,N_25313);
and U27405 (N_27405,N_24636,N_25025);
and U27406 (N_27406,N_25121,N_25661);
xnor U27407 (N_27407,N_25279,N_24125);
xnor U27408 (N_27408,N_25653,N_24547);
nor U27409 (N_27409,N_25472,N_24586);
nor U27410 (N_27410,N_24661,N_24200);
xnor U27411 (N_27411,N_24747,N_24669);
nor U27412 (N_27412,N_25763,N_24087);
nand U27413 (N_27413,N_25755,N_25706);
and U27414 (N_27414,N_24901,N_24955);
and U27415 (N_27415,N_24487,N_24451);
or U27416 (N_27416,N_24379,N_25960);
or U27417 (N_27417,N_24491,N_24140);
nor U27418 (N_27418,N_25841,N_25783);
nand U27419 (N_27419,N_25557,N_24313);
and U27420 (N_27420,N_25703,N_25014);
nor U27421 (N_27421,N_25631,N_24505);
or U27422 (N_27422,N_24703,N_25878);
nand U27423 (N_27423,N_25876,N_24757);
xnor U27424 (N_27424,N_25976,N_24102);
xor U27425 (N_27425,N_25951,N_24710);
or U27426 (N_27426,N_24570,N_25810);
xor U27427 (N_27427,N_25570,N_25414);
nor U27428 (N_27428,N_25075,N_24957);
or U27429 (N_27429,N_24940,N_25171);
nand U27430 (N_27430,N_25078,N_25020);
nand U27431 (N_27431,N_25368,N_25644);
nand U27432 (N_27432,N_25985,N_24262);
or U27433 (N_27433,N_24925,N_24554);
or U27434 (N_27434,N_24812,N_25375);
xor U27435 (N_27435,N_25022,N_24136);
nor U27436 (N_27436,N_24054,N_25874);
and U27437 (N_27437,N_24983,N_24070);
xor U27438 (N_27438,N_24145,N_24134);
xnor U27439 (N_27439,N_25168,N_25894);
nand U27440 (N_27440,N_24829,N_25205);
or U27441 (N_27441,N_24858,N_24723);
or U27442 (N_27442,N_24391,N_24981);
or U27443 (N_27443,N_25755,N_24171);
nor U27444 (N_27444,N_24279,N_24700);
nand U27445 (N_27445,N_25757,N_24512);
and U27446 (N_27446,N_25592,N_25398);
xnor U27447 (N_27447,N_25293,N_25527);
nand U27448 (N_27448,N_24587,N_24028);
or U27449 (N_27449,N_24334,N_24963);
nand U27450 (N_27450,N_24413,N_24738);
xor U27451 (N_27451,N_24323,N_25884);
nand U27452 (N_27452,N_24815,N_24269);
nand U27453 (N_27453,N_25808,N_25962);
nor U27454 (N_27454,N_25971,N_25109);
nor U27455 (N_27455,N_25667,N_24296);
nor U27456 (N_27456,N_24179,N_25364);
or U27457 (N_27457,N_24533,N_25909);
and U27458 (N_27458,N_24349,N_24764);
and U27459 (N_27459,N_25928,N_24150);
and U27460 (N_27460,N_24740,N_25287);
xnor U27461 (N_27461,N_25326,N_25265);
or U27462 (N_27462,N_25034,N_25396);
xor U27463 (N_27463,N_24837,N_24368);
nor U27464 (N_27464,N_25037,N_24631);
or U27465 (N_27465,N_25627,N_24994);
nor U27466 (N_27466,N_24352,N_24849);
nor U27467 (N_27467,N_25157,N_24826);
nand U27468 (N_27468,N_24951,N_24455);
xor U27469 (N_27469,N_24195,N_25870);
or U27470 (N_27470,N_24624,N_25364);
nor U27471 (N_27471,N_24825,N_24378);
or U27472 (N_27472,N_24108,N_25144);
xor U27473 (N_27473,N_24804,N_25153);
xnor U27474 (N_27474,N_25258,N_25949);
and U27475 (N_27475,N_24221,N_24581);
xor U27476 (N_27476,N_25948,N_24824);
xor U27477 (N_27477,N_24565,N_25877);
nor U27478 (N_27478,N_24436,N_24788);
or U27479 (N_27479,N_25375,N_25981);
and U27480 (N_27480,N_24886,N_25150);
nor U27481 (N_27481,N_25811,N_25077);
xnor U27482 (N_27482,N_25283,N_24474);
nand U27483 (N_27483,N_25683,N_24330);
nor U27484 (N_27484,N_25505,N_25232);
nand U27485 (N_27485,N_24459,N_25693);
nand U27486 (N_27486,N_24429,N_25397);
nor U27487 (N_27487,N_24146,N_24747);
xnor U27488 (N_27488,N_24377,N_25493);
and U27489 (N_27489,N_25300,N_25009);
and U27490 (N_27490,N_25609,N_24283);
and U27491 (N_27491,N_24249,N_25955);
nand U27492 (N_27492,N_24956,N_24697);
xnor U27493 (N_27493,N_25253,N_25135);
or U27494 (N_27494,N_25979,N_25050);
xor U27495 (N_27495,N_25308,N_24012);
xor U27496 (N_27496,N_25723,N_25402);
nand U27497 (N_27497,N_24861,N_24245);
xor U27498 (N_27498,N_25895,N_24392);
and U27499 (N_27499,N_25299,N_24686);
xnor U27500 (N_27500,N_25376,N_24825);
xor U27501 (N_27501,N_24619,N_25612);
and U27502 (N_27502,N_24945,N_24825);
nor U27503 (N_27503,N_25318,N_25135);
xnor U27504 (N_27504,N_25411,N_25350);
xor U27505 (N_27505,N_25241,N_25461);
and U27506 (N_27506,N_25630,N_25481);
nor U27507 (N_27507,N_24934,N_24807);
or U27508 (N_27508,N_24899,N_24260);
nand U27509 (N_27509,N_24394,N_24433);
or U27510 (N_27510,N_25520,N_25703);
and U27511 (N_27511,N_24540,N_25867);
nand U27512 (N_27512,N_24953,N_24803);
or U27513 (N_27513,N_25497,N_24220);
nand U27514 (N_27514,N_25400,N_24331);
and U27515 (N_27515,N_24042,N_24833);
xnor U27516 (N_27516,N_25770,N_25668);
and U27517 (N_27517,N_25869,N_24795);
xnor U27518 (N_27518,N_25224,N_24241);
and U27519 (N_27519,N_25933,N_25956);
nand U27520 (N_27520,N_25932,N_24013);
and U27521 (N_27521,N_24394,N_25684);
nor U27522 (N_27522,N_24891,N_25279);
nand U27523 (N_27523,N_24376,N_25128);
or U27524 (N_27524,N_24938,N_24339);
nor U27525 (N_27525,N_24325,N_24421);
or U27526 (N_27526,N_25615,N_25385);
nor U27527 (N_27527,N_25999,N_25998);
and U27528 (N_27528,N_24633,N_25159);
nor U27529 (N_27529,N_24626,N_25448);
or U27530 (N_27530,N_25228,N_24326);
xor U27531 (N_27531,N_24931,N_25221);
nor U27532 (N_27532,N_25947,N_24754);
and U27533 (N_27533,N_24213,N_25480);
nand U27534 (N_27534,N_25144,N_24785);
and U27535 (N_27535,N_24379,N_24115);
and U27536 (N_27536,N_24603,N_25562);
xnor U27537 (N_27537,N_24225,N_25536);
xor U27538 (N_27538,N_24009,N_25929);
xnor U27539 (N_27539,N_24349,N_24991);
and U27540 (N_27540,N_24048,N_24596);
or U27541 (N_27541,N_24038,N_25475);
nand U27542 (N_27542,N_24267,N_25493);
xnor U27543 (N_27543,N_24337,N_24775);
nand U27544 (N_27544,N_24454,N_24519);
or U27545 (N_27545,N_25736,N_25496);
nor U27546 (N_27546,N_25443,N_25713);
nand U27547 (N_27547,N_24231,N_24880);
nand U27548 (N_27548,N_24075,N_24415);
or U27549 (N_27549,N_24037,N_24718);
nor U27550 (N_27550,N_25812,N_25423);
and U27551 (N_27551,N_24465,N_24481);
xor U27552 (N_27552,N_25933,N_24931);
nor U27553 (N_27553,N_24966,N_24134);
or U27554 (N_27554,N_25804,N_25783);
xnor U27555 (N_27555,N_25081,N_25101);
xor U27556 (N_27556,N_24921,N_25902);
and U27557 (N_27557,N_25136,N_24795);
nand U27558 (N_27558,N_25364,N_25001);
nand U27559 (N_27559,N_24346,N_24520);
and U27560 (N_27560,N_25384,N_24874);
xor U27561 (N_27561,N_25492,N_25108);
and U27562 (N_27562,N_25652,N_24207);
nor U27563 (N_27563,N_24807,N_24256);
nor U27564 (N_27564,N_24594,N_24010);
and U27565 (N_27565,N_25031,N_25381);
xor U27566 (N_27566,N_25082,N_25642);
xor U27567 (N_27567,N_24999,N_24321);
nor U27568 (N_27568,N_25564,N_24630);
nor U27569 (N_27569,N_25718,N_24495);
xnor U27570 (N_27570,N_25741,N_25118);
xor U27571 (N_27571,N_25328,N_25641);
or U27572 (N_27572,N_24651,N_25582);
nor U27573 (N_27573,N_25288,N_24357);
nor U27574 (N_27574,N_25229,N_24785);
xnor U27575 (N_27575,N_25688,N_24012);
xnor U27576 (N_27576,N_24275,N_24148);
nand U27577 (N_27577,N_25384,N_25643);
nor U27578 (N_27578,N_25587,N_25621);
xnor U27579 (N_27579,N_25554,N_25843);
and U27580 (N_27580,N_25172,N_25585);
nor U27581 (N_27581,N_25611,N_24782);
xor U27582 (N_27582,N_25274,N_24676);
or U27583 (N_27583,N_25991,N_24948);
or U27584 (N_27584,N_25370,N_25374);
and U27585 (N_27585,N_24305,N_24459);
nand U27586 (N_27586,N_24818,N_25938);
xnor U27587 (N_27587,N_25543,N_25046);
or U27588 (N_27588,N_24127,N_25186);
and U27589 (N_27589,N_25599,N_25319);
nand U27590 (N_27590,N_25900,N_25025);
xor U27591 (N_27591,N_25608,N_24699);
nor U27592 (N_27592,N_25086,N_25484);
nor U27593 (N_27593,N_25837,N_24242);
nand U27594 (N_27594,N_25589,N_25701);
nor U27595 (N_27595,N_25408,N_24464);
xnor U27596 (N_27596,N_24105,N_24630);
or U27597 (N_27597,N_24648,N_24342);
nand U27598 (N_27598,N_25060,N_25111);
nor U27599 (N_27599,N_24212,N_24253);
nor U27600 (N_27600,N_24637,N_24115);
or U27601 (N_27601,N_25921,N_25573);
and U27602 (N_27602,N_24352,N_24130);
nand U27603 (N_27603,N_24234,N_25188);
or U27604 (N_27604,N_24087,N_24455);
nor U27605 (N_27605,N_24339,N_25377);
nor U27606 (N_27606,N_25561,N_24185);
nand U27607 (N_27607,N_25680,N_24145);
and U27608 (N_27608,N_25875,N_24917);
nand U27609 (N_27609,N_24539,N_24387);
xnor U27610 (N_27610,N_25675,N_25977);
nand U27611 (N_27611,N_24808,N_24249);
xnor U27612 (N_27612,N_24520,N_24753);
xnor U27613 (N_27613,N_25582,N_24083);
xor U27614 (N_27614,N_25314,N_24018);
nor U27615 (N_27615,N_24476,N_24977);
and U27616 (N_27616,N_24212,N_25903);
nand U27617 (N_27617,N_24747,N_25384);
or U27618 (N_27618,N_24988,N_24726);
nor U27619 (N_27619,N_25563,N_24533);
nor U27620 (N_27620,N_24828,N_25896);
or U27621 (N_27621,N_24102,N_25497);
and U27622 (N_27622,N_25818,N_25812);
nor U27623 (N_27623,N_24882,N_25063);
and U27624 (N_27624,N_25334,N_24711);
nand U27625 (N_27625,N_24584,N_25098);
or U27626 (N_27626,N_24704,N_25391);
nand U27627 (N_27627,N_25815,N_24400);
or U27628 (N_27628,N_25261,N_25939);
and U27629 (N_27629,N_25787,N_25994);
xnor U27630 (N_27630,N_25567,N_25472);
nand U27631 (N_27631,N_24283,N_24316);
nand U27632 (N_27632,N_25162,N_25167);
and U27633 (N_27633,N_24990,N_24309);
nand U27634 (N_27634,N_24847,N_25246);
xnor U27635 (N_27635,N_25693,N_24731);
nor U27636 (N_27636,N_25073,N_25926);
xnor U27637 (N_27637,N_24161,N_24464);
xnor U27638 (N_27638,N_25304,N_25244);
or U27639 (N_27639,N_24933,N_25225);
nor U27640 (N_27640,N_24016,N_24858);
nor U27641 (N_27641,N_24545,N_24194);
and U27642 (N_27642,N_25336,N_24683);
xor U27643 (N_27643,N_25747,N_24252);
nand U27644 (N_27644,N_24347,N_24535);
nand U27645 (N_27645,N_24588,N_25659);
and U27646 (N_27646,N_25608,N_24398);
nand U27647 (N_27647,N_24978,N_24005);
or U27648 (N_27648,N_24517,N_24838);
or U27649 (N_27649,N_25629,N_25686);
and U27650 (N_27650,N_25504,N_24430);
or U27651 (N_27651,N_25626,N_25218);
nor U27652 (N_27652,N_24184,N_24236);
xor U27653 (N_27653,N_25738,N_24738);
nor U27654 (N_27654,N_25981,N_24253);
or U27655 (N_27655,N_25965,N_24589);
or U27656 (N_27656,N_25359,N_24291);
xnor U27657 (N_27657,N_24679,N_24166);
nor U27658 (N_27658,N_25240,N_25443);
and U27659 (N_27659,N_24747,N_25586);
and U27660 (N_27660,N_24040,N_25397);
xor U27661 (N_27661,N_25621,N_25507);
or U27662 (N_27662,N_25850,N_24562);
or U27663 (N_27663,N_24509,N_25211);
or U27664 (N_27664,N_25612,N_24142);
nand U27665 (N_27665,N_25858,N_25164);
nor U27666 (N_27666,N_24125,N_25535);
or U27667 (N_27667,N_24562,N_24283);
or U27668 (N_27668,N_24902,N_25520);
or U27669 (N_27669,N_24605,N_25357);
and U27670 (N_27670,N_24549,N_25807);
nor U27671 (N_27671,N_25007,N_25049);
nand U27672 (N_27672,N_25442,N_24242);
nand U27673 (N_27673,N_25304,N_24501);
nand U27674 (N_27674,N_25310,N_24753);
xnor U27675 (N_27675,N_25153,N_25082);
or U27676 (N_27676,N_25704,N_25143);
or U27677 (N_27677,N_24448,N_25302);
or U27678 (N_27678,N_25033,N_24372);
xor U27679 (N_27679,N_25861,N_24013);
xnor U27680 (N_27680,N_24565,N_25055);
and U27681 (N_27681,N_25522,N_25090);
and U27682 (N_27682,N_24266,N_25841);
nand U27683 (N_27683,N_25736,N_25070);
or U27684 (N_27684,N_25226,N_24917);
nand U27685 (N_27685,N_24143,N_25951);
nor U27686 (N_27686,N_25391,N_24728);
nand U27687 (N_27687,N_25695,N_24733);
or U27688 (N_27688,N_25980,N_25566);
nand U27689 (N_27689,N_24639,N_24500);
xor U27690 (N_27690,N_24301,N_25018);
and U27691 (N_27691,N_25335,N_25201);
or U27692 (N_27692,N_24329,N_24081);
nand U27693 (N_27693,N_24291,N_24832);
nor U27694 (N_27694,N_25574,N_25352);
nand U27695 (N_27695,N_25514,N_25923);
and U27696 (N_27696,N_24204,N_24068);
nand U27697 (N_27697,N_25161,N_24642);
or U27698 (N_27698,N_24483,N_25683);
xnor U27699 (N_27699,N_24799,N_24970);
and U27700 (N_27700,N_25632,N_25995);
and U27701 (N_27701,N_25287,N_25987);
nor U27702 (N_27702,N_24963,N_25972);
and U27703 (N_27703,N_24966,N_24599);
and U27704 (N_27704,N_24088,N_24425);
or U27705 (N_27705,N_24418,N_25758);
nor U27706 (N_27706,N_24598,N_24105);
nand U27707 (N_27707,N_25514,N_24706);
nand U27708 (N_27708,N_24859,N_24860);
nor U27709 (N_27709,N_25807,N_25746);
nand U27710 (N_27710,N_24615,N_24895);
or U27711 (N_27711,N_24649,N_24047);
nand U27712 (N_27712,N_25224,N_25266);
and U27713 (N_27713,N_25988,N_25201);
nand U27714 (N_27714,N_25721,N_25850);
nand U27715 (N_27715,N_24629,N_24583);
nor U27716 (N_27716,N_25678,N_25082);
xnor U27717 (N_27717,N_24249,N_24065);
or U27718 (N_27718,N_25988,N_24211);
or U27719 (N_27719,N_24939,N_24195);
nand U27720 (N_27720,N_24524,N_24355);
nor U27721 (N_27721,N_25411,N_24145);
nand U27722 (N_27722,N_25755,N_24289);
and U27723 (N_27723,N_25619,N_25738);
nand U27724 (N_27724,N_25560,N_25520);
or U27725 (N_27725,N_25809,N_25752);
or U27726 (N_27726,N_25655,N_25733);
or U27727 (N_27727,N_25171,N_24473);
and U27728 (N_27728,N_25828,N_24661);
and U27729 (N_27729,N_25863,N_24521);
xnor U27730 (N_27730,N_24210,N_25831);
or U27731 (N_27731,N_24210,N_25559);
or U27732 (N_27732,N_24433,N_25944);
nand U27733 (N_27733,N_25532,N_24537);
and U27734 (N_27734,N_24837,N_24776);
and U27735 (N_27735,N_25021,N_25584);
nor U27736 (N_27736,N_25441,N_24698);
xor U27737 (N_27737,N_25904,N_24759);
nor U27738 (N_27738,N_24238,N_24333);
xnor U27739 (N_27739,N_24018,N_24158);
nor U27740 (N_27740,N_24173,N_24179);
and U27741 (N_27741,N_24803,N_24396);
xnor U27742 (N_27742,N_25343,N_25112);
xor U27743 (N_27743,N_25459,N_25844);
or U27744 (N_27744,N_25390,N_24192);
nor U27745 (N_27745,N_25987,N_24105);
and U27746 (N_27746,N_24011,N_25180);
nand U27747 (N_27747,N_25921,N_24885);
xor U27748 (N_27748,N_24710,N_25993);
or U27749 (N_27749,N_24983,N_24322);
xor U27750 (N_27750,N_24789,N_24795);
and U27751 (N_27751,N_25106,N_25248);
nor U27752 (N_27752,N_24733,N_24119);
or U27753 (N_27753,N_24342,N_25469);
or U27754 (N_27754,N_24414,N_24177);
nand U27755 (N_27755,N_24469,N_24055);
nor U27756 (N_27756,N_24356,N_25134);
and U27757 (N_27757,N_24666,N_25639);
nor U27758 (N_27758,N_24950,N_25743);
nand U27759 (N_27759,N_24017,N_25558);
and U27760 (N_27760,N_24742,N_24809);
or U27761 (N_27761,N_24532,N_25245);
nand U27762 (N_27762,N_25505,N_25858);
or U27763 (N_27763,N_24399,N_24028);
nand U27764 (N_27764,N_24655,N_25299);
or U27765 (N_27765,N_25802,N_24609);
or U27766 (N_27766,N_24667,N_24218);
or U27767 (N_27767,N_24383,N_25344);
xnor U27768 (N_27768,N_25714,N_24987);
xor U27769 (N_27769,N_24350,N_25487);
xnor U27770 (N_27770,N_25880,N_25580);
nand U27771 (N_27771,N_25193,N_24103);
nand U27772 (N_27772,N_25073,N_25925);
xnor U27773 (N_27773,N_25294,N_25478);
nand U27774 (N_27774,N_24548,N_24553);
and U27775 (N_27775,N_24582,N_24294);
nand U27776 (N_27776,N_24075,N_24082);
nor U27777 (N_27777,N_24780,N_24861);
xnor U27778 (N_27778,N_25305,N_24409);
or U27779 (N_27779,N_24286,N_24810);
nor U27780 (N_27780,N_25191,N_25226);
nor U27781 (N_27781,N_25878,N_25243);
nand U27782 (N_27782,N_24025,N_24980);
or U27783 (N_27783,N_25372,N_24985);
xnor U27784 (N_27784,N_24288,N_25415);
nand U27785 (N_27785,N_25376,N_25702);
nor U27786 (N_27786,N_24463,N_25828);
xnor U27787 (N_27787,N_25713,N_24229);
nor U27788 (N_27788,N_24395,N_24266);
and U27789 (N_27789,N_25415,N_25412);
xnor U27790 (N_27790,N_25666,N_24415);
nor U27791 (N_27791,N_24808,N_25000);
or U27792 (N_27792,N_25132,N_25623);
nand U27793 (N_27793,N_24933,N_24434);
xnor U27794 (N_27794,N_24675,N_25895);
xor U27795 (N_27795,N_24592,N_24485);
or U27796 (N_27796,N_24712,N_25926);
and U27797 (N_27797,N_24000,N_24948);
nor U27798 (N_27798,N_24655,N_25036);
and U27799 (N_27799,N_25593,N_24067);
nand U27800 (N_27800,N_24031,N_25688);
nand U27801 (N_27801,N_24041,N_25168);
xnor U27802 (N_27802,N_25502,N_25106);
nand U27803 (N_27803,N_24866,N_24460);
or U27804 (N_27804,N_24825,N_25600);
nand U27805 (N_27805,N_25019,N_25940);
xnor U27806 (N_27806,N_25273,N_24971);
and U27807 (N_27807,N_24129,N_24849);
nand U27808 (N_27808,N_24500,N_24369);
and U27809 (N_27809,N_25172,N_25280);
nor U27810 (N_27810,N_24340,N_24435);
nand U27811 (N_27811,N_25940,N_24405);
nand U27812 (N_27812,N_24220,N_25882);
xnor U27813 (N_27813,N_25639,N_25832);
nand U27814 (N_27814,N_25423,N_25712);
xnor U27815 (N_27815,N_25571,N_24643);
nor U27816 (N_27816,N_25219,N_24305);
nand U27817 (N_27817,N_24574,N_25559);
xor U27818 (N_27818,N_25060,N_24369);
and U27819 (N_27819,N_25267,N_24420);
nand U27820 (N_27820,N_24008,N_24374);
nor U27821 (N_27821,N_24584,N_25430);
xnor U27822 (N_27822,N_25345,N_24906);
and U27823 (N_27823,N_25701,N_25540);
and U27824 (N_27824,N_25090,N_25402);
xnor U27825 (N_27825,N_25514,N_24867);
nand U27826 (N_27826,N_25968,N_24949);
nor U27827 (N_27827,N_24880,N_25528);
and U27828 (N_27828,N_25881,N_24822);
nand U27829 (N_27829,N_24112,N_25952);
and U27830 (N_27830,N_25566,N_24001);
xnor U27831 (N_27831,N_24677,N_24202);
nor U27832 (N_27832,N_24977,N_25288);
or U27833 (N_27833,N_25601,N_24973);
nand U27834 (N_27834,N_24701,N_25085);
and U27835 (N_27835,N_25534,N_25260);
or U27836 (N_27836,N_25165,N_25858);
xnor U27837 (N_27837,N_24567,N_25543);
and U27838 (N_27838,N_25023,N_25660);
and U27839 (N_27839,N_24076,N_25863);
xnor U27840 (N_27840,N_25970,N_25412);
xnor U27841 (N_27841,N_24683,N_25116);
or U27842 (N_27842,N_25364,N_24449);
nor U27843 (N_27843,N_25857,N_24431);
and U27844 (N_27844,N_24569,N_25207);
or U27845 (N_27845,N_25365,N_25429);
or U27846 (N_27846,N_25700,N_25781);
and U27847 (N_27847,N_24515,N_24288);
or U27848 (N_27848,N_25175,N_24827);
or U27849 (N_27849,N_25382,N_25292);
xnor U27850 (N_27850,N_24593,N_25504);
nor U27851 (N_27851,N_24606,N_24874);
nor U27852 (N_27852,N_25449,N_25601);
or U27853 (N_27853,N_24708,N_24902);
nor U27854 (N_27854,N_25496,N_25754);
nand U27855 (N_27855,N_25146,N_25000);
or U27856 (N_27856,N_25861,N_25807);
xnor U27857 (N_27857,N_25395,N_25827);
or U27858 (N_27858,N_24851,N_24051);
nand U27859 (N_27859,N_24208,N_25441);
nor U27860 (N_27860,N_25474,N_24600);
nand U27861 (N_27861,N_24959,N_25908);
nor U27862 (N_27862,N_25960,N_24138);
or U27863 (N_27863,N_25760,N_24723);
xnor U27864 (N_27864,N_24030,N_24271);
nor U27865 (N_27865,N_24266,N_25450);
nand U27866 (N_27866,N_24454,N_25956);
nand U27867 (N_27867,N_24470,N_25532);
nand U27868 (N_27868,N_24225,N_25659);
nor U27869 (N_27869,N_25265,N_25501);
nor U27870 (N_27870,N_24285,N_25518);
xnor U27871 (N_27871,N_24226,N_24084);
xnor U27872 (N_27872,N_24153,N_25274);
nor U27873 (N_27873,N_25940,N_25438);
nor U27874 (N_27874,N_24848,N_24661);
xor U27875 (N_27875,N_24302,N_24246);
nor U27876 (N_27876,N_25428,N_24944);
nor U27877 (N_27877,N_24639,N_24492);
and U27878 (N_27878,N_24591,N_24771);
or U27879 (N_27879,N_24997,N_24062);
and U27880 (N_27880,N_25251,N_24677);
and U27881 (N_27881,N_24162,N_24723);
nand U27882 (N_27882,N_25063,N_24231);
and U27883 (N_27883,N_24841,N_24913);
and U27884 (N_27884,N_25327,N_25320);
nand U27885 (N_27885,N_24820,N_25173);
xor U27886 (N_27886,N_25485,N_24075);
or U27887 (N_27887,N_24403,N_24202);
xor U27888 (N_27888,N_25878,N_24873);
nand U27889 (N_27889,N_24330,N_24125);
or U27890 (N_27890,N_25280,N_25542);
and U27891 (N_27891,N_25015,N_24758);
xor U27892 (N_27892,N_25922,N_24001);
nor U27893 (N_27893,N_24243,N_25881);
xnor U27894 (N_27894,N_25663,N_25034);
xnor U27895 (N_27895,N_25787,N_25707);
or U27896 (N_27896,N_25099,N_25973);
or U27897 (N_27897,N_25142,N_24682);
nor U27898 (N_27898,N_24607,N_24465);
nor U27899 (N_27899,N_24358,N_24986);
xor U27900 (N_27900,N_24813,N_25238);
or U27901 (N_27901,N_25154,N_25146);
or U27902 (N_27902,N_24070,N_24583);
or U27903 (N_27903,N_24582,N_24081);
nand U27904 (N_27904,N_24476,N_25662);
or U27905 (N_27905,N_24734,N_24080);
or U27906 (N_27906,N_24031,N_25795);
and U27907 (N_27907,N_24219,N_25813);
nor U27908 (N_27908,N_24802,N_24689);
xor U27909 (N_27909,N_24566,N_24873);
xnor U27910 (N_27910,N_24288,N_24933);
xnor U27911 (N_27911,N_24221,N_24308);
and U27912 (N_27912,N_25367,N_25306);
or U27913 (N_27913,N_25785,N_24054);
and U27914 (N_27914,N_25957,N_25947);
xnor U27915 (N_27915,N_24334,N_25723);
xor U27916 (N_27916,N_24861,N_25515);
or U27917 (N_27917,N_25216,N_25626);
xor U27918 (N_27918,N_24792,N_24451);
and U27919 (N_27919,N_24714,N_25606);
nor U27920 (N_27920,N_24844,N_24340);
or U27921 (N_27921,N_24974,N_25557);
or U27922 (N_27922,N_24430,N_25319);
nor U27923 (N_27923,N_25143,N_25461);
nand U27924 (N_27924,N_25565,N_24585);
nand U27925 (N_27925,N_25200,N_24366);
or U27926 (N_27926,N_25202,N_25751);
nor U27927 (N_27927,N_24351,N_24680);
and U27928 (N_27928,N_25751,N_24930);
nor U27929 (N_27929,N_24466,N_24259);
xor U27930 (N_27930,N_24041,N_25044);
nor U27931 (N_27931,N_24057,N_25154);
or U27932 (N_27932,N_25932,N_24083);
nor U27933 (N_27933,N_25519,N_24954);
xor U27934 (N_27934,N_24502,N_25006);
nand U27935 (N_27935,N_24694,N_24919);
xnor U27936 (N_27936,N_24240,N_24950);
xnor U27937 (N_27937,N_25460,N_25480);
nand U27938 (N_27938,N_24675,N_24440);
and U27939 (N_27939,N_24311,N_25712);
xnor U27940 (N_27940,N_24334,N_25754);
nand U27941 (N_27941,N_25190,N_25239);
or U27942 (N_27942,N_24588,N_24828);
xnor U27943 (N_27943,N_24957,N_25166);
nand U27944 (N_27944,N_25862,N_25327);
and U27945 (N_27945,N_25351,N_24415);
nand U27946 (N_27946,N_24010,N_25005);
nor U27947 (N_27947,N_25569,N_25718);
nor U27948 (N_27948,N_24135,N_24508);
nor U27949 (N_27949,N_24179,N_25119);
or U27950 (N_27950,N_24559,N_24200);
xnor U27951 (N_27951,N_24096,N_24318);
or U27952 (N_27952,N_25578,N_25987);
nor U27953 (N_27953,N_25018,N_25389);
nand U27954 (N_27954,N_24609,N_25533);
nor U27955 (N_27955,N_24674,N_24324);
xor U27956 (N_27956,N_25123,N_24226);
nor U27957 (N_27957,N_25175,N_25548);
xnor U27958 (N_27958,N_24710,N_24374);
nand U27959 (N_27959,N_24949,N_25160);
xnor U27960 (N_27960,N_24584,N_24166);
and U27961 (N_27961,N_24331,N_25623);
nor U27962 (N_27962,N_24603,N_24889);
nand U27963 (N_27963,N_25463,N_25378);
xor U27964 (N_27964,N_25663,N_25013);
nand U27965 (N_27965,N_24622,N_24666);
nor U27966 (N_27966,N_24278,N_24392);
nor U27967 (N_27967,N_24402,N_25925);
and U27968 (N_27968,N_24208,N_24285);
or U27969 (N_27969,N_25386,N_25776);
or U27970 (N_27970,N_24987,N_25747);
and U27971 (N_27971,N_24861,N_25407);
nand U27972 (N_27972,N_24562,N_24115);
and U27973 (N_27973,N_25007,N_25456);
nand U27974 (N_27974,N_25662,N_24885);
or U27975 (N_27975,N_24065,N_24487);
or U27976 (N_27976,N_24677,N_25924);
nor U27977 (N_27977,N_24113,N_24068);
nor U27978 (N_27978,N_24903,N_25707);
and U27979 (N_27979,N_24623,N_24581);
or U27980 (N_27980,N_24299,N_24770);
and U27981 (N_27981,N_24648,N_24928);
xnor U27982 (N_27982,N_25477,N_25957);
xnor U27983 (N_27983,N_24420,N_24137);
or U27984 (N_27984,N_24222,N_24286);
and U27985 (N_27985,N_24892,N_24195);
and U27986 (N_27986,N_25595,N_25649);
xnor U27987 (N_27987,N_25812,N_24047);
and U27988 (N_27988,N_25137,N_25308);
nand U27989 (N_27989,N_24529,N_25374);
or U27990 (N_27990,N_24395,N_24340);
nand U27991 (N_27991,N_24234,N_25543);
nand U27992 (N_27992,N_24007,N_25222);
nand U27993 (N_27993,N_24482,N_24308);
and U27994 (N_27994,N_25273,N_24334);
nand U27995 (N_27995,N_25218,N_24185);
or U27996 (N_27996,N_24152,N_24850);
or U27997 (N_27997,N_24932,N_24270);
or U27998 (N_27998,N_25569,N_25373);
xnor U27999 (N_27999,N_25156,N_24044);
nand U28000 (N_28000,N_26669,N_27307);
xnor U28001 (N_28001,N_26734,N_26027);
nand U28002 (N_28002,N_26288,N_26690);
nor U28003 (N_28003,N_27206,N_27360);
nor U28004 (N_28004,N_27938,N_26930);
nand U28005 (N_28005,N_27973,N_27346);
xnor U28006 (N_28006,N_26228,N_26010);
nor U28007 (N_28007,N_27534,N_26239);
xnor U28008 (N_28008,N_27575,N_27868);
or U28009 (N_28009,N_27474,N_27131);
nand U28010 (N_28010,N_27345,N_26404);
and U28011 (N_28011,N_26525,N_26041);
and U28012 (N_28012,N_27327,N_27633);
nand U28013 (N_28013,N_26061,N_27429);
or U28014 (N_28014,N_26219,N_27304);
and U28015 (N_28015,N_26562,N_27726);
xor U28016 (N_28016,N_26092,N_26126);
nand U28017 (N_28017,N_26028,N_27324);
nand U28018 (N_28018,N_27326,N_26331);
and U28019 (N_28019,N_26012,N_27651);
and U28020 (N_28020,N_26770,N_26391);
nand U28021 (N_28021,N_26082,N_27207);
and U28022 (N_28022,N_27006,N_27836);
and U28023 (N_28023,N_27080,N_27615);
or U28024 (N_28024,N_27754,N_26718);
nor U28025 (N_28025,N_26763,N_27501);
and U28026 (N_28026,N_27662,N_26972);
xnor U28027 (N_28027,N_26801,N_27198);
or U28028 (N_28028,N_26116,N_27912);
xnor U28029 (N_28029,N_27177,N_27533);
and U28030 (N_28030,N_26354,N_26083);
nand U28031 (N_28031,N_26857,N_26453);
or U28032 (N_28032,N_26262,N_26558);
nor U28033 (N_28033,N_27775,N_26425);
xnor U28034 (N_28034,N_27433,N_27881);
xor U28035 (N_28035,N_26242,N_27136);
or U28036 (N_28036,N_27798,N_26385);
nor U28037 (N_28037,N_27144,N_26373);
nand U28038 (N_28038,N_27205,N_27719);
and U28039 (N_28039,N_26468,N_27456);
nand U28040 (N_28040,N_26475,N_26999);
nand U28041 (N_28041,N_26266,N_27493);
nor U28042 (N_28042,N_27088,N_26945);
and U28043 (N_28043,N_27190,N_26106);
or U28044 (N_28044,N_27414,N_27982);
nand U28045 (N_28045,N_26223,N_26896);
nor U28046 (N_28046,N_27029,N_27879);
nor U28047 (N_28047,N_27658,N_27491);
nor U28048 (N_28048,N_26265,N_26034);
nor U28049 (N_28049,N_27022,N_27583);
xor U28050 (N_28050,N_27368,N_27782);
nand U28051 (N_28051,N_26179,N_26470);
xnor U28052 (N_28052,N_26408,N_27652);
or U28053 (N_28053,N_27594,N_27168);
xor U28054 (N_28054,N_27259,N_26814);
and U28055 (N_28055,N_27224,N_26177);
nand U28056 (N_28056,N_26632,N_26103);
or U28057 (N_28057,N_26985,N_26026);
and U28058 (N_28058,N_27860,N_27960);
and U28059 (N_28059,N_26695,N_27415);
or U28060 (N_28060,N_27978,N_27896);
nor U28061 (N_28061,N_27680,N_27592);
and U28062 (N_28062,N_27223,N_27186);
or U28063 (N_28063,N_26381,N_26564);
and U28064 (N_28064,N_27038,N_26943);
or U28065 (N_28065,N_27567,N_26369);
or U28066 (N_28066,N_26352,N_26176);
or U28067 (N_28067,N_26273,N_27257);
xor U28068 (N_28068,N_27508,N_26346);
xnor U28069 (N_28069,N_27361,N_26359);
nor U28070 (N_28070,N_27446,N_26965);
nor U28071 (N_28071,N_26878,N_27473);
nor U28072 (N_28072,N_26893,N_26961);
and U28073 (N_28073,N_26825,N_26421);
nand U28074 (N_28074,N_27396,N_26819);
and U28075 (N_28075,N_27609,N_26949);
and U28076 (N_28076,N_26306,N_27898);
nor U28077 (N_28077,N_26710,N_26807);
xor U28078 (N_28078,N_27490,N_27556);
nand U28079 (N_28079,N_27569,N_27330);
or U28080 (N_28080,N_27820,N_27112);
nor U28081 (N_28081,N_26309,N_26668);
nor U28082 (N_28082,N_27614,N_27777);
xor U28083 (N_28083,N_26339,N_26199);
nand U28084 (N_28084,N_26606,N_26851);
or U28085 (N_28085,N_27664,N_27004);
or U28086 (N_28086,N_26534,N_26481);
xnor U28087 (N_28087,N_27760,N_27020);
or U28088 (N_28088,N_26243,N_27498);
nand U28089 (N_28089,N_27284,N_26701);
and U28090 (N_28090,N_26067,N_26233);
xnor U28091 (N_28091,N_27007,N_26004);
nand U28092 (N_28092,N_26203,N_26080);
nor U28093 (N_28093,N_27591,N_27862);
nand U28094 (N_28094,N_26571,N_27845);
xnor U28095 (N_28095,N_27027,N_26950);
nor U28096 (N_28096,N_27773,N_26341);
and U28097 (N_28097,N_27595,N_26958);
xnor U28098 (N_28098,N_27078,N_26767);
nor U28099 (N_28099,N_26245,N_26717);
xnor U28100 (N_28100,N_27031,N_26161);
or U28101 (N_28101,N_27576,N_27219);
and U28102 (N_28102,N_27215,N_26715);
nand U28103 (N_28103,N_26167,N_27788);
or U28104 (N_28104,N_27638,N_27283);
and U28105 (N_28105,N_27867,N_26058);
and U28106 (N_28106,N_27976,N_27070);
or U28107 (N_28107,N_26327,N_27821);
and U28108 (N_28108,N_27348,N_27518);
xnor U28109 (N_28109,N_27119,N_27656);
or U28110 (N_28110,N_26873,N_26900);
nor U28111 (N_28111,N_27005,N_27333);
or U28112 (N_28112,N_27395,N_26964);
xnor U28113 (N_28113,N_27837,N_26621);
nor U28114 (N_28114,N_27306,N_27099);
nor U28115 (N_28115,N_26235,N_26689);
nor U28116 (N_28116,N_26056,N_27425);
nor U28117 (N_28117,N_26638,N_26656);
or U28118 (N_28118,N_26620,N_26406);
nor U28119 (N_28119,N_27351,N_26944);
or U28120 (N_28120,N_27993,N_26711);
and U28121 (N_28121,N_26224,N_27235);
xor U28122 (N_28122,N_27959,N_26395);
and U28123 (N_28123,N_26109,N_26055);
and U28124 (N_28124,N_27994,N_27364);
and U28125 (N_28125,N_27546,N_26152);
xnor U28126 (N_28126,N_27040,N_26021);
nand U28127 (N_28127,N_27093,N_27374);
nor U28128 (N_28128,N_26051,N_27944);
and U28129 (N_28129,N_26570,N_26741);
or U28130 (N_28130,N_27663,N_26813);
nand U28131 (N_28131,N_26994,N_27786);
and U28132 (N_28132,N_27942,N_26509);
nand U28133 (N_28133,N_26646,N_27016);
nand U28134 (N_28134,N_27694,N_27013);
nand U28135 (N_28135,N_27553,N_27828);
or U28136 (N_28136,N_27890,N_26595);
xnor U28137 (N_28137,N_27061,N_27601);
and U28138 (N_28138,N_26947,N_27443);
xnor U28139 (N_28139,N_26478,N_26434);
nand U28140 (N_28140,N_27248,N_27605);
nor U28141 (N_28141,N_26146,N_26703);
xnor U28142 (N_28142,N_27157,N_26613);
nor U28143 (N_28143,N_27267,N_27757);
xor U28144 (N_28144,N_27417,N_26559);
nor U28145 (N_28145,N_26184,N_27008);
nor U28146 (N_28146,N_27204,N_26102);
nand U28147 (N_28147,N_27386,N_26450);
xnor U28148 (N_28148,N_27041,N_27162);
and U28149 (N_28149,N_27827,N_26754);
and U28150 (N_28150,N_26438,N_27412);
or U28151 (N_28151,N_26738,N_26441);
nand U28152 (N_28152,N_26025,N_27011);
nand U28153 (N_28153,N_26119,N_27671);
nand U28154 (N_28154,N_26447,N_26859);
xnor U28155 (N_28155,N_27557,N_27402);
or U28156 (N_28156,N_27289,N_27649);
nand U28157 (N_28157,N_27668,N_26956);
nor U28158 (N_28158,N_27264,N_27064);
xnor U28159 (N_28159,N_27154,N_26660);
nor U28160 (N_28160,N_26540,N_26719);
nand U28161 (N_28161,N_27627,N_26039);
nand U28162 (N_28162,N_26334,N_27953);
or U28163 (N_28163,N_26452,N_26128);
and U28164 (N_28164,N_26636,N_26072);
and U28165 (N_28165,N_26898,N_26618);
nor U28166 (N_28166,N_26993,N_27916);
or U28167 (N_28167,N_26680,N_27140);
and U28168 (N_28168,N_27126,N_26091);
nor U28169 (N_28169,N_27675,N_27794);
nor U28170 (N_28170,N_26019,N_27435);
nor U28171 (N_28171,N_27158,N_26388);
or U28172 (N_28172,N_27072,N_26508);
nand U28173 (N_28173,N_27106,N_26123);
and U28174 (N_28174,N_26410,N_26329);
nor U28175 (N_28175,N_27428,N_26370);
xnor U28176 (N_28176,N_27536,N_27081);
nor U28177 (N_28177,N_26237,N_26979);
xor U28178 (N_28178,N_27956,N_26784);
and U28179 (N_28179,N_26166,N_27923);
nand U28180 (N_28180,N_26350,N_27839);
or U28181 (N_28181,N_26557,N_27236);
and U28182 (N_28182,N_27957,N_27350);
xor U28183 (N_28183,N_27643,N_27297);
or U28184 (N_28184,N_26952,N_27104);
or U28185 (N_28185,N_27515,N_26220);
and U28186 (N_28186,N_27046,N_27288);
or U28187 (N_28187,N_26882,N_26727);
or U28188 (N_28188,N_26696,N_26845);
and U28189 (N_28189,N_27098,N_26264);
nand U28190 (N_28190,N_27657,N_26712);
xnor U28191 (N_28191,N_26476,N_26333);
nand U28192 (N_28192,N_27927,N_27111);
nand U28193 (N_28193,N_27914,N_26749);
or U28194 (N_28194,N_27679,N_26657);
xnor U28195 (N_28195,N_26778,N_26886);
xor U28196 (N_28196,N_27060,N_26629);
or U28197 (N_28197,N_26218,N_27850);
xor U28198 (N_28198,N_26572,N_27193);
xor U28199 (N_28199,N_27813,N_26008);
or U28200 (N_28200,N_27621,N_26742);
and U28201 (N_28201,N_26105,N_27066);
xor U28202 (N_28202,N_27547,N_27908);
and U28203 (N_28203,N_27571,N_27385);
xnor U28204 (N_28204,N_27139,N_26474);
nor U28205 (N_28205,N_27108,N_26609);
nand U28206 (N_28206,N_26885,N_27859);
or U28207 (N_28207,N_27150,N_26820);
xor U28208 (N_28208,N_26962,N_27378);
nand U28209 (N_28209,N_27838,N_27966);
and U28210 (N_28210,N_26420,N_27875);
and U28211 (N_28211,N_27520,N_27308);
or U28212 (N_28212,N_27573,N_27639);
or U28213 (N_28213,N_26661,N_26210);
nor U28214 (N_28214,N_26036,N_26101);
and U28215 (N_28215,N_26217,N_27199);
and U28216 (N_28216,N_26066,N_26337);
or U28217 (N_28217,N_27631,N_27612);
or U28218 (N_28218,N_27018,N_27929);
or U28219 (N_28219,N_27143,N_26533);
nor U28220 (N_28220,N_27115,N_26358);
nor U28221 (N_28221,N_27870,N_27458);
nor U28222 (N_28222,N_27053,N_26463);
or U28223 (N_28223,N_27359,N_26267);
or U28224 (N_28224,N_27864,N_26422);
xor U28225 (N_28225,N_26811,N_26673);
nand U28226 (N_28226,N_26035,N_27783);
nor U28227 (N_28227,N_27497,N_26204);
and U28228 (N_28228,N_27033,N_27389);
nor U28229 (N_28229,N_26043,N_26495);
or U28230 (N_28230,N_26976,N_26760);
xnor U28231 (N_28231,N_26249,N_26111);
xnor U28232 (N_28232,N_26650,N_27030);
nand U28233 (N_28233,N_27382,N_26589);
and U28234 (N_28234,N_27911,N_27021);
nand U28235 (N_28235,N_26926,N_27684);
nand U28236 (N_28236,N_27271,N_27634);
nand U28237 (N_28237,N_27701,N_26785);
nor U28238 (N_28238,N_26132,N_27092);
or U28239 (N_28239,N_26003,N_26662);
or U28240 (N_28240,N_26454,N_27468);
nand U28241 (N_28241,N_26097,N_27874);
nor U28242 (N_28242,N_27863,N_27347);
nor U28243 (N_28243,N_27450,N_26160);
nor U28244 (N_28244,N_27313,N_26140);
nor U28245 (N_28245,N_26577,N_26877);
and U28246 (N_28246,N_26075,N_26020);
or U28247 (N_28247,N_27921,N_26351);
nor U28248 (N_28248,N_27209,N_26290);
and U28249 (N_28249,N_26969,N_26295);
and U28250 (N_28250,N_27528,N_26940);
xor U28251 (N_28251,N_27525,N_26604);
nor U28252 (N_28252,N_26776,N_26430);
xor U28253 (N_28253,N_26340,N_27265);
xnor U28254 (N_28254,N_26681,N_27950);
nor U28255 (N_28255,N_27220,N_27165);
or U28256 (N_28256,N_27281,N_26552);
and U28257 (N_28257,N_26085,N_26183);
or U28258 (N_28258,N_27384,N_26162);
and U28259 (N_28259,N_26854,N_27105);
xnor U28260 (N_28260,N_26464,N_27065);
nand U28261 (N_28261,N_27241,N_26610);
xnor U28262 (N_28262,N_26906,N_26390);
xnor U28263 (N_28263,N_26612,N_26578);
and U28264 (N_28264,N_27856,N_27654);
or U28265 (N_28265,N_27991,N_26551);
nor U28266 (N_28266,N_27900,N_27464);
xor U28267 (N_28267,N_26221,N_27544);
and U28268 (N_28268,N_27787,N_26136);
nand U28269 (N_28269,N_26743,N_27214);
nor U28270 (N_28270,N_26207,N_27230);
or U28271 (N_28271,N_27357,N_27972);
and U28272 (N_28272,N_27660,N_26225);
nand U28273 (N_28273,N_27231,N_26556);
and U28274 (N_28274,N_27985,N_27685);
or U28275 (N_28275,N_27640,N_26174);
xnor U28276 (N_28276,N_27502,N_27507);
or U28277 (N_28277,N_26732,N_27829);
nor U28278 (N_28278,N_26922,N_27211);
nor U28279 (N_28279,N_27512,N_26448);
and U28280 (N_28280,N_26587,N_26110);
nor U28281 (N_28281,N_26512,N_27596);
nand U28282 (N_28282,N_27312,N_26586);
and U28283 (N_28283,N_26250,N_27328);
nor U28284 (N_28284,N_26403,N_26625);
and U28285 (N_28285,N_26175,N_27620);
nand U28286 (N_28286,N_27731,N_27700);
nand U28287 (N_28287,N_27965,N_26486);
or U28288 (N_28288,N_26821,N_27784);
nand U28289 (N_28289,N_27262,N_26196);
nand U28290 (N_28290,N_26460,N_27465);
nor U28291 (N_28291,N_27076,N_27320);
or U28292 (N_28292,N_27550,N_27413);
nand U28293 (N_28293,N_27800,N_27579);
nor U28294 (N_28294,N_26984,N_27954);
nor U28295 (N_28295,N_27290,N_26686);
or U28296 (N_28296,N_26550,N_27739);
or U28297 (N_28297,N_27683,N_27296);
xor U28298 (N_28298,N_26530,N_27925);
and U28299 (N_28299,N_26921,N_27311);
nand U28300 (N_28300,N_26676,N_26433);
xor U28301 (N_28301,N_26721,N_27617);
nor U28302 (N_28302,N_26929,N_27689);
nor U28303 (N_28303,N_26096,N_26757);
xnor U28304 (N_28304,N_27164,N_27260);
xor U28305 (N_28305,N_26594,N_27682);
nand U28306 (N_28306,N_27509,N_27492);
or U28307 (N_28307,N_27511,N_27762);
nand U28308 (N_28308,N_26484,N_26059);
and U28309 (N_28309,N_26674,N_27979);
nor U28310 (N_28310,N_26479,N_27125);
nor U28311 (N_28311,N_27756,N_27980);
nand U28312 (N_28312,N_26108,N_26318);
and U28313 (N_28313,N_26431,N_26321);
xnor U28314 (N_28314,N_27253,N_27009);
or U28315 (N_28315,N_26688,N_27276);
and U28316 (N_28316,N_26054,N_26465);
nand U28317 (N_28317,N_26643,N_27728);
xnor U28318 (N_28318,N_26368,N_26371);
xnor U28319 (N_28319,N_26436,N_27721);
nor U28320 (N_28320,N_26623,N_26914);
xnor U28321 (N_28321,N_27866,N_27645);
nor U28322 (N_28322,N_26649,N_27842);
nand U28323 (N_28323,N_26030,N_26153);
nor U28324 (N_28324,N_26714,N_27790);
and U28325 (N_28325,N_26605,N_27603);
or U28326 (N_28326,N_26575,N_27861);
nor U28327 (N_28327,N_27884,N_27826);
or U28328 (N_28328,N_26029,N_26678);
nor U28329 (N_28329,N_26222,N_27763);
nand U28330 (N_28330,N_27734,N_26280);
xnor U28331 (N_28331,N_26457,N_27059);
and U28332 (N_28332,N_27404,N_26156);
xnor U28333 (N_28333,N_27895,N_26378);
and U28334 (N_28334,N_27319,N_26251);
xnor U28335 (N_28335,N_27321,N_26771);
or U28336 (N_28336,N_26342,N_26942);
nand U28337 (N_28337,N_27818,N_26655);
xnor U28338 (N_28338,N_27765,N_26833);
and U28339 (N_28339,N_27750,N_27147);
xor U28340 (N_28340,N_26762,N_26169);
xor U28341 (N_28341,N_26538,N_27755);
nand U28342 (N_28342,N_27623,N_27949);
and U28343 (N_28343,N_27452,N_26302);
nor U28344 (N_28344,N_26903,N_26006);
xor U28345 (N_28345,N_26974,N_27766);
nand U28346 (N_28346,N_26442,N_27145);
or U28347 (N_28347,N_26797,N_26535);
and U28348 (N_28348,N_27709,N_27153);
or U28349 (N_28349,N_27727,N_27738);
xor U28350 (N_28350,N_26081,N_27703);
xor U28351 (N_28351,N_26279,N_27258);
nor U28352 (N_28352,N_27733,N_27607);
nor U28353 (N_28353,N_26355,N_26895);
nand U28354 (N_28354,N_27032,N_27920);
or U28355 (N_28355,N_27202,N_26305);
xor U28356 (N_28356,N_27695,N_26308);
nand U28357 (N_28357,N_26875,N_27876);
xnor U28358 (N_28358,N_26047,N_26723);
nor U28359 (N_28359,N_26752,N_26322);
and U28360 (N_28360,N_26444,N_27941);
or U28361 (N_28361,N_26393,N_26115);
nor U28362 (N_28362,N_27353,N_26642);
nand U28363 (N_28363,N_27442,N_26236);
nor U28364 (N_28364,N_27858,N_26543);
and U28365 (N_28365,N_26573,N_27341);
xor U28366 (N_28366,N_26451,N_27155);
or U28367 (N_28367,N_27432,N_26756);
nand U28368 (N_28368,N_26829,N_27272);
xor U28369 (N_28369,N_26936,N_26073);
xor U28370 (N_28370,N_26205,N_27363);
xor U28371 (N_28371,N_26170,N_27852);
and U28372 (N_28372,N_26443,N_26913);
and U28373 (N_28373,N_27940,N_26931);
xor U28374 (N_28374,N_27778,N_26528);
nand U28375 (N_28375,N_26858,N_26517);
or U28376 (N_28376,N_26848,N_27372);
and U28377 (N_28377,N_27554,N_26736);
nor U28378 (N_28378,N_26000,N_26211);
nand U28379 (N_28379,N_26198,N_27725);
nor U28380 (N_28380,N_27208,N_27323);
xnor U28381 (N_28381,N_27012,N_26614);
xor U28382 (N_28382,N_26602,N_26876);
and U28383 (N_28383,N_26315,N_26496);
xnor U28384 (N_28384,N_27977,N_27809);
nor U28385 (N_28385,N_27924,N_27463);
nor U28386 (N_28386,N_26654,N_26013);
nand U28387 (N_28387,N_26815,N_26951);
xnor U28388 (N_28388,N_27655,N_27872);
nand U28389 (N_28389,N_27928,N_27948);
xnor U28390 (N_28390,N_27537,N_26981);
and U28391 (N_28391,N_26440,N_26970);
or U28392 (N_28392,N_27134,N_26180);
nand U28393 (N_28393,N_26568,N_27411);
nor U28394 (N_28394,N_27229,N_27722);
xnor U28395 (N_28395,N_27023,N_26705);
nand U28396 (N_28396,N_26042,N_27988);
nor U28397 (N_28397,N_26720,N_26089);
xor U28398 (N_28398,N_26159,N_27124);
or U28399 (N_28399,N_26700,N_26044);
xnor U28400 (N_28400,N_26363,N_27849);
nor U28401 (N_28401,N_26399,N_26018);
or U28402 (N_28402,N_26692,N_26310);
and U28403 (N_28403,N_27201,N_27892);
or U28404 (N_28404,N_26933,N_27622);
xnor U28405 (N_28405,N_27101,N_27275);
xnor U28406 (N_28406,N_26955,N_26033);
nand U28407 (N_28407,N_27055,N_27299);
xnor U28408 (N_28408,N_26652,N_27999);
or U28409 (N_28409,N_27901,N_27251);
nor U28410 (N_28410,N_27865,N_27744);
nand U28411 (N_28411,N_26015,N_27844);
or U28412 (N_28412,N_27833,N_27650);
or U28413 (N_28413,N_27878,N_27888);
nand U28414 (N_28414,N_26675,N_27130);
xnor U28415 (N_28415,N_26255,N_26832);
or U28416 (N_28416,N_26500,N_26076);
or U28417 (N_28417,N_26232,N_26792);
nand U28418 (N_28418,N_27613,N_26432);
nand U28419 (N_28419,N_27362,N_26413);
and U28420 (N_28420,N_26397,N_27871);
and U28421 (N_28421,N_27397,N_27517);
and U28422 (N_28422,N_27522,N_27574);
or U28423 (N_28423,N_27698,N_27529);
and U28424 (N_28424,N_27071,N_26531);
or U28425 (N_28425,N_26758,N_26163);
xor U28426 (N_28426,N_27388,N_26745);
nand U28427 (N_28427,N_27217,N_27477);
nor U28428 (N_28428,N_26423,N_27172);
and U28429 (N_28429,N_27713,N_26995);
nand U28430 (N_28430,N_26835,N_27770);
nor U28431 (N_28431,N_26935,N_27799);
or U28432 (N_28432,N_27670,N_26511);
nor U28433 (N_28433,N_27095,N_26915);
nand U28434 (N_28434,N_26149,N_26488);
and U28435 (N_28435,N_27692,N_27049);
or U28436 (N_28436,N_26826,N_27527);
nor U28437 (N_28437,N_26164,N_27805);
or U28438 (N_28438,N_27880,N_27759);
and U28439 (N_28439,N_27810,N_26185);
nand U28440 (N_28440,N_27286,N_27459);
and U28441 (N_28441,N_26702,N_26640);
or U28442 (N_28442,N_26281,N_27171);
nor U28443 (N_28443,N_26287,N_27637);
nor U28444 (N_28444,N_27904,N_26987);
nor U28445 (N_28445,N_27699,N_27356);
nor U28446 (N_28446,N_26356,N_26611);
nand U28447 (N_28447,N_27048,N_26869);
or U28448 (N_28448,N_27203,N_26114);
nand U28449 (N_28449,N_26852,N_27947);
and U28450 (N_28450,N_26192,N_27636);
nor U28451 (N_28451,N_26889,N_26923);
and U28452 (N_28452,N_27624,N_27945);
or U28453 (N_28453,N_27292,N_27365);
or U28454 (N_28454,N_27376,N_26842);
or U28455 (N_28455,N_26394,N_27846);
xnor U28456 (N_28456,N_26259,N_26800);
nand U28457 (N_28457,N_26002,N_27371);
nor U28458 (N_28458,N_26565,N_26616);
or U28459 (N_28459,N_26831,N_27641);
nor U28460 (N_28460,N_27019,N_26907);
xor U28461 (N_28461,N_27398,N_26206);
and U28462 (N_28462,N_26435,N_26908);
xnor U28463 (N_28463,N_27882,N_27740);
nand U28464 (N_28464,N_27984,N_26887);
xor U28465 (N_28465,N_26840,N_26761);
nand U28466 (N_28466,N_27077,N_27975);
xor U28467 (N_28467,N_27427,N_27097);
or U28468 (N_28468,N_27513,N_27524);
nand U28469 (N_28469,N_26596,N_26986);
nor U28470 (N_28470,N_26560,N_26816);
xnor U28471 (N_28471,N_26546,N_27669);
nor U28472 (N_28472,N_26781,N_26554);
nor U28473 (N_28473,N_27934,N_26968);
or U28474 (N_28474,N_27189,N_26079);
and U28475 (N_28475,N_26338,N_26261);
nand U28476 (N_28476,N_27560,N_27337);
nand U28477 (N_28477,N_26843,N_27416);
xor U28478 (N_28478,N_27996,N_26897);
nand U28479 (N_28479,N_26181,N_27387);
or U28480 (N_28480,N_26195,N_27310);
xnor U28481 (N_28481,N_27243,N_26849);
and U28482 (N_28482,N_26467,N_27316);
xor U28483 (N_28483,N_27843,N_26585);
xor U28484 (N_28484,N_26093,N_27056);
nand U28485 (N_28485,N_26317,N_26687);
nor U28486 (N_28486,N_27226,N_27752);
nor U28487 (N_28487,N_27937,N_27221);
nand U28488 (N_28488,N_26301,N_27510);
nor U28489 (N_28489,N_26473,N_27089);
nand U28490 (N_28490,N_27291,N_27747);
or U28491 (N_28491,N_26437,N_26490);
or U28492 (N_28492,N_26014,N_26747);
and U28493 (N_28493,N_27577,N_27373);
nor U28494 (N_28494,N_27545,N_27210);
nor U28495 (N_28495,N_26418,N_27562);
and U28496 (N_28496,N_26822,N_27015);
xnor U28497 (N_28497,N_27789,N_26375);
nand U28498 (N_28498,N_27173,N_27887);
and U28499 (N_28499,N_26118,N_26284);
nor U28500 (N_28500,N_27690,N_26409);
nand U28501 (N_28501,N_27218,N_26989);
nor U28502 (N_28502,N_27822,N_26601);
and U28503 (N_28503,N_27050,N_27107);
nand U28504 (N_28504,N_27855,N_27602);
nand U28505 (N_28505,N_26412,N_26260);
and U28506 (N_28506,N_26635,N_26803);
or U28507 (N_28507,N_27516,N_26663);
and U28508 (N_28508,N_27714,N_26240);
nor U28509 (N_28509,N_26307,N_26545);
and U28510 (N_28510,N_26619,N_27303);
xor U28511 (N_28511,N_27572,N_27906);
nand U28512 (N_28512,N_26499,N_27840);
nand U28513 (N_28513,N_27399,N_26839);
or U28514 (N_28514,N_26045,N_26365);
xnor U28515 (N_28515,N_27133,N_26074);
and U28516 (N_28516,N_27903,N_27246);
nand U28517 (N_28517,N_27677,N_26173);
nor U28518 (N_28518,N_26168,N_26521);
and U28519 (N_28519,N_26874,N_26086);
nand U28520 (N_28520,N_26783,N_26729);
xnor U28521 (N_28521,N_26286,N_27628);
nand U28522 (N_28522,N_26569,N_26300);
and U28523 (N_28523,N_26855,N_26401);
and U28524 (N_28524,N_27058,N_27268);
nand U28525 (N_28525,N_27034,N_26349);
nor U28526 (N_28526,N_26155,N_27503);
or U28527 (N_28527,N_27899,N_27263);
xnor U28528 (N_28528,N_27611,N_26750);
nor U28529 (N_28529,N_27717,N_27051);
and U28530 (N_28530,N_26107,N_26542);
nor U28531 (N_28531,N_27437,N_26294);
or U28532 (N_28532,N_27256,N_26201);
and U28533 (N_28533,N_26664,N_27659);
nand U28534 (N_28534,N_26725,N_26005);
xor U28535 (N_28535,N_27405,N_26319);
nor U28536 (N_28536,N_27767,N_26501);
and U28537 (N_28537,N_26891,N_27873);
and U28538 (N_28538,N_26050,N_27819);
and U28539 (N_28539,N_26634,N_27723);
or U28540 (N_28540,N_27943,N_26384);
nand U28541 (N_28541,N_26847,N_27197);
or U28542 (N_28542,N_27295,N_27803);
nand U28543 (N_28543,N_27678,N_27600);
nand U28544 (N_28544,N_26186,N_26100);
and U28545 (N_28545,N_26130,N_27715);
or U28546 (N_28546,N_27000,N_26038);
nor U28547 (N_28547,N_27082,N_26960);
nand U28548 (N_28548,N_26812,N_27280);
nor U28549 (N_28549,N_26314,N_26275);
nor U28550 (N_28550,N_26407,N_26624);
nand U28551 (N_28551,N_27110,N_26326);
or U28552 (N_28552,N_27588,N_26780);
and U28553 (N_28553,N_27665,N_26347);
nand U28554 (N_28554,N_26890,N_26238);
xor U28555 (N_28555,N_26793,N_27377);
xor U28556 (N_28556,N_27538,N_26791);
xor U28557 (N_28557,N_27630,N_26157);
xor U28558 (N_28558,N_27806,N_27094);
and U28559 (N_28559,N_27294,N_27815);
nand U28560 (N_28560,N_26297,N_26178);
nand U28561 (N_28561,N_27245,N_26544);
xnor U28562 (N_28562,N_27393,N_27068);
and U28563 (N_28563,N_26483,N_27604);
and U28564 (N_28564,N_27952,N_27240);
and U28565 (N_28565,N_27779,N_26806);
nand U28566 (N_28566,N_26311,N_27174);
or U28567 (N_28567,N_26182,N_26805);
nand U28568 (N_28568,N_26052,N_26303);
xor U28569 (N_28569,N_26997,N_27455);
and U28570 (N_28570,N_26212,N_27768);
nor U28571 (N_28571,N_27933,N_26866);
and U28572 (N_28572,N_27551,N_26131);
and U28573 (N_28573,N_27249,N_27039);
or U28574 (N_28574,N_27394,N_27531);
or U28575 (N_28575,N_27042,N_26060);
and U28576 (N_28576,N_27519,N_26298);
or U28577 (N_28577,N_26834,N_26491);
nor U28578 (N_28578,N_27237,N_27983);
or U28579 (N_28579,N_27420,N_26292);
nand U28580 (N_28580,N_27225,N_26520);
nand U28581 (N_28581,N_27749,N_27499);
or U28582 (N_28582,N_27824,N_26285);
and U28583 (N_28583,N_27475,N_27795);
or U28584 (N_28584,N_26023,N_27057);
nor U28585 (N_28585,N_26257,N_26379);
or U28586 (N_28586,N_26017,N_27730);
xor U28587 (N_28587,N_26838,N_27269);
and U28588 (N_28588,N_26730,N_26497);
nand U28589 (N_28589,N_27370,N_27793);
xnor U28590 (N_28590,N_26117,N_26272);
nor U28591 (N_28591,N_26667,N_27802);
xor U28592 (N_28592,N_27279,N_27079);
nor U28593 (N_28593,N_27460,N_26009);
xor U28594 (N_28594,N_27073,N_27471);
xor U28595 (N_28595,N_26069,N_26104);
or U28596 (N_28596,N_27761,N_26064);
or U28597 (N_28597,N_27808,N_27687);
or U28598 (N_28598,N_26603,N_27480);
and U28599 (N_28599,N_27542,N_27122);
nor U28600 (N_28600,N_27751,N_27932);
xor U28601 (N_28601,N_26429,N_26902);
xnor U28602 (N_28602,N_26120,N_27084);
nand U28603 (N_28603,N_27024,N_26909);
xor U28604 (N_28604,N_26651,N_27247);
or U28605 (N_28605,N_27814,N_27963);
nor U28606 (N_28606,N_27392,N_27200);
or U28607 (N_28607,N_27891,N_27710);
or U28608 (N_28608,N_27159,N_26607);
nand U28609 (N_28609,N_26971,N_26597);
nor U28610 (N_28610,N_27801,N_27585);
or U28611 (N_28611,N_26622,N_27804);
nand U28612 (N_28612,N_27342,N_27811);
or U28613 (N_28613,N_27629,N_26683);
or U28614 (N_28614,N_27851,N_26948);
xor U28615 (N_28615,N_27736,N_27085);
xnor U28616 (N_28616,N_27825,N_27261);
xor U28617 (N_28617,N_27302,N_26098);
nand U28618 (N_28618,N_26522,N_26316);
xnor U28619 (N_28619,N_27135,N_27129);
nor U28620 (N_28620,N_26584,N_27010);
or U28621 (N_28621,N_26234,N_26366);
and U28622 (N_28622,N_26548,N_27449);
and U28623 (N_28623,N_26063,N_27103);
or U28624 (N_28624,N_27381,N_27113);
xor U28625 (N_28625,N_27939,N_27436);
nand U28626 (N_28626,N_27448,N_27403);
or U28627 (N_28627,N_26510,N_26916);
and U28628 (N_28628,N_26343,N_26458);
nor U28629 (N_28629,N_27278,N_26959);
nor U28630 (N_28630,N_26498,N_26647);
or U28631 (N_28631,N_26532,N_26879);
and U28632 (N_28632,N_27478,N_27044);
and U28633 (N_28633,N_26731,N_26256);
or U28634 (N_28634,N_27653,N_27543);
nand U28635 (N_28635,N_26764,N_26513);
nor U28636 (N_28636,N_27383,N_26871);
xnor U28637 (N_28637,N_26449,N_26645);
nor U28638 (N_28638,N_26946,N_27964);
nor U28639 (N_28639,N_26505,N_27191);
or U28640 (N_28640,N_26697,N_27486);
nand U28641 (N_28641,N_27329,N_26053);
and U28642 (N_28642,N_26320,N_27315);
and U28643 (N_28643,N_27505,N_27792);
and U28644 (N_28644,N_27910,N_26737);
nor U28645 (N_28645,N_26988,N_26230);
nand U28646 (N_28646,N_26046,N_27148);
nand U28647 (N_28647,N_26446,N_27841);
or U28648 (N_28648,N_27610,N_26828);
or U28649 (N_28649,N_26912,N_26924);
or U28650 (N_28650,N_26677,N_27549);
xor U28651 (N_28651,N_26514,N_27857);
nor U28652 (N_28652,N_26049,N_27325);
nor U28653 (N_28653,N_26911,N_26925);
nor U28654 (N_28654,N_26617,N_26519);
nand U28655 (N_28655,N_26990,N_27091);
or U28656 (N_28656,N_26172,N_26348);
or U28657 (N_28657,N_27581,N_27293);
and U28658 (N_28658,N_26894,N_27816);
and U28659 (N_28659,N_27674,N_26283);
xnor U28660 (N_28660,N_27180,N_26593);
xnor U28661 (N_28661,N_26837,N_26031);
xnor U28662 (N_28662,N_26576,N_26862);
xor U28663 (N_28663,N_27222,N_26065);
nand U28664 (N_28664,N_27913,N_27746);
nand U28665 (N_28665,N_27003,N_26967);
xnor U28666 (N_28666,N_27632,N_26274);
nand U28667 (N_28667,N_26229,N_26376);
or U28668 (N_28668,N_27479,N_26127);
nor U28669 (N_28669,N_27424,N_26405);
nand U28670 (N_28670,N_26860,N_26296);
nor U28671 (N_28671,N_27541,N_26555);
or U28672 (N_28672,N_27423,N_27618);
xor U28673 (N_28673,N_26753,N_27036);
and U28674 (N_28674,N_27444,N_26567);
xnor U28675 (N_28675,N_27339,N_27673);
or U28676 (N_28676,N_26057,N_26901);
nor U28677 (N_28677,N_26024,N_27274);
and U28678 (N_28678,N_26278,N_26214);
xor U28679 (N_28679,N_26599,N_26809);
xor U28680 (N_28680,N_27255,N_27232);
xnor U28681 (N_28681,N_26765,N_27183);
and U28682 (N_28682,N_26087,N_27626);
nand U28683 (N_28683,N_27409,N_27681);
or U28684 (N_28684,N_27907,N_26938);
or U28685 (N_28685,N_26466,N_27495);
or U28686 (N_28686,N_27885,N_27971);
nor U28687 (N_28687,N_27848,N_26299);
nand U28688 (N_28688,N_27379,N_26377);
and U28689 (N_28689,N_27322,N_26539);
nand U28690 (N_28690,N_26291,N_27935);
nor U28691 (N_28691,N_26480,N_26095);
nand U28692 (N_28692,N_26853,N_26150);
nor U28693 (N_28693,N_27332,N_26628);
or U28694 (N_28694,N_27213,N_27946);
or U28695 (N_28695,N_26707,N_26188);
nand U28696 (N_28696,N_27270,N_26526);
or U28697 (N_28697,N_27776,N_26637);
and U28698 (N_28698,N_26980,N_26094);
xnor U28699 (N_28699,N_26920,N_27561);
nand U28700 (N_28700,N_27354,N_26361);
xor U28701 (N_28701,N_26134,N_27149);
and U28702 (N_28702,N_27599,N_26615);
nand U28703 (N_28703,N_26827,N_26455);
and U28704 (N_28704,N_27266,N_26957);
and U28705 (N_28705,N_26864,N_26588);
or U28706 (N_28706,N_26824,N_26581);
and U28707 (N_28707,N_27758,N_26208);
nand U28708 (N_28708,N_26187,N_26367);
nand U28709 (N_28709,N_27184,N_26336);
nand U28710 (N_28710,N_27035,N_27074);
xnor U28711 (N_28711,N_27336,N_27883);
and U28712 (N_28712,N_27242,N_26641);
xnor U28713 (N_28713,N_27062,N_26398);
xnor U28714 (N_28714,N_26580,N_26716);
xor U28715 (N_28715,N_26427,N_26068);
and U28716 (N_28716,N_27711,N_27485);
xnor U28717 (N_28717,N_27028,N_27466);
xor U28718 (N_28718,N_26653,N_27096);
nor U28719 (N_28719,N_26215,N_26328);
xor U28720 (N_28720,N_27797,N_27067);
nand U28721 (N_28721,N_27285,N_26389);
nor U28722 (N_28722,N_27548,N_26563);
nor U28723 (N_28723,N_27440,N_27462);
and U28724 (N_28724,N_27566,N_26194);
nor U28725 (N_28725,N_26865,N_26518);
and U28726 (N_28726,N_27318,N_27555);
nor U28727 (N_28727,N_26934,N_26590);
and U28728 (N_28728,N_26973,N_26414);
and U28729 (N_28729,N_27422,N_27047);
or U28730 (N_28730,N_26751,N_26802);
and U28731 (N_28731,N_27457,N_26592);
xnor U28732 (N_28732,N_27743,N_27301);
nor U28733 (N_28733,N_27877,N_27791);
nand U28734 (N_28734,N_26932,N_27244);
xnor U28735 (N_28735,N_27568,N_27421);
nor U28736 (N_28736,N_27893,N_26090);
nor U28737 (N_28737,N_26277,N_27445);
nand U28738 (N_28738,N_27239,N_27451);
nand U28739 (N_28739,N_27990,N_27832);
nor U28740 (N_28740,N_26304,N_26158);
or U28741 (N_28741,N_27188,N_27407);
nor U28742 (N_28742,N_26032,N_26506);
nand U28743 (N_28743,N_27748,N_27704);
xnor U28744 (N_28744,N_26462,N_27123);
xnor U28745 (N_28745,N_26387,N_27521);
xnor U28746 (N_28746,N_26786,N_26121);
or U28747 (N_28747,N_26788,N_26227);
and U28748 (N_28748,N_26537,N_27227);
and U28749 (N_28749,N_27812,N_26818);
nand U28750 (N_28750,N_27535,N_27968);
nor U28751 (N_28751,N_27441,N_27706);
nand U28752 (N_28752,N_27598,N_27506);
xor U28753 (N_28753,N_27936,N_27915);
nor U28754 (N_28754,N_26541,N_27483);
nor U28755 (N_28755,N_26870,N_27083);
nand U28756 (N_28756,N_26529,N_26863);
nor U28757 (N_28757,N_27772,N_27305);
xnor U28758 (N_28758,N_26503,N_26561);
and U28759 (N_28759,N_26966,N_26939);
xnor U28760 (N_28760,N_26527,N_26774);
and U28761 (N_28761,N_26810,N_26639);
nor U28762 (N_28762,N_27181,N_27593);
or U28763 (N_28763,N_27166,N_26728);
nand U28764 (N_28764,N_27391,N_27228);
and U28765 (N_28765,N_27234,N_27273);
nand U28766 (N_28766,N_26790,N_27408);
nor U28767 (N_28767,N_26709,N_27358);
nand U28768 (N_28768,N_27559,N_26644);
nor U28769 (N_28769,N_27587,N_27369);
or U28770 (N_28770,N_26516,N_27063);
and U28771 (N_28771,N_26691,N_26982);
nor U28772 (N_28772,N_26088,N_26904);
or U28773 (N_28773,N_27419,N_26485);
nand U28774 (N_28774,N_27367,N_26963);
nand U28775 (N_28775,N_26954,N_27277);
nor U28776 (N_28776,N_27586,N_27484);
xnor U28777 (N_28777,N_26154,N_27995);
and U28778 (N_28778,N_27889,N_27494);
and U28779 (N_28779,N_26247,N_26372);
nor U28780 (N_28780,N_26417,N_27697);
and U28781 (N_28781,N_27334,N_26775);
nand U28782 (N_28782,N_26600,N_27514);
xor U28783 (N_28783,N_26216,N_27608);
nand U28784 (N_28784,N_26928,N_27922);
nor U28785 (N_28785,N_26658,N_26608);
nand U28786 (N_28786,N_26996,N_27335);
nand U28787 (N_28787,N_27087,N_26129);
xnor U28788 (N_28788,N_27781,N_27647);
and U28789 (N_28789,N_27905,N_27118);
xor U28790 (N_28790,N_27558,N_27539);
or U28791 (N_28791,N_27967,N_27834);
and U28792 (N_28792,N_27931,N_26553);
xor U28793 (N_28793,N_26124,N_26048);
nand U28794 (N_28794,N_27469,N_26574);
xnor U28795 (N_28795,N_26627,N_27917);
or U28796 (N_28796,N_26927,N_26953);
and U28797 (N_28797,N_27720,N_27691);
nand U28798 (N_28798,N_26746,N_26733);
and U28799 (N_28799,N_26193,N_27708);
nor U28800 (N_28800,N_27667,N_27597);
or U28801 (N_28801,N_26789,N_27926);
or U28802 (N_28802,N_27500,N_27998);
and U28803 (N_28803,N_26808,N_26415);
nor U28804 (N_28804,N_27054,N_26144);
or U28805 (N_28805,N_27981,N_26416);
or U28806 (N_28806,N_27400,N_26631);
xor U28807 (N_28807,N_26748,N_27026);
xor U28808 (N_28808,N_26293,N_26200);
xnor U28809 (N_28809,N_26844,N_27737);
xor U28810 (N_28810,N_27109,N_26536);
xnor U28811 (N_28811,N_26037,N_26489);
nand U28812 (N_28812,N_26252,N_27349);
and U28813 (N_28813,N_26492,N_26312);
and U28814 (N_28814,N_27380,N_26892);
or U28815 (N_28815,N_26330,N_26364);
nor U28816 (N_28816,N_26487,N_26910);
or U28817 (N_28817,N_27418,N_27447);
and U28818 (N_28818,N_26579,N_26011);
or U28819 (N_28819,N_26794,N_27732);
or U28820 (N_28820,N_26881,N_27461);
and U28821 (N_28821,N_26461,N_26122);
nand U28822 (N_28822,N_27309,N_27132);
or U28823 (N_28823,N_27930,N_26888);
and U28824 (N_28824,N_27902,N_26679);
xnor U28825 (N_28825,N_27196,N_26693);
nor U28826 (N_28826,N_26263,N_26226);
and U28827 (N_28827,N_27163,N_26040);
or U28828 (N_28828,N_27785,N_26566);
or U28829 (N_28829,N_26428,N_26139);
nor U28830 (N_28830,N_26143,N_26419);
nor U28831 (N_28831,N_27918,N_27406);
or U28832 (N_28832,N_27176,N_26861);
xnor U28833 (N_28833,N_26769,N_26978);
nand U28834 (N_28834,N_27317,N_27052);
nand U28835 (N_28835,N_27146,N_27482);
and U28836 (N_28836,N_26016,N_26070);
xor U28837 (N_28837,N_26884,N_27179);
nand U28838 (N_28838,N_26445,N_27152);
or U28839 (N_28839,N_27250,N_27090);
nor U28840 (N_28840,N_26872,N_26983);
xor U28841 (N_28841,N_27564,N_27120);
nor U28842 (N_28842,N_27753,N_26919);
nand U28843 (N_28843,N_26739,N_27161);
xnor U28844 (N_28844,N_27233,N_26276);
or U28845 (N_28845,N_26148,N_26850);
xor U28846 (N_28846,N_27780,N_26504);
xnor U28847 (N_28847,N_27182,N_26392);
xor U28848 (N_28848,N_27769,N_26699);
and U28849 (N_28849,N_27489,N_27823);
and U28850 (N_28850,N_27919,N_27661);
nand U28851 (N_28851,N_26804,N_26077);
nand U28852 (N_28852,N_26258,N_26502);
xnor U28853 (N_28853,N_27796,N_27958);
nand U28854 (N_28854,N_27187,N_27175);
nand U28855 (N_28855,N_26493,N_26659);
nor U28856 (N_28856,N_26231,N_27430);
nor U28857 (N_28857,N_27454,N_26469);
nor U28858 (N_28858,N_27869,N_27137);
or U28859 (N_28859,N_27344,N_26549);
nand U28860 (N_28860,N_27496,N_27635);
or U28861 (N_28861,N_26424,N_27401);
and U28862 (N_28862,N_26396,N_26357);
and U28863 (N_28863,N_26867,N_27909);
xnor U28864 (N_28864,N_27160,N_27997);
and U28865 (N_28865,N_26135,N_27114);
or U28866 (N_28866,N_27487,N_26708);
nor U28867 (N_28867,N_26759,N_27523);
xnor U28868 (N_28868,N_27470,N_27642);
or U28869 (N_28869,N_27472,N_27169);
or U28870 (N_28870,N_26202,N_27467);
or U28871 (N_28871,N_26313,N_27151);
nor U28872 (N_28872,N_27178,N_27955);
and U28873 (N_28873,N_26917,N_26941);
or U28874 (N_28874,N_26856,N_27045);
nor U28875 (N_28875,N_26062,N_26133);
nor U28876 (N_28876,N_26282,N_27043);
nor U28877 (N_28877,N_26125,N_26137);
xnor U28878 (N_28878,N_26007,N_26402);
nor U28879 (N_28879,N_26171,N_26722);
nand U28880 (N_28880,N_27619,N_26335);
xor U28881 (N_28881,N_27390,N_26323);
nor U28882 (N_28882,N_26459,N_27156);
xnor U28883 (N_28883,N_27584,N_27724);
xnor U28884 (N_28884,N_27853,N_27017);
nor U28885 (N_28885,N_27672,N_26270);
and U28886 (N_28886,N_27438,N_27565);
and U28887 (N_28887,N_26197,N_26671);
xor U28888 (N_28888,N_26724,N_26735);
xnor U28889 (N_28889,N_26766,N_27481);
or U28890 (N_28890,N_26426,N_27331);
xor U28891 (N_28891,N_27488,N_27847);
and U28892 (N_28892,N_26817,N_26684);
and U28893 (N_28893,N_26740,N_26001);
and U28894 (N_28894,N_27366,N_27526);
xor U28895 (N_28895,N_26386,N_27532);
xnor U28896 (N_28896,N_26151,N_27570);
nor U28897 (N_28897,N_26883,N_27580);
nand U28898 (N_28898,N_26268,N_26779);
and U28899 (N_28899,N_27238,N_26672);
nand U28900 (N_28900,N_26665,N_26439);
nand U28901 (N_28901,N_27606,N_27625);
and U28902 (N_28902,N_26147,N_26244);
or U28903 (N_28903,N_27986,N_27431);
and U28904 (N_28904,N_26411,N_26755);
xnor U28905 (N_28905,N_27742,N_26141);
xor U28906 (N_28906,N_27002,N_27375);
and U28907 (N_28907,N_26977,N_26382);
or U28908 (N_28908,N_26477,N_27831);
xnor U28909 (N_28909,N_26400,N_27693);
and U28910 (N_28910,N_27167,N_26113);
or U28911 (N_28911,N_27426,N_27648);
xor U28912 (N_28912,N_27530,N_27989);
xor U28913 (N_28913,N_26345,N_27764);
xnor U28914 (N_28914,N_27886,N_26191);
or U28915 (N_28915,N_27563,N_26706);
and U28916 (N_28916,N_26289,N_26841);
nor U28917 (N_28917,N_27170,N_27194);
or U28918 (N_28918,N_26772,N_27352);
or U28919 (N_28919,N_26271,N_27894);
or U28920 (N_28920,N_27582,N_27741);
or U28921 (N_28921,N_27212,N_26324);
nand U28922 (N_28922,N_26482,N_26937);
nor U28923 (N_28923,N_26836,N_27476);
or U28924 (N_28924,N_27716,N_27897);
nor U28925 (N_28925,N_26899,N_26246);
or U28926 (N_28926,N_27718,N_27578);
xor U28927 (N_28927,N_26905,N_27961);
or U28928 (N_28928,N_26248,N_26704);
nor U28929 (N_28929,N_26142,N_26022);
or U28930 (N_28930,N_27128,N_27282);
nor U28931 (N_28931,N_27001,N_26666);
nor U28932 (N_28932,N_27314,N_26472);
or U28933 (N_28933,N_27552,N_26868);
xor U28934 (N_28934,N_26209,N_26523);
and U28935 (N_28935,N_27453,N_27688);
or U28936 (N_28936,N_26798,N_27300);
nand U28937 (N_28937,N_26799,N_27616);
xnor U28938 (N_28938,N_27835,N_27141);
nor U28939 (N_28939,N_27854,N_27987);
and U28940 (N_28940,N_26269,N_26830);
xor U28941 (N_28941,N_26138,N_26583);
xnor U28942 (N_28942,N_27355,N_27086);
or U28943 (N_28943,N_27439,N_27504);
or U28944 (N_28944,N_27729,N_26084);
and U28945 (N_28945,N_27951,N_26823);
xnor U28946 (N_28946,N_26507,N_27962);
xnor U28947 (N_28947,N_26630,N_26078);
and U28948 (N_28948,N_27069,N_26726);
and U28949 (N_28949,N_26190,N_27774);
xnor U28950 (N_28950,N_26918,N_27807);
xnor U28951 (N_28951,N_26773,N_27590);
nand U28952 (N_28952,N_26880,N_26991);
or U28953 (N_28953,N_27338,N_27142);
xnor U28954 (N_28954,N_27075,N_27970);
nor U28955 (N_28955,N_27254,N_27138);
or U28956 (N_28956,N_26777,N_27771);
or U28957 (N_28957,N_26325,N_27216);
xor U28958 (N_28958,N_26992,N_26456);
xnor U28959 (N_28959,N_26782,N_26670);
and U28960 (N_28960,N_26071,N_26213);
and U28961 (N_28961,N_26380,N_26598);
nand U28962 (N_28962,N_27014,N_27712);
xnor U28963 (N_28963,N_27540,N_27735);
or U28964 (N_28964,N_27696,N_27252);
or U28965 (N_28965,N_26694,N_26344);
nand U28966 (N_28966,N_27192,N_26795);
nor U28967 (N_28967,N_27707,N_26626);
xor U28968 (N_28968,N_26998,N_26241);
or U28969 (N_28969,N_26494,N_27992);
or U28970 (N_28970,N_26685,N_27025);
and U28971 (N_28971,N_26253,N_27298);
and U28972 (N_28972,N_27702,N_26374);
xnor U28973 (N_28973,N_26189,N_26591);
and U28974 (N_28974,N_26165,N_27676);
xor U28975 (N_28975,N_27340,N_27666);
nand U28976 (N_28976,N_27037,N_26713);
and U28977 (N_28977,N_26787,N_26515);
and U28978 (N_28978,N_26648,N_26547);
xnor U28979 (N_28979,N_27434,N_27410);
xor U28980 (N_28980,N_26471,N_27974);
xor U28981 (N_28981,N_26796,N_27121);
xnor U28982 (N_28982,N_27100,N_27185);
and U28983 (N_28983,N_26846,N_26383);
xnor U28984 (N_28984,N_26975,N_27127);
and U28985 (N_28985,N_26112,N_26698);
or U28986 (N_28986,N_26362,N_27644);
or U28987 (N_28987,N_26768,N_26744);
nor U28988 (N_28988,N_27686,N_27817);
or U28989 (N_28989,N_26353,N_27969);
nand U28990 (N_28990,N_26254,N_27705);
or U28991 (N_28991,N_27745,N_27195);
xnor U28992 (N_28992,N_27102,N_27830);
nand U28993 (N_28993,N_27343,N_26582);
nand U28994 (N_28994,N_27646,N_26633);
xor U28995 (N_28995,N_27287,N_26524);
xnor U28996 (N_28996,N_27116,N_27589);
xor U28997 (N_28997,N_26682,N_26145);
nor U28998 (N_28998,N_26332,N_27117);
nand U28999 (N_28999,N_26360,N_26099);
nor U29000 (N_29000,N_27275,N_26880);
nor U29001 (N_29001,N_27651,N_27518);
and U29002 (N_29002,N_26416,N_26067);
xor U29003 (N_29003,N_26380,N_26187);
nor U29004 (N_29004,N_27897,N_26669);
nand U29005 (N_29005,N_26947,N_26752);
nand U29006 (N_29006,N_27800,N_27078);
xor U29007 (N_29007,N_26782,N_27388);
xnor U29008 (N_29008,N_27750,N_27572);
xnor U29009 (N_29009,N_26796,N_26808);
xor U29010 (N_29010,N_26984,N_26562);
or U29011 (N_29011,N_27783,N_27022);
nor U29012 (N_29012,N_27580,N_26983);
and U29013 (N_29013,N_27058,N_26878);
or U29014 (N_29014,N_27122,N_26511);
and U29015 (N_29015,N_27943,N_26166);
and U29016 (N_29016,N_27001,N_26531);
or U29017 (N_29017,N_27446,N_26924);
or U29018 (N_29018,N_26872,N_27450);
xnor U29019 (N_29019,N_26853,N_26949);
and U29020 (N_29020,N_27265,N_26769);
nor U29021 (N_29021,N_26431,N_27687);
xor U29022 (N_29022,N_26406,N_27539);
or U29023 (N_29023,N_27964,N_27179);
nand U29024 (N_29024,N_27442,N_26805);
or U29025 (N_29025,N_26423,N_26276);
nor U29026 (N_29026,N_27421,N_27998);
nor U29027 (N_29027,N_26291,N_26222);
nor U29028 (N_29028,N_27759,N_26698);
nand U29029 (N_29029,N_27039,N_26892);
nand U29030 (N_29030,N_26269,N_27029);
nor U29031 (N_29031,N_27154,N_26406);
nor U29032 (N_29032,N_27760,N_27147);
or U29033 (N_29033,N_27961,N_26660);
xor U29034 (N_29034,N_26358,N_27544);
nand U29035 (N_29035,N_27421,N_27332);
and U29036 (N_29036,N_26271,N_26106);
nand U29037 (N_29037,N_27718,N_27168);
and U29038 (N_29038,N_26347,N_26911);
xor U29039 (N_29039,N_27718,N_27311);
nand U29040 (N_29040,N_26737,N_26610);
nand U29041 (N_29041,N_27094,N_27634);
nand U29042 (N_29042,N_27810,N_26060);
nand U29043 (N_29043,N_26589,N_26376);
or U29044 (N_29044,N_26564,N_26045);
xnor U29045 (N_29045,N_26897,N_27206);
or U29046 (N_29046,N_27673,N_27776);
nand U29047 (N_29047,N_26237,N_26137);
xnor U29048 (N_29048,N_27724,N_27571);
nor U29049 (N_29049,N_27950,N_26331);
nand U29050 (N_29050,N_27132,N_26071);
xnor U29051 (N_29051,N_27755,N_26393);
nand U29052 (N_29052,N_27937,N_27703);
and U29053 (N_29053,N_26947,N_27389);
xor U29054 (N_29054,N_27770,N_26708);
nor U29055 (N_29055,N_26531,N_26343);
nand U29056 (N_29056,N_26537,N_26287);
or U29057 (N_29057,N_26618,N_27617);
and U29058 (N_29058,N_27636,N_26417);
xnor U29059 (N_29059,N_27750,N_27895);
nor U29060 (N_29060,N_26463,N_27121);
or U29061 (N_29061,N_26207,N_27267);
nor U29062 (N_29062,N_27807,N_26010);
or U29063 (N_29063,N_27139,N_27007);
and U29064 (N_29064,N_26326,N_27142);
nand U29065 (N_29065,N_26475,N_27689);
xnor U29066 (N_29066,N_26699,N_27053);
and U29067 (N_29067,N_26090,N_26084);
xor U29068 (N_29068,N_26891,N_26324);
and U29069 (N_29069,N_27192,N_26644);
or U29070 (N_29070,N_26902,N_26739);
and U29071 (N_29071,N_27497,N_27141);
xor U29072 (N_29072,N_26762,N_26753);
xor U29073 (N_29073,N_26377,N_27676);
and U29074 (N_29074,N_26905,N_27758);
nor U29075 (N_29075,N_26475,N_27799);
xor U29076 (N_29076,N_27784,N_27499);
nor U29077 (N_29077,N_26333,N_26599);
and U29078 (N_29078,N_26821,N_26620);
and U29079 (N_29079,N_27572,N_26839);
xor U29080 (N_29080,N_27586,N_27266);
nor U29081 (N_29081,N_26097,N_26115);
nor U29082 (N_29082,N_26176,N_27662);
nor U29083 (N_29083,N_27940,N_26394);
or U29084 (N_29084,N_27366,N_26876);
and U29085 (N_29085,N_26208,N_26764);
or U29086 (N_29086,N_27711,N_26291);
nand U29087 (N_29087,N_26005,N_27921);
nand U29088 (N_29088,N_26738,N_26501);
xor U29089 (N_29089,N_26104,N_27476);
xor U29090 (N_29090,N_26032,N_26141);
xor U29091 (N_29091,N_26875,N_26483);
or U29092 (N_29092,N_27616,N_26735);
xnor U29093 (N_29093,N_26069,N_27862);
or U29094 (N_29094,N_27636,N_27704);
and U29095 (N_29095,N_27567,N_27601);
or U29096 (N_29096,N_27450,N_27486);
xnor U29097 (N_29097,N_26872,N_26559);
xnor U29098 (N_29098,N_26745,N_27144);
nor U29099 (N_29099,N_26731,N_27776);
xor U29100 (N_29100,N_26665,N_26607);
nand U29101 (N_29101,N_27767,N_27237);
and U29102 (N_29102,N_26536,N_26039);
nand U29103 (N_29103,N_26873,N_26126);
nand U29104 (N_29104,N_27107,N_26321);
nor U29105 (N_29105,N_27558,N_27696);
nor U29106 (N_29106,N_26321,N_26492);
nor U29107 (N_29107,N_27843,N_27461);
xnor U29108 (N_29108,N_26729,N_26451);
xnor U29109 (N_29109,N_27187,N_27477);
or U29110 (N_29110,N_26389,N_27699);
nor U29111 (N_29111,N_27226,N_27197);
xor U29112 (N_29112,N_26855,N_27328);
xnor U29113 (N_29113,N_27211,N_26266);
and U29114 (N_29114,N_26052,N_26185);
or U29115 (N_29115,N_27063,N_26765);
and U29116 (N_29116,N_26876,N_26700);
nor U29117 (N_29117,N_27627,N_27953);
xor U29118 (N_29118,N_27842,N_27924);
or U29119 (N_29119,N_27231,N_26312);
nand U29120 (N_29120,N_27989,N_26430);
or U29121 (N_29121,N_26285,N_26967);
xnor U29122 (N_29122,N_27971,N_27340);
nor U29123 (N_29123,N_26408,N_27656);
nand U29124 (N_29124,N_26034,N_27550);
xor U29125 (N_29125,N_27597,N_27108);
and U29126 (N_29126,N_27369,N_26076);
nor U29127 (N_29127,N_27433,N_26916);
nor U29128 (N_29128,N_26491,N_26912);
nor U29129 (N_29129,N_26923,N_26324);
nand U29130 (N_29130,N_27329,N_27376);
or U29131 (N_29131,N_26582,N_27518);
or U29132 (N_29132,N_27373,N_26232);
xor U29133 (N_29133,N_27331,N_27769);
and U29134 (N_29134,N_26888,N_26615);
or U29135 (N_29135,N_27052,N_27091);
nor U29136 (N_29136,N_27718,N_26017);
or U29137 (N_29137,N_26059,N_27718);
or U29138 (N_29138,N_26513,N_27056);
or U29139 (N_29139,N_27686,N_26167);
or U29140 (N_29140,N_27490,N_26173);
nor U29141 (N_29141,N_26416,N_27244);
nor U29142 (N_29142,N_27387,N_27917);
nand U29143 (N_29143,N_26008,N_27906);
xor U29144 (N_29144,N_26307,N_26704);
or U29145 (N_29145,N_26355,N_26776);
and U29146 (N_29146,N_26974,N_27668);
xor U29147 (N_29147,N_27022,N_27651);
and U29148 (N_29148,N_27048,N_27369);
nor U29149 (N_29149,N_26268,N_27543);
xor U29150 (N_29150,N_27332,N_27391);
nand U29151 (N_29151,N_26272,N_27952);
or U29152 (N_29152,N_26826,N_27037);
nand U29153 (N_29153,N_27952,N_26987);
and U29154 (N_29154,N_27030,N_27516);
nand U29155 (N_29155,N_27914,N_26593);
or U29156 (N_29156,N_26248,N_27165);
and U29157 (N_29157,N_27859,N_27026);
xor U29158 (N_29158,N_27200,N_26462);
or U29159 (N_29159,N_26006,N_27844);
or U29160 (N_29160,N_27268,N_26506);
nand U29161 (N_29161,N_27459,N_27564);
xnor U29162 (N_29162,N_27051,N_26147);
and U29163 (N_29163,N_27754,N_26748);
nor U29164 (N_29164,N_27832,N_27247);
and U29165 (N_29165,N_26235,N_27063);
nor U29166 (N_29166,N_26688,N_26264);
or U29167 (N_29167,N_26657,N_27775);
and U29168 (N_29168,N_26373,N_27089);
or U29169 (N_29169,N_26026,N_27007);
or U29170 (N_29170,N_27398,N_26655);
or U29171 (N_29171,N_26904,N_26962);
xnor U29172 (N_29172,N_26958,N_26214);
nand U29173 (N_29173,N_26406,N_27609);
nor U29174 (N_29174,N_27204,N_27063);
nor U29175 (N_29175,N_26414,N_26575);
and U29176 (N_29176,N_27745,N_26819);
nand U29177 (N_29177,N_27666,N_27800);
nand U29178 (N_29178,N_26485,N_27963);
nor U29179 (N_29179,N_26523,N_27187);
and U29180 (N_29180,N_27227,N_26495);
nor U29181 (N_29181,N_26036,N_26173);
nand U29182 (N_29182,N_26344,N_27112);
nand U29183 (N_29183,N_27853,N_27996);
nand U29184 (N_29184,N_27798,N_27029);
and U29185 (N_29185,N_26502,N_26520);
and U29186 (N_29186,N_26918,N_26552);
xor U29187 (N_29187,N_26489,N_26138);
and U29188 (N_29188,N_26020,N_26616);
and U29189 (N_29189,N_27378,N_26663);
and U29190 (N_29190,N_27931,N_27687);
nor U29191 (N_29191,N_27318,N_27547);
nor U29192 (N_29192,N_26050,N_26661);
or U29193 (N_29193,N_27877,N_27283);
nor U29194 (N_29194,N_26684,N_26767);
xor U29195 (N_29195,N_27083,N_26442);
nor U29196 (N_29196,N_27619,N_27925);
xnor U29197 (N_29197,N_26883,N_26133);
and U29198 (N_29198,N_26828,N_26819);
nor U29199 (N_29199,N_26425,N_26361);
xnor U29200 (N_29200,N_26374,N_26512);
nor U29201 (N_29201,N_26642,N_26839);
or U29202 (N_29202,N_27019,N_27033);
nor U29203 (N_29203,N_26807,N_27970);
or U29204 (N_29204,N_26411,N_26417);
nor U29205 (N_29205,N_27445,N_27326);
and U29206 (N_29206,N_26334,N_26388);
xnor U29207 (N_29207,N_26133,N_27610);
or U29208 (N_29208,N_27234,N_27328);
xor U29209 (N_29209,N_26307,N_26478);
or U29210 (N_29210,N_27114,N_27384);
or U29211 (N_29211,N_27181,N_26808);
or U29212 (N_29212,N_26532,N_26851);
or U29213 (N_29213,N_27217,N_26252);
nor U29214 (N_29214,N_26738,N_26687);
and U29215 (N_29215,N_26715,N_26706);
nand U29216 (N_29216,N_26719,N_26081);
nor U29217 (N_29217,N_26778,N_26124);
nand U29218 (N_29218,N_27595,N_27823);
xnor U29219 (N_29219,N_26773,N_26891);
or U29220 (N_29220,N_27040,N_27278);
nor U29221 (N_29221,N_27699,N_27817);
nor U29222 (N_29222,N_26951,N_26055);
nand U29223 (N_29223,N_27052,N_26714);
xnor U29224 (N_29224,N_26671,N_27940);
xor U29225 (N_29225,N_26226,N_26264);
or U29226 (N_29226,N_26867,N_26434);
and U29227 (N_29227,N_27963,N_26421);
or U29228 (N_29228,N_26573,N_26322);
or U29229 (N_29229,N_26044,N_26220);
nand U29230 (N_29230,N_26099,N_27190);
and U29231 (N_29231,N_27780,N_26480);
nand U29232 (N_29232,N_26783,N_26737);
or U29233 (N_29233,N_27257,N_27753);
and U29234 (N_29234,N_26630,N_26758);
and U29235 (N_29235,N_26189,N_27113);
xor U29236 (N_29236,N_27407,N_27017);
nand U29237 (N_29237,N_27981,N_26271);
xor U29238 (N_29238,N_26120,N_27258);
nand U29239 (N_29239,N_27143,N_27353);
nor U29240 (N_29240,N_27349,N_27552);
or U29241 (N_29241,N_27019,N_26540);
xor U29242 (N_29242,N_26144,N_26723);
or U29243 (N_29243,N_26126,N_27738);
xor U29244 (N_29244,N_27973,N_27586);
or U29245 (N_29245,N_26764,N_27116);
or U29246 (N_29246,N_27968,N_27345);
and U29247 (N_29247,N_27819,N_27135);
and U29248 (N_29248,N_26763,N_27540);
and U29249 (N_29249,N_27631,N_26427);
and U29250 (N_29250,N_26332,N_26066);
nor U29251 (N_29251,N_27035,N_26091);
xor U29252 (N_29252,N_27247,N_26208);
or U29253 (N_29253,N_27978,N_26035);
nand U29254 (N_29254,N_26586,N_26177);
nand U29255 (N_29255,N_27823,N_26517);
and U29256 (N_29256,N_27274,N_26470);
xnor U29257 (N_29257,N_27164,N_27314);
or U29258 (N_29258,N_27668,N_27907);
xor U29259 (N_29259,N_26496,N_26526);
or U29260 (N_29260,N_27466,N_26539);
nor U29261 (N_29261,N_26376,N_26109);
nand U29262 (N_29262,N_27603,N_26466);
nand U29263 (N_29263,N_27465,N_26332);
nand U29264 (N_29264,N_27568,N_27354);
nor U29265 (N_29265,N_27976,N_27141);
nor U29266 (N_29266,N_27097,N_27193);
or U29267 (N_29267,N_27863,N_27380);
nand U29268 (N_29268,N_27201,N_26033);
nor U29269 (N_29269,N_27330,N_27990);
xnor U29270 (N_29270,N_27260,N_26695);
nor U29271 (N_29271,N_27671,N_26517);
nand U29272 (N_29272,N_27203,N_26009);
nand U29273 (N_29273,N_26520,N_26946);
nand U29274 (N_29274,N_26842,N_27593);
nor U29275 (N_29275,N_27142,N_26392);
nor U29276 (N_29276,N_27996,N_26351);
nand U29277 (N_29277,N_27058,N_26359);
nor U29278 (N_29278,N_26056,N_27418);
or U29279 (N_29279,N_26070,N_27595);
xor U29280 (N_29280,N_26722,N_26191);
or U29281 (N_29281,N_26295,N_26799);
xnor U29282 (N_29282,N_26131,N_26813);
or U29283 (N_29283,N_26943,N_27664);
nor U29284 (N_29284,N_26666,N_26877);
and U29285 (N_29285,N_27402,N_26678);
or U29286 (N_29286,N_26012,N_27032);
nor U29287 (N_29287,N_27102,N_26900);
or U29288 (N_29288,N_26405,N_27660);
or U29289 (N_29289,N_26527,N_27774);
nand U29290 (N_29290,N_26836,N_27413);
or U29291 (N_29291,N_27446,N_27976);
nand U29292 (N_29292,N_27647,N_27857);
xor U29293 (N_29293,N_27879,N_26945);
xnor U29294 (N_29294,N_27139,N_27161);
nor U29295 (N_29295,N_27650,N_26062);
and U29296 (N_29296,N_26833,N_26818);
nor U29297 (N_29297,N_27070,N_26703);
or U29298 (N_29298,N_27372,N_27241);
xnor U29299 (N_29299,N_27631,N_27594);
xnor U29300 (N_29300,N_26489,N_26464);
xnor U29301 (N_29301,N_26286,N_26469);
nand U29302 (N_29302,N_26355,N_27964);
and U29303 (N_29303,N_26604,N_27766);
or U29304 (N_29304,N_26846,N_26103);
and U29305 (N_29305,N_27339,N_27495);
xnor U29306 (N_29306,N_27559,N_26329);
xnor U29307 (N_29307,N_27782,N_26128);
and U29308 (N_29308,N_26345,N_26700);
or U29309 (N_29309,N_26640,N_26047);
xnor U29310 (N_29310,N_26698,N_26592);
and U29311 (N_29311,N_26072,N_26215);
and U29312 (N_29312,N_27717,N_27010);
nand U29313 (N_29313,N_26409,N_27913);
or U29314 (N_29314,N_26097,N_27468);
xor U29315 (N_29315,N_27838,N_26728);
nand U29316 (N_29316,N_26534,N_27714);
nand U29317 (N_29317,N_27951,N_27630);
or U29318 (N_29318,N_26564,N_27798);
and U29319 (N_29319,N_26185,N_26753);
and U29320 (N_29320,N_27063,N_26322);
nand U29321 (N_29321,N_27408,N_26558);
or U29322 (N_29322,N_26750,N_27564);
xor U29323 (N_29323,N_26812,N_27505);
nand U29324 (N_29324,N_26255,N_27073);
nand U29325 (N_29325,N_26798,N_27204);
nor U29326 (N_29326,N_27516,N_26513);
and U29327 (N_29327,N_27730,N_26051);
or U29328 (N_29328,N_26927,N_26935);
nand U29329 (N_29329,N_26213,N_26667);
nand U29330 (N_29330,N_27301,N_27427);
xor U29331 (N_29331,N_26482,N_26725);
xnor U29332 (N_29332,N_27722,N_27055);
and U29333 (N_29333,N_26022,N_26084);
or U29334 (N_29334,N_27514,N_27390);
and U29335 (N_29335,N_27199,N_26287);
nor U29336 (N_29336,N_26506,N_26699);
and U29337 (N_29337,N_27871,N_26824);
xnor U29338 (N_29338,N_26047,N_26853);
nand U29339 (N_29339,N_26132,N_26232);
or U29340 (N_29340,N_27979,N_27449);
or U29341 (N_29341,N_26782,N_26041);
nand U29342 (N_29342,N_26425,N_26143);
xor U29343 (N_29343,N_27681,N_27645);
and U29344 (N_29344,N_26095,N_26503);
nand U29345 (N_29345,N_26216,N_26669);
or U29346 (N_29346,N_27778,N_27499);
xnor U29347 (N_29347,N_26270,N_27759);
nand U29348 (N_29348,N_26706,N_27008);
and U29349 (N_29349,N_27275,N_27504);
or U29350 (N_29350,N_26360,N_27705);
nor U29351 (N_29351,N_26080,N_27739);
or U29352 (N_29352,N_27580,N_27554);
xor U29353 (N_29353,N_27750,N_27904);
or U29354 (N_29354,N_27668,N_27877);
and U29355 (N_29355,N_27013,N_27097);
xnor U29356 (N_29356,N_26162,N_27712);
xor U29357 (N_29357,N_27402,N_27682);
and U29358 (N_29358,N_26965,N_26089);
xnor U29359 (N_29359,N_26569,N_27661);
nor U29360 (N_29360,N_26982,N_27502);
nand U29361 (N_29361,N_27695,N_26920);
or U29362 (N_29362,N_27732,N_27357);
or U29363 (N_29363,N_27877,N_27715);
xnor U29364 (N_29364,N_27552,N_26709);
and U29365 (N_29365,N_26804,N_26928);
or U29366 (N_29366,N_27175,N_27941);
nor U29367 (N_29367,N_27389,N_27283);
nor U29368 (N_29368,N_26487,N_27868);
nand U29369 (N_29369,N_26418,N_27589);
and U29370 (N_29370,N_27897,N_26043);
xnor U29371 (N_29371,N_27940,N_26337);
nor U29372 (N_29372,N_27047,N_27379);
and U29373 (N_29373,N_26802,N_27568);
xor U29374 (N_29374,N_27673,N_26059);
or U29375 (N_29375,N_27943,N_27064);
or U29376 (N_29376,N_26326,N_26859);
nand U29377 (N_29377,N_26621,N_26827);
or U29378 (N_29378,N_27633,N_27376);
or U29379 (N_29379,N_27916,N_26817);
nor U29380 (N_29380,N_27627,N_26911);
xnor U29381 (N_29381,N_26555,N_26092);
nor U29382 (N_29382,N_27746,N_26963);
nand U29383 (N_29383,N_27351,N_27848);
nor U29384 (N_29384,N_27659,N_26768);
xnor U29385 (N_29385,N_26684,N_26323);
nor U29386 (N_29386,N_26459,N_26234);
and U29387 (N_29387,N_27076,N_26506);
nor U29388 (N_29388,N_27922,N_26663);
and U29389 (N_29389,N_27389,N_27741);
nand U29390 (N_29390,N_26758,N_26870);
and U29391 (N_29391,N_26371,N_26071);
nor U29392 (N_29392,N_27493,N_26855);
or U29393 (N_29393,N_27724,N_27974);
xor U29394 (N_29394,N_27733,N_26832);
xnor U29395 (N_29395,N_26491,N_27011);
nor U29396 (N_29396,N_26506,N_27548);
or U29397 (N_29397,N_27772,N_27714);
or U29398 (N_29398,N_26587,N_26283);
nand U29399 (N_29399,N_26997,N_27075);
nor U29400 (N_29400,N_26961,N_26643);
xor U29401 (N_29401,N_26404,N_27681);
and U29402 (N_29402,N_27633,N_27978);
or U29403 (N_29403,N_26714,N_27903);
nand U29404 (N_29404,N_27905,N_27233);
or U29405 (N_29405,N_26799,N_26409);
and U29406 (N_29406,N_27625,N_26858);
nor U29407 (N_29407,N_26402,N_26036);
nor U29408 (N_29408,N_27599,N_27312);
nor U29409 (N_29409,N_26008,N_27809);
or U29410 (N_29410,N_27039,N_27759);
nor U29411 (N_29411,N_26520,N_27879);
nor U29412 (N_29412,N_27981,N_27270);
xor U29413 (N_29413,N_26872,N_26048);
nor U29414 (N_29414,N_26231,N_27778);
nand U29415 (N_29415,N_26744,N_26501);
nand U29416 (N_29416,N_26723,N_27842);
xnor U29417 (N_29417,N_27160,N_27755);
nor U29418 (N_29418,N_26646,N_26542);
or U29419 (N_29419,N_27888,N_27667);
and U29420 (N_29420,N_26412,N_26170);
or U29421 (N_29421,N_27120,N_27082);
nor U29422 (N_29422,N_26952,N_27582);
xor U29423 (N_29423,N_27418,N_26664);
and U29424 (N_29424,N_27232,N_26101);
xnor U29425 (N_29425,N_27541,N_26558);
and U29426 (N_29426,N_27688,N_26460);
xor U29427 (N_29427,N_26706,N_27232);
and U29428 (N_29428,N_26689,N_27322);
xor U29429 (N_29429,N_27872,N_27979);
xor U29430 (N_29430,N_26251,N_26141);
nand U29431 (N_29431,N_26805,N_27411);
and U29432 (N_29432,N_26763,N_27272);
and U29433 (N_29433,N_27939,N_27208);
xnor U29434 (N_29434,N_27377,N_27718);
and U29435 (N_29435,N_27424,N_26070);
and U29436 (N_29436,N_26105,N_27464);
or U29437 (N_29437,N_27343,N_27325);
xnor U29438 (N_29438,N_27660,N_26398);
nand U29439 (N_29439,N_26323,N_26478);
nor U29440 (N_29440,N_27171,N_26135);
xnor U29441 (N_29441,N_27523,N_26334);
xor U29442 (N_29442,N_26410,N_27802);
nand U29443 (N_29443,N_27080,N_26097);
and U29444 (N_29444,N_27327,N_27767);
xnor U29445 (N_29445,N_27391,N_26028);
nand U29446 (N_29446,N_27928,N_26751);
xnor U29447 (N_29447,N_27945,N_27497);
xor U29448 (N_29448,N_26842,N_27065);
nor U29449 (N_29449,N_26020,N_27106);
and U29450 (N_29450,N_26902,N_26359);
nor U29451 (N_29451,N_26190,N_26207);
nand U29452 (N_29452,N_27631,N_26629);
and U29453 (N_29453,N_26839,N_26975);
and U29454 (N_29454,N_26204,N_27294);
and U29455 (N_29455,N_27130,N_27951);
and U29456 (N_29456,N_27506,N_27821);
nand U29457 (N_29457,N_26018,N_27916);
and U29458 (N_29458,N_27862,N_26797);
or U29459 (N_29459,N_26186,N_27606);
and U29460 (N_29460,N_27510,N_27619);
nand U29461 (N_29461,N_26529,N_27163);
nand U29462 (N_29462,N_26046,N_27887);
xnor U29463 (N_29463,N_26054,N_26062);
xor U29464 (N_29464,N_27685,N_26587);
and U29465 (N_29465,N_27784,N_27513);
xnor U29466 (N_29466,N_26776,N_27719);
nand U29467 (N_29467,N_27595,N_27115);
and U29468 (N_29468,N_26824,N_27346);
or U29469 (N_29469,N_26578,N_26226);
nor U29470 (N_29470,N_26197,N_26191);
and U29471 (N_29471,N_26054,N_26688);
nor U29472 (N_29472,N_27227,N_26046);
and U29473 (N_29473,N_27517,N_27444);
nand U29474 (N_29474,N_27096,N_27601);
nor U29475 (N_29475,N_26030,N_27452);
or U29476 (N_29476,N_26938,N_27652);
and U29477 (N_29477,N_26729,N_26164);
nor U29478 (N_29478,N_26163,N_27129);
and U29479 (N_29479,N_27807,N_27540);
xnor U29480 (N_29480,N_27766,N_26588);
and U29481 (N_29481,N_26451,N_27093);
nor U29482 (N_29482,N_27953,N_27645);
nor U29483 (N_29483,N_27134,N_27851);
nor U29484 (N_29484,N_27700,N_27114);
nand U29485 (N_29485,N_26940,N_27661);
or U29486 (N_29486,N_27268,N_27705);
xnor U29487 (N_29487,N_26910,N_26744);
or U29488 (N_29488,N_27778,N_26514);
or U29489 (N_29489,N_27936,N_26115);
nor U29490 (N_29490,N_26779,N_27150);
nand U29491 (N_29491,N_27341,N_27883);
xnor U29492 (N_29492,N_26320,N_27980);
nand U29493 (N_29493,N_26057,N_26602);
nor U29494 (N_29494,N_26029,N_26736);
nand U29495 (N_29495,N_27942,N_26686);
or U29496 (N_29496,N_26695,N_27471);
nand U29497 (N_29497,N_27715,N_27964);
nand U29498 (N_29498,N_27766,N_26082);
and U29499 (N_29499,N_26045,N_26321);
nand U29500 (N_29500,N_27472,N_27198);
and U29501 (N_29501,N_26513,N_26950);
or U29502 (N_29502,N_26008,N_26617);
and U29503 (N_29503,N_26546,N_26819);
xor U29504 (N_29504,N_27245,N_27017);
nor U29505 (N_29505,N_26052,N_26986);
xor U29506 (N_29506,N_27852,N_27878);
nor U29507 (N_29507,N_27793,N_27175);
nand U29508 (N_29508,N_27712,N_27838);
or U29509 (N_29509,N_27923,N_27159);
nand U29510 (N_29510,N_27512,N_26078);
nand U29511 (N_29511,N_26156,N_27398);
nor U29512 (N_29512,N_26466,N_26471);
nor U29513 (N_29513,N_26868,N_27574);
or U29514 (N_29514,N_26281,N_27271);
or U29515 (N_29515,N_26215,N_27285);
xnor U29516 (N_29516,N_26410,N_26300);
xor U29517 (N_29517,N_26714,N_27945);
and U29518 (N_29518,N_27677,N_26103);
and U29519 (N_29519,N_26999,N_27821);
xnor U29520 (N_29520,N_26320,N_27320);
nor U29521 (N_29521,N_27986,N_27616);
or U29522 (N_29522,N_26695,N_27246);
xor U29523 (N_29523,N_27980,N_26742);
and U29524 (N_29524,N_26389,N_27139);
nor U29525 (N_29525,N_26986,N_27732);
or U29526 (N_29526,N_27200,N_26159);
xor U29527 (N_29527,N_26211,N_26106);
or U29528 (N_29528,N_26509,N_27892);
or U29529 (N_29529,N_26259,N_27497);
or U29530 (N_29530,N_27387,N_27429);
nand U29531 (N_29531,N_27278,N_27026);
or U29532 (N_29532,N_26737,N_26790);
and U29533 (N_29533,N_27502,N_26622);
nand U29534 (N_29534,N_26545,N_27034);
nand U29535 (N_29535,N_26872,N_26100);
nand U29536 (N_29536,N_26058,N_27924);
nand U29537 (N_29537,N_26345,N_27435);
nor U29538 (N_29538,N_26741,N_27175);
xor U29539 (N_29539,N_27976,N_26624);
or U29540 (N_29540,N_27740,N_27091);
nand U29541 (N_29541,N_26699,N_26899);
xnor U29542 (N_29542,N_26086,N_26042);
nor U29543 (N_29543,N_26603,N_27472);
nand U29544 (N_29544,N_26573,N_27450);
nor U29545 (N_29545,N_26364,N_26649);
xnor U29546 (N_29546,N_26945,N_27549);
nor U29547 (N_29547,N_26767,N_27829);
or U29548 (N_29548,N_26194,N_26146);
and U29549 (N_29549,N_27349,N_27816);
nor U29550 (N_29550,N_26334,N_26121);
and U29551 (N_29551,N_26209,N_26631);
nand U29552 (N_29552,N_26457,N_27027);
nor U29553 (N_29553,N_27824,N_26620);
xnor U29554 (N_29554,N_27608,N_26724);
and U29555 (N_29555,N_26509,N_27908);
xnor U29556 (N_29556,N_27889,N_26461);
nor U29557 (N_29557,N_27067,N_26155);
nand U29558 (N_29558,N_26112,N_27493);
xnor U29559 (N_29559,N_27030,N_27138);
nand U29560 (N_29560,N_26504,N_27345);
or U29561 (N_29561,N_27649,N_26121);
and U29562 (N_29562,N_27973,N_26313);
or U29563 (N_29563,N_27774,N_27454);
nand U29564 (N_29564,N_26734,N_27287);
and U29565 (N_29565,N_26474,N_26291);
and U29566 (N_29566,N_27611,N_27874);
and U29567 (N_29567,N_27047,N_26902);
and U29568 (N_29568,N_27369,N_27097);
or U29569 (N_29569,N_26218,N_26698);
xor U29570 (N_29570,N_26385,N_27081);
nor U29571 (N_29571,N_27908,N_26960);
or U29572 (N_29572,N_27147,N_26242);
xnor U29573 (N_29573,N_26544,N_27225);
and U29574 (N_29574,N_26913,N_26453);
xor U29575 (N_29575,N_27877,N_26706);
or U29576 (N_29576,N_27436,N_27274);
nand U29577 (N_29577,N_26990,N_26402);
nand U29578 (N_29578,N_27789,N_26350);
xor U29579 (N_29579,N_27244,N_27636);
nand U29580 (N_29580,N_26634,N_26032);
xor U29581 (N_29581,N_27233,N_26338);
xnor U29582 (N_29582,N_27862,N_27062);
xnor U29583 (N_29583,N_26572,N_27121);
nor U29584 (N_29584,N_27925,N_27945);
nor U29585 (N_29585,N_27319,N_27713);
xor U29586 (N_29586,N_27538,N_26798);
xnor U29587 (N_29587,N_26981,N_27120);
nand U29588 (N_29588,N_27827,N_26593);
xor U29589 (N_29589,N_27791,N_26564);
xor U29590 (N_29590,N_26835,N_26936);
nor U29591 (N_29591,N_27095,N_27674);
nand U29592 (N_29592,N_26693,N_26433);
nor U29593 (N_29593,N_26813,N_27048);
nand U29594 (N_29594,N_26693,N_26295);
and U29595 (N_29595,N_26545,N_26484);
and U29596 (N_29596,N_26451,N_27044);
nand U29597 (N_29597,N_26247,N_26145);
nor U29598 (N_29598,N_26877,N_26770);
and U29599 (N_29599,N_27347,N_27314);
xor U29600 (N_29600,N_26949,N_27250);
and U29601 (N_29601,N_26455,N_27200);
and U29602 (N_29602,N_26040,N_27796);
nand U29603 (N_29603,N_27351,N_26514);
xnor U29604 (N_29604,N_26892,N_26088);
and U29605 (N_29605,N_26402,N_26340);
nand U29606 (N_29606,N_26376,N_27859);
xor U29607 (N_29607,N_26806,N_27305);
xor U29608 (N_29608,N_26768,N_27109);
and U29609 (N_29609,N_27608,N_27662);
and U29610 (N_29610,N_27492,N_26748);
or U29611 (N_29611,N_27208,N_27481);
or U29612 (N_29612,N_26580,N_26874);
or U29613 (N_29613,N_27251,N_26270);
or U29614 (N_29614,N_26420,N_26315);
nor U29615 (N_29615,N_27132,N_27208);
xor U29616 (N_29616,N_26515,N_26638);
xor U29617 (N_29617,N_26981,N_27692);
or U29618 (N_29618,N_26574,N_26671);
nor U29619 (N_29619,N_27359,N_27966);
and U29620 (N_29620,N_27614,N_27137);
or U29621 (N_29621,N_27448,N_27777);
or U29622 (N_29622,N_26483,N_26100);
xnor U29623 (N_29623,N_27023,N_26538);
nand U29624 (N_29624,N_26207,N_27672);
nand U29625 (N_29625,N_27804,N_26802);
and U29626 (N_29626,N_27332,N_26600);
nor U29627 (N_29627,N_27729,N_27801);
nand U29628 (N_29628,N_26671,N_26338);
xor U29629 (N_29629,N_27975,N_27632);
xor U29630 (N_29630,N_26361,N_26269);
and U29631 (N_29631,N_27508,N_27165);
xor U29632 (N_29632,N_26143,N_26628);
xor U29633 (N_29633,N_26576,N_27901);
and U29634 (N_29634,N_26460,N_27899);
and U29635 (N_29635,N_26632,N_27728);
and U29636 (N_29636,N_26610,N_27190);
and U29637 (N_29637,N_27466,N_27785);
or U29638 (N_29638,N_26109,N_26258);
nor U29639 (N_29639,N_26065,N_26398);
nand U29640 (N_29640,N_27028,N_26200);
nand U29641 (N_29641,N_26940,N_26243);
nor U29642 (N_29642,N_27046,N_27744);
nor U29643 (N_29643,N_26062,N_27231);
and U29644 (N_29644,N_26444,N_26649);
or U29645 (N_29645,N_27386,N_27106);
and U29646 (N_29646,N_27267,N_26550);
xnor U29647 (N_29647,N_27721,N_27677);
or U29648 (N_29648,N_26865,N_27190);
or U29649 (N_29649,N_27277,N_27219);
nor U29650 (N_29650,N_27178,N_27341);
xnor U29651 (N_29651,N_26515,N_27659);
and U29652 (N_29652,N_27527,N_26320);
or U29653 (N_29653,N_27212,N_26833);
or U29654 (N_29654,N_26787,N_27605);
and U29655 (N_29655,N_26988,N_27531);
xnor U29656 (N_29656,N_26866,N_26910);
or U29657 (N_29657,N_27448,N_26651);
xor U29658 (N_29658,N_27366,N_26577);
nand U29659 (N_29659,N_27390,N_27406);
or U29660 (N_29660,N_27157,N_26288);
nor U29661 (N_29661,N_27436,N_27664);
or U29662 (N_29662,N_26279,N_27517);
xor U29663 (N_29663,N_26152,N_27543);
nor U29664 (N_29664,N_26956,N_26848);
nand U29665 (N_29665,N_27787,N_26483);
nand U29666 (N_29666,N_26283,N_26728);
xor U29667 (N_29667,N_26583,N_26577);
and U29668 (N_29668,N_27271,N_27412);
and U29669 (N_29669,N_26794,N_27290);
and U29670 (N_29670,N_27356,N_27841);
xnor U29671 (N_29671,N_27838,N_27967);
xor U29672 (N_29672,N_26997,N_27065);
nand U29673 (N_29673,N_26955,N_26240);
and U29674 (N_29674,N_26582,N_27152);
nand U29675 (N_29675,N_27990,N_27128);
xor U29676 (N_29676,N_27677,N_27161);
and U29677 (N_29677,N_27129,N_26433);
nand U29678 (N_29678,N_27465,N_26860);
nand U29679 (N_29679,N_26585,N_27153);
or U29680 (N_29680,N_27461,N_26219);
xnor U29681 (N_29681,N_27329,N_26960);
xnor U29682 (N_29682,N_27507,N_26336);
nand U29683 (N_29683,N_26507,N_26888);
and U29684 (N_29684,N_27559,N_26863);
xnor U29685 (N_29685,N_26184,N_26474);
and U29686 (N_29686,N_26777,N_26122);
nor U29687 (N_29687,N_27564,N_26483);
or U29688 (N_29688,N_26291,N_26980);
or U29689 (N_29689,N_27504,N_27632);
nor U29690 (N_29690,N_27139,N_27029);
and U29691 (N_29691,N_27123,N_26961);
xnor U29692 (N_29692,N_27365,N_26259);
and U29693 (N_29693,N_26379,N_26274);
and U29694 (N_29694,N_26680,N_27465);
xnor U29695 (N_29695,N_26606,N_27522);
nand U29696 (N_29696,N_27413,N_26903);
or U29697 (N_29697,N_27716,N_27411);
nand U29698 (N_29698,N_26833,N_27517);
and U29699 (N_29699,N_27400,N_27640);
and U29700 (N_29700,N_27674,N_26822);
or U29701 (N_29701,N_27518,N_27468);
xnor U29702 (N_29702,N_26389,N_27594);
xnor U29703 (N_29703,N_27402,N_27713);
xnor U29704 (N_29704,N_27915,N_26653);
or U29705 (N_29705,N_27055,N_26348);
or U29706 (N_29706,N_27798,N_26482);
nor U29707 (N_29707,N_27939,N_26751);
or U29708 (N_29708,N_27974,N_26092);
xor U29709 (N_29709,N_27270,N_27900);
nand U29710 (N_29710,N_26328,N_27526);
or U29711 (N_29711,N_27757,N_26834);
xor U29712 (N_29712,N_26609,N_26487);
and U29713 (N_29713,N_26662,N_27802);
and U29714 (N_29714,N_27141,N_26740);
and U29715 (N_29715,N_26279,N_27743);
xor U29716 (N_29716,N_26829,N_27349);
nand U29717 (N_29717,N_26262,N_26562);
and U29718 (N_29718,N_26288,N_26727);
or U29719 (N_29719,N_26076,N_26941);
xnor U29720 (N_29720,N_27288,N_27413);
nand U29721 (N_29721,N_26682,N_27268);
and U29722 (N_29722,N_27328,N_26487);
xor U29723 (N_29723,N_27377,N_27519);
and U29724 (N_29724,N_26382,N_26330);
nor U29725 (N_29725,N_26896,N_26091);
nor U29726 (N_29726,N_27237,N_26330);
nand U29727 (N_29727,N_26585,N_26589);
nor U29728 (N_29728,N_27507,N_26571);
xnor U29729 (N_29729,N_26610,N_27210);
and U29730 (N_29730,N_26058,N_27307);
nand U29731 (N_29731,N_26765,N_27734);
xnor U29732 (N_29732,N_26271,N_26427);
xor U29733 (N_29733,N_27136,N_26052);
nand U29734 (N_29734,N_27357,N_26387);
or U29735 (N_29735,N_27121,N_26434);
nor U29736 (N_29736,N_26006,N_27908);
or U29737 (N_29737,N_26404,N_26382);
nor U29738 (N_29738,N_26212,N_27062);
or U29739 (N_29739,N_26650,N_27285);
nor U29740 (N_29740,N_26759,N_26134);
nor U29741 (N_29741,N_26580,N_26282);
nand U29742 (N_29742,N_26180,N_27494);
or U29743 (N_29743,N_26061,N_27301);
xor U29744 (N_29744,N_26857,N_26808);
nor U29745 (N_29745,N_26123,N_27783);
nor U29746 (N_29746,N_27059,N_27017);
or U29747 (N_29747,N_26435,N_26438);
nand U29748 (N_29748,N_26125,N_26539);
xnor U29749 (N_29749,N_27476,N_27139);
xnor U29750 (N_29750,N_27237,N_26294);
and U29751 (N_29751,N_27273,N_26804);
xor U29752 (N_29752,N_26543,N_27688);
xnor U29753 (N_29753,N_26576,N_26944);
nor U29754 (N_29754,N_27689,N_27820);
or U29755 (N_29755,N_26982,N_27027);
nor U29756 (N_29756,N_26410,N_27893);
or U29757 (N_29757,N_27283,N_27041);
and U29758 (N_29758,N_26913,N_27345);
nand U29759 (N_29759,N_26812,N_26623);
nor U29760 (N_29760,N_27193,N_27980);
xnor U29761 (N_29761,N_26523,N_26902);
nand U29762 (N_29762,N_26573,N_26938);
xnor U29763 (N_29763,N_27325,N_27206);
nor U29764 (N_29764,N_27687,N_27696);
or U29765 (N_29765,N_26705,N_27801);
or U29766 (N_29766,N_26703,N_27892);
and U29767 (N_29767,N_27962,N_26559);
or U29768 (N_29768,N_26981,N_27720);
or U29769 (N_29769,N_26315,N_27931);
nor U29770 (N_29770,N_26390,N_26308);
nand U29771 (N_29771,N_27498,N_26003);
or U29772 (N_29772,N_26369,N_26321);
and U29773 (N_29773,N_27673,N_27826);
nand U29774 (N_29774,N_27226,N_26190);
xor U29775 (N_29775,N_27080,N_27658);
or U29776 (N_29776,N_26011,N_27270);
nand U29777 (N_29777,N_26139,N_26615);
and U29778 (N_29778,N_27473,N_27740);
or U29779 (N_29779,N_26034,N_26970);
xnor U29780 (N_29780,N_26673,N_27940);
nor U29781 (N_29781,N_26491,N_27962);
and U29782 (N_29782,N_26853,N_27624);
xor U29783 (N_29783,N_26971,N_26291);
or U29784 (N_29784,N_26528,N_26109);
nand U29785 (N_29785,N_26355,N_27181);
and U29786 (N_29786,N_26402,N_27587);
nor U29787 (N_29787,N_27710,N_26577);
or U29788 (N_29788,N_26657,N_27345);
nor U29789 (N_29789,N_27457,N_27383);
xor U29790 (N_29790,N_26337,N_26359);
and U29791 (N_29791,N_26627,N_26325);
or U29792 (N_29792,N_27984,N_27044);
xor U29793 (N_29793,N_27006,N_27187);
nand U29794 (N_29794,N_26985,N_26997);
and U29795 (N_29795,N_26598,N_27729);
nor U29796 (N_29796,N_26120,N_26233);
nor U29797 (N_29797,N_27749,N_27996);
nand U29798 (N_29798,N_26378,N_27168);
xor U29799 (N_29799,N_27408,N_27457);
or U29800 (N_29800,N_26451,N_27313);
nand U29801 (N_29801,N_26552,N_26793);
xnor U29802 (N_29802,N_27535,N_27041);
nor U29803 (N_29803,N_26740,N_27716);
or U29804 (N_29804,N_26152,N_27706);
and U29805 (N_29805,N_27769,N_26306);
and U29806 (N_29806,N_26364,N_26505);
nand U29807 (N_29807,N_27882,N_27938);
xnor U29808 (N_29808,N_26018,N_27300);
nor U29809 (N_29809,N_26976,N_26802);
nand U29810 (N_29810,N_27164,N_27528);
nand U29811 (N_29811,N_27916,N_27514);
xnor U29812 (N_29812,N_26750,N_26802);
nor U29813 (N_29813,N_27376,N_27441);
nor U29814 (N_29814,N_26399,N_27831);
nand U29815 (N_29815,N_27849,N_27684);
or U29816 (N_29816,N_27816,N_26701);
nand U29817 (N_29817,N_27713,N_27581);
nand U29818 (N_29818,N_26692,N_26236);
nand U29819 (N_29819,N_27412,N_27252);
xnor U29820 (N_29820,N_27113,N_27019);
nand U29821 (N_29821,N_26934,N_27437);
xnor U29822 (N_29822,N_26767,N_26770);
or U29823 (N_29823,N_26095,N_26890);
or U29824 (N_29824,N_26209,N_26332);
or U29825 (N_29825,N_26289,N_27133);
xor U29826 (N_29826,N_26499,N_27957);
or U29827 (N_29827,N_27601,N_27299);
nand U29828 (N_29828,N_27069,N_27121);
xnor U29829 (N_29829,N_26323,N_26368);
nor U29830 (N_29830,N_26271,N_26875);
nor U29831 (N_29831,N_27391,N_27050);
nor U29832 (N_29832,N_27628,N_27077);
nor U29833 (N_29833,N_26555,N_27187);
xnor U29834 (N_29834,N_26657,N_27896);
nor U29835 (N_29835,N_27904,N_26428);
xor U29836 (N_29836,N_27023,N_27301);
xor U29837 (N_29837,N_27915,N_26486);
nor U29838 (N_29838,N_26041,N_27426);
nand U29839 (N_29839,N_26925,N_26503);
or U29840 (N_29840,N_27807,N_27186);
nor U29841 (N_29841,N_27684,N_27042);
nor U29842 (N_29842,N_26584,N_26159);
nand U29843 (N_29843,N_26848,N_27364);
xnor U29844 (N_29844,N_27079,N_27387);
nand U29845 (N_29845,N_26545,N_27379);
xor U29846 (N_29846,N_26705,N_27412);
or U29847 (N_29847,N_26786,N_27144);
or U29848 (N_29848,N_26748,N_27193);
or U29849 (N_29849,N_26013,N_27875);
and U29850 (N_29850,N_26540,N_27978);
xor U29851 (N_29851,N_27105,N_26280);
or U29852 (N_29852,N_27619,N_27412);
or U29853 (N_29853,N_26675,N_27958);
and U29854 (N_29854,N_26305,N_27315);
nand U29855 (N_29855,N_26776,N_26521);
nor U29856 (N_29856,N_26943,N_26238);
or U29857 (N_29857,N_27095,N_27905);
nor U29858 (N_29858,N_26778,N_27007);
or U29859 (N_29859,N_27805,N_27806);
nor U29860 (N_29860,N_27339,N_27443);
xnor U29861 (N_29861,N_27413,N_27108);
and U29862 (N_29862,N_27094,N_27637);
nor U29863 (N_29863,N_27210,N_26723);
nor U29864 (N_29864,N_26572,N_26553);
xnor U29865 (N_29865,N_27755,N_26253);
or U29866 (N_29866,N_27050,N_27703);
nand U29867 (N_29867,N_26865,N_27847);
and U29868 (N_29868,N_27081,N_26892);
nand U29869 (N_29869,N_27991,N_26085);
nor U29870 (N_29870,N_27281,N_26381);
and U29871 (N_29871,N_26589,N_26519);
nor U29872 (N_29872,N_26900,N_26034);
nand U29873 (N_29873,N_27507,N_27434);
xor U29874 (N_29874,N_26595,N_27141);
xnor U29875 (N_29875,N_27566,N_27713);
and U29876 (N_29876,N_27476,N_26883);
xnor U29877 (N_29877,N_26989,N_27763);
and U29878 (N_29878,N_27945,N_27360);
or U29879 (N_29879,N_27548,N_26218);
nand U29880 (N_29880,N_27347,N_26340);
or U29881 (N_29881,N_27985,N_26703);
nor U29882 (N_29882,N_26479,N_26807);
nor U29883 (N_29883,N_27023,N_26732);
or U29884 (N_29884,N_27072,N_27428);
and U29885 (N_29885,N_26572,N_27170);
nor U29886 (N_29886,N_26142,N_26272);
nor U29887 (N_29887,N_27491,N_26245);
nor U29888 (N_29888,N_27032,N_26979);
nand U29889 (N_29889,N_26837,N_26680);
xor U29890 (N_29890,N_27461,N_26214);
nand U29891 (N_29891,N_26107,N_27758);
nand U29892 (N_29892,N_27196,N_27511);
xnor U29893 (N_29893,N_27474,N_26822);
nand U29894 (N_29894,N_27391,N_26929);
or U29895 (N_29895,N_26830,N_26410);
nand U29896 (N_29896,N_26799,N_26546);
or U29897 (N_29897,N_26395,N_26706);
or U29898 (N_29898,N_26766,N_27277);
xnor U29899 (N_29899,N_26090,N_26214);
nor U29900 (N_29900,N_26893,N_26379);
or U29901 (N_29901,N_27971,N_26239);
nor U29902 (N_29902,N_26263,N_27041);
nand U29903 (N_29903,N_26533,N_26129);
xnor U29904 (N_29904,N_26674,N_26452);
xnor U29905 (N_29905,N_27645,N_26006);
nand U29906 (N_29906,N_26082,N_27676);
or U29907 (N_29907,N_27819,N_27662);
nand U29908 (N_29908,N_27169,N_27646);
xnor U29909 (N_29909,N_27383,N_27372);
xnor U29910 (N_29910,N_27576,N_27372);
and U29911 (N_29911,N_27772,N_26979);
or U29912 (N_29912,N_26960,N_26157);
xor U29913 (N_29913,N_27849,N_27658);
xor U29914 (N_29914,N_27719,N_27152);
or U29915 (N_29915,N_27141,N_27083);
and U29916 (N_29916,N_27472,N_26994);
and U29917 (N_29917,N_26039,N_26544);
or U29918 (N_29918,N_27846,N_26521);
and U29919 (N_29919,N_27317,N_27865);
nor U29920 (N_29920,N_27098,N_27451);
nor U29921 (N_29921,N_27748,N_26542);
xor U29922 (N_29922,N_27244,N_27856);
nor U29923 (N_29923,N_26895,N_26329);
and U29924 (N_29924,N_26666,N_26696);
nand U29925 (N_29925,N_27718,N_26643);
nand U29926 (N_29926,N_26626,N_26177);
and U29927 (N_29927,N_26570,N_26882);
xor U29928 (N_29928,N_27702,N_26002);
nor U29929 (N_29929,N_27569,N_26538);
nand U29930 (N_29930,N_27446,N_27898);
nand U29931 (N_29931,N_27717,N_26375);
and U29932 (N_29932,N_26316,N_27005);
and U29933 (N_29933,N_27251,N_26361);
and U29934 (N_29934,N_27940,N_27811);
nand U29935 (N_29935,N_27567,N_26654);
or U29936 (N_29936,N_27773,N_26730);
nor U29937 (N_29937,N_26279,N_26917);
nand U29938 (N_29938,N_27067,N_26338);
nand U29939 (N_29939,N_27464,N_26789);
and U29940 (N_29940,N_27890,N_26833);
or U29941 (N_29941,N_26902,N_26504);
xnor U29942 (N_29942,N_26360,N_26542);
xnor U29943 (N_29943,N_27335,N_26740);
nand U29944 (N_29944,N_26802,N_27947);
xor U29945 (N_29945,N_27810,N_26057);
or U29946 (N_29946,N_27488,N_27237);
nor U29947 (N_29947,N_26734,N_27794);
and U29948 (N_29948,N_27099,N_26535);
nand U29949 (N_29949,N_26785,N_27579);
or U29950 (N_29950,N_27354,N_26228);
nand U29951 (N_29951,N_26048,N_27843);
nor U29952 (N_29952,N_27268,N_27470);
and U29953 (N_29953,N_27077,N_27056);
or U29954 (N_29954,N_26634,N_26974);
nand U29955 (N_29955,N_27356,N_26269);
nor U29956 (N_29956,N_27129,N_26496);
and U29957 (N_29957,N_27261,N_27891);
or U29958 (N_29958,N_26773,N_27540);
nor U29959 (N_29959,N_26915,N_27608);
or U29960 (N_29960,N_26804,N_26160);
nor U29961 (N_29961,N_27249,N_27737);
or U29962 (N_29962,N_26524,N_26596);
nand U29963 (N_29963,N_26314,N_27400);
xor U29964 (N_29964,N_27881,N_27887);
and U29965 (N_29965,N_26553,N_26999);
nor U29966 (N_29966,N_26300,N_27252);
and U29967 (N_29967,N_27266,N_27855);
nand U29968 (N_29968,N_26654,N_26474);
xor U29969 (N_29969,N_27037,N_27560);
and U29970 (N_29970,N_26878,N_27363);
nand U29971 (N_29971,N_26428,N_27381);
and U29972 (N_29972,N_26074,N_26134);
nor U29973 (N_29973,N_27450,N_27094);
nor U29974 (N_29974,N_26771,N_26563);
nor U29975 (N_29975,N_26392,N_26613);
nand U29976 (N_29976,N_27613,N_26799);
xnor U29977 (N_29977,N_27431,N_27659);
xor U29978 (N_29978,N_26902,N_26430);
nand U29979 (N_29979,N_26197,N_27511);
nand U29980 (N_29980,N_27883,N_26674);
or U29981 (N_29981,N_27545,N_26390);
or U29982 (N_29982,N_27598,N_27714);
xnor U29983 (N_29983,N_26375,N_27193);
nand U29984 (N_29984,N_27722,N_26164);
nor U29985 (N_29985,N_26946,N_26884);
nand U29986 (N_29986,N_27609,N_26990);
nand U29987 (N_29987,N_26674,N_27182);
and U29988 (N_29988,N_27194,N_26152);
nand U29989 (N_29989,N_26678,N_26708);
or U29990 (N_29990,N_26191,N_27843);
xor U29991 (N_29991,N_26441,N_27725);
nor U29992 (N_29992,N_27751,N_26212);
and U29993 (N_29993,N_27344,N_27290);
and U29994 (N_29994,N_26490,N_26017);
and U29995 (N_29995,N_27021,N_27166);
or U29996 (N_29996,N_26714,N_26018);
and U29997 (N_29997,N_26343,N_26227);
nor U29998 (N_29998,N_26061,N_26435);
and U29999 (N_29999,N_26427,N_26202);
nand UO_0 (O_0,N_29856,N_28031);
and UO_1 (O_1,N_29771,N_28890);
and UO_2 (O_2,N_28300,N_29366);
or UO_3 (O_3,N_28313,N_29910);
xor UO_4 (O_4,N_29852,N_29136);
and UO_5 (O_5,N_29499,N_29898);
or UO_6 (O_6,N_28563,N_29644);
xor UO_7 (O_7,N_28649,N_28228);
xnor UO_8 (O_8,N_28298,N_28693);
nor UO_9 (O_9,N_29020,N_28501);
nor UO_10 (O_10,N_29601,N_28554);
and UO_11 (O_11,N_29507,N_28381);
xor UO_12 (O_12,N_29867,N_28422);
nand UO_13 (O_13,N_29440,N_29751);
xnor UO_14 (O_14,N_28665,N_29805);
nor UO_15 (O_15,N_29205,N_28541);
nand UO_16 (O_16,N_29840,N_28608);
nand UO_17 (O_17,N_28136,N_28118);
nor UO_18 (O_18,N_28833,N_28186);
or UO_19 (O_19,N_28323,N_29139);
nor UO_20 (O_20,N_29168,N_28721);
nor UO_21 (O_21,N_28002,N_29464);
xor UO_22 (O_22,N_29900,N_29713);
or UO_23 (O_23,N_29978,N_28847);
and UO_24 (O_24,N_29091,N_28653);
nor UO_25 (O_25,N_28112,N_29110);
nand UO_26 (O_26,N_28322,N_29930);
nand UO_27 (O_27,N_29480,N_29591);
and UO_28 (O_28,N_29768,N_29195);
and UO_29 (O_29,N_29680,N_29879);
and UO_30 (O_30,N_29718,N_29230);
nor UO_31 (O_31,N_28899,N_28285);
nand UO_32 (O_32,N_28971,N_29066);
nor UO_33 (O_33,N_28060,N_29203);
nand UO_34 (O_34,N_29769,N_28761);
nand UO_35 (O_35,N_28707,N_28142);
xnor UO_36 (O_36,N_29465,N_29542);
nand UO_37 (O_37,N_28138,N_29620);
or UO_38 (O_38,N_29524,N_29027);
nand UO_39 (O_39,N_29980,N_29748);
nor UO_40 (O_40,N_29054,N_28929);
nor UO_41 (O_41,N_29976,N_28044);
and UO_42 (O_42,N_28294,N_29035);
nand UO_43 (O_43,N_28543,N_28542);
or UO_44 (O_44,N_29134,N_29806);
and UO_45 (O_45,N_29154,N_28902);
or UO_46 (O_46,N_29551,N_28640);
or UO_47 (O_47,N_29624,N_29165);
nor UO_48 (O_48,N_28612,N_28567);
and UO_49 (O_49,N_29240,N_29038);
or UO_50 (O_50,N_28836,N_29371);
nor UO_51 (O_51,N_29181,N_29942);
and UO_52 (O_52,N_28454,N_28908);
or UO_53 (O_53,N_29323,N_28686);
or UO_54 (O_54,N_28279,N_28914);
nand UO_55 (O_55,N_29354,N_28708);
and UO_56 (O_56,N_29526,N_28759);
or UO_57 (O_57,N_29794,N_28276);
xnor UO_58 (O_58,N_29398,N_28360);
xor UO_59 (O_59,N_29523,N_29362);
or UO_60 (O_60,N_28507,N_28208);
nand UO_61 (O_61,N_29690,N_29302);
or UO_62 (O_62,N_28844,N_29498);
or UO_63 (O_63,N_29972,N_28973);
and UO_64 (O_64,N_29698,N_29204);
nand UO_65 (O_65,N_29741,N_29039);
nor UO_66 (O_66,N_28842,N_29073);
nand UO_67 (O_67,N_28858,N_29272);
or UO_68 (O_68,N_29825,N_28756);
and UO_69 (O_69,N_29904,N_29599);
or UO_70 (O_70,N_29519,N_28077);
and UO_71 (O_71,N_29937,N_28078);
nor UO_72 (O_72,N_29209,N_29701);
xor UO_73 (O_73,N_29504,N_28968);
or UO_74 (O_74,N_28366,N_29176);
nand UO_75 (O_75,N_28273,N_28943);
nor UO_76 (O_76,N_28898,N_28132);
and UO_77 (O_77,N_28714,N_29691);
xor UO_78 (O_78,N_28473,N_29030);
nor UO_79 (O_79,N_29408,N_29126);
nand UO_80 (O_80,N_29502,N_28675);
nand UO_81 (O_81,N_28951,N_29512);
nor UO_82 (O_82,N_28616,N_29000);
nand UO_83 (O_83,N_29872,N_29400);
xnor UO_84 (O_84,N_28198,N_28987);
and UO_85 (O_85,N_29822,N_29076);
xnor UO_86 (O_86,N_29372,N_29034);
or UO_87 (O_87,N_28210,N_29380);
nand UO_88 (O_88,N_29579,N_29202);
or UO_89 (O_89,N_29429,N_29926);
nor UO_90 (O_90,N_28872,N_28846);
nor UO_91 (O_91,N_29311,N_28015);
nand UO_92 (O_92,N_29839,N_28339);
xnor UO_93 (O_93,N_28853,N_29723);
nand UO_94 (O_94,N_29527,N_29901);
xor UO_95 (O_95,N_29662,N_29656);
xnor UO_96 (O_96,N_29486,N_29142);
nand UO_97 (O_97,N_28436,N_28026);
xnor UO_98 (O_98,N_28682,N_28578);
nor UO_99 (O_99,N_28318,N_29534);
and UO_100 (O_100,N_28103,N_29836);
xor UO_101 (O_101,N_28755,N_29052);
nand UO_102 (O_102,N_29044,N_28676);
nor UO_103 (O_103,N_28217,N_29053);
xnor UO_104 (O_104,N_28931,N_29515);
nor UO_105 (O_105,N_29638,N_28412);
nor UO_106 (O_106,N_29358,N_29614);
nor UO_107 (O_107,N_28011,N_28086);
nand UO_108 (O_108,N_28382,N_28762);
nand UO_109 (O_109,N_28822,N_29037);
xnor UO_110 (O_110,N_28358,N_28281);
xor UO_111 (O_111,N_29316,N_29835);
xor UO_112 (O_112,N_29497,N_28962);
nand UO_113 (O_113,N_28362,N_28128);
nor UO_114 (O_114,N_29161,N_29753);
and UO_115 (O_115,N_29317,N_28841);
or UO_116 (O_116,N_28202,N_29006);
nand UO_117 (O_117,N_29549,N_28239);
or UO_118 (O_118,N_28718,N_28697);
xnor UO_119 (O_119,N_28798,N_28260);
or UO_120 (O_120,N_29897,N_29873);
xnor UO_121 (O_121,N_28195,N_29984);
xor UO_122 (O_122,N_29944,N_29736);
xnor UO_123 (O_123,N_29231,N_28831);
and UO_124 (O_124,N_28233,N_29494);
and UO_125 (O_125,N_29212,N_29538);
nand UO_126 (O_126,N_28857,N_29047);
nand UO_127 (O_127,N_29708,N_28089);
xor UO_128 (O_128,N_28625,N_29508);
xnor UO_129 (O_129,N_28711,N_28367);
nand UO_130 (O_130,N_29284,N_28049);
or UO_131 (O_131,N_29724,N_28059);
xor UO_132 (O_132,N_28614,N_29016);
xor UO_133 (O_133,N_28516,N_29153);
and UO_134 (O_134,N_28662,N_29818);
nand UO_135 (O_135,N_29629,N_29552);
nor UO_136 (O_136,N_29124,N_29145);
nand UO_137 (O_137,N_28532,N_29580);
nor UO_138 (O_138,N_28437,N_28188);
nand UO_139 (O_139,N_28915,N_29781);
and UO_140 (O_140,N_28215,N_28944);
nor UO_141 (O_141,N_29556,N_28737);
nand UO_142 (O_142,N_28181,N_29503);
nand UO_143 (O_143,N_28865,N_29612);
nor UO_144 (O_144,N_28861,N_28304);
or UO_145 (O_145,N_28776,N_28778);
and UO_146 (O_146,N_28054,N_29807);
xnor UO_147 (O_147,N_29925,N_29437);
nand UO_148 (O_148,N_28775,N_29721);
nand UO_149 (O_149,N_28528,N_28005);
xnor UO_150 (O_150,N_29761,N_28355);
or UO_151 (O_151,N_29948,N_29678);
and UO_152 (O_152,N_29619,N_29903);
nand UO_153 (O_153,N_28140,N_29774);
nand UO_154 (O_154,N_29249,N_28334);
xnor UO_155 (O_155,N_28311,N_28591);
and UO_156 (O_156,N_28124,N_28634);
nor UO_157 (O_157,N_28832,N_28960);
and UO_158 (O_158,N_29776,N_29637);
nand UO_159 (O_159,N_28348,N_29611);
xnor UO_160 (O_160,N_28874,N_29773);
nand UO_161 (O_161,N_28975,N_28674);
and UO_162 (O_162,N_28234,N_29716);
nand UO_163 (O_163,N_29533,N_28664);
xor UO_164 (O_164,N_28327,N_29151);
and UO_165 (O_165,N_28760,N_28061);
xor UO_166 (O_166,N_28869,N_29892);
or UO_167 (O_167,N_28731,N_28540);
and UO_168 (O_168,N_29863,N_28411);
or UO_169 (O_169,N_28785,N_29522);
and UO_170 (O_170,N_29148,N_28629);
nand UO_171 (O_171,N_29379,N_29859);
or UO_172 (O_172,N_28288,N_28115);
xor UO_173 (O_173,N_28074,N_28854);
and UO_174 (O_174,N_29567,N_28657);
nor UO_175 (O_175,N_28699,N_28428);
nor UO_176 (O_176,N_29957,N_28976);
nor UO_177 (O_177,N_29529,N_29633);
xor UO_178 (O_178,N_29762,N_29965);
xor UO_179 (O_179,N_28619,N_29179);
nand UO_180 (O_180,N_28748,N_28647);
xnor UO_181 (O_181,N_29282,N_28372);
and UO_182 (O_182,N_28840,N_28400);
xnor UO_183 (O_183,N_28918,N_29014);
xnor UO_184 (O_184,N_29132,N_29888);
and UO_185 (O_185,N_28741,N_28162);
and UO_186 (O_186,N_29247,N_28802);
and UO_187 (O_187,N_28661,N_29639);
nor UO_188 (O_188,N_29578,N_28896);
nand UO_189 (O_189,N_29729,N_28200);
and UO_190 (O_190,N_29012,N_28804);
or UO_191 (O_191,N_29383,N_28409);
xnor UO_192 (O_192,N_29869,N_29089);
nor UO_193 (O_193,N_28864,N_29460);
and UO_194 (O_194,N_29878,N_28644);
xor UO_195 (O_195,N_28338,N_28749);
xnor UO_196 (O_196,N_28232,N_29953);
or UO_197 (O_197,N_28497,N_28303);
and UO_198 (O_198,N_28314,N_29501);
xor UO_199 (O_199,N_29293,N_28559);
nor UO_200 (O_200,N_28287,N_28316);
nor UO_201 (O_201,N_29597,N_29295);
nand UO_202 (O_202,N_29386,N_29575);
and UO_203 (O_203,N_29844,N_28105);
or UO_204 (O_204,N_29495,N_29059);
and UO_205 (O_205,N_29439,N_29402);
nor UO_206 (O_206,N_29565,N_29245);
or UO_207 (O_207,N_28248,N_29422);
nand UO_208 (O_208,N_28550,N_29631);
nand UO_209 (O_209,N_28242,N_28211);
nand UO_210 (O_210,N_29651,N_29222);
nand UO_211 (O_211,N_29539,N_28726);
nand UO_212 (O_212,N_29283,N_28130);
or UO_213 (O_213,N_29998,N_29180);
xnor UO_214 (O_214,N_28191,N_29048);
and UO_215 (O_215,N_29259,N_28763);
nand UO_216 (O_216,N_29555,N_28064);
nor UO_217 (O_217,N_28692,N_28702);
nor UO_218 (O_218,N_28556,N_29933);
or UO_219 (O_219,N_28383,N_29349);
nor UO_220 (O_220,N_28109,N_28593);
nor UO_221 (O_221,N_29845,N_29322);
nor UO_222 (O_222,N_29392,N_29274);
nand UO_223 (O_223,N_29988,N_29028);
nand UO_224 (O_224,N_29094,N_28326);
and UO_225 (O_225,N_29674,N_28293);
and UO_226 (O_226,N_29609,N_28149);
nor UO_227 (O_227,N_28937,N_29021);
or UO_228 (O_228,N_29419,N_28380);
or UO_229 (O_229,N_29671,N_28803);
or UO_230 (O_230,N_28827,N_28911);
nor UO_231 (O_231,N_29796,N_29820);
nand UO_232 (O_232,N_29384,N_29833);
xor UO_233 (O_233,N_29017,N_28672);
or UO_234 (O_234,N_28565,N_29418);
xor UO_235 (O_235,N_28536,N_28570);
xor UO_236 (O_236,N_28863,N_29610);
or UO_237 (O_237,N_29974,N_28517);
nor UO_238 (O_238,N_29628,N_29598);
nand UO_239 (O_239,N_29144,N_28666);
nor UO_240 (O_240,N_28835,N_28399);
xor UO_241 (O_241,N_28292,N_29650);
or UO_242 (O_242,N_29686,N_29615);
and UO_243 (O_243,N_28772,N_29868);
nand UO_244 (O_244,N_28585,N_29080);
xnor UO_245 (O_245,N_29061,N_28265);
and UO_246 (O_246,N_29968,N_28196);
and UO_247 (O_247,N_29009,N_28212);
xor UO_248 (O_248,N_28753,N_28179);
and UO_249 (O_249,N_28880,N_29381);
nand UO_250 (O_250,N_28480,N_29636);
xnor UO_251 (O_251,N_28405,N_28558);
xor UO_252 (O_252,N_29434,N_29561);
xnor UO_253 (O_253,N_28888,N_28493);
nor UO_254 (O_254,N_28793,N_29887);
and UO_255 (O_255,N_28247,N_29286);
or UO_256 (O_256,N_28343,N_28901);
and UO_257 (O_257,N_28855,N_29956);
or UO_258 (O_258,N_28946,N_29074);
xor UO_259 (O_259,N_28354,N_28096);
nand UO_260 (O_260,N_29003,N_29468);
nand UO_261 (O_261,N_29743,N_28678);
nor UO_262 (O_262,N_28254,N_29416);
nor UO_263 (O_263,N_29025,N_28733);
nand UO_264 (O_264,N_29278,N_28237);
or UO_265 (O_265,N_29592,N_28081);
or UO_266 (O_266,N_29778,N_29780);
nand UO_267 (O_267,N_29234,N_28098);
xor UO_268 (O_268,N_28168,N_28642);
or UO_269 (O_269,N_28996,N_29786);
xor UO_270 (O_270,N_29617,N_28679);
xor UO_271 (O_271,N_28867,N_28113);
and UO_272 (O_272,N_28499,N_29253);
nand UO_273 (O_273,N_28402,N_29344);
nand UO_274 (O_274,N_28894,N_28114);
and UO_275 (O_275,N_29966,N_28922);
nand UO_276 (O_276,N_29788,N_29606);
nand UO_277 (O_277,N_28983,N_28020);
nand UO_278 (O_278,N_28650,N_29934);
xor UO_279 (O_279,N_28335,N_29476);
and UO_280 (O_280,N_29216,N_29816);
nand UO_281 (O_281,N_29239,N_28154);
nand UO_282 (O_282,N_28754,N_29725);
or UO_283 (O_283,N_29623,N_29129);
xor UO_284 (O_284,N_29544,N_29919);
and UO_285 (O_285,N_28361,N_28161);
or UO_286 (O_286,N_29432,N_29397);
nand UO_287 (O_287,N_28241,N_29233);
and UO_288 (O_288,N_29206,N_29070);
xnor UO_289 (O_289,N_29455,N_29276);
xnor UO_290 (O_290,N_29351,N_29564);
nand UO_291 (O_291,N_28445,N_29532);
nand UO_292 (O_292,N_29950,N_29023);
nor UO_293 (O_293,N_28144,N_29826);
or UO_294 (O_294,N_28691,N_28312);
and UO_295 (O_295,N_28342,N_28371);
and UO_296 (O_296,N_29352,N_28477);
nand UO_297 (O_297,N_28615,N_29814);
xnor UO_298 (O_298,N_28732,N_29441);
xor UO_299 (O_299,N_28427,N_29586);
nand UO_300 (O_300,N_29127,N_28701);
and UO_301 (O_301,N_29160,N_29128);
nand UO_302 (O_302,N_28302,N_29902);
xor UO_303 (O_303,N_28134,N_29433);
or UO_304 (O_304,N_28843,N_28838);
nor UO_305 (O_305,N_28909,N_28799);
nor UO_306 (O_306,N_29373,N_28457);
nand UO_307 (O_307,N_28900,N_29307);
nand UO_308 (O_308,N_28618,N_29102);
and UO_309 (O_309,N_28997,N_29008);
nand UO_310 (O_310,N_28980,N_28576);
nand UO_311 (O_311,N_28582,N_29189);
nor UO_312 (O_312,N_29471,N_28801);
nand UO_313 (O_313,N_28189,N_28222);
xnor UO_314 (O_314,N_28373,N_29866);
xnor UO_315 (O_315,N_29287,N_28546);
xnor UO_316 (O_316,N_28547,N_29280);
nor UO_317 (O_317,N_29467,N_28496);
or UO_318 (O_318,N_28491,N_29196);
nand UO_319 (O_319,N_29135,N_29141);
nor UO_320 (O_320,N_28163,N_28083);
xor UO_321 (O_321,N_28735,N_28272);
nand UO_322 (O_322,N_29928,N_29535);
nand UO_323 (O_323,N_28277,N_28458);
nand UO_324 (O_324,N_28949,N_28449);
nand UO_325 (O_325,N_29895,N_28255);
nand UO_326 (O_326,N_29993,N_28368);
and UO_327 (O_327,N_28527,N_29331);
and UO_328 (O_328,N_28815,N_28876);
and UO_329 (O_329,N_29057,N_28966);
xnor UO_330 (O_330,N_28413,N_28484);
nor UO_331 (O_331,N_29103,N_28448);
and UO_332 (O_332,N_29105,N_28921);
or UO_333 (O_333,N_28000,N_28809);
nand UO_334 (O_334,N_28253,N_29961);
or UO_335 (O_335,N_29388,N_29117);
nand UO_336 (O_336,N_29120,N_28752);
and UO_337 (O_337,N_28021,N_29224);
nand UO_338 (O_338,N_29960,N_29042);
nand UO_339 (O_339,N_29746,N_28116);
and UO_340 (O_340,N_28624,N_28845);
xor UO_341 (O_341,N_28283,N_29913);
xor UO_342 (O_342,N_29767,N_28597);
or UO_343 (O_343,N_28447,N_29568);
nor UO_344 (O_344,N_28429,N_29649);
nand UO_345 (O_345,N_29370,N_28167);
and UO_346 (O_346,N_28638,N_29583);
or UO_347 (O_347,N_28385,N_29051);
nor UO_348 (O_348,N_28606,N_29920);
xor UO_349 (O_349,N_28299,N_29257);
nand UO_350 (O_350,N_28525,N_28414);
nand UO_351 (O_351,N_29613,N_29604);
nor UO_352 (O_352,N_29453,N_28301);
nand UO_353 (O_353,N_29213,N_29423);
nor UO_354 (O_354,N_28487,N_28187);
xnor UO_355 (O_355,N_29100,N_28820);
nand UO_356 (O_356,N_29755,N_28455);
nand UO_357 (O_357,N_29595,N_29608);
or UO_358 (O_358,N_28014,N_28668);
and UO_359 (O_359,N_28159,N_29041);
and UO_360 (O_360,N_29645,N_29147);
or UO_361 (O_361,N_29346,N_28461);
and UO_362 (O_362,N_29810,N_29880);
xor UO_363 (O_363,N_28331,N_28267);
nand UO_364 (O_364,N_28476,N_29332);
xnor UO_365 (O_365,N_29977,N_29634);
and UO_366 (O_366,N_29226,N_29795);
nor UO_367 (O_367,N_29210,N_28648);
xnor UO_368 (O_368,N_29749,N_28621);
nor UO_369 (O_369,N_29116,N_29026);
nor UO_370 (O_370,N_28472,N_29273);
xor UO_371 (O_371,N_29712,N_29324);
nand UO_372 (O_372,N_29492,N_28177);
or UO_373 (O_373,N_28819,N_28376);
or UO_374 (O_374,N_28403,N_28590);
nand UO_375 (O_375,N_29837,N_28829);
and UO_376 (O_376,N_28645,N_28961);
and UO_377 (O_377,N_29082,N_28421);
xnor UO_378 (O_378,N_28782,N_29720);
nand UO_379 (O_379,N_29469,N_28280);
nor UO_380 (O_380,N_29236,N_29908);
nand UO_381 (O_381,N_28522,N_29955);
nand UO_382 (O_382,N_28143,N_28719);
nand UO_383 (O_383,N_29485,N_29987);
and UO_384 (O_384,N_28690,N_28029);
nor UO_385 (O_385,N_28218,N_28694);
or UO_386 (O_386,N_28505,N_28093);
nand UO_387 (O_387,N_29197,N_29970);
or UO_388 (O_388,N_28347,N_29447);
or UO_389 (O_389,N_28652,N_28641);
nor UO_390 (O_390,N_29420,N_29269);
xnor UO_391 (O_391,N_29391,N_28417);
and UO_392 (O_392,N_29336,N_28193);
and UO_393 (O_393,N_28295,N_28521);
and UO_394 (O_394,N_28340,N_28800);
and UO_395 (O_395,N_29765,N_29394);
nor UO_396 (O_396,N_28063,N_29406);
nor UO_397 (O_397,N_29943,N_29275);
and UO_398 (O_398,N_28336,N_28940);
nor UO_399 (O_399,N_29952,N_28510);
nor UO_400 (O_400,N_29266,N_29451);
and UO_401 (O_401,N_28950,N_29548);
or UO_402 (O_402,N_28566,N_28249);
nor UO_403 (O_403,N_28069,N_28630);
nor UO_404 (O_404,N_28720,N_29097);
nor UO_405 (O_405,N_29800,N_29137);
and UO_406 (O_406,N_29939,N_28219);
and UO_407 (O_407,N_29758,N_28626);
and UO_408 (O_408,N_29002,N_28765);
nor UO_409 (O_409,N_29854,N_28956);
nand UO_410 (O_410,N_28278,N_28529);
or UO_411 (O_411,N_29581,N_28194);
nor UO_412 (O_412,N_28740,N_29764);
nand UO_413 (O_413,N_28953,N_29894);
nand UO_414 (O_414,N_29990,N_29164);
xnor UO_415 (O_415,N_28062,N_28110);
and UO_416 (O_416,N_28004,N_28147);
nand UO_417 (O_417,N_28165,N_29475);
and UO_418 (O_418,N_28553,N_28999);
and UO_419 (O_419,N_29511,N_29681);
nor UO_420 (O_420,N_28043,N_29829);
or UO_421 (O_421,N_28356,N_28724);
xnor UO_422 (O_422,N_29294,N_28920);
or UO_423 (O_423,N_29715,N_28526);
nor UO_424 (O_424,N_29647,N_29005);
nand UO_425 (O_425,N_28099,N_28916);
nor UO_426 (O_426,N_29109,N_29188);
or UO_427 (O_427,N_29679,N_28817);
and UO_428 (O_428,N_29264,N_29355);
and UO_429 (O_429,N_29752,N_29013);
nor UO_430 (O_430,N_29463,N_29265);
nand UO_431 (O_431,N_29646,N_28851);
xor UO_432 (O_432,N_28426,N_28344);
or UO_433 (O_433,N_29367,N_28581);
and UO_434 (O_434,N_28418,N_29593);
nor UO_435 (O_435,N_28750,N_29999);
nand UO_436 (O_436,N_28157,N_29228);
nor UO_437 (O_437,N_28523,N_28231);
or UO_438 (O_438,N_28531,N_29461);
or UO_439 (O_439,N_28329,N_29396);
and UO_440 (O_440,N_28780,N_29215);
or UO_441 (O_441,N_29403,N_29341);
nor UO_442 (O_442,N_29490,N_29032);
or UO_443 (O_443,N_28141,N_28082);
or UO_444 (O_444,N_28126,N_29121);
nand UO_445 (O_445,N_29882,N_29857);
or UO_446 (O_446,N_28577,N_29365);
and UO_447 (O_447,N_28611,N_28271);
and UO_448 (O_448,N_28032,N_29312);
nor UO_449 (O_449,N_29940,N_28715);
or UO_450 (O_450,N_29803,N_28407);
nor UO_451 (O_451,N_29850,N_28917);
nand UO_452 (O_452,N_28164,N_29547);
nand UO_453 (O_453,N_28848,N_29348);
nor UO_454 (O_454,N_29889,N_29558);
and UO_455 (O_455,N_28932,N_28036);
nand UO_456 (O_456,N_28057,N_29347);
or UO_457 (O_457,N_28744,N_29454);
and UO_458 (O_458,N_29959,N_29360);
nand UO_459 (O_459,N_28259,N_28101);
or UO_460 (O_460,N_29938,N_29665);
and UO_461 (O_461,N_29877,N_28037);
nor UO_462 (O_462,N_29301,N_28862);
and UO_463 (O_463,N_29242,N_28613);
or UO_464 (O_464,N_29941,N_28470);
nor UO_465 (O_465,N_28518,N_29707);
xnor UO_466 (O_466,N_28238,N_29574);
nand UO_467 (O_467,N_28274,N_29802);
and UO_468 (O_468,N_29260,N_29177);
nor UO_469 (O_469,N_29306,N_29169);
and UO_470 (O_470,N_29150,N_28310);
or UO_471 (O_471,N_29525,N_29830);
or UO_472 (O_472,N_29875,N_29760);
or UO_473 (O_473,N_29906,N_28425);
nor UO_474 (O_474,N_29757,N_29675);
nor UO_475 (O_475,N_28464,N_29572);
nand UO_476 (O_476,N_28991,N_29178);
and UO_477 (O_477,N_29149,N_28736);
or UO_478 (O_478,N_28882,N_28884);
and UO_479 (O_479,N_29983,N_29848);
or UO_480 (O_480,N_29256,N_28463);
or UO_481 (O_481,N_28746,N_28148);
or UO_482 (O_482,N_28220,N_28758);
and UO_483 (O_483,N_29364,N_29812);
nand UO_484 (O_484,N_28628,N_29670);
or UO_485 (O_485,N_28513,N_29409);
xnor UO_486 (O_486,N_28622,N_28795);
nand UO_487 (O_487,N_28075,N_28509);
nand UO_488 (O_488,N_29573,N_28654);
and UO_489 (O_489,N_28180,N_29911);
nor UO_490 (O_490,N_29119,N_28533);
nor UO_491 (O_491,N_28879,N_28927);
nor UO_492 (O_492,N_28430,N_28174);
nand UO_493 (O_493,N_28646,N_29885);
nand UO_494 (O_494,N_28135,N_28107);
nor UO_495 (O_495,N_29194,N_29248);
and UO_496 (O_496,N_29208,N_28388);
and UO_497 (O_497,N_29717,N_28813);
and UO_498 (O_498,N_28419,N_29589);
nor UO_499 (O_499,N_29214,N_28467);
nand UO_500 (O_500,N_29096,N_29945);
nand UO_501 (O_501,N_28038,N_28045);
xor UO_502 (O_502,N_28315,N_28695);
and UO_503 (O_503,N_29982,N_28739);
and UO_504 (O_504,N_29115,N_28537);
nand UO_505 (O_505,N_29683,N_28607);
or UO_506 (O_506,N_28067,N_28046);
or UO_507 (O_507,N_28401,N_28291);
nor UO_508 (O_508,N_29479,N_29326);
nand UO_509 (O_509,N_29779,N_29255);
nand UO_510 (O_510,N_29669,N_28459);
xnor UO_511 (O_511,N_28866,N_29841);
nor UO_512 (O_512,N_29602,N_28985);
and UO_513 (O_513,N_29672,N_28805);
and UO_514 (O_514,N_28913,N_28111);
and UO_515 (O_515,N_28252,N_29123);
and UO_516 (O_516,N_28609,N_28544);
nand UO_517 (O_517,N_29218,N_28839);
and UO_518 (O_518,N_28013,N_29865);
xnor UO_519 (O_519,N_29731,N_28268);
or UO_520 (O_520,N_29050,N_28512);
xor UO_521 (O_521,N_28881,N_29513);
xor UO_522 (O_522,N_29550,N_28050);
nor UO_523 (O_523,N_28673,N_28284);
nand UO_524 (O_524,N_28660,N_29157);
nor UO_525 (O_525,N_29049,N_29912);
and UO_526 (O_526,N_28623,N_28564);
or UO_527 (O_527,N_29577,N_28025);
xor UO_528 (O_528,N_29664,N_29060);
or UO_529 (O_529,N_29530,N_29193);
nand UO_530 (O_530,N_28768,N_28936);
xnor UO_531 (O_531,N_28016,N_29155);
nand UO_532 (O_532,N_29167,N_28893);
or UO_533 (O_533,N_28886,N_29314);
xor UO_534 (O_534,N_28588,N_28589);
or UO_535 (O_535,N_28555,N_28035);
xnor UO_536 (O_536,N_28538,N_28369);
or UO_537 (O_537,N_28769,N_29340);
or UO_538 (O_538,N_29431,N_29086);
nor UO_539 (O_539,N_29143,N_29684);
or UO_540 (O_540,N_29745,N_29443);
and UO_541 (O_541,N_29517,N_29470);
nor UO_542 (O_542,N_28967,N_28955);
nand UO_543 (O_543,N_28824,N_29677);
nor UO_544 (O_544,N_29954,N_29378);
and UO_545 (O_545,N_29072,N_29084);
nand UO_546 (O_546,N_28201,N_29981);
or UO_547 (O_547,N_28456,N_29079);
nand UO_548 (O_548,N_28790,N_29616);
and UO_549 (O_549,N_28003,N_28655);
nor UO_550 (O_550,N_29905,N_28689);
or UO_551 (O_551,N_28153,N_29390);
and UO_552 (O_552,N_29241,N_29744);
and UO_553 (O_553,N_28197,N_28595);
nor UO_554 (O_554,N_29727,N_29688);
xor UO_555 (O_555,N_28905,N_29404);
or UO_556 (O_556,N_29756,N_29566);
or UO_557 (O_557,N_29466,N_28122);
nor UO_558 (O_558,N_29946,N_28151);
nand UO_559 (O_559,N_29413,N_28988);
nor UO_560 (O_560,N_28090,N_28912);
nor UO_561 (O_561,N_29831,N_28859);
xnor UO_562 (O_562,N_28977,N_28658);
xnor UO_563 (O_563,N_29085,N_29095);
and UO_564 (O_564,N_28723,N_28321);
nor UO_565 (O_565,N_28444,N_28441);
nor UO_566 (O_566,N_28830,N_28535);
xnor UO_567 (O_567,N_28071,N_29909);
nand UO_568 (O_568,N_28465,N_29310);
or UO_569 (O_569,N_28225,N_29296);
nor UO_570 (O_570,N_28432,N_29838);
nand UO_571 (O_571,N_28906,N_29281);
and UO_572 (O_572,N_29935,N_28246);
xor UO_573 (O_573,N_28007,N_28969);
xor UO_574 (O_574,N_28710,N_28959);
xnor UO_575 (O_575,N_29986,N_29330);
xor UO_576 (O_576,N_29927,N_28370);
and UO_577 (O_577,N_28156,N_28561);
xnor UO_578 (O_578,N_29417,N_29254);
xnor UO_579 (O_579,N_28954,N_28392);
xor UO_580 (O_580,N_28424,N_29162);
and UO_581 (O_581,N_29438,N_29232);
and UO_582 (O_582,N_28637,N_28023);
and UO_583 (O_583,N_28781,N_29198);
and UO_584 (O_584,N_28635,N_29985);
and UO_585 (O_585,N_29363,N_28072);
nor UO_586 (O_586,N_29329,N_29682);
nor UO_587 (O_587,N_29130,N_28221);
xor UO_588 (O_588,N_29090,N_28080);
nor UO_589 (O_589,N_28981,N_29319);
xnor UO_590 (O_590,N_29907,N_29184);
xnor UO_591 (O_591,N_29223,N_28681);
or UO_592 (O_592,N_29518,N_28552);
nand UO_593 (O_593,N_28040,N_29170);
nand UO_594 (O_594,N_28745,N_28269);
nand UO_595 (O_595,N_28172,N_29797);
nand UO_596 (O_596,N_29704,N_29971);
xor UO_597 (O_597,N_28131,N_28317);
or UO_598 (O_598,N_28928,N_28774);
or UO_599 (O_599,N_28685,N_29183);
nand UO_600 (O_600,N_29740,N_28257);
or UO_601 (O_601,N_29932,N_28094);
nor UO_602 (O_602,N_29742,N_29687);
and UO_603 (O_603,N_29063,N_29697);
xnor UO_604 (O_604,N_28479,N_29799);
and UO_605 (O_605,N_28022,N_29456);
xnor UO_606 (O_606,N_28818,N_28452);
and UO_607 (O_607,N_29313,N_29531);
nor UO_608 (O_608,N_28942,N_29401);
nand UO_609 (O_609,N_29673,N_29393);
or UO_610 (O_610,N_29237,N_28363);
nand UO_611 (O_611,N_28903,N_28433);
nor UO_612 (O_612,N_28214,N_28514);
and UO_613 (O_613,N_28730,N_28982);
or UO_614 (O_614,N_28575,N_28012);
nand UO_615 (O_615,N_28481,N_28305);
or UO_616 (O_616,N_28856,N_29449);
and UO_617 (O_617,N_29015,N_29361);
xnor UO_618 (O_618,N_29819,N_29676);
nor UO_619 (O_619,N_29412,N_29004);
or UO_620 (O_620,N_29728,N_29557);
nand UO_621 (O_621,N_28308,N_28264);
nand UO_622 (O_622,N_28341,N_28992);
nand UO_623 (O_623,N_28435,N_28097);
or UO_624 (O_624,N_29827,N_29131);
nand UO_625 (O_625,N_29493,N_28783);
nor UO_626 (O_626,N_28065,N_28216);
nand UO_627 (O_627,N_29415,N_29220);
nand UO_628 (O_628,N_28387,N_28592);
and UO_629 (O_629,N_29784,N_28398);
xor UO_630 (O_630,N_28812,N_29484);
nand UO_631 (O_631,N_28438,N_29922);
nand UO_632 (O_632,N_29536,N_28777);
xor UO_633 (O_633,N_29385,N_28738);
xnor UO_634 (O_634,N_28571,N_29375);
or UO_635 (O_635,N_29969,N_28506);
and UO_636 (O_636,N_29864,N_29874);
or UO_637 (O_637,N_28519,N_29267);
xor UO_638 (O_638,N_28825,N_29576);
and UO_639 (O_639,N_29268,N_29472);
nor UO_640 (O_640,N_29702,N_29787);
or UO_641 (O_641,N_29270,N_29125);
nand UO_642 (O_642,N_28670,N_29711);
nand UO_643 (O_643,N_29345,N_29657);
xor UO_644 (O_644,N_28703,N_29929);
or UO_645 (O_645,N_29734,N_28352);
nand UO_646 (O_646,N_28494,N_29733);
and UO_647 (O_647,N_28712,N_29621);
nand UO_648 (O_648,N_29750,N_28446);
or UO_649 (O_649,N_28713,N_29289);
xnor UO_650 (O_650,N_29685,N_28757);
and UO_651 (O_651,N_29989,N_29353);
or UO_652 (O_652,N_28883,N_28223);
or UO_653 (O_653,N_28182,N_29040);
nor UO_654 (O_654,N_29763,N_29019);
and UO_655 (O_655,N_29395,N_28796);
nand UO_656 (O_656,N_29187,N_28227);
and UO_657 (O_657,N_28993,N_28133);
nor UO_658 (O_658,N_28478,N_29399);
xnor UO_659 (O_659,N_29338,N_28791);
or UO_660 (O_660,N_28704,N_28282);
nand UO_661 (O_661,N_29732,N_28053);
or UO_662 (O_662,N_29847,N_29064);
nand UO_663 (O_663,N_29101,N_28604);
nor UO_664 (O_664,N_28137,N_28667);
nand UO_665 (O_665,N_29007,N_29849);
xnor UO_666 (O_666,N_28979,N_29588);
xor UO_667 (O_667,N_29092,N_29596);
and UO_668 (O_668,N_28471,N_28379);
or UO_669 (O_669,N_29159,N_28834);
nand UO_670 (O_670,N_28423,N_28150);
nor UO_671 (O_671,N_29436,N_28926);
nor UO_672 (O_672,N_29305,N_28307);
nor UO_673 (O_673,N_28474,N_28207);
nand UO_674 (O_674,N_29630,N_28008);
or UO_675 (O_675,N_28633,N_29923);
or UO_676 (O_676,N_28572,N_28010);
and UO_677 (O_677,N_29133,N_28594);
or UO_678 (O_678,N_28410,N_29158);
nand UO_679 (O_679,N_28586,N_28792);
and UO_680 (O_680,N_29936,N_29045);
or UO_681 (O_681,N_28717,N_28209);
xnor UO_682 (O_682,N_29335,N_29714);
or UO_683 (O_683,N_28503,N_29114);
or UO_684 (O_684,N_29792,N_28889);
or UO_685 (O_685,N_28378,N_28251);
and UO_686 (O_686,N_28243,N_28823);
nor UO_687 (O_687,N_29478,N_28669);
and UO_688 (O_688,N_29915,N_28404);
and UO_689 (O_689,N_28203,N_28048);
and UO_690 (O_690,N_29545,N_28384);
nor UO_691 (O_691,N_29914,N_29022);
and UO_692 (O_692,N_29029,N_29288);
nand UO_693 (O_693,N_28687,N_28828);
or UO_694 (O_694,N_29088,N_28175);
and UO_695 (O_695,N_29992,N_28958);
nand UO_696 (O_696,N_28860,N_29071);
or UO_697 (O_697,N_28100,N_29166);
nand UO_698 (O_698,N_29846,N_28659);
nand UO_699 (O_699,N_28390,N_28394);
or UO_700 (O_700,N_28158,N_29011);
or UO_701 (O_701,N_29947,N_29709);
xor UO_702 (O_702,N_28947,N_29747);
nand UO_703 (O_703,N_28562,N_28056);
xnor UO_704 (O_704,N_28039,N_28989);
nor UO_705 (O_705,N_29425,N_29808);
nor UO_706 (O_706,N_28807,N_28364);
xnor UO_707 (O_707,N_29140,N_29387);
nand UO_708 (O_708,N_28963,N_28486);
or UO_709 (O_709,N_28337,N_29112);
or UO_710 (O_710,N_29916,N_28127);
nand UO_711 (O_711,N_28598,N_28286);
or UO_712 (O_712,N_28125,N_29046);
and UO_713 (O_713,N_28850,N_28871);
or UO_714 (O_714,N_28579,N_29766);
xor UO_715 (O_715,N_28891,N_29661);
nand UO_716 (O_716,N_29350,N_28152);
or UO_717 (O_717,N_28986,N_28068);
nor UO_718 (O_718,N_29554,N_29790);
nor UO_719 (O_719,N_29327,N_28770);
nand UO_720 (O_720,N_29815,N_28837);
nor UO_721 (O_721,N_29065,N_28974);
and UO_722 (O_722,N_29093,N_29668);
nand UO_723 (O_723,N_28236,N_29540);
xor UO_724 (O_724,N_28601,N_28306);
xnor UO_725 (O_725,N_29730,N_28490);
nor UO_726 (O_726,N_28945,N_29654);
xor UO_727 (O_727,N_29446,N_28088);
or UO_728 (O_728,N_29722,N_28030);
xor UO_729 (O_729,N_28995,N_29077);
or UO_730 (O_730,N_29261,N_28206);
or UO_731 (O_731,N_28873,N_28079);
xor UO_732 (O_732,N_29809,N_29113);
xor UO_733 (O_733,N_28683,N_29457);
nor UO_734 (O_734,N_29191,N_29299);
or UO_735 (O_735,N_28930,N_29543);
and UO_736 (O_736,N_28545,N_28171);
nand UO_737 (O_737,N_29871,N_29893);
or UO_738 (O_738,N_29481,N_28984);
or UO_739 (O_739,N_29884,N_29410);
or UO_740 (O_740,N_28018,N_29357);
nor UO_741 (O_741,N_28475,N_28808);
nor UO_742 (O_742,N_28450,N_28957);
nand UO_743 (O_743,N_28705,N_29426);
nand UO_744 (O_744,N_29081,N_28706);
nand UO_745 (O_745,N_29368,N_28240);
nand UO_746 (O_746,N_29182,N_29359);
or UO_747 (O_747,N_29024,N_29693);
and UO_748 (O_748,N_29376,N_29921);
xnor UO_749 (O_749,N_28192,N_28617);
nand UO_750 (O_750,N_28178,N_29924);
xor UO_751 (O_751,N_29421,N_28548);
nor UO_752 (O_752,N_29277,N_29655);
or UO_753 (O_753,N_28258,N_28121);
nor UO_754 (O_754,N_29201,N_29791);
or UO_755 (O_755,N_29315,N_28250);
nand UO_756 (O_756,N_29860,N_29828);
xnor UO_757 (O_757,N_29735,N_29660);
nand UO_758 (O_758,N_28393,N_29069);
xnor UO_759 (O_759,N_29635,N_28696);
nand UO_760 (O_760,N_29500,N_28878);
nand UO_761 (O_761,N_29862,N_28453);
nand UO_762 (O_762,N_28087,N_28024);
nor UO_763 (O_763,N_28434,N_29477);
or UO_764 (O_764,N_29843,N_28226);
or UO_765 (O_765,N_29424,N_28263);
xor UO_766 (O_766,N_28786,N_28729);
and UO_767 (O_767,N_28875,N_29428);
nor UO_768 (O_768,N_28330,N_29243);
xor UO_769 (O_769,N_28395,N_28084);
or UO_770 (O_770,N_29377,N_28102);
xor UO_771 (O_771,N_29785,N_29798);
nor UO_772 (O_772,N_29300,N_29739);
nor UO_773 (O_773,N_29018,N_28938);
and UO_774 (O_774,N_28027,N_29285);
xnor UO_775 (O_775,N_28391,N_28047);
xor UO_776 (O_776,N_29632,N_28166);
and UO_777 (O_777,N_29605,N_29321);
nor UO_778 (O_778,N_29356,N_28145);
and UO_779 (O_779,N_28155,N_28204);
nand UO_780 (O_780,N_29343,N_29823);
xnor UO_781 (O_781,N_28119,N_28469);
nor UO_782 (O_782,N_28184,N_29759);
nand UO_783 (O_783,N_29473,N_28205);
or UO_784 (O_784,N_28332,N_29448);
nand UO_785 (O_785,N_29252,N_29516);
and UO_786 (O_786,N_29445,N_29514);
xnor UO_787 (O_787,N_28656,N_29754);
xor UO_788 (O_788,N_28256,N_28511);
nand UO_789 (O_789,N_29949,N_28767);
xor UO_790 (O_790,N_29694,N_29250);
nand UO_791 (O_791,N_28001,N_28345);
and UO_792 (O_792,N_29570,N_28764);
nand UO_793 (O_793,N_29099,N_29692);
xnor UO_794 (O_794,N_29834,N_29118);
xnor UO_795 (O_795,N_28743,N_28389);
nor UO_796 (O_796,N_28034,N_29411);
nor UO_797 (O_797,N_28123,N_28129);
nor UO_798 (O_798,N_29618,N_29033);
nand UO_799 (O_799,N_29876,N_29339);
xor UO_800 (O_800,N_28910,N_29689);
or UO_801 (O_801,N_28006,N_29666);
nand UO_802 (O_802,N_29546,N_29001);
nor UO_803 (O_803,N_28076,N_29304);
nor UO_804 (O_804,N_29653,N_29663);
nand UO_805 (O_805,N_28998,N_29056);
or UO_806 (O_806,N_29087,N_29207);
nand UO_807 (O_807,N_28431,N_29290);
xnor UO_808 (O_808,N_28408,N_28440);
xor UO_809 (O_809,N_29967,N_29997);
and UO_810 (O_810,N_29156,N_28146);
nand UO_811 (O_811,N_29483,N_28573);
xor UO_812 (O_812,N_28771,N_29560);
xnor UO_813 (O_813,N_28524,N_29738);
nor UO_814 (O_814,N_28374,N_29309);
xnor UO_815 (O_815,N_28751,N_29200);
nor UO_816 (O_816,N_29271,N_28797);
and UO_817 (O_817,N_28466,N_29462);
nand UO_818 (O_818,N_29559,N_28952);
nand UO_819 (O_819,N_29186,N_28468);
nand UO_820 (O_820,N_29793,N_29010);
nor UO_821 (O_821,N_28639,N_29104);
nand UO_822 (O_822,N_29458,N_28406);
nor UO_823 (O_823,N_28092,N_29973);
nand UO_824 (O_824,N_29870,N_28375);
and UO_825 (O_825,N_28091,N_29777);
nand UO_826 (O_826,N_29505,N_28627);
or UO_827 (O_827,N_29528,N_28972);
nor UO_828 (O_828,N_28349,N_29217);
or UO_829 (O_829,N_28700,N_29899);
and UO_830 (O_830,N_28557,N_29333);
nor UO_831 (O_831,N_28169,N_28492);
nor UO_832 (O_832,N_28320,N_29043);
and UO_833 (O_833,N_29521,N_28887);
nor UO_834 (O_834,N_28709,N_29963);
xnor UO_835 (O_835,N_28877,N_29227);
xnor UO_836 (O_836,N_29861,N_29891);
and UO_837 (O_837,N_28948,N_29107);
nor UO_838 (O_838,N_29726,N_28568);
nand UO_839 (O_839,N_29964,N_29851);
and UO_840 (O_840,N_28643,N_28574);
and UO_841 (O_841,N_28605,N_29083);
xor UO_842 (O_842,N_28319,N_29958);
and UO_843 (O_843,N_29450,N_28734);
or UO_844 (O_844,N_28631,N_28041);
nor UO_845 (O_845,N_29667,N_29171);
and UO_846 (O_846,N_29488,N_29832);
xnor UO_847 (O_847,N_28261,N_28350);
nand UO_848 (O_848,N_28170,N_28651);
and UO_849 (O_849,N_29067,N_29407);
nand UO_850 (O_850,N_29238,N_28964);
and UO_851 (O_851,N_29185,N_28680);
xor UO_852 (O_852,N_29487,N_29703);
xnor UO_853 (O_853,N_28885,N_29298);
or UO_854 (O_854,N_28482,N_29643);
nand UO_855 (O_855,N_28199,N_29648);
nand UO_856 (O_856,N_28502,N_29098);
nand UO_857 (O_857,N_29699,N_29444);
xnor UO_858 (O_858,N_28500,N_28620);
nand UO_859 (O_859,N_29122,N_28534);
nand UO_860 (O_860,N_28925,N_29853);
or UO_861 (O_861,N_29775,N_28120);
xor UO_862 (O_862,N_28033,N_29995);
nand UO_863 (O_863,N_28632,N_29626);
nand UO_864 (O_864,N_29627,N_28990);
xnor UO_865 (O_865,N_28266,N_28584);
nor UO_866 (O_866,N_28462,N_28810);
or UO_867 (O_867,N_28907,N_28747);
nor UO_868 (O_868,N_28333,N_28052);
and UO_869 (O_869,N_28017,N_29640);
nand UO_870 (O_870,N_28042,N_29318);
nor UO_871 (O_871,N_28173,N_28275);
xnor UO_872 (O_872,N_28919,N_28821);
or UO_873 (O_873,N_29813,N_29520);
and UO_874 (O_874,N_29435,N_28583);
or UO_875 (O_875,N_29152,N_28489);
nand UO_876 (O_876,N_28727,N_28442);
or UO_877 (O_877,N_28019,N_29821);
xnor UO_878 (O_878,N_29334,N_29031);
nor UO_879 (O_879,N_28814,N_28244);
nand UO_880 (O_880,N_29600,N_29642);
xor UO_881 (O_881,N_28245,N_28587);
or UO_882 (O_882,N_29811,N_29192);
nand UO_883 (O_883,N_28224,N_29174);
xor UO_884 (O_884,N_29695,N_29569);
or UO_885 (O_885,N_28779,N_29369);
nor UO_886 (O_886,N_29325,N_29962);
nand UO_887 (O_887,N_28070,N_28028);
xor UO_888 (O_888,N_28009,N_28934);
and UO_889 (O_889,N_28725,N_28904);
nand UO_890 (O_890,N_29607,N_29506);
nor UO_891 (O_891,N_28270,N_29931);
nand UO_892 (O_892,N_29279,N_29442);
or UO_893 (O_893,N_29172,N_28698);
or UO_894 (O_894,N_29414,N_28055);
xnor UO_895 (O_895,N_29584,N_28386);
nand UO_896 (O_896,N_29146,N_28108);
or UO_897 (O_897,N_28722,N_29991);
nand UO_898 (O_898,N_28420,N_29622);
nor UO_899 (O_899,N_29225,N_28636);
xor UO_900 (O_900,N_29246,N_28994);
and UO_901 (O_901,N_28530,N_28610);
nand UO_902 (O_902,N_29190,N_28970);
and UO_903 (O_903,N_28811,N_28443);
nand UO_904 (O_904,N_29244,N_29111);
nand UO_905 (O_905,N_29427,N_28935);
xnor UO_906 (O_906,N_28359,N_29883);
xnor UO_907 (O_907,N_29824,N_28515);
xor UO_908 (O_908,N_28965,N_29075);
and UO_909 (O_909,N_29262,N_29263);
xnor UO_910 (O_910,N_29308,N_29173);
or UO_911 (O_911,N_28602,N_28262);
nor UO_912 (O_912,N_29585,N_28377);
nor UO_913 (O_913,N_28852,N_29625);
xnor UO_914 (O_914,N_28139,N_29337);
nand UO_915 (O_915,N_29890,N_29858);
or UO_916 (O_916,N_29817,N_28766);
nand UO_917 (O_917,N_28058,N_28495);
or UO_918 (O_918,N_29509,N_29199);
or UO_919 (O_919,N_29055,N_28868);
nor UO_920 (O_920,N_28870,N_28728);
nand UO_921 (O_921,N_29563,N_29896);
or UO_922 (O_922,N_28580,N_29211);
or UO_923 (O_923,N_28600,N_28788);
xor UO_924 (O_924,N_29496,N_29801);
nand UO_925 (O_925,N_28213,N_28185);
xnor UO_926 (O_926,N_28560,N_28106);
or UO_927 (O_927,N_29163,N_28229);
nand UO_928 (O_928,N_29782,N_29594);
xnor UO_929 (O_929,N_29710,N_29996);
xor UO_930 (O_930,N_29062,N_29068);
or UO_931 (O_931,N_29459,N_28508);
nor UO_932 (O_932,N_29562,N_29108);
or UO_933 (O_933,N_28324,N_28397);
and UO_934 (O_934,N_28924,N_28230);
xor UO_935 (O_935,N_29719,N_28551);
xnor UO_936 (O_936,N_28684,N_29235);
and UO_937 (O_937,N_29881,N_29994);
xor UO_938 (O_938,N_28806,N_28663);
or UO_939 (O_939,N_29175,N_29292);
or UO_940 (O_940,N_28095,N_29855);
xor UO_941 (O_941,N_29320,N_28978);
or UO_942 (O_942,N_29789,N_28895);
and UO_943 (O_943,N_29491,N_28923);
xor UO_944 (O_944,N_29770,N_29582);
nand UO_945 (O_945,N_28603,N_29553);
or UO_946 (O_946,N_29804,N_28104);
nor UO_947 (O_947,N_28520,N_29510);
xnor UO_948 (O_948,N_28296,N_28549);
nor UO_949 (O_949,N_28190,N_29917);
xor UO_950 (O_950,N_29541,N_28939);
or UO_951 (O_951,N_29658,N_28289);
xor UO_952 (O_952,N_29106,N_29342);
nand UO_953 (O_953,N_29783,N_29979);
nor UO_954 (O_954,N_28351,N_28849);
xnor UO_955 (O_955,N_29975,N_29641);
or UO_956 (O_956,N_29737,N_28085);
nor UO_957 (O_957,N_29138,N_28784);
nand UO_958 (O_958,N_28599,N_28504);
nand UO_959 (O_959,N_28671,N_28488);
xor UO_960 (O_960,N_29078,N_29374);
and UO_961 (O_961,N_28415,N_29382);
nor UO_962 (O_962,N_28365,N_28742);
and UO_963 (O_963,N_28826,N_29430);
and UO_964 (O_964,N_28297,N_28160);
xor UO_965 (O_965,N_28787,N_29659);
or UO_966 (O_966,N_28933,N_29590);
and UO_967 (O_967,N_28309,N_29603);
and UO_968 (O_968,N_28325,N_28483);
nor UO_969 (O_969,N_28117,N_28596);
nand UO_970 (O_970,N_28073,N_28451);
nor UO_971 (O_971,N_29706,N_28892);
nor UO_972 (O_972,N_29258,N_28941);
xnor UO_973 (O_973,N_28416,N_29219);
or UO_974 (O_974,N_28773,N_29221);
and UO_975 (O_975,N_29587,N_28328);
nand UO_976 (O_976,N_28794,N_28677);
or UO_977 (O_977,N_29700,N_28051);
nand UO_978 (O_978,N_29571,N_28439);
and UO_979 (O_979,N_29251,N_28460);
xnor UO_980 (O_980,N_29303,N_29489);
nand UO_981 (O_981,N_28346,N_28539);
and UO_982 (O_982,N_28357,N_29537);
or UO_983 (O_983,N_28897,N_28183);
or UO_984 (O_984,N_29482,N_29389);
and UO_985 (O_985,N_29705,N_29229);
nor UO_986 (O_986,N_29918,N_29405);
nor UO_987 (O_987,N_28569,N_29474);
xor UO_988 (O_988,N_28485,N_29291);
xor UO_989 (O_989,N_29452,N_29652);
and UO_990 (O_990,N_29328,N_28176);
and UO_991 (O_991,N_28716,N_28066);
nand UO_992 (O_992,N_29696,N_28353);
nand UO_993 (O_993,N_28396,N_29842);
and UO_994 (O_994,N_28816,N_28290);
xnor UO_995 (O_995,N_28789,N_29772);
and UO_996 (O_996,N_28688,N_28235);
nor UO_997 (O_997,N_29297,N_29951);
nor UO_998 (O_998,N_29886,N_29058);
nand UO_999 (O_999,N_28498,N_29036);
and UO_1000 (O_1000,N_28901,N_28056);
nand UO_1001 (O_1001,N_29266,N_29676);
or UO_1002 (O_1002,N_29717,N_28090);
xor UO_1003 (O_1003,N_28755,N_29864);
nand UO_1004 (O_1004,N_28618,N_29552);
or UO_1005 (O_1005,N_28049,N_28183);
xnor UO_1006 (O_1006,N_29059,N_29563);
xnor UO_1007 (O_1007,N_29697,N_29135);
and UO_1008 (O_1008,N_29682,N_28405);
and UO_1009 (O_1009,N_29854,N_28704);
nand UO_1010 (O_1010,N_29286,N_28842);
nand UO_1011 (O_1011,N_29065,N_28905);
xor UO_1012 (O_1012,N_29564,N_28748);
and UO_1013 (O_1013,N_28235,N_29878);
or UO_1014 (O_1014,N_28835,N_28725);
and UO_1015 (O_1015,N_28164,N_29856);
nor UO_1016 (O_1016,N_29497,N_28416);
or UO_1017 (O_1017,N_28029,N_29151);
xnor UO_1018 (O_1018,N_29391,N_28145);
xor UO_1019 (O_1019,N_29221,N_29337);
nor UO_1020 (O_1020,N_28663,N_28279);
nor UO_1021 (O_1021,N_28871,N_29964);
and UO_1022 (O_1022,N_28432,N_29248);
and UO_1023 (O_1023,N_28727,N_29408);
or UO_1024 (O_1024,N_28975,N_28366);
or UO_1025 (O_1025,N_29602,N_28443);
nor UO_1026 (O_1026,N_28323,N_29885);
or UO_1027 (O_1027,N_29920,N_28274);
xor UO_1028 (O_1028,N_29005,N_28118);
nand UO_1029 (O_1029,N_28240,N_29805);
xor UO_1030 (O_1030,N_28213,N_29654);
nand UO_1031 (O_1031,N_28020,N_28204);
nor UO_1032 (O_1032,N_28492,N_28422);
and UO_1033 (O_1033,N_28291,N_28228);
or UO_1034 (O_1034,N_29811,N_29922);
nand UO_1035 (O_1035,N_28833,N_29321);
xnor UO_1036 (O_1036,N_29057,N_29028);
nor UO_1037 (O_1037,N_29732,N_28798);
xor UO_1038 (O_1038,N_29691,N_28491);
xnor UO_1039 (O_1039,N_29074,N_29536);
xor UO_1040 (O_1040,N_29940,N_29663);
nand UO_1041 (O_1041,N_28927,N_28774);
nand UO_1042 (O_1042,N_28785,N_28636);
xor UO_1043 (O_1043,N_29066,N_28529);
and UO_1044 (O_1044,N_28284,N_29075);
nand UO_1045 (O_1045,N_28710,N_28900);
nand UO_1046 (O_1046,N_29230,N_28318);
xnor UO_1047 (O_1047,N_28418,N_28534);
xor UO_1048 (O_1048,N_28867,N_29322);
or UO_1049 (O_1049,N_29166,N_28851);
and UO_1050 (O_1050,N_28389,N_29009);
nand UO_1051 (O_1051,N_29432,N_29952);
nand UO_1052 (O_1052,N_28421,N_28356);
nand UO_1053 (O_1053,N_28796,N_28042);
xor UO_1054 (O_1054,N_28973,N_29673);
nor UO_1055 (O_1055,N_28048,N_29274);
nand UO_1056 (O_1056,N_29296,N_28071);
nand UO_1057 (O_1057,N_29237,N_28831);
and UO_1058 (O_1058,N_29940,N_28918);
xnor UO_1059 (O_1059,N_28777,N_28378);
and UO_1060 (O_1060,N_29164,N_28892);
xor UO_1061 (O_1061,N_28722,N_28332);
or UO_1062 (O_1062,N_28287,N_28953);
or UO_1063 (O_1063,N_28970,N_29283);
xnor UO_1064 (O_1064,N_29080,N_29467);
and UO_1065 (O_1065,N_29437,N_29537);
nand UO_1066 (O_1066,N_29287,N_29506);
nor UO_1067 (O_1067,N_28545,N_28451);
xor UO_1068 (O_1068,N_28666,N_29012);
and UO_1069 (O_1069,N_29319,N_29616);
nand UO_1070 (O_1070,N_29764,N_28567);
and UO_1071 (O_1071,N_28046,N_28320);
nand UO_1072 (O_1072,N_28674,N_28257);
and UO_1073 (O_1073,N_28840,N_29761);
xnor UO_1074 (O_1074,N_29610,N_28854);
or UO_1075 (O_1075,N_29618,N_29315);
and UO_1076 (O_1076,N_29447,N_28624);
nand UO_1077 (O_1077,N_28968,N_29931);
or UO_1078 (O_1078,N_29861,N_29039);
nor UO_1079 (O_1079,N_29866,N_29066);
nand UO_1080 (O_1080,N_28691,N_29565);
and UO_1081 (O_1081,N_29734,N_29128);
and UO_1082 (O_1082,N_28104,N_29934);
nand UO_1083 (O_1083,N_28486,N_28067);
nor UO_1084 (O_1084,N_28526,N_28196);
or UO_1085 (O_1085,N_28557,N_29074);
or UO_1086 (O_1086,N_28031,N_28114);
nand UO_1087 (O_1087,N_28750,N_28887);
nand UO_1088 (O_1088,N_28455,N_28956);
or UO_1089 (O_1089,N_28038,N_28435);
nand UO_1090 (O_1090,N_28723,N_28959);
nor UO_1091 (O_1091,N_28268,N_28569);
xnor UO_1092 (O_1092,N_29776,N_29304);
xnor UO_1093 (O_1093,N_28371,N_28333);
or UO_1094 (O_1094,N_28618,N_29995);
and UO_1095 (O_1095,N_28150,N_28661);
or UO_1096 (O_1096,N_28936,N_29893);
nor UO_1097 (O_1097,N_28897,N_28575);
or UO_1098 (O_1098,N_28362,N_29203);
and UO_1099 (O_1099,N_29785,N_29276);
or UO_1100 (O_1100,N_28374,N_28865);
and UO_1101 (O_1101,N_28211,N_28673);
nor UO_1102 (O_1102,N_29332,N_29556);
or UO_1103 (O_1103,N_28145,N_29316);
nor UO_1104 (O_1104,N_28971,N_28667);
xnor UO_1105 (O_1105,N_28406,N_28135);
nor UO_1106 (O_1106,N_29874,N_28055);
or UO_1107 (O_1107,N_29625,N_29467);
and UO_1108 (O_1108,N_28657,N_28681);
and UO_1109 (O_1109,N_28496,N_29607);
nor UO_1110 (O_1110,N_29786,N_29643);
xor UO_1111 (O_1111,N_28659,N_29216);
nor UO_1112 (O_1112,N_29549,N_28397);
and UO_1113 (O_1113,N_28776,N_29446);
or UO_1114 (O_1114,N_28893,N_28533);
and UO_1115 (O_1115,N_29249,N_29206);
xor UO_1116 (O_1116,N_28743,N_29293);
nor UO_1117 (O_1117,N_29521,N_28076);
or UO_1118 (O_1118,N_28421,N_29355);
or UO_1119 (O_1119,N_29858,N_28663);
or UO_1120 (O_1120,N_28119,N_28467);
xor UO_1121 (O_1121,N_28712,N_29311);
or UO_1122 (O_1122,N_29943,N_28995);
or UO_1123 (O_1123,N_29179,N_28040);
xor UO_1124 (O_1124,N_29983,N_28388);
or UO_1125 (O_1125,N_29239,N_29063);
and UO_1126 (O_1126,N_28434,N_28915);
and UO_1127 (O_1127,N_28132,N_29986);
nand UO_1128 (O_1128,N_29736,N_29314);
and UO_1129 (O_1129,N_28783,N_28654);
or UO_1130 (O_1130,N_28232,N_28174);
xnor UO_1131 (O_1131,N_29396,N_28406);
xor UO_1132 (O_1132,N_28136,N_28444);
and UO_1133 (O_1133,N_29026,N_28114);
nand UO_1134 (O_1134,N_28662,N_28010);
nor UO_1135 (O_1135,N_29044,N_29448);
and UO_1136 (O_1136,N_28616,N_29031);
and UO_1137 (O_1137,N_29878,N_29843);
and UO_1138 (O_1138,N_29461,N_28883);
xnor UO_1139 (O_1139,N_28764,N_28863);
and UO_1140 (O_1140,N_29655,N_29019);
or UO_1141 (O_1141,N_28774,N_28689);
nor UO_1142 (O_1142,N_28236,N_28163);
xnor UO_1143 (O_1143,N_28403,N_28575);
or UO_1144 (O_1144,N_28271,N_29806);
and UO_1145 (O_1145,N_29517,N_28187);
or UO_1146 (O_1146,N_28322,N_29413);
nor UO_1147 (O_1147,N_29874,N_29492);
nand UO_1148 (O_1148,N_28174,N_28409);
xor UO_1149 (O_1149,N_29308,N_28871);
or UO_1150 (O_1150,N_29700,N_29376);
xnor UO_1151 (O_1151,N_29698,N_28626);
xnor UO_1152 (O_1152,N_28954,N_28650);
or UO_1153 (O_1153,N_29370,N_28375);
nand UO_1154 (O_1154,N_29714,N_28985);
nand UO_1155 (O_1155,N_28110,N_28198);
or UO_1156 (O_1156,N_29376,N_29153);
xor UO_1157 (O_1157,N_29124,N_29921);
or UO_1158 (O_1158,N_29381,N_29243);
and UO_1159 (O_1159,N_28697,N_28866);
and UO_1160 (O_1160,N_28743,N_29923);
nor UO_1161 (O_1161,N_28580,N_29997);
nand UO_1162 (O_1162,N_28499,N_29691);
xor UO_1163 (O_1163,N_29550,N_29671);
nor UO_1164 (O_1164,N_28948,N_28705);
nand UO_1165 (O_1165,N_28879,N_28261);
nor UO_1166 (O_1166,N_28289,N_29999);
nor UO_1167 (O_1167,N_29795,N_28394);
nand UO_1168 (O_1168,N_29110,N_28514);
and UO_1169 (O_1169,N_28963,N_28232);
or UO_1170 (O_1170,N_28822,N_28089);
or UO_1171 (O_1171,N_29734,N_28237);
nand UO_1172 (O_1172,N_28940,N_29107);
xor UO_1173 (O_1173,N_29498,N_28286);
and UO_1174 (O_1174,N_28970,N_28586);
nor UO_1175 (O_1175,N_29013,N_29718);
nand UO_1176 (O_1176,N_28731,N_28706);
and UO_1177 (O_1177,N_28083,N_29888);
and UO_1178 (O_1178,N_28230,N_28504);
or UO_1179 (O_1179,N_28409,N_28154);
nor UO_1180 (O_1180,N_28629,N_29073);
or UO_1181 (O_1181,N_29982,N_29684);
or UO_1182 (O_1182,N_29627,N_28920);
nand UO_1183 (O_1183,N_29206,N_29221);
or UO_1184 (O_1184,N_29759,N_28453);
xor UO_1185 (O_1185,N_29059,N_29417);
and UO_1186 (O_1186,N_28173,N_28017);
xor UO_1187 (O_1187,N_29446,N_28995);
and UO_1188 (O_1188,N_28036,N_29668);
nand UO_1189 (O_1189,N_28718,N_28827);
nor UO_1190 (O_1190,N_29636,N_28524);
and UO_1191 (O_1191,N_29942,N_28029);
xor UO_1192 (O_1192,N_28539,N_28068);
nand UO_1193 (O_1193,N_29739,N_29468);
nor UO_1194 (O_1194,N_28263,N_29976);
nor UO_1195 (O_1195,N_28480,N_29907);
and UO_1196 (O_1196,N_29640,N_29958);
and UO_1197 (O_1197,N_28010,N_28406);
or UO_1198 (O_1198,N_28704,N_29643);
or UO_1199 (O_1199,N_28282,N_29511);
and UO_1200 (O_1200,N_29566,N_28250);
or UO_1201 (O_1201,N_29835,N_28696);
and UO_1202 (O_1202,N_29692,N_29515);
nand UO_1203 (O_1203,N_28599,N_28978);
nor UO_1204 (O_1204,N_29978,N_29692);
nor UO_1205 (O_1205,N_29257,N_28750);
and UO_1206 (O_1206,N_28930,N_28874);
xnor UO_1207 (O_1207,N_28690,N_29532);
and UO_1208 (O_1208,N_29455,N_28749);
xor UO_1209 (O_1209,N_29710,N_29846);
nor UO_1210 (O_1210,N_29618,N_29344);
nand UO_1211 (O_1211,N_29315,N_29666);
or UO_1212 (O_1212,N_28574,N_28722);
xor UO_1213 (O_1213,N_28523,N_29520);
or UO_1214 (O_1214,N_29278,N_29539);
and UO_1215 (O_1215,N_29722,N_29480);
nand UO_1216 (O_1216,N_28668,N_28916);
nor UO_1217 (O_1217,N_28682,N_29864);
xnor UO_1218 (O_1218,N_29588,N_29438);
or UO_1219 (O_1219,N_28840,N_28791);
or UO_1220 (O_1220,N_29427,N_28342);
nor UO_1221 (O_1221,N_29212,N_29187);
or UO_1222 (O_1222,N_29516,N_28305);
or UO_1223 (O_1223,N_28245,N_28700);
nand UO_1224 (O_1224,N_28521,N_28657);
xnor UO_1225 (O_1225,N_28846,N_29313);
nand UO_1226 (O_1226,N_28243,N_28882);
nand UO_1227 (O_1227,N_28164,N_28388);
nor UO_1228 (O_1228,N_28120,N_28825);
nor UO_1229 (O_1229,N_28521,N_28413);
nand UO_1230 (O_1230,N_28572,N_28761);
or UO_1231 (O_1231,N_29362,N_28913);
nand UO_1232 (O_1232,N_28646,N_29393);
and UO_1233 (O_1233,N_29064,N_29094);
nand UO_1234 (O_1234,N_28608,N_28108);
nor UO_1235 (O_1235,N_29309,N_28493);
xnor UO_1236 (O_1236,N_28896,N_29771);
nand UO_1237 (O_1237,N_28631,N_28107);
xor UO_1238 (O_1238,N_29033,N_28974);
nand UO_1239 (O_1239,N_28110,N_29417);
or UO_1240 (O_1240,N_29793,N_29921);
or UO_1241 (O_1241,N_29585,N_28176);
nand UO_1242 (O_1242,N_28477,N_28623);
or UO_1243 (O_1243,N_28805,N_29350);
xor UO_1244 (O_1244,N_29486,N_28335);
and UO_1245 (O_1245,N_28708,N_28269);
nor UO_1246 (O_1246,N_29903,N_29233);
nor UO_1247 (O_1247,N_28814,N_28802);
and UO_1248 (O_1248,N_29771,N_28161);
nor UO_1249 (O_1249,N_29665,N_28495);
and UO_1250 (O_1250,N_29680,N_28151);
nor UO_1251 (O_1251,N_29966,N_28678);
xor UO_1252 (O_1252,N_28036,N_29517);
nor UO_1253 (O_1253,N_28142,N_28250);
nor UO_1254 (O_1254,N_28398,N_28624);
nor UO_1255 (O_1255,N_29091,N_29459);
or UO_1256 (O_1256,N_28401,N_28066);
xor UO_1257 (O_1257,N_28866,N_28628);
nor UO_1258 (O_1258,N_29250,N_28493);
or UO_1259 (O_1259,N_28921,N_29908);
and UO_1260 (O_1260,N_28887,N_28922);
or UO_1261 (O_1261,N_29751,N_28775);
and UO_1262 (O_1262,N_28278,N_28686);
nand UO_1263 (O_1263,N_29399,N_28519);
nand UO_1264 (O_1264,N_28966,N_28264);
xor UO_1265 (O_1265,N_29854,N_28616);
xor UO_1266 (O_1266,N_29814,N_29562);
nand UO_1267 (O_1267,N_29728,N_28629);
nand UO_1268 (O_1268,N_29256,N_28468);
xor UO_1269 (O_1269,N_29178,N_29995);
and UO_1270 (O_1270,N_28011,N_28861);
or UO_1271 (O_1271,N_29375,N_28492);
nand UO_1272 (O_1272,N_28523,N_28641);
xor UO_1273 (O_1273,N_28307,N_28470);
nand UO_1274 (O_1274,N_28512,N_28711);
nand UO_1275 (O_1275,N_28037,N_29824);
and UO_1276 (O_1276,N_29678,N_28651);
or UO_1277 (O_1277,N_29084,N_29374);
and UO_1278 (O_1278,N_28510,N_29964);
nor UO_1279 (O_1279,N_29836,N_28136);
nor UO_1280 (O_1280,N_28329,N_28407);
or UO_1281 (O_1281,N_28417,N_29073);
and UO_1282 (O_1282,N_28180,N_28349);
nand UO_1283 (O_1283,N_28197,N_29812);
nand UO_1284 (O_1284,N_29108,N_29125);
xnor UO_1285 (O_1285,N_28369,N_28325);
and UO_1286 (O_1286,N_28172,N_29926);
nand UO_1287 (O_1287,N_28951,N_29210);
nand UO_1288 (O_1288,N_29080,N_28762);
xor UO_1289 (O_1289,N_29830,N_29295);
xor UO_1290 (O_1290,N_29378,N_28326);
nor UO_1291 (O_1291,N_28707,N_28693);
nor UO_1292 (O_1292,N_29093,N_29468);
xor UO_1293 (O_1293,N_28722,N_29062);
nand UO_1294 (O_1294,N_28819,N_28794);
nor UO_1295 (O_1295,N_28646,N_29073);
nor UO_1296 (O_1296,N_28725,N_29791);
or UO_1297 (O_1297,N_29948,N_29838);
xor UO_1298 (O_1298,N_28654,N_29008);
or UO_1299 (O_1299,N_28641,N_28180);
nand UO_1300 (O_1300,N_29005,N_29488);
nand UO_1301 (O_1301,N_28788,N_29392);
or UO_1302 (O_1302,N_29800,N_29817);
nor UO_1303 (O_1303,N_29167,N_29750);
nor UO_1304 (O_1304,N_28577,N_29114);
nand UO_1305 (O_1305,N_28572,N_29583);
nand UO_1306 (O_1306,N_28613,N_29034);
or UO_1307 (O_1307,N_28393,N_28250);
or UO_1308 (O_1308,N_28658,N_28524);
and UO_1309 (O_1309,N_29394,N_28339);
and UO_1310 (O_1310,N_29917,N_28908);
and UO_1311 (O_1311,N_29722,N_29697);
nor UO_1312 (O_1312,N_29965,N_29928);
or UO_1313 (O_1313,N_29698,N_28522);
nand UO_1314 (O_1314,N_28268,N_28043);
nor UO_1315 (O_1315,N_29640,N_28718);
xor UO_1316 (O_1316,N_28589,N_28737);
nand UO_1317 (O_1317,N_29625,N_28521);
nor UO_1318 (O_1318,N_28816,N_29709);
nor UO_1319 (O_1319,N_29628,N_29029);
or UO_1320 (O_1320,N_29857,N_29567);
nor UO_1321 (O_1321,N_28847,N_28347);
nor UO_1322 (O_1322,N_28527,N_28281);
or UO_1323 (O_1323,N_29009,N_28948);
or UO_1324 (O_1324,N_29995,N_29647);
nand UO_1325 (O_1325,N_29916,N_28239);
nor UO_1326 (O_1326,N_28463,N_29837);
xor UO_1327 (O_1327,N_29785,N_29200);
xor UO_1328 (O_1328,N_28007,N_28820);
or UO_1329 (O_1329,N_28758,N_28827);
or UO_1330 (O_1330,N_29582,N_29565);
xnor UO_1331 (O_1331,N_29917,N_29907);
xnor UO_1332 (O_1332,N_28865,N_29880);
nor UO_1333 (O_1333,N_28750,N_28124);
nor UO_1334 (O_1334,N_28661,N_29362);
nand UO_1335 (O_1335,N_28995,N_29804);
nor UO_1336 (O_1336,N_29919,N_29293);
and UO_1337 (O_1337,N_28278,N_28276);
or UO_1338 (O_1338,N_28699,N_28787);
nor UO_1339 (O_1339,N_28737,N_28002);
or UO_1340 (O_1340,N_28414,N_29460);
nand UO_1341 (O_1341,N_28082,N_28163);
nand UO_1342 (O_1342,N_29606,N_29002);
and UO_1343 (O_1343,N_28677,N_29222);
xor UO_1344 (O_1344,N_29405,N_29813);
nand UO_1345 (O_1345,N_29232,N_29001);
nor UO_1346 (O_1346,N_28578,N_29431);
xor UO_1347 (O_1347,N_28256,N_29806);
nand UO_1348 (O_1348,N_28660,N_28733);
xnor UO_1349 (O_1349,N_29649,N_29445);
or UO_1350 (O_1350,N_29793,N_28339);
or UO_1351 (O_1351,N_28464,N_28186);
nor UO_1352 (O_1352,N_29062,N_28487);
and UO_1353 (O_1353,N_29536,N_28215);
xor UO_1354 (O_1354,N_28033,N_28906);
or UO_1355 (O_1355,N_28422,N_28522);
xnor UO_1356 (O_1356,N_28651,N_29633);
xor UO_1357 (O_1357,N_29770,N_28667);
or UO_1358 (O_1358,N_28165,N_29900);
nand UO_1359 (O_1359,N_29490,N_29081);
or UO_1360 (O_1360,N_29873,N_29787);
xor UO_1361 (O_1361,N_28366,N_28169);
nand UO_1362 (O_1362,N_28964,N_29075);
xnor UO_1363 (O_1363,N_28399,N_29629);
or UO_1364 (O_1364,N_28195,N_28035);
and UO_1365 (O_1365,N_28065,N_29378);
or UO_1366 (O_1366,N_29328,N_29679);
nor UO_1367 (O_1367,N_29048,N_28948);
or UO_1368 (O_1368,N_28522,N_29748);
nor UO_1369 (O_1369,N_29880,N_29418);
and UO_1370 (O_1370,N_28904,N_29058);
nand UO_1371 (O_1371,N_29917,N_28625);
xor UO_1372 (O_1372,N_28215,N_28011);
nand UO_1373 (O_1373,N_28206,N_28693);
xnor UO_1374 (O_1374,N_28925,N_29701);
and UO_1375 (O_1375,N_29554,N_29417);
or UO_1376 (O_1376,N_29834,N_28232);
or UO_1377 (O_1377,N_28932,N_29591);
nand UO_1378 (O_1378,N_29857,N_28269);
nand UO_1379 (O_1379,N_29720,N_29030);
xnor UO_1380 (O_1380,N_28344,N_29934);
or UO_1381 (O_1381,N_28916,N_29609);
nor UO_1382 (O_1382,N_29642,N_29468);
xnor UO_1383 (O_1383,N_28836,N_29846);
or UO_1384 (O_1384,N_28242,N_28523);
or UO_1385 (O_1385,N_29049,N_29323);
or UO_1386 (O_1386,N_28522,N_29411);
nor UO_1387 (O_1387,N_29013,N_28148);
or UO_1388 (O_1388,N_29064,N_28247);
and UO_1389 (O_1389,N_29602,N_29233);
nor UO_1390 (O_1390,N_29879,N_29779);
or UO_1391 (O_1391,N_29242,N_29437);
xnor UO_1392 (O_1392,N_29709,N_28223);
nor UO_1393 (O_1393,N_28397,N_29129);
nor UO_1394 (O_1394,N_29747,N_28277);
nand UO_1395 (O_1395,N_29222,N_29987);
nor UO_1396 (O_1396,N_28980,N_29711);
xnor UO_1397 (O_1397,N_28399,N_28988);
or UO_1398 (O_1398,N_28976,N_28931);
nand UO_1399 (O_1399,N_28991,N_28298);
and UO_1400 (O_1400,N_29988,N_29667);
xor UO_1401 (O_1401,N_29333,N_28139);
or UO_1402 (O_1402,N_28098,N_29138);
and UO_1403 (O_1403,N_29560,N_29419);
or UO_1404 (O_1404,N_28900,N_29708);
xor UO_1405 (O_1405,N_29442,N_28244);
and UO_1406 (O_1406,N_28631,N_28487);
xor UO_1407 (O_1407,N_29245,N_28136);
xor UO_1408 (O_1408,N_29826,N_29162);
nor UO_1409 (O_1409,N_29915,N_28936);
xor UO_1410 (O_1410,N_28682,N_29061);
or UO_1411 (O_1411,N_29925,N_28275);
or UO_1412 (O_1412,N_29491,N_28242);
xnor UO_1413 (O_1413,N_29731,N_29974);
xor UO_1414 (O_1414,N_29888,N_29399);
nand UO_1415 (O_1415,N_29029,N_28003);
nand UO_1416 (O_1416,N_29296,N_29418);
nor UO_1417 (O_1417,N_29940,N_29470);
nor UO_1418 (O_1418,N_28066,N_29882);
and UO_1419 (O_1419,N_28186,N_29231);
xor UO_1420 (O_1420,N_28701,N_28414);
nor UO_1421 (O_1421,N_29964,N_28262);
xor UO_1422 (O_1422,N_28482,N_28896);
xnor UO_1423 (O_1423,N_29069,N_29968);
xor UO_1424 (O_1424,N_29231,N_29690);
nand UO_1425 (O_1425,N_29498,N_29848);
xor UO_1426 (O_1426,N_28878,N_28957);
xor UO_1427 (O_1427,N_29823,N_29476);
and UO_1428 (O_1428,N_28317,N_29596);
and UO_1429 (O_1429,N_29411,N_28345);
xor UO_1430 (O_1430,N_28506,N_29663);
nand UO_1431 (O_1431,N_28145,N_28657);
xnor UO_1432 (O_1432,N_29042,N_28589);
nand UO_1433 (O_1433,N_29754,N_28446);
nor UO_1434 (O_1434,N_28571,N_29388);
nand UO_1435 (O_1435,N_28166,N_29417);
and UO_1436 (O_1436,N_28661,N_29911);
nor UO_1437 (O_1437,N_29117,N_28342);
nor UO_1438 (O_1438,N_29888,N_29218);
nand UO_1439 (O_1439,N_28758,N_28592);
or UO_1440 (O_1440,N_29821,N_29283);
or UO_1441 (O_1441,N_28032,N_29484);
nor UO_1442 (O_1442,N_28274,N_28244);
and UO_1443 (O_1443,N_29938,N_28919);
xnor UO_1444 (O_1444,N_28715,N_28892);
and UO_1445 (O_1445,N_28788,N_29234);
and UO_1446 (O_1446,N_29180,N_29968);
or UO_1447 (O_1447,N_29556,N_29314);
xnor UO_1448 (O_1448,N_28548,N_29226);
nand UO_1449 (O_1449,N_29718,N_29981);
nor UO_1450 (O_1450,N_28089,N_28065);
or UO_1451 (O_1451,N_29956,N_28823);
nand UO_1452 (O_1452,N_28816,N_28831);
and UO_1453 (O_1453,N_29039,N_29589);
or UO_1454 (O_1454,N_29682,N_29570);
nand UO_1455 (O_1455,N_28428,N_29199);
or UO_1456 (O_1456,N_28175,N_28443);
xor UO_1457 (O_1457,N_28043,N_28649);
nor UO_1458 (O_1458,N_28193,N_28887);
nand UO_1459 (O_1459,N_29825,N_29571);
or UO_1460 (O_1460,N_28512,N_28768);
xnor UO_1461 (O_1461,N_28819,N_28358);
xor UO_1462 (O_1462,N_29513,N_29026);
or UO_1463 (O_1463,N_29739,N_28714);
nor UO_1464 (O_1464,N_29768,N_29808);
or UO_1465 (O_1465,N_28190,N_29264);
nor UO_1466 (O_1466,N_29977,N_28789);
and UO_1467 (O_1467,N_29587,N_29621);
and UO_1468 (O_1468,N_29772,N_29350);
and UO_1469 (O_1469,N_29932,N_28980);
or UO_1470 (O_1470,N_28149,N_28111);
nor UO_1471 (O_1471,N_28334,N_28192);
xor UO_1472 (O_1472,N_28774,N_28377);
and UO_1473 (O_1473,N_29615,N_28437);
nand UO_1474 (O_1474,N_29570,N_28039);
nand UO_1475 (O_1475,N_29884,N_29577);
nor UO_1476 (O_1476,N_29234,N_29110);
nand UO_1477 (O_1477,N_28572,N_28297);
and UO_1478 (O_1478,N_29378,N_28268);
xor UO_1479 (O_1479,N_28556,N_29046);
and UO_1480 (O_1480,N_29327,N_29445);
or UO_1481 (O_1481,N_29534,N_28861);
nor UO_1482 (O_1482,N_29595,N_28697);
nor UO_1483 (O_1483,N_29625,N_28301);
nand UO_1484 (O_1484,N_28664,N_28884);
and UO_1485 (O_1485,N_29938,N_28315);
and UO_1486 (O_1486,N_29752,N_29210);
and UO_1487 (O_1487,N_28605,N_29490);
nand UO_1488 (O_1488,N_29916,N_29971);
nand UO_1489 (O_1489,N_29601,N_28746);
xnor UO_1490 (O_1490,N_28302,N_29841);
nor UO_1491 (O_1491,N_28187,N_29660);
or UO_1492 (O_1492,N_28426,N_29587);
or UO_1493 (O_1493,N_28949,N_29888);
xor UO_1494 (O_1494,N_29252,N_28517);
nand UO_1495 (O_1495,N_29859,N_28284);
nor UO_1496 (O_1496,N_28015,N_29420);
or UO_1497 (O_1497,N_28737,N_29813);
xor UO_1498 (O_1498,N_28282,N_28350);
nor UO_1499 (O_1499,N_29356,N_28283);
and UO_1500 (O_1500,N_28846,N_29467);
and UO_1501 (O_1501,N_28283,N_28907);
xor UO_1502 (O_1502,N_29067,N_29249);
or UO_1503 (O_1503,N_29323,N_28602);
nor UO_1504 (O_1504,N_28774,N_29702);
xnor UO_1505 (O_1505,N_28510,N_28025);
nand UO_1506 (O_1506,N_28213,N_28318);
nor UO_1507 (O_1507,N_29707,N_29270);
nand UO_1508 (O_1508,N_28436,N_29335);
and UO_1509 (O_1509,N_28091,N_28419);
nor UO_1510 (O_1510,N_29490,N_28616);
xor UO_1511 (O_1511,N_28592,N_29090);
nand UO_1512 (O_1512,N_28837,N_29180);
or UO_1513 (O_1513,N_29514,N_29859);
nor UO_1514 (O_1514,N_29750,N_29297);
or UO_1515 (O_1515,N_29820,N_29982);
nor UO_1516 (O_1516,N_29191,N_29111);
or UO_1517 (O_1517,N_28982,N_28036);
nand UO_1518 (O_1518,N_29834,N_29114);
or UO_1519 (O_1519,N_28072,N_29530);
xnor UO_1520 (O_1520,N_28991,N_29625);
nand UO_1521 (O_1521,N_28406,N_28720);
and UO_1522 (O_1522,N_28923,N_28436);
nor UO_1523 (O_1523,N_28072,N_28248);
xnor UO_1524 (O_1524,N_28403,N_29456);
nor UO_1525 (O_1525,N_29035,N_29754);
and UO_1526 (O_1526,N_29269,N_29193);
xnor UO_1527 (O_1527,N_28081,N_28890);
or UO_1528 (O_1528,N_29364,N_28936);
nor UO_1529 (O_1529,N_28860,N_29532);
xor UO_1530 (O_1530,N_29989,N_29520);
xor UO_1531 (O_1531,N_29556,N_28013);
or UO_1532 (O_1532,N_28667,N_29968);
or UO_1533 (O_1533,N_29743,N_29484);
or UO_1534 (O_1534,N_29730,N_28539);
and UO_1535 (O_1535,N_28867,N_28710);
xor UO_1536 (O_1536,N_29044,N_29734);
nand UO_1537 (O_1537,N_29795,N_28989);
xor UO_1538 (O_1538,N_29031,N_29471);
or UO_1539 (O_1539,N_29496,N_28542);
nand UO_1540 (O_1540,N_28638,N_28434);
and UO_1541 (O_1541,N_29266,N_29406);
and UO_1542 (O_1542,N_29582,N_28714);
nor UO_1543 (O_1543,N_28393,N_29283);
or UO_1544 (O_1544,N_29054,N_28116);
or UO_1545 (O_1545,N_28954,N_29960);
nor UO_1546 (O_1546,N_29099,N_29258);
nor UO_1547 (O_1547,N_28381,N_29391);
or UO_1548 (O_1548,N_28917,N_29100);
or UO_1549 (O_1549,N_29832,N_28818);
and UO_1550 (O_1550,N_28413,N_29300);
nor UO_1551 (O_1551,N_29846,N_28088);
or UO_1552 (O_1552,N_28942,N_28971);
and UO_1553 (O_1553,N_29351,N_28963);
nor UO_1554 (O_1554,N_29041,N_28271);
nand UO_1555 (O_1555,N_29159,N_28736);
xor UO_1556 (O_1556,N_28944,N_29791);
or UO_1557 (O_1557,N_28515,N_29734);
nand UO_1558 (O_1558,N_29477,N_28159);
nor UO_1559 (O_1559,N_29745,N_29432);
and UO_1560 (O_1560,N_29125,N_29012);
xor UO_1561 (O_1561,N_28819,N_29045);
nor UO_1562 (O_1562,N_28726,N_28529);
nand UO_1563 (O_1563,N_28119,N_28260);
nand UO_1564 (O_1564,N_28294,N_29917);
nand UO_1565 (O_1565,N_28299,N_29918);
xor UO_1566 (O_1566,N_29845,N_29380);
xor UO_1567 (O_1567,N_28330,N_29988);
and UO_1568 (O_1568,N_28176,N_28910);
or UO_1569 (O_1569,N_28117,N_28280);
or UO_1570 (O_1570,N_28448,N_28307);
and UO_1571 (O_1571,N_28359,N_28981);
nor UO_1572 (O_1572,N_28008,N_29096);
or UO_1573 (O_1573,N_29425,N_28296);
and UO_1574 (O_1574,N_29627,N_28605);
xnor UO_1575 (O_1575,N_28227,N_28632);
or UO_1576 (O_1576,N_28314,N_28870);
nand UO_1577 (O_1577,N_29357,N_28110);
xor UO_1578 (O_1578,N_29072,N_29161);
nand UO_1579 (O_1579,N_29896,N_28622);
xor UO_1580 (O_1580,N_29975,N_29063);
nor UO_1581 (O_1581,N_28415,N_29075);
nor UO_1582 (O_1582,N_29631,N_28105);
nand UO_1583 (O_1583,N_28287,N_29544);
or UO_1584 (O_1584,N_28849,N_28210);
xor UO_1585 (O_1585,N_28728,N_29072);
or UO_1586 (O_1586,N_28504,N_28795);
nand UO_1587 (O_1587,N_28486,N_28833);
nand UO_1588 (O_1588,N_28541,N_29405);
or UO_1589 (O_1589,N_28027,N_28072);
or UO_1590 (O_1590,N_29851,N_28141);
xor UO_1591 (O_1591,N_28025,N_28571);
nor UO_1592 (O_1592,N_29058,N_29901);
nand UO_1593 (O_1593,N_29367,N_28497);
or UO_1594 (O_1594,N_28559,N_29538);
nor UO_1595 (O_1595,N_28801,N_29440);
xor UO_1596 (O_1596,N_28816,N_28964);
nor UO_1597 (O_1597,N_28312,N_28189);
nor UO_1598 (O_1598,N_28984,N_29120);
and UO_1599 (O_1599,N_29579,N_28684);
or UO_1600 (O_1600,N_28286,N_28004);
and UO_1601 (O_1601,N_28896,N_28886);
and UO_1602 (O_1602,N_28254,N_29279);
nor UO_1603 (O_1603,N_29547,N_28241);
nor UO_1604 (O_1604,N_28839,N_28628);
and UO_1605 (O_1605,N_29717,N_29934);
nor UO_1606 (O_1606,N_29374,N_29314);
xnor UO_1607 (O_1607,N_28437,N_28839);
or UO_1608 (O_1608,N_29119,N_28199);
or UO_1609 (O_1609,N_28773,N_28750);
and UO_1610 (O_1610,N_29558,N_28134);
or UO_1611 (O_1611,N_28721,N_28266);
xor UO_1612 (O_1612,N_28729,N_28320);
xor UO_1613 (O_1613,N_29291,N_28140);
nand UO_1614 (O_1614,N_29284,N_28337);
or UO_1615 (O_1615,N_29337,N_28773);
nand UO_1616 (O_1616,N_29320,N_28652);
or UO_1617 (O_1617,N_28155,N_28783);
nor UO_1618 (O_1618,N_28307,N_28941);
xnor UO_1619 (O_1619,N_28293,N_28304);
nor UO_1620 (O_1620,N_28468,N_29178);
and UO_1621 (O_1621,N_29097,N_29020);
xnor UO_1622 (O_1622,N_28281,N_28317);
and UO_1623 (O_1623,N_28420,N_29319);
nand UO_1624 (O_1624,N_29203,N_28701);
or UO_1625 (O_1625,N_29868,N_29381);
nor UO_1626 (O_1626,N_29603,N_28432);
and UO_1627 (O_1627,N_29097,N_28996);
and UO_1628 (O_1628,N_29361,N_29306);
or UO_1629 (O_1629,N_28646,N_29870);
or UO_1630 (O_1630,N_29154,N_28934);
xor UO_1631 (O_1631,N_29836,N_28675);
xnor UO_1632 (O_1632,N_28880,N_28363);
or UO_1633 (O_1633,N_29908,N_29225);
nand UO_1634 (O_1634,N_28473,N_28087);
xor UO_1635 (O_1635,N_29756,N_29030);
xnor UO_1636 (O_1636,N_29550,N_29961);
nand UO_1637 (O_1637,N_29805,N_28831);
nor UO_1638 (O_1638,N_29989,N_29029);
and UO_1639 (O_1639,N_28946,N_29830);
or UO_1640 (O_1640,N_28556,N_29494);
nand UO_1641 (O_1641,N_29342,N_29967);
nor UO_1642 (O_1642,N_28180,N_28291);
and UO_1643 (O_1643,N_28121,N_29828);
xnor UO_1644 (O_1644,N_28329,N_28432);
or UO_1645 (O_1645,N_28771,N_28474);
nand UO_1646 (O_1646,N_28328,N_28180);
nor UO_1647 (O_1647,N_29766,N_28741);
nand UO_1648 (O_1648,N_29441,N_29206);
nand UO_1649 (O_1649,N_28167,N_28717);
nor UO_1650 (O_1650,N_28054,N_28567);
nand UO_1651 (O_1651,N_29401,N_28424);
nor UO_1652 (O_1652,N_29144,N_28656);
nor UO_1653 (O_1653,N_29778,N_29122);
and UO_1654 (O_1654,N_29162,N_29632);
or UO_1655 (O_1655,N_29684,N_29035);
xnor UO_1656 (O_1656,N_28265,N_28043);
nand UO_1657 (O_1657,N_29265,N_29567);
nand UO_1658 (O_1658,N_29653,N_28278);
nor UO_1659 (O_1659,N_28101,N_29856);
or UO_1660 (O_1660,N_28486,N_29532);
xor UO_1661 (O_1661,N_28317,N_29586);
xnor UO_1662 (O_1662,N_29021,N_28230);
xor UO_1663 (O_1663,N_29786,N_28468);
or UO_1664 (O_1664,N_28341,N_29590);
nor UO_1665 (O_1665,N_29605,N_28161);
nor UO_1666 (O_1666,N_28187,N_28389);
xnor UO_1667 (O_1667,N_29288,N_29357);
xor UO_1668 (O_1668,N_28621,N_29747);
or UO_1669 (O_1669,N_28485,N_29204);
xor UO_1670 (O_1670,N_28604,N_28577);
nand UO_1671 (O_1671,N_28270,N_29790);
nor UO_1672 (O_1672,N_29398,N_29351);
and UO_1673 (O_1673,N_29737,N_28207);
xor UO_1674 (O_1674,N_29087,N_29968);
xor UO_1675 (O_1675,N_28809,N_29605);
and UO_1676 (O_1676,N_29459,N_29538);
nand UO_1677 (O_1677,N_28652,N_29392);
and UO_1678 (O_1678,N_28022,N_29365);
xnor UO_1679 (O_1679,N_29880,N_28950);
and UO_1680 (O_1680,N_28392,N_28604);
or UO_1681 (O_1681,N_29556,N_29656);
and UO_1682 (O_1682,N_29340,N_28698);
nor UO_1683 (O_1683,N_29079,N_28517);
nor UO_1684 (O_1684,N_29024,N_28431);
or UO_1685 (O_1685,N_29495,N_28055);
and UO_1686 (O_1686,N_29183,N_28492);
or UO_1687 (O_1687,N_28599,N_28724);
or UO_1688 (O_1688,N_29568,N_28983);
nor UO_1689 (O_1689,N_29150,N_29800);
xor UO_1690 (O_1690,N_29993,N_29177);
or UO_1691 (O_1691,N_28306,N_29613);
nand UO_1692 (O_1692,N_28072,N_29708);
xnor UO_1693 (O_1693,N_28258,N_29031);
nor UO_1694 (O_1694,N_28162,N_29539);
nor UO_1695 (O_1695,N_29139,N_28357);
nor UO_1696 (O_1696,N_28641,N_28049);
nand UO_1697 (O_1697,N_29871,N_29296);
and UO_1698 (O_1698,N_28893,N_28756);
and UO_1699 (O_1699,N_28979,N_29365);
or UO_1700 (O_1700,N_28414,N_29447);
nor UO_1701 (O_1701,N_28890,N_29268);
xor UO_1702 (O_1702,N_28343,N_29286);
xnor UO_1703 (O_1703,N_29332,N_29184);
nand UO_1704 (O_1704,N_28345,N_28678);
and UO_1705 (O_1705,N_28519,N_28556);
and UO_1706 (O_1706,N_28984,N_29197);
nor UO_1707 (O_1707,N_29033,N_29345);
xor UO_1708 (O_1708,N_28637,N_28073);
nor UO_1709 (O_1709,N_28767,N_28193);
nor UO_1710 (O_1710,N_28068,N_29387);
or UO_1711 (O_1711,N_29787,N_29972);
nor UO_1712 (O_1712,N_29588,N_29570);
nand UO_1713 (O_1713,N_28886,N_29150);
nor UO_1714 (O_1714,N_29432,N_29545);
or UO_1715 (O_1715,N_29561,N_29694);
and UO_1716 (O_1716,N_29728,N_29815);
nor UO_1717 (O_1717,N_28016,N_28646);
nor UO_1718 (O_1718,N_28648,N_29292);
xor UO_1719 (O_1719,N_28465,N_29376);
xor UO_1720 (O_1720,N_29167,N_29324);
and UO_1721 (O_1721,N_28583,N_28751);
xor UO_1722 (O_1722,N_28644,N_29173);
or UO_1723 (O_1723,N_29116,N_28598);
xnor UO_1724 (O_1724,N_28479,N_28628);
xor UO_1725 (O_1725,N_28562,N_28040);
nand UO_1726 (O_1726,N_29380,N_29735);
and UO_1727 (O_1727,N_29194,N_29058);
or UO_1728 (O_1728,N_29159,N_28832);
nand UO_1729 (O_1729,N_29057,N_28363);
or UO_1730 (O_1730,N_29821,N_29525);
nand UO_1731 (O_1731,N_28704,N_28411);
and UO_1732 (O_1732,N_28977,N_29362);
xor UO_1733 (O_1733,N_28631,N_28663);
nand UO_1734 (O_1734,N_29425,N_28523);
nand UO_1735 (O_1735,N_29202,N_28493);
nand UO_1736 (O_1736,N_29495,N_29757);
xnor UO_1737 (O_1737,N_28017,N_29473);
nor UO_1738 (O_1738,N_29251,N_28143);
xor UO_1739 (O_1739,N_28743,N_28074);
or UO_1740 (O_1740,N_29112,N_28393);
nor UO_1741 (O_1741,N_29394,N_29435);
or UO_1742 (O_1742,N_29090,N_29250);
or UO_1743 (O_1743,N_29820,N_29029);
and UO_1744 (O_1744,N_29513,N_28269);
or UO_1745 (O_1745,N_28696,N_28943);
xnor UO_1746 (O_1746,N_28312,N_28815);
nand UO_1747 (O_1747,N_28418,N_29054);
and UO_1748 (O_1748,N_28867,N_28209);
or UO_1749 (O_1749,N_28152,N_28715);
or UO_1750 (O_1750,N_29218,N_29902);
nand UO_1751 (O_1751,N_29106,N_29985);
nor UO_1752 (O_1752,N_28691,N_29040);
nor UO_1753 (O_1753,N_29185,N_28707);
xor UO_1754 (O_1754,N_29717,N_28890);
xnor UO_1755 (O_1755,N_28531,N_28608);
or UO_1756 (O_1756,N_28129,N_29747);
nand UO_1757 (O_1757,N_28891,N_28756);
nand UO_1758 (O_1758,N_28951,N_28465);
nand UO_1759 (O_1759,N_29289,N_28167);
xor UO_1760 (O_1760,N_28823,N_28960);
and UO_1761 (O_1761,N_28722,N_28831);
xnor UO_1762 (O_1762,N_29086,N_29880);
and UO_1763 (O_1763,N_29606,N_29896);
or UO_1764 (O_1764,N_29437,N_29228);
or UO_1765 (O_1765,N_28062,N_28725);
nor UO_1766 (O_1766,N_29700,N_29016);
or UO_1767 (O_1767,N_28067,N_28727);
and UO_1768 (O_1768,N_28586,N_29934);
nand UO_1769 (O_1769,N_29161,N_28881);
or UO_1770 (O_1770,N_28327,N_28381);
nand UO_1771 (O_1771,N_29398,N_29453);
nand UO_1772 (O_1772,N_29552,N_29033);
and UO_1773 (O_1773,N_29240,N_29250);
and UO_1774 (O_1774,N_28243,N_28755);
and UO_1775 (O_1775,N_28637,N_28511);
xor UO_1776 (O_1776,N_28939,N_29285);
xor UO_1777 (O_1777,N_28875,N_29296);
nor UO_1778 (O_1778,N_29925,N_29118);
xnor UO_1779 (O_1779,N_28281,N_28394);
xor UO_1780 (O_1780,N_29486,N_29854);
and UO_1781 (O_1781,N_29298,N_29078);
nand UO_1782 (O_1782,N_28539,N_29868);
nand UO_1783 (O_1783,N_28531,N_28248);
nor UO_1784 (O_1784,N_29564,N_28775);
and UO_1785 (O_1785,N_28704,N_29762);
and UO_1786 (O_1786,N_28850,N_29754);
and UO_1787 (O_1787,N_28869,N_28594);
nor UO_1788 (O_1788,N_29419,N_28520);
nand UO_1789 (O_1789,N_28016,N_29279);
xor UO_1790 (O_1790,N_29700,N_29302);
or UO_1791 (O_1791,N_29389,N_29907);
and UO_1792 (O_1792,N_28272,N_28955);
and UO_1793 (O_1793,N_28288,N_28195);
and UO_1794 (O_1794,N_28529,N_29090);
nand UO_1795 (O_1795,N_29665,N_28166);
xor UO_1796 (O_1796,N_29223,N_29718);
xor UO_1797 (O_1797,N_29874,N_29212);
xnor UO_1798 (O_1798,N_29480,N_29585);
xor UO_1799 (O_1799,N_28215,N_29755);
nor UO_1800 (O_1800,N_28786,N_28980);
and UO_1801 (O_1801,N_28085,N_29643);
nand UO_1802 (O_1802,N_28595,N_28500);
and UO_1803 (O_1803,N_28290,N_29547);
and UO_1804 (O_1804,N_28836,N_29564);
nand UO_1805 (O_1805,N_29701,N_28058);
xor UO_1806 (O_1806,N_28339,N_28983);
or UO_1807 (O_1807,N_29786,N_29340);
nor UO_1808 (O_1808,N_28129,N_29011);
nand UO_1809 (O_1809,N_29549,N_28914);
xnor UO_1810 (O_1810,N_28129,N_29408);
and UO_1811 (O_1811,N_29686,N_29803);
nand UO_1812 (O_1812,N_28678,N_29370);
nor UO_1813 (O_1813,N_29567,N_28455);
xor UO_1814 (O_1814,N_28420,N_28649);
xor UO_1815 (O_1815,N_29347,N_29941);
nand UO_1816 (O_1816,N_29038,N_28443);
and UO_1817 (O_1817,N_29548,N_29024);
and UO_1818 (O_1818,N_28901,N_29267);
or UO_1819 (O_1819,N_29285,N_29396);
nand UO_1820 (O_1820,N_29088,N_29276);
xor UO_1821 (O_1821,N_29538,N_29976);
nor UO_1822 (O_1822,N_29109,N_29200);
nor UO_1823 (O_1823,N_29823,N_29725);
xor UO_1824 (O_1824,N_28432,N_29767);
xor UO_1825 (O_1825,N_28803,N_28269);
and UO_1826 (O_1826,N_29652,N_29179);
and UO_1827 (O_1827,N_29019,N_29469);
nand UO_1828 (O_1828,N_28824,N_28393);
or UO_1829 (O_1829,N_29392,N_29990);
and UO_1830 (O_1830,N_29063,N_29820);
or UO_1831 (O_1831,N_28950,N_29482);
or UO_1832 (O_1832,N_28676,N_29156);
nand UO_1833 (O_1833,N_29492,N_29068);
or UO_1834 (O_1834,N_29840,N_28186);
or UO_1835 (O_1835,N_28873,N_29326);
nand UO_1836 (O_1836,N_28478,N_28873);
and UO_1837 (O_1837,N_28980,N_29621);
or UO_1838 (O_1838,N_28652,N_28601);
nand UO_1839 (O_1839,N_29136,N_29375);
and UO_1840 (O_1840,N_28464,N_29100);
and UO_1841 (O_1841,N_29090,N_28806);
xnor UO_1842 (O_1842,N_28051,N_29580);
nand UO_1843 (O_1843,N_28388,N_28733);
or UO_1844 (O_1844,N_29574,N_29217);
or UO_1845 (O_1845,N_29876,N_28258);
nor UO_1846 (O_1846,N_28204,N_29036);
and UO_1847 (O_1847,N_28824,N_29554);
or UO_1848 (O_1848,N_28623,N_29907);
xor UO_1849 (O_1849,N_29922,N_29544);
or UO_1850 (O_1850,N_28315,N_29374);
and UO_1851 (O_1851,N_29814,N_28448);
and UO_1852 (O_1852,N_28895,N_28410);
or UO_1853 (O_1853,N_29685,N_29053);
nand UO_1854 (O_1854,N_28612,N_29644);
and UO_1855 (O_1855,N_29583,N_28055);
nand UO_1856 (O_1856,N_28957,N_28431);
nand UO_1857 (O_1857,N_28988,N_28068);
and UO_1858 (O_1858,N_28980,N_28755);
nand UO_1859 (O_1859,N_28164,N_29636);
nand UO_1860 (O_1860,N_28737,N_29714);
xnor UO_1861 (O_1861,N_28989,N_28304);
nor UO_1862 (O_1862,N_29424,N_28196);
xnor UO_1863 (O_1863,N_28554,N_29262);
nor UO_1864 (O_1864,N_29587,N_29475);
and UO_1865 (O_1865,N_29338,N_28268);
nand UO_1866 (O_1866,N_29018,N_28420);
nor UO_1867 (O_1867,N_29819,N_28694);
xnor UO_1868 (O_1868,N_28825,N_28396);
xnor UO_1869 (O_1869,N_29161,N_29020);
or UO_1870 (O_1870,N_28166,N_29198);
or UO_1871 (O_1871,N_29859,N_29278);
xnor UO_1872 (O_1872,N_29230,N_28205);
or UO_1873 (O_1873,N_28665,N_29907);
or UO_1874 (O_1874,N_29845,N_28698);
and UO_1875 (O_1875,N_29335,N_29176);
or UO_1876 (O_1876,N_29065,N_28607);
or UO_1877 (O_1877,N_28461,N_29400);
xnor UO_1878 (O_1878,N_29766,N_28876);
nor UO_1879 (O_1879,N_29667,N_28981);
and UO_1880 (O_1880,N_28189,N_28536);
nand UO_1881 (O_1881,N_28643,N_28326);
and UO_1882 (O_1882,N_29091,N_28426);
nor UO_1883 (O_1883,N_28921,N_28215);
and UO_1884 (O_1884,N_28976,N_29682);
and UO_1885 (O_1885,N_29407,N_29827);
nor UO_1886 (O_1886,N_28155,N_28690);
or UO_1887 (O_1887,N_28190,N_28069);
nor UO_1888 (O_1888,N_28362,N_29204);
nand UO_1889 (O_1889,N_28733,N_29492);
nor UO_1890 (O_1890,N_28336,N_28765);
and UO_1891 (O_1891,N_29286,N_29184);
nand UO_1892 (O_1892,N_29249,N_29593);
nor UO_1893 (O_1893,N_29086,N_28614);
or UO_1894 (O_1894,N_29480,N_29331);
xor UO_1895 (O_1895,N_29332,N_29250);
and UO_1896 (O_1896,N_28884,N_28637);
nor UO_1897 (O_1897,N_29313,N_29514);
or UO_1898 (O_1898,N_28355,N_29739);
nor UO_1899 (O_1899,N_28167,N_28175);
or UO_1900 (O_1900,N_29774,N_29023);
and UO_1901 (O_1901,N_28539,N_28336);
and UO_1902 (O_1902,N_28762,N_29206);
nand UO_1903 (O_1903,N_29853,N_28665);
nand UO_1904 (O_1904,N_29621,N_28209);
nor UO_1905 (O_1905,N_29995,N_29694);
xor UO_1906 (O_1906,N_29531,N_28101);
nor UO_1907 (O_1907,N_28949,N_28115);
and UO_1908 (O_1908,N_28902,N_29753);
and UO_1909 (O_1909,N_28643,N_29931);
or UO_1910 (O_1910,N_29182,N_29436);
nor UO_1911 (O_1911,N_29767,N_29330);
xor UO_1912 (O_1912,N_28497,N_29728);
nand UO_1913 (O_1913,N_28457,N_28451);
and UO_1914 (O_1914,N_28391,N_29261);
xor UO_1915 (O_1915,N_28194,N_28921);
nor UO_1916 (O_1916,N_28090,N_28996);
and UO_1917 (O_1917,N_29992,N_28225);
and UO_1918 (O_1918,N_29830,N_28642);
nor UO_1919 (O_1919,N_29930,N_29552);
nor UO_1920 (O_1920,N_29662,N_28367);
nor UO_1921 (O_1921,N_28931,N_29565);
nand UO_1922 (O_1922,N_29428,N_29946);
and UO_1923 (O_1923,N_28664,N_29514);
or UO_1924 (O_1924,N_29483,N_29348);
xnor UO_1925 (O_1925,N_29685,N_29468);
or UO_1926 (O_1926,N_28525,N_28111);
nand UO_1927 (O_1927,N_28535,N_28855);
and UO_1928 (O_1928,N_28950,N_28303);
and UO_1929 (O_1929,N_29829,N_29435);
nor UO_1930 (O_1930,N_29992,N_29729);
xnor UO_1931 (O_1931,N_28179,N_29349);
and UO_1932 (O_1932,N_28241,N_28543);
or UO_1933 (O_1933,N_28375,N_28351);
nor UO_1934 (O_1934,N_29321,N_28143);
nand UO_1935 (O_1935,N_28100,N_29697);
and UO_1936 (O_1936,N_28410,N_29434);
and UO_1937 (O_1937,N_28712,N_28893);
nand UO_1938 (O_1938,N_29308,N_28432);
or UO_1939 (O_1939,N_29264,N_29906);
nor UO_1940 (O_1940,N_29899,N_28440);
xnor UO_1941 (O_1941,N_28553,N_28173);
or UO_1942 (O_1942,N_29057,N_29188);
and UO_1943 (O_1943,N_29143,N_28769);
xnor UO_1944 (O_1944,N_29572,N_29361);
nand UO_1945 (O_1945,N_28281,N_28425);
or UO_1946 (O_1946,N_29904,N_29017);
or UO_1947 (O_1947,N_28482,N_28802);
nor UO_1948 (O_1948,N_29612,N_29732);
xor UO_1949 (O_1949,N_28633,N_29024);
or UO_1950 (O_1950,N_29161,N_28275);
nor UO_1951 (O_1951,N_29598,N_29722);
xnor UO_1952 (O_1952,N_28135,N_28849);
nor UO_1953 (O_1953,N_28772,N_28262);
or UO_1954 (O_1954,N_29287,N_29331);
or UO_1955 (O_1955,N_28810,N_28740);
and UO_1956 (O_1956,N_28962,N_29372);
and UO_1957 (O_1957,N_28194,N_28089);
and UO_1958 (O_1958,N_29285,N_29204);
and UO_1959 (O_1959,N_28031,N_29332);
nor UO_1960 (O_1960,N_29277,N_29712);
nand UO_1961 (O_1961,N_29352,N_28725);
nor UO_1962 (O_1962,N_29233,N_28556);
nor UO_1963 (O_1963,N_29821,N_28881);
or UO_1964 (O_1964,N_29607,N_29156);
and UO_1965 (O_1965,N_28383,N_28024);
xnor UO_1966 (O_1966,N_28001,N_29046);
nor UO_1967 (O_1967,N_28278,N_28791);
and UO_1968 (O_1968,N_28538,N_28717);
or UO_1969 (O_1969,N_28507,N_29866);
nand UO_1970 (O_1970,N_28053,N_29113);
and UO_1971 (O_1971,N_28123,N_29208);
xor UO_1972 (O_1972,N_28613,N_28344);
or UO_1973 (O_1973,N_29932,N_28864);
or UO_1974 (O_1974,N_28773,N_28244);
xor UO_1975 (O_1975,N_29446,N_28621);
and UO_1976 (O_1976,N_29740,N_29340);
and UO_1977 (O_1977,N_29071,N_29637);
xnor UO_1978 (O_1978,N_28158,N_29798);
xor UO_1979 (O_1979,N_29403,N_29047);
xor UO_1980 (O_1980,N_29685,N_29658);
nand UO_1981 (O_1981,N_28961,N_29330);
nor UO_1982 (O_1982,N_28301,N_28238);
xnor UO_1983 (O_1983,N_29950,N_29792);
and UO_1984 (O_1984,N_29845,N_29324);
nand UO_1985 (O_1985,N_28645,N_29490);
nand UO_1986 (O_1986,N_28505,N_28063);
xnor UO_1987 (O_1987,N_29892,N_28652);
nor UO_1988 (O_1988,N_28775,N_28589);
xnor UO_1989 (O_1989,N_28161,N_28254);
xnor UO_1990 (O_1990,N_29446,N_28185);
nand UO_1991 (O_1991,N_28341,N_29003);
or UO_1992 (O_1992,N_28143,N_29182);
nand UO_1993 (O_1993,N_28434,N_28760);
xor UO_1994 (O_1994,N_28068,N_28076);
nor UO_1995 (O_1995,N_28140,N_28243);
xor UO_1996 (O_1996,N_29859,N_28768);
or UO_1997 (O_1997,N_28477,N_29273);
and UO_1998 (O_1998,N_29418,N_28692);
or UO_1999 (O_1999,N_29705,N_29731);
xor UO_2000 (O_2000,N_29970,N_28005);
nor UO_2001 (O_2001,N_28311,N_29217);
nor UO_2002 (O_2002,N_28948,N_28388);
nand UO_2003 (O_2003,N_28971,N_29948);
nand UO_2004 (O_2004,N_29567,N_29209);
xnor UO_2005 (O_2005,N_28453,N_29906);
nor UO_2006 (O_2006,N_29496,N_28267);
nand UO_2007 (O_2007,N_28460,N_28909);
nand UO_2008 (O_2008,N_28898,N_29315);
nand UO_2009 (O_2009,N_29654,N_28283);
or UO_2010 (O_2010,N_28412,N_28394);
xor UO_2011 (O_2011,N_28035,N_29467);
nand UO_2012 (O_2012,N_28358,N_28730);
and UO_2013 (O_2013,N_28058,N_29773);
xnor UO_2014 (O_2014,N_28183,N_29625);
nand UO_2015 (O_2015,N_29459,N_28694);
nand UO_2016 (O_2016,N_28159,N_29347);
nor UO_2017 (O_2017,N_29885,N_28856);
nand UO_2018 (O_2018,N_28617,N_29724);
nor UO_2019 (O_2019,N_28751,N_29612);
and UO_2020 (O_2020,N_29212,N_28769);
or UO_2021 (O_2021,N_29829,N_28158);
or UO_2022 (O_2022,N_29924,N_29927);
nand UO_2023 (O_2023,N_28127,N_29833);
nand UO_2024 (O_2024,N_28481,N_29471);
and UO_2025 (O_2025,N_28941,N_29461);
and UO_2026 (O_2026,N_28873,N_28706);
nand UO_2027 (O_2027,N_29348,N_29195);
nor UO_2028 (O_2028,N_28999,N_28496);
xor UO_2029 (O_2029,N_28009,N_28492);
nand UO_2030 (O_2030,N_29456,N_29914);
nand UO_2031 (O_2031,N_28397,N_29359);
xnor UO_2032 (O_2032,N_28037,N_28828);
nor UO_2033 (O_2033,N_29107,N_28342);
nor UO_2034 (O_2034,N_29935,N_29838);
nor UO_2035 (O_2035,N_28228,N_28730);
nand UO_2036 (O_2036,N_29876,N_29163);
nand UO_2037 (O_2037,N_29593,N_28264);
or UO_2038 (O_2038,N_29566,N_29065);
nand UO_2039 (O_2039,N_28843,N_29372);
nand UO_2040 (O_2040,N_29670,N_29277);
or UO_2041 (O_2041,N_29549,N_28200);
nand UO_2042 (O_2042,N_28025,N_29645);
nor UO_2043 (O_2043,N_28939,N_28643);
and UO_2044 (O_2044,N_29351,N_28115);
or UO_2045 (O_2045,N_28128,N_29798);
nor UO_2046 (O_2046,N_28137,N_28201);
xnor UO_2047 (O_2047,N_28468,N_28024);
and UO_2048 (O_2048,N_29209,N_29829);
nand UO_2049 (O_2049,N_29346,N_29839);
xor UO_2050 (O_2050,N_28732,N_29573);
nand UO_2051 (O_2051,N_29480,N_29112);
and UO_2052 (O_2052,N_29333,N_28684);
and UO_2053 (O_2053,N_29522,N_28826);
xor UO_2054 (O_2054,N_29638,N_28781);
xnor UO_2055 (O_2055,N_29879,N_29973);
or UO_2056 (O_2056,N_28612,N_29910);
or UO_2057 (O_2057,N_28187,N_28825);
xor UO_2058 (O_2058,N_28203,N_28722);
nor UO_2059 (O_2059,N_28425,N_28535);
or UO_2060 (O_2060,N_29388,N_29096);
xnor UO_2061 (O_2061,N_29121,N_29365);
nand UO_2062 (O_2062,N_29574,N_29378);
or UO_2063 (O_2063,N_28382,N_29990);
nand UO_2064 (O_2064,N_28418,N_29494);
xnor UO_2065 (O_2065,N_29640,N_29311);
nand UO_2066 (O_2066,N_28999,N_29949);
xnor UO_2067 (O_2067,N_28527,N_28050);
nand UO_2068 (O_2068,N_29385,N_28285);
xnor UO_2069 (O_2069,N_28957,N_28718);
or UO_2070 (O_2070,N_28483,N_29844);
or UO_2071 (O_2071,N_28554,N_29327);
nor UO_2072 (O_2072,N_28203,N_28261);
or UO_2073 (O_2073,N_28045,N_28729);
xor UO_2074 (O_2074,N_29735,N_28351);
nor UO_2075 (O_2075,N_28575,N_29821);
xor UO_2076 (O_2076,N_29922,N_28264);
or UO_2077 (O_2077,N_29014,N_29028);
and UO_2078 (O_2078,N_28946,N_28065);
xor UO_2079 (O_2079,N_28245,N_29380);
and UO_2080 (O_2080,N_28597,N_29197);
nor UO_2081 (O_2081,N_29875,N_28838);
or UO_2082 (O_2082,N_29061,N_28341);
nor UO_2083 (O_2083,N_29225,N_28917);
nand UO_2084 (O_2084,N_29780,N_29444);
xnor UO_2085 (O_2085,N_29332,N_28302);
xnor UO_2086 (O_2086,N_28940,N_29908);
nor UO_2087 (O_2087,N_29785,N_29583);
nand UO_2088 (O_2088,N_28030,N_28359);
or UO_2089 (O_2089,N_29875,N_29975);
or UO_2090 (O_2090,N_28052,N_29171);
and UO_2091 (O_2091,N_28075,N_29825);
nand UO_2092 (O_2092,N_29966,N_29424);
nand UO_2093 (O_2093,N_29950,N_29673);
xnor UO_2094 (O_2094,N_29751,N_28694);
nor UO_2095 (O_2095,N_28395,N_29791);
xor UO_2096 (O_2096,N_29486,N_28319);
and UO_2097 (O_2097,N_28357,N_29886);
or UO_2098 (O_2098,N_28969,N_29152);
nand UO_2099 (O_2099,N_28298,N_29550);
nand UO_2100 (O_2100,N_28071,N_29413);
nand UO_2101 (O_2101,N_29742,N_28255);
nand UO_2102 (O_2102,N_28457,N_28770);
nand UO_2103 (O_2103,N_28484,N_29039);
xnor UO_2104 (O_2104,N_28819,N_29896);
or UO_2105 (O_2105,N_29311,N_28110);
xor UO_2106 (O_2106,N_28621,N_28443);
or UO_2107 (O_2107,N_28367,N_28208);
nor UO_2108 (O_2108,N_29928,N_28975);
nand UO_2109 (O_2109,N_29637,N_28963);
nand UO_2110 (O_2110,N_29894,N_28874);
nor UO_2111 (O_2111,N_28534,N_29051);
xor UO_2112 (O_2112,N_29694,N_28406);
nor UO_2113 (O_2113,N_29426,N_28540);
xor UO_2114 (O_2114,N_28796,N_28849);
or UO_2115 (O_2115,N_29350,N_28594);
nand UO_2116 (O_2116,N_29621,N_29359);
xnor UO_2117 (O_2117,N_28590,N_28759);
xor UO_2118 (O_2118,N_28466,N_29839);
nand UO_2119 (O_2119,N_29231,N_29185);
xnor UO_2120 (O_2120,N_29362,N_29116);
xnor UO_2121 (O_2121,N_28079,N_28689);
xnor UO_2122 (O_2122,N_29821,N_28282);
or UO_2123 (O_2123,N_29955,N_28714);
nand UO_2124 (O_2124,N_28137,N_29698);
and UO_2125 (O_2125,N_28187,N_29034);
or UO_2126 (O_2126,N_28535,N_28789);
or UO_2127 (O_2127,N_28169,N_28243);
nor UO_2128 (O_2128,N_29856,N_29534);
xor UO_2129 (O_2129,N_29925,N_28567);
or UO_2130 (O_2130,N_28020,N_28804);
nand UO_2131 (O_2131,N_29837,N_28336);
nor UO_2132 (O_2132,N_28766,N_28376);
or UO_2133 (O_2133,N_28097,N_29139);
nand UO_2134 (O_2134,N_28648,N_29843);
xnor UO_2135 (O_2135,N_28492,N_28577);
xnor UO_2136 (O_2136,N_28866,N_29124);
nand UO_2137 (O_2137,N_28212,N_29959);
and UO_2138 (O_2138,N_28703,N_28068);
nor UO_2139 (O_2139,N_29391,N_28749);
nor UO_2140 (O_2140,N_29131,N_29604);
xnor UO_2141 (O_2141,N_28817,N_28922);
and UO_2142 (O_2142,N_29743,N_29110);
or UO_2143 (O_2143,N_29685,N_29379);
xor UO_2144 (O_2144,N_28216,N_29946);
xnor UO_2145 (O_2145,N_29209,N_28991);
nand UO_2146 (O_2146,N_29543,N_28269);
nor UO_2147 (O_2147,N_29176,N_28025);
and UO_2148 (O_2148,N_28466,N_29344);
nand UO_2149 (O_2149,N_28798,N_28729);
or UO_2150 (O_2150,N_28330,N_28018);
xor UO_2151 (O_2151,N_28083,N_29830);
nand UO_2152 (O_2152,N_28782,N_29946);
and UO_2153 (O_2153,N_28146,N_28507);
nand UO_2154 (O_2154,N_28335,N_29715);
nand UO_2155 (O_2155,N_28479,N_29534);
nand UO_2156 (O_2156,N_29890,N_28472);
and UO_2157 (O_2157,N_29875,N_28128);
or UO_2158 (O_2158,N_28250,N_28105);
xor UO_2159 (O_2159,N_29220,N_28257);
and UO_2160 (O_2160,N_28639,N_28267);
xnor UO_2161 (O_2161,N_28706,N_29816);
or UO_2162 (O_2162,N_29431,N_28798);
and UO_2163 (O_2163,N_29766,N_29258);
or UO_2164 (O_2164,N_29380,N_29922);
nand UO_2165 (O_2165,N_28771,N_29640);
or UO_2166 (O_2166,N_28326,N_29749);
nand UO_2167 (O_2167,N_29594,N_29445);
or UO_2168 (O_2168,N_29483,N_29304);
nor UO_2169 (O_2169,N_28331,N_28297);
nand UO_2170 (O_2170,N_28860,N_28032);
nand UO_2171 (O_2171,N_29844,N_28620);
xnor UO_2172 (O_2172,N_28191,N_29081);
or UO_2173 (O_2173,N_29235,N_28002);
xnor UO_2174 (O_2174,N_28829,N_29037);
and UO_2175 (O_2175,N_28300,N_29964);
or UO_2176 (O_2176,N_29074,N_29888);
nor UO_2177 (O_2177,N_28803,N_29011);
xnor UO_2178 (O_2178,N_28981,N_29020);
nand UO_2179 (O_2179,N_29586,N_28744);
and UO_2180 (O_2180,N_29571,N_29548);
xnor UO_2181 (O_2181,N_28363,N_28641);
or UO_2182 (O_2182,N_28887,N_28242);
nand UO_2183 (O_2183,N_29094,N_28825);
or UO_2184 (O_2184,N_28973,N_28145);
nor UO_2185 (O_2185,N_28364,N_28232);
or UO_2186 (O_2186,N_29976,N_29511);
nor UO_2187 (O_2187,N_28192,N_28359);
nand UO_2188 (O_2188,N_28178,N_28984);
nand UO_2189 (O_2189,N_28468,N_29191);
nand UO_2190 (O_2190,N_29578,N_28928);
or UO_2191 (O_2191,N_29178,N_29602);
and UO_2192 (O_2192,N_29449,N_28139);
nand UO_2193 (O_2193,N_29203,N_28233);
xor UO_2194 (O_2194,N_28596,N_28265);
and UO_2195 (O_2195,N_29580,N_28428);
xnor UO_2196 (O_2196,N_29282,N_29724);
xnor UO_2197 (O_2197,N_28725,N_28839);
or UO_2198 (O_2198,N_28908,N_29722);
xor UO_2199 (O_2199,N_28472,N_28393);
nand UO_2200 (O_2200,N_29932,N_29588);
or UO_2201 (O_2201,N_29250,N_29972);
nor UO_2202 (O_2202,N_29364,N_28536);
xor UO_2203 (O_2203,N_28111,N_29070);
nor UO_2204 (O_2204,N_28187,N_29832);
or UO_2205 (O_2205,N_28435,N_29351);
and UO_2206 (O_2206,N_29494,N_29927);
xor UO_2207 (O_2207,N_29277,N_29118);
nand UO_2208 (O_2208,N_29729,N_29015);
nand UO_2209 (O_2209,N_29727,N_29380);
xor UO_2210 (O_2210,N_28167,N_29095);
and UO_2211 (O_2211,N_29611,N_29160);
nor UO_2212 (O_2212,N_29245,N_28391);
nor UO_2213 (O_2213,N_29428,N_29467);
or UO_2214 (O_2214,N_28560,N_29766);
nor UO_2215 (O_2215,N_29820,N_29892);
or UO_2216 (O_2216,N_29706,N_28368);
or UO_2217 (O_2217,N_28112,N_29759);
or UO_2218 (O_2218,N_29207,N_29790);
nand UO_2219 (O_2219,N_29276,N_29002);
or UO_2220 (O_2220,N_28032,N_28631);
and UO_2221 (O_2221,N_28933,N_29296);
nand UO_2222 (O_2222,N_28231,N_28009);
xor UO_2223 (O_2223,N_29755,N_28135);
or UO_2224 (O_2224,N_28223,N_29966);
and UO_2225 (O_2225,N_28621,N_28844);
nand UO_2226 (O_2226,N_29171,N_28372);
or UO_2227 (O_2227,N_29910,N_28678);
and UO_2228 (O_2228,N_29348,N_29696);
nor UO_2229 (O_2229,N_29392,N_29409);
nand UO_2230 (O_2230,N_29558,N_28054);
nand UO_2231 (O_2231,N_28974,N_28910);
and UO_2232 (O_2232,N_28514,N_29916);
nor UO_2233 (O_2233,N_29992,N_28710);
or UO_2234 (O_2234,N_29425,N_28847);
xnor UO_2235 (O_2235,N_29718,N_29481);
and UO_2236 (O_2236,N_29231,N_29563);
nor UO_2237 (O_2237,N_29995,N_28586);
or UO_2238 (O_2238,N_29217,N_28875);
and UO_2239 (O_2239,N_29425,N_28041);
or UO_2240 (O_2240,N_28175,N_28076);
and UO_2241 (O_2241,N_29211,N_28985);
and UO_2242 (O_2242,N_28678,N_28457);
or UO_2243 (O_2243,N_28407,N_29173);
and UO_2244 (O_2244,N_29416,N_29905);
nand UO_2245 (O_2245,N_29042,N_28757);
xnor UO_2246 (O_2246,N_28525,N_29965);
or UO_2247 (O_2247,N_29009,N_29926);
nor UO_2248 (O_2248,N_29807,N_28841);
xnor UO_2249 (O_2249,N_29766,N_29616);
and UO_2250 (O_2250,N_28055,N_29836);
xor UO_2251 (O_2251,N_29026,N_28857);
nand UO_2252 (O_2252,N_29000,N_29941);
nor UO_2253 (O_2253,N_29474,N_28459);
xor UO_2254 (O_2254,N_28966,N_29872);
nor UO_2255 (O_2255,N_28317,N_28012);
xor UO_2256 (O_2256,N_28096,N_28297);
and UO_2257 (O_2257,N_28470,N_28861);
nand UO_2258 (O_2258,N_29526,N_28302);
and UO_2259 (O_2259,N_28337,N_28013);
nand UO_2260 (O_2260,N_28537,N_28511);
nor UO_2261 (O_2261,N_29200,N_28615);
or UO_2262 (O_2262,N_29367,N_29743);
or UO_2263 (O_2263,N_28113,N_29727);
or UO_2264 (O_2264,N_29455,N_28344);
nand UO_2265 (O_2265,N_29090,N_29421);
or UO_2266 (O_2266,N_29730,N_28898);
nor UO_2267 (O_2267,N_29853,N_28766);
xor UO_2268 (O_2268,N_29868,N_28519);
and UO_2269 (O_2269,N_28129,N_29739);
or UO_2270 (O_2270,N_28979,N_29654);
xor UO_2271 (O_2271,N_28142,N_28392);
and UO_2272 (O_2272,N_29687,N_28555);
nor UO_2273 (O_2273,N_28042,N_28217);
and UO_2274 (O_2274,N_29940,N_28887);
or UO_2275 (O_2275,N_28841,N_29458);
nor UO_2276 (O_2276,N_29233,N_28645);
nor UO_2277 (O_2277,N_28428,N_28637);
xor UO_2278 (O_2278,N_28191,N_29583);
nand UO_2279 (O_2279,N_28078,N_29311);
nand UO_2280 (O_2280,N_28130,N_29675);
and UO_2281 (O_2281,N_28963,N_28848);
and UO_2282 (O_2282,N_29970,N_29094);
or UO_2283 (O_2283,N_28067,N_28443);
xnor UO_2284 (O_2284,N_29845,N_28465);
nand UO_2285 (O_2285,N_28925,N_29557);
or UO_2286 (O_2286,N_28420,N_28037);
nand UO_2287 (O_2287,N_28303,N_28302);
and UO_2288 (O_2288,N_29460,N_28862);
or UO_2289 (O_2289,N_29693,N_28859);
and UO_2290 (O_2290,N_28059,N_29913);
or UO_2291 (O_2291,N_29200,N_29567);
xor UO_2292 (O_2292,N_28525,N_29351);
or UO_2293 (O_2293,N_28924,N_29878);
xor UO_2294 (O_2294,N_29284,N_28163);
or UO_2295 (O_2295,N_29251,N_29232);
nor UO_2296 (O_2296,N_28027,N_29016);
xor UO_2297 (O_2297,N_28174,N_28208);
or UO_2298 (O_2298,N_29733,N_28401);
nand UO_2299 (O_2299,N_29238,N_28160);
xnor UO_2300 (O_2300,N_28315,N_28153);
xnor UO_2301 (O_2301,N_28267,N_29006);
xor UO_2302 (O_2302,N_28774,N_28169);
or UO_2303 (O_2303,N_29145,N_29817);
nand UO_2304 (O_2304,N_28118,N_29609);
and UO_2305 (O_2305,N_28051,N_29798);
nand UO_2306 (O_2306,N_28387,N_29869);
nand UO_2307 (O_2307,N_28020,N_29771);
or UO_2308 (O_2308,N_28076,N_29199);
xnor UO_2309 (O_2309,N_28071,N_29225);
and UO_2310 (O_2310,N_28081,N_29053);
xnor UO_2311 (O_2311,N_28667,N_29648);
nand UO_2312 (O_2312,N_28080,N_28060);
xor UO_2313 (O_2313,N_29047,N_29740);
nor UO_2314 (O_2314,N_29203,N_29441);
xor UO_2315 (O_2315,N_29991,N_28768);
xnor UO_2316 (O_2316,N_29754,N_29224);
and UO_2317 (O_2317,N_28006,N_29065);
or UO_2318 (O_2318,N_28345,N_29723);
xnor UO_2319 (O_2319,N_29782,N_29633);
and UO_2320 (O_2320,N_29848,N_29204);
xnor UO_2321 (O_2321,N_29648,N_28712);
or UO_2322 (O_2322,N_29518,N_28344);
or UO_2323 (O_2323,N_28874,N_29073);
nand UO_2324 (O_2324,N_28297,N_29679);
nor UO_2325 (O_2325,N_28459,N_28691);
nand UO_2326 (O_2326,N_29597,N_28471);
or UO_2327 (O_2327,N_28570,N_28357);
and UO_2328 (O_2328,N_29411,N_29033);
or UO_2329 (O_2329,N_28693,N_29084);
nor UO_2330 (O_2330,N_28213,N_29798);
xor UO_2331 (O_2331,N_28907,N_29934);
nor UO_2332 (O_2332,N_28400,N_28237);
or UO_2333 (O_2333,N_28728,N_28752);
nand UO_2334 (O_2334,N_28719,N_28195);
or UO_2335 (O_2335,N_28137,N_28053);
or UO_2336 (O_2336,N_28323,N_28698);
and UO_2337 (O_2337,N_28434,N_29424);
and UO_2338 (O_2338,N_28125,N_29639);
nand UO_2339 (O_2339,N_28534,N_28222);
xor UO_2340 (O_2340,N_29922,N_29169);
or UO_2341 (O_2341,N_29518,N_28788);
nor UO_2342 (O_2342,N_29793,N_28318);
nor UO_2343 (O_2343,N_29539,N_29344);
xnor UO_2344 (O_2344,N_28956,N_29449);
or UO_2345 (O_2345,N_28722,N_28592);
nor UO_2346 (O_2346,N_29119,N_28968);
nor UO_2347 (O_2347,N_29265,N_28909);
and UO_2348 (O_2348,N_28392,N_29828);
nand UO_2349 (O_2349,N_29832,N_28108);
and UO_2350 (O_2350,N_28804,N_28161);
or UO_2351 (O_2351,N_28756,N_29094);
nand UO_2352 (O_2352,N_29311,N_28473);
or UO_2353 (O_2353,N_29584,N_28799);
and UO_2354 (O_2354,N_29387,N_28954);
or UO_2355 (O_2355,N_28706,N_28604);
or UO_2356 (O_2356,N_28192,N_29736);
and UO_2357 (O_2357,N_29291,N_28980);
nand UO_2358 (O_2358,N_29737,N_28250);
nand UO_2359 (O_2359,N_29501,N_28422);
xor UO_2360 (O_2360,N_29904,N_28305);
or UO_2361 (O_2361,N_28254,N_28213);
xor UO_2362 (O_2362,N_29331,N_28426);
nor UO_2363 (O_2363,N_28096,N_29224);
and UO_2364 (O_2364,N_28284,N_29110);
nor UO_2365 (O_2365,N_28964,N_28536);
nor UO_2366 (O_2366,N_29247,N_28161);
nor UO_2367 (O_2367,N_29645,N_28468);
nor UO_2368 (O_2368,N_28817,N_28070);
nand UO_2369 (O_2369,N_29901,N_29589);
xor UO_2370 (O_2370,N_29802,N_28901);
and UO_2371 (O_2371,N_29956,N_28944);
and UO_2372 (O_2372,N_29289,N_28257);
or UO_2373 (O_2373,N_28440,N_28937);
and UO_2374 (O_2374,N_29802,N_28994);
or UO_2375 (O_2375,N_29064,N_28657);
nor UO_2376 (O_2376,N_28850,N_28664);
or UO_2377 (O_2377,N_29409,N_28122);
and UO_2378 (O_2378,N_28598,N_28565);
and UO_2379 (O_2379,N_29977,N_29867);
xor UO_2380 (O_2380,N_29062,N_28973);
and UO_2381 (O_2381,N_29355,N_29047);
nor UO_2382 (O_2382,N_28206,N_29363);
nand UO_2383 (O_2383,N_28640,N_29676);
nor UO_2384 (O_2384,N_29606,N_29841);
or UO_2385 (O_2385,N_28194,N_29093);
nor UO_2386 (O_2386,N_29594,N_28674);
and UO_2387 (O_2387,N_29314,N_29031);
and UO_2388 (O_2388,N_28823,N_29790);
xor UO_2389 (O_2389,N_28348,N_28319);
xnor UO_2390 (O_2390,N_28800,N_29766);
nand UO_2391 (O_2391,N_28646,N_29089);
nand UO_2392 (O_2392,N_28316,N_28389);
nor UO_2393 (O_2393,N_29065,N_29702);
xnor UO_2394 (O_2394,N_29160,N_28335);
xnor UO_2395 (O_2395,N_29005,N_29331);
xnor UO_2396 (O_2396,N_28916,N_28550);
and UO_2397 (O_2397,N_28325,N_28365);
nor UO_2398 (O_2398,N_29041,N_29805);
and UO_2399 (O_2399,N_28911,N_28286);
nand UO_2400 (O_2400,N_28498,N_28832);
or UO_2401 (O_2401,N_29407,N_29424);
xor UO_2402 (O_2402,N_28724,N_29775);
or UO_2403 (O_2403,N_28664,N_28701);
nand UO_2404 (O_2404,N_29508,N_29047);
and UO_2405 (O_2405,N_28157,N_28171);
xnor UO_2406 (O_2406,N_28214,N_28098);
nor UO_2407 (O_2407,N_28083,N_28508);
or UO_2408 (O_2408,N_29174,N_28682);
nor UO_2409 (O_2409,N_29100,N_28459);
xnor UO_2410 (O_2410,N_28066,N_28387);
and UO_2411 (O_2411,N_29661,N_28479);
or UO_2412 (O_2412,N_28440,N_29525);
nor UO_2413 (O_2413,N_29095,N_28944);
nand UO_2414 (O_2414,N_29494,N_29154);
or UO_2415 (O_2415,N_29374,N_28147);
and UO_2416 (O_2416,N_29769,N_28090);
and UO_2417 (O_2417,N_28798,N_29457);
nor UO_2418 (O_2418,N_29682,N_28896);
or UO_2419 (O_2419,N_28928,N_28895);
and UO_2420 (O_2420,N_29227,N_29812);
nor UO_2421 (O_2421,N_28142,N_29425);
nand UO_2422 (O_2422,N_28848,N_29385);
xor UO_2423 (O_2423,N_29472,N_28625);
and UO_2424 (O_2424,N_28078,N_29339);
xnor UO_2425 (O_2425,N_29852,N_29438);
nand UO_2426 (O_2426,N_28789,N_28292);
nor UO_2427 (O_2427,N_28550,N_28463);
nor UO_2428 (O_2428,N_29543,N_28985);
nand UO_2429 (O_2429,N_28655,N_28793);
xnor UO_2430 (O_2430,N_28418,N_29067);
or UO_2431 (O_2431,N_28842,N_29783);
or UO_2432 (O_2432,N_29703,N_28010);
nor UO_2433 (O_2433,N_29386,N_28554);
or UO_2434 (O_2434,N_29351,N_28844);
nand UO_2435 (O_2435,N_29008,N_28216);
and UO_2436 (O_2436,N_29160,N_28823);
and UO_2437 (O_2437,N_29508,N_29299);
and UO_2438 (O_2438,N_28063,N_28630);
and UO_2439 (O_2439,N_28292,N_28727);
nor UO_2440 (O_2440,N_29120,N_29770);
nor UO_2441 (O_2441,N_29661,N_28356);
nor UO_2442 (O_2442,N_28698,N_29648);
and UO_2443 (O_2443,N_28444,N_29303);
nor UO_2444 (O_2444,N_29324,N_28986);
or UO_2445 (O_2445,N_29850,N_28926);
and UO_2446 (O_2446,N_29459,N_29722);
nor UO_2447 (O_2447,N_28454,N_29123);
nor UO_2448 (O_2448,N_29047,N_28712);
nor UO_2449 (O_2449,N_29013,N_28210);
and UO_2450 (O_2450,N_28217,N_28895);
nor UO_2451 (O_2451,N_28952,N_28280);
or UO_2452 (O_2452,N_29976,N_29697);
xor UO_2453 (O_2453,N_29063,N_29247);
and UO_2454 (O_2454,N_28307,N_28812);
and UO_2455 (O_2455,N_29607,N_28834);
xnor UO_2456 (O_2456,N_29797,N_29155);
nor UO_2457 (O_2457,N_28934,N_28482);
nor UO_2458 (O_2458,N_29616,N_29186);
nand UO_2459 (O_2459,N_29086,N_28965);
xnor UO_2460 (O_2460,N_29470,N_29706);
and UO_2461 (O_2461,N_28297,N_28699);
and UO_2462 (O_2462,N_29516,N_28048);
and UO_2463 (O_2463,N_29720,N_29360);
or UO_2464 (O_2464,N_28785,N_28118);
nand UO_2465 (O_2465,N_28259,N_28613);
or UO_2466 (O_2466,N_28236,N_29558);
or UO_2467 (O_2467,N_29303,N_29316);
and UO_2468 (O_2468,N_29838,N_28862);
and UO_2469 (O_2469,N_29309,N_29072);
and UO_2470 (O_2470,N_28895,N_28584);
xor UO_2471 (O_2471,N_29665,N_28991);
nor UO_2472 (O_2472,N_29146,N_29489);
nor UO_2473 (O_2473,N_28893,N_28422);
xnor UO_2474 (O_2474,N_28396,N_29298);
xnor UO_2475 (O_2475,N_28110,N_28272);
and UO_2476 (O_2476,N_28064,N_29498);
nor UO_2477 (O_2477,N_29426,N_28376);
and UO_2478 (O_2478,N_28945,N_29388);
nor UO_2479 (O_2479,N_28277,N_28370);
and UO_2480 (O_2480,N_28115,N_29571);
nor UO_2481 (O_2481,N_29407,N_29154);
nor UO_2482 (O_2482,N_29325,N_28099);
xnor UO_2483 (O_2483,N_28677,N_28838);
and UO_2484 (O_2484,N_28040,N_28737);
and UO_2485 (O_2485,N_28794,N_29198);
or UO_2486 (O_2486,N_29112,N_29645);
and UO_2487 (O_2487,N_28692,N_28572);
or UO_2488 (O_2488,N_28091,N_28267);
nor UO_2489 (O_2489,N_29511,N_28824);
xnor UO_2490 (O_2490,N_28470,N_29848);
nand UO_2491 (O_2491,N_28475,N_28521);
nor UO_2492 (O_2492,N_29422,N_28620);
xnor UO_2493 (O_2493,N_29954,N_28146);
nand UO_2494 (O_2494,N_28920,N_28872);
nand UO_2495 (O_2495,N_29188,N_28321);
xor UO_2496 (O_2496,N_28000,N_28209);
xnor UO_2497 (O_2497,N_28923,N_28550);
nand UO_2498 (O_2498,N_29471,N_28934);
or UO_2499 (O_2499,N_28050,N_29179);
xor UO_2500 (O_2500,N_29001,N_29865);
nand UO_2501 (O_2501,N_29964,N_28408);
and UO_2502 (O_2502,N_29253,N_29411);
xor UO_2503 (O_2503,N_28274,N_29465);
nor UO_2504 (O_2504,N_29395,N_29773);
nor UO_2505 (O_2505,N_28299,N_29978);
or UO_2506 (O_2506,N_28405,N_28174);
nand UO_2507 (O_2507,N_28735,N_29842);
nor UO_2508 (O_2508,N_29966,N_28050);
nand UO_2509 (O_2509,N_28206,N_28548);
nor UO_2510 (O_2510,N_28844,N_29686);
nor UO_2511 (O_2511,N_28819,N_28790);
and UO_2512 (O_2512,N_29561,N_28911);
nor UO_2513 (O_2513,N_28905,N_29247);
or UO_2514 (O_2514,N_29749,N_28943);
and UO_2515 (O_2515,N_28342,N_29508);
nor UO_2516 (O_2516,N_29451,N_29937);
xnor UO_2517 (O_2517,N_29514,N_28513);
nand UO_2518 (O_2518,N_29636,N_29916);
and UO_2519 (O_2519,N_29279,N_29060);
and UO_2520 (O_2520,N_29714,N_28109);
or UO_2521 (O_2521,N_28426,N_29302);
nor UO_2522 (O_2522,N_28899,N_28005);
nor UO_2523 (O_2523,N_29440,N_28512);
nor UO_2524 (O_2524,N_28566,N_28461);
or UO_2525 (O_2525,N_29722,N_28993);
nand UO_2526 (O_2526,N_29208,N_29929);
nand UO_2527 (O_2527,N_28346,N_29276);
xor UO_2528 (O_2528,N_28101,N_29493);
xor UO_2529 (O_2529,N_28764,N_29889);
or UO_2530 (O_2530,N_29302,N_29864);
nor UO_2531 (O_2531,N_28912,N_29732);
xor UO_2532 (O_2532,N_28935,N_29342);
or UO_2533 (O_2533,N_29685,N_29917);
or UO_2534 (O_2534,N_29301,N_29972);
nand UO_2535 (O_2535,N_29751,N_28216);
nand UO_2536 (O_2536,N_29693,N_29528);
xnor UO_2537 (O_2537,N_29417,N_28916);
or UO_2538 (O_2538,N_29568,N_29690);
xnor UO_2539 (O_2539,N_29811,N_29868);
nand UO_2540 (O_2540,N_29211,N_29659);
xor UO_2541 (O_2541,N_28578,N_28367);
nand UO_2542 (O_2542,N_28761,N_28576);
nand UO_2543 (O_2543,N_28057,N_29611);
xor UO_2544 (O_2544,N_28981,N_28305);
nand UO_2545 (O_2545,N_28885,N_29714);
xor UO_2546 (O_2546,N_29755,N_29029);
nor UO_2547 (O_2547,N_28870,N_29716);
or UO_2548 (O_2548,N_29929,N_29872);
nor UO_2549 (O_2549,N_29739,N_29655);
nand UO_2550 (O_2550,N_28749,N_29343);
xnor UO_2551 (O_2551,N_28624,N_29426);
or UO_2552 (O_2552,N_29487,N_29802);
or UO_2553 (O_2553,N_29214,N_29587);
and UO_2554 (O_2554,N_29826,N_29703);
or UO_2555 (O_2555,N_28256,N_28053);
and UO_2556 (O_2556,N_28985,N_29829);
nor UO_2557 (O_2557,N_29806,N_28776);
nor UO_2558 (O_2558,N_29339,N_28479);
nor UO_2559 (O_2559,N_29375,N_29028);
xnor UO_2560 (O_2560,N_29730,N_28995);
nor UO_2561 (O_2561,N_28743,N_28932);
nor UO_2562 (O_2562,N_28126,N_28700);
xor UO_2563 (O_2563,N_29072,N_29905);
nor UO_2564 (O_2564,N_29243,N_28635);
or UO_2565 (O_2565,N_28741,N_28192);
nor UO_2566 (O_2566,N_28519,N_29220);
or UO_2567 (O_2567,N_28072,N_29732);
xnor UO_2568 (O_2568,N_29002,N_28604);
or UO_2569 (O_2569,N_29060,N_28717);
xor UO_2570 (O_2570,N_28260,N_28608);
xnor UO_2571 (O_2571,N_29059,N_28180);
xor UO_2572 (O_2572,N_29971,N_29038);
nand UO_2573 (O_2573,N_28207,N_28076);
and UO_2574 (O_2574,N_28956,N_28836);
nand UO_2575 (O_2575,N_28797,N_28879);
and UO_2576 (O_2576,N_29422,N_29205);
xor UO_2577 (O_2577,N_29499,N_29183);
nand UO_2578 (O_2578,N_29364,N_29056);
or UO_2579 (O_2579,N_28442,N_29422);
nand UO_2580 (O_2580,N_28938,N_29821);
nand UO_2581 (O_2581,N_28605,N_28639);
and UO_2582 (O_2582,N_29309,N_28952);
or UO_2583 (O_2583,N_29589,N_29547);
nand UO_2584 (O_2584,N_28689,N_29942);
xor UO_2585 (O_2585,N_29469,N_28729);
and UO_2586 (O_2586,N_28169,N_28602);
xor UO_2587 (O_2587,N_29118,N_28150);
xnor UO_2588 (O_2588,N_29771,N_28743);
and UO_2589 (O_2589,N_29373,N_29485);
or UO_2590 (O_2590,N_29125,N_29386);
nor UO_2591 (O_2591,N_28567,N_28285);
nand UO_2592 (O_2592,N_29719,N_28379);
or UO_2593 (O_2593,N_29247,N_28440);
or UO_2594 (O_2594,N_28508,N_28838);
or UO_2595 (O_2595,N_29209,N_29338);
and UO_2596 (O_2596,N_28666,N_29011);
nand UO_2597 (O_2597,N_29842,N_28539);
nand UO_2598 (O_2598,N_29352,N_29409);
nor UO_2599 (O_2599,N_29903,N_28566);
nand UO_2600 (O_2600,N_28569,N_29110);
or UO_2601 (O_2601,N_29292,N_28533);
or UO_2602 (O_2602,N_28544,N_28976);
and UO_2603 (O_2603,N_28078,N_29249);
xnor UO_2604 (O_2604,N_29364,N_29560);
nand UO_2605 (O_2605,N_28858,N_29281);
nor UO_2606 (O_2606,N_29790,N_28144);
or UO_2607 (O_2607,N_28366,N_29536);
nand UO_2608 (O_2608,N_28242,N_28579);
or UO_2609 (O_2609,N_28638,N_28842);
xnor UO_2610 (O_2610,N_29751,N_29002);
and UO_2611 (O_2611,N_29982,N_29365);
nand UO_2612 (O_2612,N_29106,N_28696);
and UO_2613 (O_2613,N_29940,N_29287);
nand UO_2614 (O_2614,N_29044,N_29447);
xor UO_2615 (O_2615,N_28208,N_29100);
nor UO_2616 (O_2616,N_28763,N_29264);
nand UO_2617 (O_2617,N_29098,N_28394);
nand UO_2618 (O_2618,N_29391,N_28778);
nor UO_2619 (O_2619,N_29374,N_29582);
and UO_2620 (O_2620,N_29132,N_29775);
xnor UO_2621 (O_2621,N_28063,N_29436);
xnor UO_2622 (O_2622,N_29755,N_29672);
or UO_2623 (O_2623,N_29525,N_28020);
xnor UO_2624 (O_2624,N_28902,N_29985);
and UO_2625 (O_2625,N_29572,N_29203);
nor UO_2626 (O_2626,N_28072,N_28488);
and UO_2627 (O_2627,N_28026,N_29690);
and UO_2628 (O_2628,N_28385,N_28097);
xnor UO_2629 (O_2629,N_28344,N_28452);
xnor UO_2630 (O_2630,N_28516,N_28680);
and UO_2631 (O_2631,N_29068,N_28304);
nor UO_2632 (O_2632,N_29444,N_28941);
nand UO_2633 (O_2633,N_29837,N_29038);
xor UO_2634 (O_2634,N_29885,N_29946);
nand UO_2635 (O_2635,N_29027,N_29655);
nand UO_2636 (O_2636,N_29258,N_29889);
or UO_2637 (O_2637,N_28125,N_29841);
nand UO_2638 (O_2638,N_29999,N_28335);
nor UO_2639 (O_2639,N_29574,N_29755);
xnor UO_2640 (O_2640,N_29195,N_29870);
nand UO_2641 (O_2641,N_28594,N_29410);
or UO_2642 (O_2642,N_28999,N_28280);
or UO_2643 (O_2643,N_28398,N_29370);
and UO_2644 (O_2644,N_29699,N_29989);
xnor UO_2645 (O_2645,N_28830,N_29534);
or UO_2646 (O_2646,N_28564,N_29073);
and UO_2647 (O_2647,N_29117,N_29008);
nand UO_2648 (O_2648,N_29108,N_28705);
nor UO_2649 (O_2649,N_29385,N_28422);
xor UO_2650 (O_2650,N_29803,N_29163);
and UO_2651 (O_2651,N_29476,N_28362);
xor UO_2652 (O_2652,N_28461,N_28722);
or UO_2653 (O_2653,N_29850,N_28766);
and UO_2654 (O_2654,N_28164,N_28536);
nor UO_2655 (O_2655,N_28538,N_29225);
or UO_2656 (O_2656,N_29133,N_29575);
nand UO_2657 (O_2657,N_28844,N_28601);
and UO_2658 (O_2658,N_28182,N_28586);
xnor UO_2659 (O_2659,N_29199,N_28971);
nor UO_2660 (O_2660,N_29391,N_29113);
and UO_2661 (O_2661,N_29636,N_29768);
nand UO_2662 (O_2662,N_29836,N_28801);
nor UO_2663 (O_2663,N_28862,N_28674);
nor UO_2664 (O_2664,N_28708,N_29045);
or UO_2665 (O_2665,N_28673,N_29955);
or UO_2666 (O_2666,N_29556,N_29707);
nor UO_2667 (O_2667,N_29717,N_29258);
nor UO_2668 (O_2668,N_28041,N_28447);
nor UO_2669 (O_2669,N_28739,N_28339);
or UO_2670 (O_2670,N_29969,N_28262);
nor UO_2671 (O_2671,N_29317,N_28119);
and UO_2672 (O_2672,N_28946,N_28268);
and UO_2673 (O_2673,N_28791,N_28736);
nor UO_2674 (O_2674,N_28341,N_29429);
and UO_2675 (O_2675,N_28080,N_28057);
and UO_2676 (O_2676,N_29912,N_28815);
nand UO_2677 (O_2677,N_28846,N_29635);
nand UO_2678 (O_2678,N_29203,N_29059);
nand UO_2679 (O_2679,N_29856,N_29207);
nand UO_2680 (O_2680,N_28326,N_29971);
nand UO_2681 (O_2681,N_29847,N_28140);
nor UO_2682 (O_2682,N_28867,N_28360);
xnor UO_2683 (O_2683,N_28468,N_28731);
and UO_2684 (O_2684,N_29663,N_29581);
and UO_2685 (O_2685,N_29226,N_29555);
nand UO_2686 (O_2686,N_28755,N_28456);
or UO_2687 (O_2687,N_29835,N_29141);
xor UO_2688 (O_2688,N_28504,N_29857);
xnor UO_2689 (O_2689,N_28546,N_29427);
and UO_2690 (O_2690,N_28137,N_29996);
and UO_2691 (O_2691,N_29251,N_29767);
or UO_2692 (O_2692,N_29855,N_29287);
nor UO_2693 (O_2693,N_28611,N_29723);
or UO_2694 (O_2694,N_29208,N_28810);
or UO_2695 (O_2695,N_28523,N_29959);
nand UO_2696 (O_2696,N_29236,N_29350);
or UO_2697 (O_2697,N_28802,N_28841);
xor UO_2698 (O_2698,N_28644,N_29314);
nor UO_2699 (O_2699,N_28402,N_29108);
xor UO_2700 (O_2700,N_28017,N_28065);
and UO_2701 (O_2701,N_29759,N_28349);
and UO_2702 (O_2702,N_29592,N_29090);
and UO_2703 (O_2703,N_28608,N_28115);
nor UO_2704 (O_2704,N_28520,N_29736);
xor UO_2705 (O_2705,N_29735,N_28933);
xnor UO_2706 (O_2706,N_29617,N_29287);
and UO_2707 (O_2707,N_29927,N_29920);
nand UO_2708 (O_2708,N_29884,N_29562);
nand UO_2709 (O_2709,N_28342,N_28780);
nand UO_2710 (O_2710,N_29686,N_28056);
and UO_2711 (O_2711,N_28156,N_28525);
xor UO_2712 (O_2712,N_28968,N_28498);
xor UO_2713 (O_2713,N_28387,N_28650);
nand UO_2714 (O_2714,N_28998,N_29985);
and UO_2715 (O_2715,N_28516,N_29897);
and UO_2716 (O_2716,N_28008,N_29129);
nand UO_2717 (O_2717,N_29045,N_29256);
nor UO_2718 (O_2718,N_29014,N_28867);
xor UO_2719 (O_2719,N_28510,N_29578);
and UO_2720 (O_2720,N_29909,N_29125);
or UO_2721 (O_2721,N_28186,N_29164);
or UO_2722 (O_2722,N_28112,N_29892);
nor UO_2723 (O_2723,N_29245,N_28584);
nor UO_2724 (O_2724,N_29155,N_28982);
nand UO_2725 (O_2725,N_28184,N_29195);
nand UO_2726 (O_2726,N_29465,N_29214);
xor UO_2727 (O_2727,N_29479,N_29521);
or UO_2728 (O_2728,N_29823,N_28701);
xnor UO_2729 (O_2729,N_29252,N_29364);
nand UO_2730 (O_2730,N_28740,N_28764);
nand UO_2731 (O_2731,N_28250,N_29093);
and UO_2732 (O_2732,N_29236,N_29239);
and UO_2733 (O_2733,N_29419,N_28393);
nand UO_2734 (O_2734,N_28750,N_28631);
nor UO_2735 (O_2735,N_28505,N_29368);
or UO_2736 (O_2736,N_29638,N_29083);
and UO_2737 (O_2737,N_28067,N_29399);
and UO_2738 (O_2738,N_29340,N_29484);
nand UO_2739 (O_2739,N_29030,N_28027);
and UO_2740 (O_2740,N_29274,N_29220);
nand UO_2741 (O_2741,N_29925,N_28190);
nor UO_2742 (O_2742,N_28737,N_29153);
or UO_2743 (O_2743,N_28873,N_29056);
xnor UO_2744 (O_2744,N_29072,N_28661);
xor UO_2745 (O_2745,N_28736,N_28794);
and UO_2746 (O_2746,N_28146,N_28895);
or UO_2747 (O_2747,N_28792,N_29259);
xor UO_2748 (O_2748,N_29075,N_29094);
or UO_2749 (O_2749,N_29928,N_28104);
or UO_2750 (O_2750,N_29841,N_28074);
or UO_2751 (O_2751,N_29929,N_29482);
nor UO_2752 (O_2752,N_29053,N_28534);
nand UO_2753 (O_2753,N_28070,N_29989);
or UO_2754 (O_2754,N_29293,N_29119);
and UO_2755 (O_2755,N_29261,N_28053);
or UO_2756 (O_2756,N_28773,N_29696);
nand UO_2757 (O_2757,N_28425,N_29454);
nor UO_2758 (O_2758,N_28704,N_29447);
xnor UO_2759 (O_2759,N_29430,N_29106);
and UO_2760 (O_2760,N_29037,N_29034);
nor UO_2761 (O_2761,N_28255,N_29726);
or UO_2762 (O_2762,N_28320,N_28656);
and UO_2763 (O_2763,N_28417,N_29525);
xnor UO_2764 (O_2764,N_29225,N_28884);
nor UO_2765 (O_2765,N_28545,N_29043);
nand UO_2766 (O_2766,N_29871,N_28717);
xnor UO_2767 (O_2767,N_29435,N_29832);
nand UO_2768 (O_2768,N_29157,N_28618);
and UO_2769 (O_2769,N_29389,N_28617);
nand UO_2770 (O_2770,N_29127,N_29968);
and UO_2771 (O_2771,N_28603,N_29661);
or UO_2772 (O_2772,N_29063,N_28984);
or UO_2773 (O_2773,N_28717,N_29956);
or UO_2774 (O_2774,N_28263,N_29848);
nor UO_2775 (O_2775,N_28715,N_28189);
or UO_2776 (O_2776,N_29684,N_28872);
nand UO_2777 (O_2777,N_29186,N_28230);
nor UO_2778 (O_2778,N_28224,N_29416);
and UO_2779 (O_2779,N_29502,N_29762);
xnor UO_2780 (O_2780,N_29182,N_28532);
nor UO_2781 (O_2781,N_28829,N_28567);
nand UO_2782 (O_2782,N_29676,N_28353);
nand UO_2783 (O_2783,N_28224,N_29586);
or UO_2784 (O_2784,N_29310,N_29587);
and UO_2785 (O_2785,N_28908,N_28148);
xnor UO_2786 (O_2786,N_29322,N_29708);
and UO_2787 (O_2787,N_29855,N_29632);
or UO_2788 (O_2788,N_28059,N_29768);
xor UO_2789 (O_2789,N_28680,N_28817);
nand UO_2790 (O_2790,N_29634,N_29970);
nand UO_2791 (O_2791,N_29301,N_29401);
nand UO_2792 (O_2792,N_29875,N_28348);
or UO_2793 (O_2793,N_29032,N_29793);
xor UO_2794 (O_2794,N_29134,N_28928);
and UO_2795 (O_2795,N_28627,N_29149);
nand UO_2796 (O_2796,N_29696,N_29877);
xnor UO_2797 (O_2797,N_28158,N_28796);
xnor UO_2798 (O_2798,N_29199,N_28283);
nand UO_2799 (O_2799,N_28664,N_29387);
xor UO_2800 (O_2800,N_28397,N_29396);
xnor UO_2801 (O_2801,N_29165,N_28528);
or UO_2802 (O_2802,N_28905,N_29564);
or UO_2803 (O_2803,N_29569,N_28163);
and UO_2804 (O_2804,N_28952,N_29609);
xor UO_2805 (O_2805,N_28490,N_28102);
and UO_2806 (O_2806,N_28740,N_28162);
and UO_2807 (O_2807,N_28923,N_28904);
nand UO_2808 (O_2808,N_28134,N_29845);
xnor UO_2809 (O_2809,N_29923,N_29424);
nor UO_2810 (O_2810,N_29238,N_29990);
nand UO_2811 (O_2811,N_29941,N_29760);
and UO_2812 (O_2812,N_28068,N_28519);
xor UO_2813 (O_2813,N_29575,N_28927);
xor UO_2814 (O_2814,N_28095,N_28422);
nor UO_2815 (O_2815,N_29591,N_28941);
nand UO_2816 (O_2816,N_29964,N_28791);
nor UO_2817 (O_2817,N_29986,N_28896);
nor UO_2818 (O_2818,N_29411,N_28105);
xnor UO_2819 (O_2819,N_28840,N_28804);
and UO_2820 (O_2820,N_28939,N_28978);
and UO_2821 (O_2821,N_28882,N_29671);
nor UO_2822 (O_2822,N_29828,N_29289);
nor UO_2823 (O_2823,N_28364,N_29853);
or UO_2824 (O_2824,N_29503,N_28113);
xnor UO_2825 (O_2825,N_28546,N_29722);
nand UO_2826 (O_2826,N_29366,N_28951);
nor UO_2827 (O_2827,N_28907,N_28081);
or UO_2828 (O_2828,N_28209,N_29786);
nor UO_2829 (O_2829,N_29343,N_29966);
nand UO_2830 (O_2830,N_29896,N_29494);
nand UO_2831 (O_2831,N_28320,N_29430);
nor UO_2832 (O_2832,N_29709,N_29539);
nor UO_2833 (O_2833,N_28048,N_29410);
nor UO_2834 (O_2834,N_29961,N_29568);
xnor UO_2835 (O_2835,N_28703,N_28040);
nor UO_2836 (O_2836,N_29344,N_28238);
and UO_2837 (O_2837,N_29829,N_29786);
nand UO_2838 (O_2838,N_28701,N_29125);
and UO_2839 (O_2839,N_29260,N_29145);
nor UO_2840 (O_2840,N_29599,N_29738);
nand UO_2841 (O_2841,N_29608,N_29964);
or UO_2842 (O_2842,N_29924,N_29849);
and UO_2843 (O_2843,N_29014,N_28681);
and UO_2844 (O_2844,N_28141,N_29064);
nand UO_2845 (O_2845,N_28731,N_29162);
nor UO_2846 (O_2846,N_29776,N_29073);
or UO_2847 (O_2847,N_29860,N_28735);
or UO_2848 (O_2848,N_28803,N_29001);
nor UO_2849 (O_2849,N_29636,N_29973);
nand UO_2850 (O_2850,N_28451,N_28528);
xnor UO_2851 (O_2851,N_29154,N_29319);
nand UO_2852 (O_2852,N_29928,N_28429);
nor UO_2853 (O_2853,N_28560,N_29596);
xnor UO_2854 (O_2854,N_28399,N_29008);
nor UO_2855 (O_2855,N_28247,N_28062);
xnor UO_2856 (O_2856,N_28229,N_28882);
nand UO_2857 (O_2857,N_28413,N_29656);
nand UO_2858 (O_2858,N_28974,N_28987);
nor UO_2859 (O_2859,N_29108,N_29582);
nor UO_2860 (O_2860,N_28072,N_28711);
nand UO_2861 (O_2861,N_28093,N_29031);
or UO_2862 (O_2862,N_28087,N_28374);
xor UO_2863 (O_2863,N_29047,N_28210);
or UO_2864 (O_2864,N_28949,N_29998);
and UO_2865 (O_2865,N_28138,N_29380);
and UO_2866 (O_2866,N_29566,N_28115);
nor UO_2867 (O_2867,N_29072,N_29140);
and UO_2868 (O_2868,N_29842,N_29611);
and UO_2869 (O_2869,N_29498,N_28939);
xnor UO_2870 (O_2870,N_28529,N_29957);
nor UO_2871 (O_2871,N_28283,N_28028);
xnor UO_2872 (O_2872,N_28504,N_28669);
xor UO_2873 (O_2873,N_28270,N_29672);
or UO_2874 (O_2874,N_29901,N_28897);
xor UO_2875 (O_2875,N_28570,N_29917);
and UO_2876 (O_2876,N_29822,N_28493);
nand UO_2877 (O_2877,N_28667,N_28123);
nor UO_2878 (O_2878,N_28266,N_29661);
xor UO_2879 (O_2879,N_28092,N_28405);
xnor UO_2880 (O_2880,N_29238,N_29831);
xnor UO_2881 (O_2881,N_28073,N_29304);
xor UO_2882 (O_2882,N_29585,N_28054);
xor UO_2883 (O_2883,N_28417,N_29204);
and UO_2884 (O_2884,N_29198,N_28732);
nand UO_2885 (O_2885,N_28048,N_28762);
nor UO_2886 (O_2886,N_28642,N_28338);
xnor UO_2887 (O_2887,N_29115,N_28346);
or UO_2888 (O_2888,N_29545,N_29964);
nor UO_2889 (O_2889,N_29540,N_28474);
nand UO_2890 (O_2890,N_29788,N_29037);
xnor UO_2891 (O_2891,N_28922,N_29603);
nor UO_2892 (O_2892,N_29129,N_29815);
xor UO_2893 (O_2893,N_28766,N_28199);
or UO_2894 (O_2894,N_28977,N_29348);
xor UO_2895 (O_2895,N_29483,N_28021);
nand UO_2896 (O_2896,N_28912,N_28963);
nand UO_2897 (O_2897,N_29730,N_29399);
and UO_2898 (O_2898,N_29287,N_29367);
and UO_2899 (O_2899,N_29522,N_28565);
or UO_2900 (O_2900,N_29301,N_29693);
xnor UO_2901 (O_2901,N_29080,N_29261);
nand UO_2902 (O_2902,N_28695,N_28430);
nor UO_2903 (O_2903,N_29267,N_29916);
nand UO_2904 (O_2904,N_29873,N_28913);
nor UO_2905 (O_2905,N_29257,N_29666);
and UO_2906 (O_2906,N_28867,N_28130);
xnor UO_2907 (O_2907,N_29770,N_28599);
xor UO_2908 (O_2908,N_29590,N_28460);
nand UO_2909 (O_2909,N_29710,N_28650);
nand UO_2910 (O_2910,N_29806,N_29550);
nor UO_2911 (O_2911,N_29267,N_28685);
or UO_2912 (O_2912,N_28940,N_29133);
nor UO_2913 (O_2913,N_29551,N_28043);
or UO_2914 (O_2914,N_29370,N_29489);
nand UO_2915 (O_2915,N_29047,N_29700);
nand UO_2916 (O_2916,N_28099,N_28257);
or UO_2917 (O_2917,N_28258,N_29289);
or UO_2918 (O_2918,N_28980,N_29873);
xnor UO_2919 (O_2919,N_28158,N_29381);
nand UO_2920 (O_2920,N_28990,N_28769);
xor UO_2921 (O_2921,N_28439,N_29522);
xor UO_2922 (O_2922,N_28849,N_28644);
and UO_2923 (O_2923,N_29104,N_29999);
or UO_2924 (O_2924,N_29465,N_28593);
nor UO_2925 (O_2925,N_29123,N_29472);
nor UO_2926 (O_2926,N_29343,N_28894);
nor UO_2927 (O_2927,N_29488,N_29229);
nor UO_2928 (O_2928,N_29750,N_29622);
nor UO_2929 (O_2929,N_28788,N_29015);
xor UO_2930 (O_2930,N_29688,N_28575);
nor UO_2931 (O_2931,N_29878,N_28945);
and UO_2932 (O_2932,N_29254,N_29066);
and UO_2933 (O_2933,N_29139,N_29402);
nand UO_2934 (O_2934,N_28434,N_29805);
xnor UO_2935 (O_2935,N_28374,N_29720);
nor UO_2936 (O_2936,N_29253,N_28263);
or UO_2937 (O_2937,N_29412,N_29075);
nor UO_2938 (O_2938,N_28475,N_28251);
xor UO_2939 (O_2939,N_28674,N_28391);
xnor UO_2940 (O_2940,N_29512,N_28715);
nand UO_2941 (O_2941,N_29603,N_28663);
nor UO_2942 (O_2942,N_28073,N_29975);
or UO_2943 (O_2943,N_28380,N_29340);
xor UO_2944 (O_2944,N_29335,N_28086);
xnor UO_2945 (O_2945,N_28609,N_29784);
or UO_2946 (O_2946,N_29938,N_29428);
xnor UO_2947 (O_2947,N_29844,N_28369);
nor UO_2948 (O_2948,N_29291,N_29712);
or UO_2949 (O_2949,N_29310,N_29533);
and UO_2950 (O_2950,N_29049,N_28735);
xnor UO_2951 (O_2951,N_29530,N_28523);
nor UO_2952 (O_2952,N_28226,N_28928);
or UO_2953 (O_2953,N_28908,N_28727);
nand UO_2954 (O_2954,N_28677,N_28182);
xor UO_2955 (O_2955,N_28980,N_28185);
and UO_2956 (O_2956,N_28195,N_28351);
nand UO_2957 (O_2957,N_28102,N_29849);
or UO_2958 (O_2958,N_28409,N_29255);
or UO_2959 (O_2959,N_28806,N_28280);
or UO_2960 (O_2960,N_29094,N_28892);
xor UO_2961 (O_2961,N_29478,N_28135);
xor UO_2962 (O_2962,N_28625,N_29291);
or UO_2963 (O_2963,N_28089,N_29258);
and UO_2964 (O_2964,N_29882,N_28720);
and UO_2965 (O_2965,N_29352,N_28632);
and UO_2966 (O_2966,N_28438,N_28059);
nand UO_2967 (O_2967,N_29168,N_29937);
and UO_2968 (O_2968,N_29681,N_28343);
xnor UO_2969 (O_2969,N_28620,N_29049);
or UO_2970 (O_2970,N_29352,N_28656);
and UO_2971 (O_2971,N_28579,N_29910);
or UO_2972 (O_2972,N_29059,N_29212);
and UO_2973 (O_2973,N_29800,N_28485);
nand UO_2974 (O_2974,N_28298,N_28494);
and UO_2975 (O_2975,N_28824,N_28360);
nand UO_2976 (O_2976,N_29203,N_28623);
nand UO_2977 (O_2977,N_29770,N_28244);
or UO_2978 (O_2978,N_29700,N_28542);
or UO_2979 (O_2979,N_29590,N_28407);
nor UO_2980 (O_2980,N_29859,N_29698);
nand UO_2981 (O_2981,N_29518,N_29336);
or UO_2982 (O_2982,N_28556,N_29155);
nand UO_2983 (O_2983,N_28552,N_29462);
and UO_2984 (O_2984,N_28188,N_29783);
and UO_2985 (O_2985,N_28665,N_28629);
nor UO_2986 (O_2986,N_29426,N_29565);
or UO_2987 (O_2987,N_29665,N_29343);
and UO_2988 (O_2988,N_28550,N_29342);
nand UO_2989 (O_2989,N_28832,N_29582);
and UO_2990 (O_2990,N_28889,N_29404);
and UO_2991 (O_2991,N_29686,N_28197);
nand UO_2992 (O_2992,N_29759,N_29156);
and UO_2993 (O_2993,N_28427,N_29442);
and UO_2994 (O_2994,N_29093,N_29714);
nor UO_2995 (O_2995,N_28762,N_28740);
xor UO_2996 (O_2996,N_29315,N_28497);
nand UO_2997 (O_2997,N_28502,N_29756);
nor UO_2998 (O_2998,N_28783,N_29450);
xnor UO_2999 (O_2999,N_29737,N_29728);
nor UO_3000 (O_3000,N_29588,N_28202);
or UO_3001 (O_3001,N_29221,N_29941);
nor UO_3002 (O_3002,N_28280,N_28980);
or UO_3003 (O_3003,N_28531,N_29807);
or UO_3004 (O_3004,N_28917,N_28042);
nor UO_3005 (O_3005,N_28984,N_29065);
nor UO_3006 (O_3006,N_29161,N_28735);
nor UO_3007 (O_3007,N_29865,N_29941);
or UO_3008 (O_3008,N_29194,N_29793);
or UO_3009 (O_3009,N_28182,N_28567);
or UO_3010 (O_3010,N_29025,N_28986);
nor UO_3011 (O_3011,N_29331,N_28983);
nand UO_3012 (O_3012,N_28789,N_28595);
and UO_3013 (O_3013,N_29334,N_28180);
nand UO_3014 (O_3014,N_29399,N_28504);
xor UO_3015 (O_3015,N_29154,N_29931);
and UO_3016 (O_3016,N_28570,N_29888);
nor UO_3017 (O_3017,N_28399,N_29052);
nor UO_3018 (O_3018,N_29810,N_29683);
or UO_3019 (O_3019,N_29821,N_29056);
nor UO_3020 (O_3020,N_28981,N_29907);
nand UO_3021 (O_3021,N_28812,N_28378);
nor UO_3022 (O_3022,N_29533,N_28155);
or UO_3023 (O_3023,N_28418,N_28213);
nor UO_3024 (O_3024,N_29831,N_28830);
xor UO_3025 (O_3025,N_28796,N_29308);
and UO_3026 (O_3026,N_28499,N_29019);
nand UO_3027 (O_3027,N_28506,N_29868);
nand UO_3028 (O_3028,N_28882,N_28622);
and UO_3029 (O_3029,N_29517,N_29629);
or UO_3030 (O_3030,N_29641,N_28853);
nand UO_3031 (O_3031,N_29425,N_29874);
nor UO_3032 (O_3032,N_29354,N_29184);
nor UO_3033 (O_3033,N_28698,N_29336);
xor UO_3034 (O_3034,N_28423,N_29820);
xnor UO_3035 (O_3035,N_28157,N_29169);
and UO_3036 (O_3036,N_29266,N_29491);
nand UO_3037 (O_3037,N_29341,N_29677);
or UO_3038 (O_3038,N_29079,N_29519);
and UO_3039 (O_3039,N_28713,N_29719);
and UO_3040 (O_3040,N_29974,N_28291);
or UO_3041 (O_3041,N_29917,N_28280);
xor UO_3042 (O_3042,N_28296,N_29366);
and UO_3043 (O_3043,N_29330,N_28258);
or UO_3044 (O_3044,N_28864,N_28091);
nor UO_3045 (O_3045,N_29621,N_28399);
and UO_3046 (O_3046,N_28862,N_29714);
nor UO_3047 (O_3047,N_29640,N_28077);
or UO_3048 (O_3048,N_28787,N_29043);
nand UO_3049 (O_3049,N_28535,N_29636);
and UO_3050 (O_3050,N_29929,N_29120);
and UO_3051 (O_3051,N_28732,N_29469);
xor UO_3052 (O_3052,N_28653,N_29446);
nand UO_3053 (O_3053,N_28358,N_29162);
or UO_3054 (O_3054,N_29545,N_29092);
nand UO_3055 (O_3055,N_28071,N_28218);
nor UO_3056 (O_3056,N_29119,N_28650);
xnor UO_3057 (O_3057,N_29740,N_29978);
xor UO_3058 (O_3058,N_29073,N_29638);
or UO_3059 (O_3059,N_29386,N_29479);
or UO_3060 (O_3060,N_28040,N_29913);
nand UO_3061 (O_3061,N_29563,N_29909);
nor UO_3062 (O_3062,N_29475,N_29230);
nor UO_3063 (O_3063,N_28008,N_28558);
nor UO_3064 (O_3064,N_29430,N_29996);
or UO_3065 (O_3065,N_28584,N_28135);
nand UO_3066 (O_3066,N_28225,N_29256);
nand UO_3067 (O_3067,N_29362,N_28418);
and UO_3068 (O_3068,N_28629,N_29721);
xnor UO_3069 (O_3069,N_28995,N_29092);
or UO_3070 (O_3070,N_28264,N_28925);
or UO_3071 (O_3071,N_29932,N_28680);
xor UO_3072 (O_3072,N_29038,N_28575);
or UO_3073 (O_3073,N_29574,N_28839);
nand UO_3074 (O_3074,N_29251,N_29529);
xor UO_3075 (O_3075,N_28863,N_29890);
xnor UO_3076 (O_3076,N_29403,N_28106);
nor UO_3077 (O_3077,N_28834,N_29193);
nand UO_3078 (O_3078,N_29313,N_28273);
and UO_3079 (O_3079,N_29123,N_28097);
nor UO_3080 (O_3080,N_28883,N_29539);
nand UO_3081 (O_3081,N_28495,N_29549);
or UO_3082 (O_3082,N_28345,N_29711);
xor UO_3083 (O_3083,N_29235,N_28326);
or UO_3084 (O_3084,N_28693,N_28197);
and UO_3085 (O_3085,N_28764,N_29141);
and UO_3086 (O_3086,N_28423,N_29444);
nand UO_3087 (O_3087,N_29754,N_29610);
and UO_3088 (O_3088,N_28595,N_28780);
xnor UO_3089 (O_3089,N_28135,N_28124);
nor UO_3090 (O_3090,N_29843,N_28122);
xor UO_3091 (O_3091,N_29265,N_28355);
and UO_3092 (O_3092,N_29322,N_28265);
nor UO_3093 (O_3093,N_29957,N_29246);
or UO_3094 (O_3094,N_28912,N_29775);
or UO_3095 (O_3095,N_29024,N_29422);
or UO_3096 (O_3096,N_28459,N_29362);
and UO_3097 (O_3097,N_29574,N_28537);
nand UO_3098 (O_3098,N_29008,N_29602);
xor UO_3099 (O_3099,N_28427,N_28259);
xor UO_3100 (O_3100,N_29604,N_29506);
nor UO_3101 (O_3101,N_29839,N_28445);
nand UO_3102 (O_3102,N_28013,N_29817);
nand UO_3103 (O_3103,N_29825,N_29045);
xnor UO_3104 (O_3104,N_28392,N_28323);
and UO_3105 (O_3105,N_28575,N_28528);
nand UO_3106 (O_3106,N_28545,N_29149);
xnor UO_3107 (O_3107,N_29485,N_28260);
nor UO_3108 (O_3108,N_29454,N_28658);
and UO_3109 (O_3109,N_29006,N_29487);
and UO_3110 (O_3110,N_28805,N_28448);
nor UO_3111 (O_3111,N_28215,N_29496);
and UO_3112 (O_3112,N_28223,N_28321);
and UO_3113 (O_3113,N_28066,N_29832);
nand UO_3114 (O_3114,N_28763,N_29964);
and UO_3115 (O_3115,N_28736,N_29645);
nand UO_3116 (O_3116,N_28585,N_28359);
nand UO_3117 (O_3117,N_28229,N_29904);
and UO_3118 (O_3118,N_29844,N_29572);
nand UO_3119 (O_3119,N_29605,N_29706);
or UO_3120 (O_3120,N_29326,N_28894);
and UO_3121 (O_3121,N_29688,N_29537);
or UO_3122 (O_3122,N_29615,N_29108);
or UO_3123 (O_3123,N_28964,N_28444);
or UO_3124 (O_3124,N_28200,N_28416);
nand UO_3125 (O_3125,N_29168,N_29664);
and UO_3126 (O_3126,N_28701,N_28200);
nor UO_3127 (O_3127,N_29357,N_29922);
or UO_3128 (O_3128,N_28771,N_28846);
xor UO_3129 (O_3129,N_28878,N_29096);
nand UO_3130 (O_3130,N_29820,N_29371);
and UO_3131 (O_3131,N_29850,N_28114);
xnor UO_3132 (O_3132,N_28486,N_29459);
nor UO_3133 (O_3133,N_29597,N_29065);
and UO_3134 (O_3134,N_28361,N_28590);
or UO_3135 (O_3135,N_29723,N_29077);
or UO_3136 (O_3136,N_29582,N_29010);
or UO_3137 (O_3137,N_29034,N_28035);
or UO_3138 (O_3138,N_28506,N_29131);
or UO_3139 (O_3139,N_28304,N_28255);
xor UO_3140 (O_3140,N_29558,N_29303);
and UO_3141 (O_3141,N_28096,N_29378);
nand UO_3142 (O_3142,N_28692,N_28674);
nand UO_3143 (O_3143,N_28603,N_29977);
and UO_3144 (O_3144,N_29412,N_29454);
or UO_3145 (O_3145,N_28667,N_29506);
or UO_3146 (O_3146,N_29779,N_29618);
xnor UO_3147 (O_3147,N_28191,N_29476);
and UO_3148 (O_3148,N_28331,N_29351);
nor UO_3149 (O_3149,N_28486,N_29981);
xor UO_3150 (O_3150,N_28139,N_29785);
nand UO_3151 (O_3151,N_28567,N_29745);
and UO_3152 (O_3152,N_29035,N_29489);
or UO_3153 (O_3153,N_28791,N_29987);
or UO_3154 (O_3154,N_29798,N_29403);
and UO_3155 (O_3155,N_28558,N_28640);
xnor UO_3156 (O_3156,N_28628,N_29292);
xor UO_3157 (O_3157,N_29854,N_28199);
nor UO_3158 (O_3158,N_28765,N_28665);
xor UO_3159 (O_3159,N_29946,N_29691);
xnor UO_3160 (O_3160,N_29691,N_29763);
nand UO_3161 (O_3161,N_28513,N_28016);
nor UO_3162 (O_3162,N_29627,N_29982);
or UO_3163 (O_3163,N_28629,N_29437);
and UO_3164 (O_3164,N_29412,N_29998);
and UO_3165 (O_3165,N_29321,N_29428);
nand UO_3166 (O_3166,N_29307,N_28615);
and UO_3167 (O_3167,N_29861,N_29585);
xnor UO_3168 (O_3168,N_29788,N_28633);
xor UO_3169 (O_3169,N_28003,N_28662);
or UO_3170 (O_3170,N_28212,N_28983);
nand UO_3171 (O_3171,N_28179,N_28614);
xnor UO_3172 (O_3172,N_29831,N_28848);
nand UO_3173 (O_3173,N_28092,N_29122);
and UO_3174 (O_3174,N_28564,N_28363);
nand UO_3175 (O_3175,N_29161,N_28147);
xor UO_3176 (O_3176,N_29080,N_29543);
nand UO_3177 (O_3177,N_28875,N_28405);
and UO_3178 (O_3178,N_29588,N_29004);
and UO_3179 (O_3179,N_28525,N_29380);
xnor UO_3180 (O_3180,N_29900,N_28475);
xnor UO_3181 (O_3181,N_29286,N_28628);
nor UO_3182 (O_3182,N_29196,N_29038);
or UO_3183 (O_3183,N_28382,N_28605);
and UO_3184 (O_3184,N_28812,N_29997);
and UO_3185 (O_3185,N_28880,N_29519);
xor UO_3186 (O_3186,N_29745,N_29674);
or UO_3187 (O_3187,N_28750,N_29403);
xnor UO_3188 (O_3188,N_28239,N_29371);
nand UO_3189 (O_3189,N_28033,N_28119);
nand UO_3190 (O_3190,N_29795,N_28056);
nor UO_3191 (O_3191,N_28712,N_28266);
nand UO_3192 (O_3192,N_28649,N_28512);
nor UO_3193 (O_3193,N_28208,N_28398);
nand UO_3194 (O_3194,N_28316,N_29835);
or UO_3195 (O_3195,N_29221,N_29082);
nor UO_3196 (O_3196,N_28490,N_28819);
xor UO_3197 (O_3197,N_29093,N_29457);
nor UO_3198 (O_3198,N_28107,N_28457);
xor UO_3199 (O_3199,N_28773,N_28440);
nand UO_3200 (O_3200,N_28230,N_29062);
and UO_3201 (O_3201,N_29804,N_29519);
and UO_3202 (O_3202,N_29868,N_28365);
xor UO_3203 (O_3203,N_29538,N_29066);
nand UO_3204 (O_3204,N_29343,N_28609);
or UO_3205 (O_3205,N_28154,N_29710);
or UO_3206 (O_3206,N_29080,N_28598);
and UO_3207 (O_3207,N_28902,N_28023);
and UO_3208 (O_3208,N_28104,N_28456);
nand UO_3209 (O_3209,N_29345,N_28461);
or UO_3210 (O_3210,N_29555,N_29847);
xor UO_3211 (O_3211,N_28913,N_29565);
xor UO_3212 (O_3212,N_29775,N_28154);
and UO_3213 (O_3213,N_28446,N_28703);
or UO_3214 (O_3214,N_29909,N_29074);
or UO_3215 (O_3215,N_28085,N_28299);
or UO_3216 (O_3216,N_28482,N_29464);
and UO_3217 (O_3217,N_29448,N_29178);
nor UO_3218 (O_3218,N_29325,N_29547);
and UO_3219 (O_3219,N_29486,N_29066);
or UO_3220 (O_3220,N_29062,N_28492);
and UO_3221 (O_3221,N_28210,N_29069);
and UO_3222 (O_3222,N_29870,N_28675);
xnor UO_3223 (O_3223,N_28014,N_29891);
nor UO_3224 (O_3224,N_29335,N_29641);
nor UO_3225 (O_3225,N_28722,N_28951);
and UO_3226 (O_3226,N_29658,N_28087);
xnor UO_3227 (O_3227,N_29536,N_29998);
xnor UO_3228 (O_3228,N_28024,N_29883);
nor UO_3229 (O_3229,N_29065,N_29884);
or UO_3230 (O_3230,N_29781,N_28499);
and UO_3231 (O_3231,N_28972,N_28971);
or UO_3232 (O_3232,N_29892,N_29866);
nor UO_3233 (O_3233,N_29686,N_28964);
nand UO_3234 (O_3234,N_29910,N_28746);
nor UO_3235 (O_3235,N_28887,N_28986);
nand UO_3236 (O_3236,N_29173,N_29346);
and UO_3237 (O_3237,N_28120,N_28952);
nor UO_3238 (O_3238,N_28077,N_28934);
and UO_3239 (O_3239,N_28820,N_29832);
nand UO_3240 (O_3240,N_29117,N_29411);
and UO_3241 (O_3241,N_29527,N_29089);
nor UO_3242 (O_3242,N_29503,N_28543);
nand UO_3243 (O_3243,N_29120,N_28387);
nor UO_3244 (O_3244,N_28455,N_28682);
nor UO_3245 (O_3245,N_28480,N_28215);
xnor UO_3246 (O_3246,N_28064,N_29020);
xnor UO_3247 (O_3247,N_28488,N_29546);
nand UO_3248 (O_3248,N_28286,N_28363);
nor UO_3249 (O_3249,N_28989,N_29401);
nand UO_3250 (O_3250,N_29126,N_28213);
or UO_3251 (O_3251,N_29412,N_29821);
or UO_3252 (O_3252,N_28694,N_28035);
nor UO_3253 (O_3253,N_29730,N_29208);
and UO_3254 (O_3254,N_28637,N_28426);
or UO_3255 (O_3255,N_29926,N_28119);
and UO_3256 (O_3256,N_29673,N_29325);
and UO_3257 (O_3257,N_28062,N_29356);
xor UO_3258 (O_3258,N_28228,N_29525);
nand UO_3259 (O_3259,N_29531,N_29714);
xnor UO_3260 (O_3260,N_29848,N_29910);
nor UO_3261 (O_3261,N_29616,N_28695);
or UO_3262 (O_3262,N_28622,N_29114);
nand UO_3263 (O_3263,N_28766,N_29261);
nor UO_3264 (O_3264,N_28646,N_29898);
or UO_3265 (O_3265,N_28200,N_28315);
nor UO_3266 (O_3266,N_29707,N_29854);
xnor UO_3267 (O_3267,N_28885,N_28047);
and UO_3268 (O_3268,N_28654,N_29208);
and UO_3269 (O_3269,N_28658,N_28051);
and UO_3270 (O_3270,N_29376,N_29432);
xor UO_3271 (O_3271,N_29831,N_29501);
and UO_3272 (O_3272,N_29530,N_29897);
nand UO_3273 (O_3273,N_28929,N_29348);
nand UO_3274 (O_3274,N_28227,N_29883);
or UO_3275 (O_3275,N_28347,N_28837);
and UO_3276 (O_3276,N_28531,N_29234);
and UO_3277 (O_3277,N_29513,N_28632);
xor UO_3278 (O_3278,N_29435,N_29347);
or UO_3279 (O_3279,N_29638,N_28859);
nand UO_3280 (O_3280,N_29240,N_28354);
and UO_3281 (O_3281,N_28062,N_28552);
xnor UO_3282 (O_3282,N_28557,N_28511);
or UO_3283 (O_3283,N_29948,N_29830);
or UO_3284 (O_3284,N_29914,N_29144);
and UO_3285 (O_3285,N_28843,N_28249);
xor UO_3286 (O_3286,N_28562,N_29924);
nor UO_3287 (O_3287,N_28685,N_29016);
and UO_3288 (O_3288,N_28704,N_29715);
and UO_3289 (O_3289,N_28545,N_29188);
or UO_3290 (O_3290,N_29387,N_28257);
xnor UO_3291 (O_3291,N_28801,N_28370);
nor UO_3292 (O_3292,N_29827,N_29336);
xnor UO_3293 (O_3293,N_29447,N_29298);
or UO_3294 (O_3294,N_28725,N_28166);
nor UO_3295 (O_3295,N_28240,N_28575);
nor UO_3296 (O_3296,N_28870,N_29134);
and UO_3297 (O_3297,N_28784,N_28785);
nand UO_3298 (O_3298,N_29726,N_28316);
and UO_3299 (O_3299,N_29103,N_28958);
nor UO_3300 (O_3300,N_29448,N_29713);
nand UO_3301 (O_3301,N_28502,N_28604);
nor UO_3302 (O_3302,N_29562,N_29351);
nand UO_3303 (O_3303,N_29129,N_28831);
nor UO_3304 (O_3304,N_29175,N_29749);
or UO_3305 (O_3305,N_28502,N_29105);
or UO_3306 (O_3306,N_28528,N_28714);
nand UO_3307 (O_3307,N_29866,N_29344);
nor UO_3308 (O_3308,N_29065,N_28438);
nor UO_3309 (O_3309,N_29961,N_28914);
and UO_3310 (O_3310,N_28009,N_29745);
xor UO_3311 (O_3311,N_28099,N_29783);
xnor UO_3312 (O_3312,N_29662,N_28450);
and UO_3313 (O_3313,N_28352,N_28032);
xor UO_3314 (O_3314,N_28586,N_29163);
and UO_3315 (O_3315,N_28494,N_28915);
nor UO_3316 (O_3316,N_28913,N_29464);
nand UO_3317 (O_3317,N_29087,N_29986);
and UO_3318 (O_3318,N_29735,N_29193);
xnor UO_3319 (O_3319,N_28029,N_29294);
xnor UO_3320 (O_3320,N_28586,N_28176);
nor UO_3321 (O_3321,N_28468,N_29328);
xor UO_3322 (O_3322,N_28194,N_29942);
nor UO_3323 (O_3323,N_28118,N_29286);
nand UO_3324 (O_3324,N_29558,N_28841);
nand UO_3325 (O_3325,N_29894,N_28468);
xnor UO_3326 (O_3326,N_28107,N_28229);
xor UO_3327 (O_3327,N_28688,N_29856);
nand UO_3328 (O_3328,N_29682,N_28986);
xor UO_3329 (O_3329,N_28144,N_29990);
or UO_3330 (O_3330,N_28197,N_28858);
nand UO_3331 (O_3331,N_28544,N_29653);
nand UO_3332 (O_3332,N_28636,N_28737);
xor UO_3333 (O_3333,N_28120,N_28303);
and UO_3334 (O_3334,N_29238,N_28161);
nor UO_3335 (O_3335,N_29398,N_29342);
and UO_3336 (O_3336,N_28118,N_29250);
or UO_3337 (O_3337,N_29716,N_29124);
or UO_3338 (O_3338,N_29072,N_29272);
nor UO_3339 (O_3339,N_28290,N_28494);
nand UO_3340 (O_3340,N_29882,N_29266);
or UO_3341 (O_3341,N_29201,N_29177);
or UO_3342 (O_3342,N_29559,N_29291);
xnor UO_3343 (O_3343,N_28900,N_29793);
nor UO_3344 (O_3344,N_28397,N_29663);
nor UO_3345 (O_3345,N_29756,N_28764);
and UO_3346 (O_3346,N_28338,N_29992);
and UO_3347 (O_3347,N_29286,N_28238);
and UO_3348 (O_3348,N_29946,N_28570);
xnor UO_3349 (O_3349,N_28276,N_28911);
and UO_3350 (O_3350,N_28058,N_28907);
nand UO_3351 (O_3351,N_29047,N_29692);
nor UO_3352 (O_3352,N_28338,N_29321);
xor UO_3353 (O_3353,N_29763,N_29263);
and UO_3354 (O_3354,N_29444,N_29253);
nand UO_3355 (O_3355,N_28290,N_28502);
and UO_3356 (O_3356,N_29383,N_28656);
nand UO_3357 (O_3357,N_29346,N_28075);
and UO_3358 (O_3358,N_28200,N_28864);
and UO_3359 (O_3359,N_28310,N_28763);
and UO_3360 (O_3360,N_29621,N_29781);
xnor UO_3361 (O_3361,N_28278,N_28579);
or UO_3362 (O_3362,N_29279,N_29911);
nor UO_3363 (O_3363,N_28026,N_29078);
and UO_3364 (O_3364,N_28739,N_29068);
or UO_3365 (O_3365,N_28021,N_28027);
or UO_3366 (O_3366,N_29527,N_28176);
or UO_3367 (O_3367,N_28508,N_29294);
nand UO_3368 (O_3368,N_28606,N_28264);
nor UO_3369 (O_3369,N_29157,N_28254);
nand UO_3370 (O_3370,N_28420,N_28784);
nand UO_3371 (O_3371,N_29428,N_29345);
nor UO_3372 (O_3372,N_28262,N_28194);
and UO_3373 (O_3373,N_28142,N_29294);
or UO_3374 (O_3374,N_28672,N_29578);
and UO_3375 (O_3375,N_28575,N_28173);
xnor UO_3376 (O_3376,N_29685,N_29160);
and UO_3377 (O_3377,N_29010,N_29006);
and UO_3378 (O_3378,N_29656,N_29593);
xnor UO_3379 (O_3379,N_29371,N_29376);
nand UO_3380 (O_3380,N_28291,N_28769);
or UO_3381 (O_3381,N_28298,N_29888);
nand UO_3382 (O_3382,N_28885,N_29465);
nand UO_3383 (O_3383,N_28672,N_29060);
xor UO_3384 (O_3384,N_29954,N_28669);
nand UO_3385 (O_3385,N_28527,N_29780);
nor UO_3386 (O_3386,N_29271,N_28557);
nand UO_3387 (O_3387,N_28654,N_28640);
xor UO_3388 (O_3388,N_29961,N_29729);
and UO_3389 (O_3389,N_28455,N_28576);
or UO_3390 (O_3390,N_28301,N_28748);
and UO_3391 (O_3391,N_28054,N_29660);
and UO_3392 (O_3392,N_29922,N_29492);
nand UO_3393 (O_3393,N_29928,N_29172);
nand UO_3394 (O_3394,N_29647,N_28475);
and UO_3395 (O_3395,N_29111,N_29574);
or UO_3396 (O_3396,N_29931,N_28387);
xor UO_3397 (O_3397,N_29553,N_28021);
or UO_3398 (O_3398,N_29687,N_28389);
nor UO_3399 (O_3399,N_28110,N_28046);
nand UO_3400 (O_3400,N_28436,N_29368);
and UO_3401 (O_3401,N_28416,N_29709);
nand UO_3402 (O_3402,N_29172,N_28219);
nand UO_3403 (O_3403,N_29052,N_29339);
and UO_3404 (O_3404,N_29406,N_28691);
nor UO_3405 (O_3405,N_29576,N_29850);
xor UO_3406 (O_3406,N_29174,N_28606);
nor UO_3407 (O_3407,N_29759,N_29774);
nor UO_3408 (O_3408,N_29489,N_28654);
nand UO_3409 (O_3409,N_29600,N_28111);
nor UO_3410 (O_3410,N_28432,N_29690);
nor UO_3411 (O_3411,N_29808,N_29085);
xnor UO_3412 (O_3412,N_29957,N_28078);
xor UO_3413 (O_3413,N_29915,N_29115);
nand UO_3414 (O_3414,N_29405,N_28706);
xor UO_3415 (O_3415,N_28447,N_29226);
or UO_3416 (O_3416,N_29965,N_29418);
nor UO_3417 (O_3417,N_28370,N_29515);
nand UO_3418 (O_3418,N_28983,N_29834);
xnor UO_3419 (O_3419,N_28095,N_28160);
and UO_3420 (O_3420,N_28164,N_28400);
nor UO_3421 (O_3421,N_29154,N_29564);
or UO_3422 (O_3422,N_28297,N_29422);
and UO_3423 (O_3423,N_28024,N_29326);
xnor UO_3424 (O_3424,N_29514,N_28220);
or UO_3425 (O_3425,N_28844,N_29064);
nor UO_3426 (O_3426,N_28950,N_29750);
xnor UO_3427 (O_3427,N_29839,N_29668);
nor UO_3428 (O_3428,N_28922,N_29740);
and UO_3429 (O_3429,N_29020,N_29657);
or UO_3430 (O_3430,N_29922,N_28043);
nor UO_3431 (O_3431,N_29142,N_29583);
or UO_3432 (O_3432,N_29095,N_29439);
nor UO_3433 (O_3433,N_28628,N_29907);
nor UO_3434 (O_3434,N_29721,N_29457);
nor UO_3435 (O_3435,N_29367,N_29338);
nand UO_3436 (O_3436,N_28169,N_29165);
or UO_3437 (O_3437,N_29983,N_29823);
and UO_3438 (O_3438,N_28736,N_28607);
and UO_3439 (O_3439,N_28379,N_29217);
nand UO_3440 (O_3440,N_28517,N_29777);
or UO_3441 (O_3441,N_29650,N_29178);
or UO_3442 (O_3442,N_28900,N_28274);
xnor UO_3443 (O_3443,N_28952,N_28418);
nand UO_3444 (O_3444,N_28815,N_29322);
or UO_3445 (O_3445,N_29410,N_29760);
xnor UO_3446 (O_3446,N_29587,N_29224);
xor UO_3447 (O_3447,N_28269,N_28139);
nor UO_3448 (O_3448,N_29121,N_29334);
or UO_3449 (O_3449,N_28361,N_28745);
and UO_3450 (O_3450,N_28543,N_28085);
and UO_3451 (O_3451,N_29607,N_29046);
xor UO_3452 (O_3452,N_29516,N_29888);
and UO_3453 (O_3453,N_28428,N_28321);
nor UO_3454 (O_3454,N_28841,N_29757);
and UO_3455 (O_3455,N_28830,N_29518);
nand UO_3456 (O_3456,N_29764,N_28221);
nand UO_3457 (O_3457,N_28448,N_28092);
and UO_3458 (O_3458,N_29876,N_29684);
nor UO_3459 (O_3459,N_28155,N_28597);
xnor UO_3460 (O_3460,N_29161,N_28208);
nand UO_3461 (O_3461,N_28498,N_28035);
xor UO_3462 (O_3462,N_29611,N_29621);
or UO_3463 (O_3463,N_28987,N_28233);
or UO_3464 (O_3464,N_29545,N_29200);
nand UO_3465 (O_3465,N_29087,N_28133);
xor UO_3466 (O_3466,N_28945,N_28191);
or UO_3467 (O_3467,N_28580,N_29741);
and UO_3468 (O_3468,N_29718,N_29819);
nor UO_3469 (O_3469,N_28971,N_29994);
or UO_3470 (O_3470,N_29615,N_29017);
and UO_3471 (O_3471,N_29860,N_29999);
nand UO_3472 (O_3472,N_28802,N_28418);
or UO_3473 (O_3473,N_28864,N_28749);
nand UO_3474 (O_3474,N_28530,N_28510);
or UO_3475 (O_3475,N_29779,N_28989);
and UO_3476 (O_3476,N_28720,N_28175);
xor UO_3477 (O_3477,N_28075,N_29555);
or UO_3478 (O_3478,N_28857,N_29564);
and UO_3479 (O_3479,N_29728,N_29252);
nor UO_3480 (O_3480,N_28749,N_29576);
nor UO_3481 (O_3481,N_29205,N_28454);
and UO_3482 (O_3482,N_28151,N_29142);
nor UO_3483 (O_3483,N_29841,N_28728);
nor UO_3484 (O_3484,N_28580,N_29181);
nand UO_3485 (O_3485,N_28140,N_29226);
or UO_3486 (O_3486,N_28178,N_29603);
nor UO_3487 (O_3487,N_28877,N_29647);
and UO_3488 (O_3488,N_29435,N_28261);
and UO_3489 (O_3489,N_29560,N_29853);
nand UO_3490 (O_3490,N_28859,N_29323);
and UO_3491 (O_3491,N_29880,N_29804);
or UO_3492 (O_3492,N_29100,N_28311);
and UO_3493 (O_3493,N_29147,N_29924);
nand UO_3494 (O_3494,N_28669,N_28567);
nor UO_3495 (O_3495,N_29106,N_28188);
xnor UO_3496 (O_3496,N_29912,N_28180);
nand UO_3497 (O_3497,N_29727,N_28292);
and UO_3498 (O_3498,N_28852,N_29092);
nand UO_3499 (O_3499,N_29178,N_28122);
endmodule