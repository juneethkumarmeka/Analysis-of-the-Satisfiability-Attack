module basic_1000_10000_1500_10_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_624,In_458);
and U1 (N_1,In_536,In_745);
and U2 (N_2,In_617,In_658);
nand U3 (N_3,In_893,In_453);
nor U4 (N_4,In_887,In_852);
nand U5 (N_5,In_335,In_396);
nor U6 (N_6,In_25,In_984);
nor U7 (N_7,In_585,In_939);
and U8 (N_8,In_107,In_651);
or U9 (N_9,In_549,In_227);
nand U10 (N_10,In_293,In_460);
or U11 (N_11,In_730,In_118);
and U12 (N_12,In_388,In_265);
nor U13 (N_13,In_260,In_389);
or U14 (N_14,In_591,In_773);
and U15 (N_15,In_85,In_18);
nor U16 (N_16,In_59,In_461);
nand U17 (N_17,In_73,In_271);
and U18 (N_18,In_646,In_524);
nand U19 (N_19,In_661,In_614);
nand U20 (N_20,In_662,In_900);
nor U21 (N_21,In_580,In_343);
nor U22 (N_22,In_578,In_344);
and U23 (N_23,In_256,In_161);
nand U24 (N_24,In_503,In_204);
nor U25 (N_25,In_245,In_237);
xnor U26 (N_26,In_55,In_378);
or U27 (N_27,In_990,In_569);
and U28 (N_28,In_598,In_75);
xnor U29 (N_29,In_270,In_123);
or U30 (N_30,In_373,In_427);
nand U31 (N_31,In_716,In_446);
and U32 (N_32,In_249,In_201);
nand U33 (N_33,In_821,In_493);
nand U34 (N_34,In_57,In_626);
nor U35 (N_35,In_680,In_240);
or U36 (N_36,In_760,In_211);
and U37 (N_37,In_183,In_637);
or U38 (N_38,In_202,In_106);
or U39 (N_39,In_142,In_21);
or U40 (N_40,In_842,In_883);
and U41 (N_41,In_197,In_307);
nor U42 (N_42,In_330,In_896);
nand U43 (N_43,In_456,In_496);
nor U44 (N_44,In_704,In_384);
or U45 (N_45,In_792,In_944);
or U46 (N_46,In_380,In_922);
and U47 (N_47,In_188,In_250);
or U48 (N_48,In_949,In_766);
nand U49 (N_49,In_403,In_826);
and U50 (N_50,In_191,In_746);
or U51 (N_51,In_119,In_909);
nor U52 (N_52,In_606,In_234);
or U53 (N_53,In_868,In_394);
nand U54 (N_54,In_988,In_339);
or U55 (N_55,In_708,In_914);
and U56 (N_56,In_799,In_4);
nand U57 (N_57,In_855,In_608);
nor U58 (N_58,In_711,In_807);
nand U59 (N_59,In_565,In_630);
or U60 (N_60,In_919,In_80);
nand U61 (N_61,In_400,In_395);
nor U62 (N_62,In_146,In_751);
nand U63 (N_63,In_596,In_438);
or U64 (N_64,In_647,In_114);
and U65 (N_65,In_952,In_487);
and U66 (N_66,In_7,In_537);
nand U67 (N_67,In_153,In_720);
nand U68 (N_68,In_528,In_797);
nor U69 (N_69,In_193,In_212);
nand U70 (N_70,In_444,In_800);
nor U71 (N_71,In_15,In_513);
nor U72 (N_72,In_361,In_758);
and U73 (N_73,In_87,In_172);
and U74 (N_74,In_543,In_712);
nor U75 (N_75,In_982,In_482);
or U76 (N_76,In_89,In_466);
nand U77 (N_77,In_672,In_124);
nor U78 (N_78,In_295,In_121);
nor U79 (N_79,In_276,In_872);
and U80 (N_80,In_207,In_638);
nand U81 (N_81,In_586,In_471);
or U82 (N_82,In_304,In_835);
nand U83 (N_83,In_701,In_786);
or U84 (N_84,In_404,In_383);
nand U85 (N_85,In_457,In_664);
xor U86 (N_86,In_554,In_744);
nand U87 (N_87,In_429,In_2);
nor U88 (N_88,In_721,In_734);
nor U89 (N_89,In_911,In_521);
xnor U90 (N_90,In_441,In_527);
nand U91 (N_91,In_523,In_477);
and U92 (N_92,In_686,In_607);
or U93 (N_93,In_534,In_152);
xnor U94 (N_94,In_406,In_26);
or U95 (N_95,In_597,In_130);
nor U96 (N_96,In_350,In_185);
nor U97 (N_97,In_874,In_722);
or U98 (N_98,In_653,In_829);
nand U99 (N_99,In_309,In_865);
and U100 (N_100,In_961,In_88);
and U101 (N_101,In_138,In_115);
and U102 (N_102,In_987,In_362);
nand U103 (N_103,In_31,In_345);
nor U104 (N_104,In_945,In_723);
or U105 (N_105,In_951,In_184);
and U106 (N_106,In_558,In_878);
nor U107 (N_107,In_219,In_353);
and U108 (N_108,In_377,In_439);
or U109 (N_109,In_289,In_168);
nor U110 (N_110,In_871,In_62);
or U111 (N_111,In_431,In_510);
xor U112 (N_112,In_450,In_684);
and U113 (N_113,In_870,In_160);
and U114 (N_114,In_217,In_315);
or U115 (N_115,In_666,In_690);
nor U116 (N_116,In_538,In_170);
nor U117 (N_117,In_135,In_332);
nor U118 (N_118,In_425,In_508);
or U119 (N_119,In_100,In_673);
nor U120 (N_120,In_742,In_419);
nor U121 (N_121,In_678,In_82);
or U122 (N_122,In_341,In_516);
nand U123 (N_123,In_418,In_703);
and U124 (N_124,In_539,In_297);
or U125 (N_125,In_314,In_137);
or U126 (N_126,In_851,In_925);
or U127 (N_127,In_519,In_0);
and U128 (N_128,In_622,In_834);
and U129 (N_129,In_950,In_53);
nor U130 (N_130,In_175,In_422);
or U131 (N_131,In_485,In_469);
nand U132 (N_132,In_136,In_99);
and U133 (N_133,In_975,In_858);
nand U134 (N_134,In_426,In_13);
or U135 (N_135,In_974,In_648);
nor U136 (N_136,In_958,In_301);
nand U137 (N_137,In_902,In_1);
xor U138 (N_138,In_897,In_410);
and U139 (N_139,In_447,In_837);
nand U140 (N_140,In_72,In_986);
or U141 (N_141,In_873,In_58);
or U142 (N_142,In_924,In_507);
xor U143 (N_143,In_640,In_236);
nor U144 (N_144,In_903,In_102);
nand U145 (N_145,In_134,In_215);
and U146 (N_146,In_994,In_143);
nor U147 (N_147,In_767,In_601);
or U148 (N_148,In_724,In_805);
nor U149 (N_149,In_81,In_557);
nor U150 (N_150,In_368,In_583);
or U151 (N_151,In_973,In_398);
nand U152 (N_152,In_451,In_252);
nor U153 (N_153,In_750,In_509);
or U154 (N_154,In_150,In_908);
and U155 (N_155,In_28,In_23);
and U156 (N_156,In_41,In_79);
nand U157 (N_157,In_32,In_983);
nand U158 (N_158,In_719,In_752);
nand U159 (N_159,In_228,In_970);
or U160 (N_160,In_687,In_194);
and U161 (N_161,In_242,In_525);
nor U162 (N_162,In_162,In_199);
and U163 (N_163,In_27,In_595);
nor U164 (N_164,In_259,In_869);
or U165 (N_165,In_235,In_111);
or U166 (N_166,In_544,In_39);
and U167 (N_167,In_402,In_880);
xnor U168 (N_168,In_346,In_784);
nand U169 (N_169,In_247,In_104);
nor U170 (N_170,In_101,In_37);
and U171 (N_171,In_670,In_824);
nand U172 (N_172,In_381,In_713);
and U173 (N_173,In_693,In_47);
or U174 (N_174,In_652,In_348);
or U175 (N_175,In_480,In_189);
and U176 (N_176,In_502,In_229);
or U177 (N_177,In_738,In_725);
and U178 (N_178,In_290,In_809);
or U179 (N_179,In_782,In_299);
nand U180 (N_180,In_553,In_291);
and U181 (N_181,In_220,In_501);
nand U182 (N_182,In_483,In_167);
nor U183 (N_183,In_899,In_552);
xnor U184 (N_184,In_603,In_531);
or U185 (N_185,In_24,In_840);
nand U186 (N_186,In_506,In_756);
or U187 (N_187,In_650,In_127);
or U188 (N_188,In_743,In_582);
nor U189 (N_189,In_891,In_495);
xnor U190 (N_190,In_803,In_709);
or U191 (N_191,In_955,In_665);
nand U192 (N_192,In_688,In_882);
or U193 (N_193,In_649,In_187);
and U194 (N_194,In_845,In_52);
xor U195 (N_195,In_546,In_755);
nand U196 (N_196,In_435,In_86);
and U197 (N_197,In_946,In_915);
nor U198 (N_198,In_997,In_927);
nor U199 (N_199,In_407,In_541);
and U200 (N_200,In_611,In_555);
and U201 (N_201,In_841,In_556);
and U202 (N_202,In_238,In_904);
or U203 (N_203,In_963,In_359);
nor U204 (N_204,In_338,In_604);
nand U205 (N_205,In_620,In_486);
and U206 (N_206,In_937,In_414);
nand U207 (N_207,In_46,In_186);
and U208 (N_208,In_989,In_551);
nor U209 (N_209,In_639,In_22);
nand U210 (N_210,In_679,In_205);
or U211 (N_211,In_685,In_329);
or U212 (N_212,In_529,In_996);
and U213 (N_213,In_497,In_642);
nand U214 (N_214,In_374,In_462);
or U215 (N_215,In_491,In_190);
nand U216 (N_216,In_780,In_563);
nand U217 (N_217,In_500,In_935);
or U218 (N_218,In_791,In_218);
and U219 (N_219,In_843,In_328);
xnor U220 (N_220,In_629,In_365);
nor U221 (N_221,In_820,In_459);
nor U222 (N_222,In_264,In_567);
nand U223 (N_223,In_960,In_93);
or U224 (N_224,In_154,In_736);
or U225 (N_225,In_609,In_408);
nor U226 (N_226,In_68,In_584);
nand U227 (N_227,In_375,In_993);
xor U228 (N_228,In_333,In_610);
or U229 (N_229,In_676,In_279);
or U230 (N_230,In_17,In_827);
nand U231 (N_231,In_443,In_321);
nand U232 (N_232,In_494,In_209);
or U233 (N_233,In_258,In_163);
nand U234 (N_234,In_540,In_397);
and U235 (N_235,In_222,In_412);
or U236 (N_236,In_421,In_886);
and U237 (N_237,In_367,In_139);
nor U238 (N_238,In_895,In_644);
and U239 (N_239,In_737,In_933);
nand U240 (N_240,In_566,In_174);
and U241 (N_241,In_434,In_273);
or U242 (N_242,In_342,In_463);
nand U243 (N_243,In_112,In_748);
and U244 (N_244,In_790,In_850);
or U245 (N_245,In_633,In_63);
and U246 (N_246,In_305,In_56);
nor U247 (N_247,In_173,In_940);
nand U248 (N_248,In_726,In_436);
nand U249 (N_249,In_262,In_581);
nand U250 (N_250,In_200,In_787);
or U251 (N_251,In_511,In_371);
nand U252 (N_252,In_96,In_717);
nand U253 (N_253,In_832,In_122);
and U254 (N_254,In_753,In_117);
and U255 (N_255,In_43,In_409);
nand U256 (N_256,In_277,In_269);
or U257 (N_257,In_147,In_317);
or U258 (N_258,In_979,In_731);
or U259 (N_259,In_433,In_817);
and U260 (N_260,In_244,In_966);
or U261 (N_261,In_968,In_454);
nand U262 (N_262,In_517,In_828);
nand U263 (N_263,In_798,In_856);
or U264 (N_264,In_390,In_464);
or U265 (N_265,In_941,In_133);
xor U266 (N_266,In_452,In_991);
and U267 (N_267,In_533,In_683);
nor U268 (N_268,In_593,In_877);
or U269 (N_269,In_449,In_921);
nand U270 (N_270,In_929,In_702);
or U271 (N_271,In_707,In_785);
and U272 (N_272,In_38,In_19);
and U273 (N_273,In_54,In_326);
nor U274 (N_274,In_579,In_232);
nand U275 (N_275,In_733,In_814);
and U276 (N_276,In_420,In_283);
nand U277 (N_277,In_674,In_774);
nand U278 (N_278,In_77,In_8);
and U279 (N_279,In_303,In_148);
and U280 (N_280,In_165,In_74);
nor U281 (N_281,In_61,In_490);
nand U282 (N_282,In_621,In_777);
nor U283 (N_283,In_816,In_934);
nand U284 (N_284,In_947,In_386);
and U285 (N_285,In_370,In_10);
nand U286 (N_286,In_178,In_867);
nor U287 (N_287,In_357,In_718);
xnor U288 (N_288,In_729,In_387);
and U289 (N_289,In_340,In_772);
nor U290 (N_290,In_324,In_655);
and U291 (N_291,In_66,In_978);
or U292 (N_292,In_254,In_831);
nor U293 (N_293,In_623,In_660);
nor U294 (N_294,In_864,In_512);
nand U295 (N_295,In_128,In_715);
nand U296 (N_296,In_892,In_60);
and U297 (N_297,In_612,In_920);
xnor U298 (N_298,In_196,In_455);
or U299 (N_299,In_468,In_268);
or U300 (N_300,In_592,In_802);
and U301 (N_301,In_475,In_67);
nor U302 (N_302,In_225,In_956);
nor U303 (N_303,In_931,In_284);
and U304 (N_304,In_696,In_881);
and U305 (N_305,In_795,In_263);
nor U306 (N_306,In_42,In_972);
nor U307 (N_307,In_337,In_589);
and U308 (N_308,In_92,In_568);
and U309 (N_309,In_530,In_839);
or U310 (N_310,In_577,In_51);
nand U311 (N_311,In_532,In_659);
and U312 (N_312,In_794,In_778);
nor U313 (N_313,In_964,In_876);
and U314 (N_314,In_518,In_311);
or U315 (N_315,In_405,In_239);
nor U316 (N_316,In_616,In_628);
nor U317 (N_317,In_962,In_515);
and U318 (N_318,In_999,In_815);
nor U319 (N_319,In_765,In_559);
nor U320 (N_320,In_282,In_923);
or U321 (N_321,In_417,In_64);
xor U322 (N_322,In_657,In_274);
and U323 (N_323,In_12,In_120);
or U324 (N_324,In_411,In_894);
nor U325 (N_325,In_29,In_230);
or U326 (N_326,In_48,In_995);
nor U327 (N_327,In_912,In_266);
nor U328 (N_328,In_484,In_833);
nor U329 (N_329,In_587,In_706);
or U330 (N_330,In_36,In_600);
or U331 (N_331,In_334,In_627);
or U332 (N_332,In_985,In_11);
and U333 (N_333,In_980,In_618);
or U334 (N_334,In_822,In_306);
nor U335 (N_335,In_84,In_705);
nor U336 (N_336,In_393,In_906);
and U337 (N_337,In_967,In_499);
nor U338 (N_338,In_879,In_50);
nand U339 (N_339,In_20,In_632);
nor U340 (N_340,In_913,In_572);
and U341 (N_341,In_331,In_322);
and U342 (N_342,In_938,In_957);
and U343 (N_343,In_861,In_221);
or U344 (N_344,In_599,In_885);
nand U345 (N_345,In_695,In_192);
nor U346 (N_346,In_233,In_261);
nand U347 (N_347,In_602,In_129);
and U348 (N_348,In_166,In_930);
nor U349 (N_349,In_203,In_16);
and U350 (N_350,In_369,In_520);
nor U351 (N_351,In_916,In_489);
nand U352 (N_352,In_472,In_49);
nand U353 (N_353,In_789,In_294);
nor U354 (N_354,In_976,In_643);
nand U355 (N_355,In_700,In_936);
nor U356 (N_356,In_34,In_171);
nand U357 (N_357,In_116,In_108);
and U358 (N_358,In_35,In_248);
or U359 (N_359,In_257,In_849);
or U360 (N_360,In_594,In_157);
nand U361 (N_361,In_465,In_70);
or U362 (N_362,In_208,In_176);
and U363 (N_363,In_575,In_360);
and U364 (N_364,In_327,In_764);
or U365 (N_365,In_347,In_698);
nand U366 (N_366,In_846,In_522);
and U367 (N_367,In_308,In_363);
and U368 (N_368,In_625,In_103);
and U369 (N_369,In_195,In_689);
nand U370 (N_370,In_866,In_747);
nor U371 (N_371,In_884,In_198);
nor U372 (N_372,In_739,In_862);
nand U373 (N_373,In_918,In_574);
and U374 (N_374,In_440,In_180);
xor U375 (N_375,In_366,In_83);
nand U376 (N_376,In_351,In_992);
nand U377 (N_377,In_998,In_6);
nand U378 (N_378,In_78,In_488);
nand U379 (N_379,In_216,In_292);
nand U380 (N_380,In_818,In_391);
or U381 (N_381,In_65,In_355);
nor U382 (N_382,In_354,In_844);
xor U383 (N_383,In_573,In_323);
and U384 (N_384,In_231,In_741);
and U385 (N_385,In_109,In_863);
nand U386 (N_386,In_562,In_156);
nand U387 (N_387,In_898,In_164);
and U388 (N_388,In_761,In_954);
nor U389 (N_389,In_3,In_470);
nor U390 (N_390,In_645,In_131);
nor U391 (N_391,In_71,In_910);
and U392 (N_392,In_663,In_560);
and U393 (N_393,In_793,In_675);
and U394 (N_394,In_727,In_430);
nand U395 (N_395,In_770,In_888);
nor U396 (N_396,In_325,In_179);
and U397 (N_397,In_771,In_182);
nand U398 (N_398,In_810,In_498);
nand U399 (N_399,In_977,In_9);
nor U400 (N_400,In_825,In_382);
nand U401 (N_401,In_779,In_634);
and U402 (N_402,In_467,In_281);
or U403 (N_403,In_481,In_423);
and U404 (N_404,In_125,In_413);
or U405 (N_405,In_631,In_953);
nand U406 (N_406,In_571,In_749);
and U407 (N_407,In_206,In_775);
and U408 (N_408,In_514,In_668);
or U409 (N_409,In_588,In_932);
nand U410 (N_410,In_267,In_319);
and U411 (N_411,In_728,In_853);
and U412 (N_412,In_769,In_788);
nor U413 (N_413,In_547,In_302);
nor U414 (N_414,In_300,In_768);
nand U415 (N_415,In_246,In_545);
nor U416 (N_416,In_619,In_5);
nand U417 (N_417,In_95,In_358);
or U418 (N_418,In_442,In_364);
nand U419 (N_419,In_223,In_318);
or U420 (N_420,In_14,In_90);
and U421 (N_421,In_310,In_275);
or U422 (N_422,In_437,In_492);
nor U423 (N_423,In_313,In_969);
nor U424 (N_424,In_372,In_697);
nor U425 (N_425,In_590,In_399);
and U426 (N_426,In_812,In_349);
and U427 (N_427,In_759,In_505);
or U428 (N_428,In_45,In_177);
or U429 (N_429,In_356,In_401);
nand U430 (N_430,In_682,In_917);
nor U431 (N_431,In_213,In_763);
or U432 (N_432,In_416,In_905);
nor U433 (N_433,In_141,In_875);
nand U434 (N_434,In_819,In_943);
nor U435 (N_435,In_285,In_635);
or U436 (N_436,In_243,In_928);
nand U437 (N_437,In_241,In_615);
and U438 (N_438,In_226,In_811);
or U439 (N_439,In_838,In_76);
and U440 (N_440,In_570,In_714);
and U441 (N_441,In_847,In_526);
and U442 (N_442,In_801,In_432);
xnor U443 (N_443,In_255,In_140);
and U444 (N_444,In_474,In_40);
and U445 (N_445,In_113,In_479);
and U446 (N_446,In_691,In_796);
nand U447 (N_447,In_576,In_613);
or U448 (N_448,In_251,In_144);
and U449 (N_449,In_859,In_287);
nor U450 (N_450,In_30,In_836);
nand U451 (N_451,In_681,In_735);
nand U452 (N_452,In_890,In_278);
or U453 (N_453,In_316,In_667);
or U454 (N_454,In_699,In_654);
and U455 (N_455,In_776,In_854);
or U456 (N_456,In_889,In_352);
or U457 (N_457,In_110,In_948);
and U458 (N_458,In_415,In_145);
nand U459 (N_459,In_677,In_379);
nand U460 (N_460,In_542,In_907);
nand U461 (N_461,In_224,In_105);
nor U462 (N_462,In_808,In_385);
or U463 (N_463,In_312,In_320);
nor U464 (N_464,In_830,In_149);
nor U465 (N_465,In_69,In_860);
xnor U466 (N_466,In_669,In_561);
nor U467 (N_467,In_424,In_159);
nand U468 (N_468,In_813,In_169);
nor U469 (N_469,In_965,In_762);
nand U470 (N_470,In_94,In_781);
nand U471 (N_471,In_641,In_298);
and U472 (N_472,In_288,In_97);
or U473 (N_473,In_126,In_376);
and U474 (N_474,In_981,In_710);
nand U475 (N_475,In_296,In_478);
and U476 (N_476,In_806,In_91);
and U477 (N_477,In_392,In_942);
or U478 (N_478,In_694,In_286);
or U479 (N_479,In_732,In_857);
or U480 (N_480,In_636,In_473);
nor U481 (N_481,In_44,In_656);
nor U482 (N_482,In_132,In_550);
and U483 (N_483,In_504,In_210);
and U484 (N_484,In_98,In_155);
and U485 (N_485,In_971,In_445);
or U486 (N_486,In_564,In_428);
or U487 (N_487,In_823,In_214);
nor U488 (N_488,In_848,In_754);
and U489 (N_489,In_926,In_740);
nor U490 (N_490,In_692,In_605);
nor U491 (N_491,In_253,In_181);
nor U492 (N_492,In_448,In_959);
nor U493 (N_493,In_151,In_804);
and U494 (N_494,In_280,In_783);
nand U495 (N_495,In_671,In_901);
nor U496 (N_496,In_757,In_158);
nor U497 (N_497,In_476,In_33);
and U498 (N_498,In_548,In_272);
nor U499 (N_499,In_535,In_336);
nor U500 (N_500,In_828,In_949);
nand U501 (N_501,In_855,In_862);
and U502 (N_502,In_73,In_537);
and U503 (N_503,In_943,In_217);
or U504 (N_504,In_756,In_719);
and U505 (N_505,In_376,In_612);
nor U506 (N_506,In_881,In_289);
and U507 (N_507,In_546,In_465);
nand U508 (N_508,In_952,In_522);
and U509 (N_509,In_520,In_109);
nor U510 (N_510,In_501,In_603);
nor U511 (N_511,In_691,In_585);
nor U512 (N_512,In_144,In_130);
or U513 (N_513,In_165,In_420);
or U514 (N_514,In_528,In_869);
and U515 (N_515,In_841,In_963);
and U516 (N_516,In_458,In_527);
nor U517 (N_517,In_507,In_107);
nand U518 (N_518,In_292,In_614);
or U519 (N_519,In_265,In_242);
or U520 (N_520,In_532,In_937);
and U521 (N_521,In_757,In_498);
nor U522 (N_522,In_684,In_902);
nand U523 (N_523,In_890,In_434);
and U524 (N_524,In_694,In_293);
and U525 (N_525,In_990,In_979);
nor U526 (N_526,In_134,In_358);
nor U527 (N_527,In_412,In_475);
or U528 (N_528,In_976,In_967);
or U529 (N_529,In_179,In_938);
nand U530 (N_530,In_747,In_459);
nand U531 (N_531,In_903,In_145);
nand U532 (N_532,In_946,In_140);
and U533 (N_533,In_999,In_425);
or U534 (N_534,In_931,In_706);
nand U535 (N_535,In_885,In_24);
nand U536 (N_536,In_263,In_113);
and U537 (N_537,In_727,In_863);
nand U538 (N_538,In_734,In_807);
nand U539 (N_539,In_187,In_269);
nand U540 (N_540,In_774,In_183);
nor U541 (N_541,In_906,In_369);
nand U542 (N_542,In_140,In_597);
and U543 (N_543,In_601,In_765);
or U544 (N_544,In_295,In_278);
nand U545 (N_545,In_790,In_746);
nand U546 (N_546,In_519,In_174);
nor U547 (N_547,In_517,In_775);
and U548 (N_548,In_377,In_623);
nand U549 (N_549,In_413,In_802);
and U550 (N_550,In_63,In_574);
nand U551 (N_551,In_625,In_84);
or U552 (N_552,In_520,In_831);
nor U553 (N_553,In_474,In_434);
and U554 (N_554,In_260,In_285);
and U555 (N_555,In_610,In_128);
nor U556 (N_556,In_909,In_51);
nand U557 (N_557,In_789,In_609);
xor U558 (N_558,In_814,In_26);
nor U559 (N_559,In_304,In_823);
nand U560 (N_560,In_698,In_564);
and U561 (N_561,In_382,In_812);
xor U562 (N_562,In_594,In_811);
and U563 (N_563,In_586,In_998);
nand U564 (N_564,In_439,In_233);
nand U565 (N_565,In_959,In_165);
nand U566 (N_566,In_945,In_619);
or U567 (N_567,In_329,In_879);
and U568 (N_568,In_909,In_467);
and U569 (N_569,In_643,In_191);
and U570 (N_570,In_675,In_256);
nand U571 (N_571,In_606,In_153);
or U572 (N_572,In_861,In_343);
nor U573 (N_573,In_274,In_447);
nor U574 (N_574,In_275,In_527);
nor U575 (N_575,In_81,In_891);
nand U576 (N_576,In_421,In_265);
and U577 (N_577,In_485,In_462);
or U578 (N_578,In_60,In_181);
or U579 (N_579,In_858,In_621);
nor U580 (N_580,In_680,In_685);
nor U581 (N_581,In_596,In_126);
nand U582 (N_582,In_734,In_289);
and U583 (N_583,In_153,In_497);
and U584 (N_584,In_538,In_98);
nand U585 (N_585,In_914,In_267);
or U586 (N_586,In_459,In_119);
nor U587 (N_587,In_324,In_373);
nand U588 (N_588,In_691,In_276);
nor U589 (N_589,In_60,In_434);
and U590 (N_590,In_289,In_740);
nand U591 (N_591,In_115,In_928);
or U592 (N_592,In_663,In_882);
or U593 (N_593,In_930,In_38);
and U594 (N_594,In_2,In_979);
or U595 (N_595,In_205,In_549);
nand U596 (N_596,In_745,In_862);
nor U597 (N_597,In_647,In_515);
and U598 (N_598,In_537,In_798);
and U599 (N_599,In_585,In_174);
and U600 (N_600,In_102,In_660);
nor U601 (N_601,In_47,In_604);
nand U602 (N_602,In_288,In_616);
xor U603 (N_603,In_892,In_101);
nand U604 (N_604,In_150,In_588);
xor U605 (N_605,In_293,In_298);
nand U606 (N_606,In_931,In_66);
or U607 (N_607,In_532,In_23);
nor U608 (N_608,In_774,In_293);
nand U609 (N_609,In_385,In_321);
nand U610 (N_610,In_283,In_61);
and U611 (N_611,In_992,In_240);
and U612 (N_612,In_154,In_638);
nor U613 (N_613,In_836,In_401);
or U614 (N_614,In_36,In_855);
nand U615 (N_615,In_424,In_75);
nor U616 (N_616,In_544,In_652);
nand U617 (N_617,In_591,In_901);
nand U618 (N_618,In_867,In_773);
nand U619 (N_619,In_617,In_759);
or U620 (N_620,In_3,In_995);
or U621 (N_621,In_690,In_963);
and U622 (N_622,In_372,In_101);
and U623 (N_623,In_625,In_593);
nand U624 (N_624,In_399,In_568);
nand U625 (N_625,In_627,In_335);
nand U626 (N_626,In_226,In_903);
nor U627 (N_627,In_444,In_185);
or U628 (N_628,In_402,In_705);
nand U629 (N_629,In_472,In_142);
or U630 (N_630,In_547,In_430);
xor U631 (N_631,In_390,In_753);
nand U632 (N_632,In_367,In_178);
and U633 (N_633,In_825,In_774);
nor U634 (N_634,In_499,In_674);
nand U635 (N_635,In_97,In_820);
nand U636 (N_636,In_686,In_401);
and U637 (N_637,In_220,In_936);
or U638 (N_638,In_874,In_131);
and U639 (N_639,In_591,In_483);
xor U640 (N_640,In_707,In_425);
or U641 (N_641,In_72,In_50);
nor U642 (N_642,In_525,In_207);
and U643 (N_643,In_540,In_750);
and U644 (N_644,In_90,In_514);
xnor U645 (N_645,In_877,In_313);
nor U646 (N_646,In_509,In_567);
nor U647 (N_647,In_675,In_82);
nand U648 (N_648,In_728,In_685);
and U649 (N_649,In_434,In_506);
nand U650 (N_650,In_687,In_785);
nor U651 (N_651,In_68,In_353);
nor U652 (N_652,In_279,In_797);
nor U653 (N_653,In_569,In_821);
nor U654 (N_654,In_274,In_24);
and U655 (N_655,In_159,In_317);
nor U656 (N_656,In_268,In_886);
and U657 (N_657,In_57,In_639);
or U658 (N_658,In_545,In_834);
nor U659 (N_659,In_529,In_958);
nor U660 (N_660,In_566,In_332);
nor U661 (N_661,In_684,In_894);
nor U662 (N_662,In_553,In_300);
or U663 (N_663,In_542,In_75);
nor U664 (N_664,In_749,In_739);
and U665 (N_665,In_689,In_805);
or U666 (N_666,In_592,In_174);
or U667 (N_667,In_401,In_277);
and U668 (N_668,In_534,In_689);
nor U669 (N_669,In_79,In_17);
nor U670 (N_670,In_85,In_590);
nand U671 (N_671,In_971,In_823);
or U672 (N_672,In_332,In_81);
and U673 (N_673,In_383,In_630);
or U674 (N_674,In_921,In_23);
or U675 (N_675,In_779,In_33);
nand U676 (N_676,In_736,In_834);
or U677 (N_677,In_421,In_20);
or U678 (N_678,In_722,In_293);
and U679 (N_679,In_936,In_2);
or U680 (N_680,In_201,In_641);
and U681 (N_681,In_530,In_730);
nor U682 (N_682,In_680,In_130);
and U683 (N_683,In_20,In_898);
nand U684 (N_684,In_234,In_102);
nand U685 (N_685,In_906,In_253);
nor U686 (N_686,In_323,In_904);
nand U687 (N_687,In_535,In_355);
and U688 (N_688,In_703,In_135);
nor U689 (N_689,In_520,In_791);
xor U690 (N_690,In_7,In_248);
and U691 (N_691,In_85,In_149);
nor U692 (N_692,In_274,In_895);
and U693 (N_693,In_61,In_52);
and U694 (N_694,In_962,In_954);
nand U695 (N_695,In_790,In_216);
nand U696 (N_696,In_660,In_857);
or U697 (N_697,In_501,In_205);
or U698 (N_698,In_474,In_684);
nor U699 (N_699,In_883,In_732);
and U700 (N_700,In_748,In_974);
nor U701 (N_701,In_553,In_117);
and U702 (N_702,In_777,In_188);
xor U703 (N_703,In_823,In_961);
nor U704 (N_704,In_84,In_101);
or U705 (N_705,In_745,In_837);
or U706 (N_706,In_336,In_736);
and U707 (N_707,In_321,In_841);
nor U708 (N_708,In_28,In_269);
nor U709 (N_709,In_738,In_776);
or U710 (N_710,In_546,In_98);
xnor U711 (N_711,In_588,In_707);
nand U712 (N_712,In_552,In_848);
nand U713 (N_713,In_676,In_363);
and U714 (N_714,In_501,In_464);
nand U715 (N_715,In_418,In_211);
and U716 (N_716,In_336,In_265);
nor U717 (N_717,In_388,In_116);
nand U718 (N_718,In_875,In_357);
and U719 (N_719,In_254,In_169);
and U720 (N_720,In_990,In_216);
or U721 (N_721,In_565,In_216);
and U722 (N_722,In_653,In_203);
or U723 (N_723,In_408,In_828);
nand U724 (N_724,In_87,In_65);
nand U725 (N_725,In_645,In_141);
and U726 (N_726,In_57,In_622);
and U727 (N_727,In_574,In_186);
and U728 (N_728,In_277,In_132);
or U729 (N_729,In_248,In_939);
or U730 (N_730,In_815,In_198);
nor U731 (N_731,In_304,In_229);
nand U732 (N_732,In_357,In_797);
nand U733 (N_733,In_761,In_864);
and U734 (N_734,In_314,In_633);
and U735 (N_735,In_117,In_487);
or U736 (N_736,In_792,In_380);
nand U737 (N_737,In_942,In_449);
nand U738 (N_738,In_245,In_800);
and U739 (N_739,In_165,In_903);
and U740 (N_740,In_161,In_365);
nand U741 (N_741,In_215,In_993);
nand U742 (N_742,In_259,In_492);
or U743 (N_743,In_490,In_537);
and U744 (N_744,In_773,In_37);
or U745 (N_745,In_117,In_639);
xor U746 (N_746,In_197,In_54);
and U747 (N_747,In_208,In_122);
or U748 (N_748,In_285,In_388);
nand U749 (N_749,In_375,In_43);
nor U750 (N_750,In_256,In_110);
and U751 (N_751,In_151,In_636);
and U752 (N_752,In_705,In_332);
nor U753 (N_753,In_890,In_109);
nor U754 (N_754,In_15,In_190);
nor U755 (N_755,In_138,In_646);
nor U756 (N_756,In_822,In_58);
and U757 (N_757,In_853,In_513);
or U758 (N_758,In_771,In_913);
nand U759 (N_759,In_546,In_478);
and U760 (N_760,In_767,In_528);
and U761 (N_761,In_450,In_99);
or U762 (N_762,In_296,In_968);
and U763 (N_763,In_569,In_656);
and U764 (N_764,In_589,In_676);
nor U765 (N_765,In_631,In_311);
nand U766 (N_766,In_160,In_805);
or U767 (N_767,In_396,In_739);
nor U768 (N_768,In_400,In_17);
nand U769 (N_769,In_571,In_800);
nor U770 (N_770,In_578,In_550);
nand U771 (N_771,In_478,In_946);
xnor U772 (N_772,In_550,In_593);
or U773 (N_773,In_561,In_951);
xnor U774 (N_774,In_551,In_914);
nor U775 (N_775,In_918,In_305);
and U776 (N_776,In_291,In_688);
nand U777 (N_777,In_372,In_436);
nand U778 (N_778,In_373,In_525);
nand U779 (N_779,In_588,In_576);
and U780 (N_780,In_135,In_706);
and U781 (N_781,In_893,In_667);
nor U782 (N_782,In_636,In_155);
nand U783 (N_783,In_488,In_226);
or U784 (N_784,In_928,In_504);
nor U785 (N_785,In_805,In_281);
or U786 (N_786,In_555,In_689);
and U787 (N_787,In_124,In_254);
nand U788 (N_788,In_216,In_741);
or U789 (N_789,In_410,In_299);
nor U790 (N_790,In_307,In_62);
and U791 (N_791,In_680,In_88);
nand U792 (N_792,In_354,In_600);
nand U793 (N_793,In_947,In_588);
or U794 (N_794,In_513,In_543);
xor U795 (N_795,In_414,In_631);
nor U796 (N_796,In_640,In_650);
nor U797 (N_797,In_691,In_679);
nor U798 (N_798,In_732,In_337);
and U799 (N_799,In_809,In_322);
or U800 (N_800,In_611,In_301);
nor U801 (N_801,In_599,In_134);
and U802 (N_802,In_553,In_337);
nand U803 (N_803,In_459,In_200);
or U804 (N_804,In_388,In_437);
or U805 (N_805,In_566,In_996);
nor U806 (N_806,In_172,In_899);
nand U807 (N_807,In_999,In_993);
nand U808 (N_808,In_836,In_734);
nand U809 (N_809,In_422,In_289);
nor U810 (N_810,In_71,In_410);
and U811 (N_811,In_545,In_311);
nor U812 (N_812,In_31,In_226);
and U813 (N_813,In_131,In_954);
or U814 (N_814,In_256,In_757);
and U815 (N_815,In_235,In_137);
or U816 (N_816,In_467,In_877);
nand U817 (N_817,In_718,In_456);
and U818 (N_818,In_852,In_855);
nand U819 (N_819,In_501,In_743);
and U820 (N_820,In_472,In_739);
and U821 (N_821,In_990,In_161);
nor U822 (N_822,In_915,In_424);
nand U823 (N_823,In_652,In_58);
nor U824 (N_824,In_568,In_280);
nor U825 (N_825,In_72,In_281);
nor U826 (N_826,In_119,In_943);
nor U827 (N_827,In_848,In_717);
xor U828 (N_828,In_441,In_943);
nand U829 (N_829,In_613,In_294);
or U830 (N_830,In_489,In_239);
and U831 (N_831,In_338,In_815);
nand U832 (N_832,In_498,In_412);
nand U833 (N_833,In_954,In_550);
nor U834 (N_834,In_27,In_372);
nand U835 (N_835,In_387,In_893);
and U836 (N_836,In_422,In_31);
and U837 (N_837,In_917,In_645);
nor U838 (N_838,In_563,In_32);
and U839 (N_839,In_921,In_197);
and U840 (N_840,In_970,In_961);
xnor U841 (N_841,In_424,In_289);
nor U842 (N_842,In_574,In_441);
nand U843 (N_843,In_398,In_76);
and U844 (N_844,In_9,In_158);
and U845 (N_845,In_160,In_30);
nor U846 (N_846,In_927,In_658);
and U847 (N_847,In_335,In_508);
nor U848 (N_848,In_687,In_868);
xnor U849 (N_849,In_782,In_296);
nor U850 (N_850,In_814,In_534);
nand U851 (N_851,In_221,In_452);
and U852 (N_852,In_175,In_764);
nor U853 (N_853,In_288,In_933);
or U854 (N_854,In_610,In_214);
and U855 (N_855,In_993,In_274);
nand U856 (N_856,In_922,In_74);
nand U857 (N_857,In_306,In_580);
and U858 (N_858,In_648,In_164);
nand U859 (N_859,In_522,In_151);
or U860 (N_860,In_4,In_713);
or U861 (N_861,In_981,In_417);
nand U862 (N_862,In_255,In_274);
nor U863 (N_863,In_33,In_91);
nor U864 (N_864,In_167,In_183);
or U865 (N_865,In_859,In_421);
or U866 (N_866,In_402,In_362);
nand U867 (N_867,In_623,In_914);
nand U868 (N_868,In_592,In_819);
or U869 (N_869,In_390,In_921);
nand U870 (N_870,In_689,In_65);
and U871 (N_871,In_421,In_94);
nor U872 (N_872,In_583,In_359);
nand U873 (N_873,In_127,In_915);
or U874 (N_874,In_348,In_994);
nand U875 (N_875,In_279,In_452);
nor U876 (N_876,In_87,In_232);
nand U877 (N_877,In_755,In_697);
nor U878 (N_878,In_272,In_759);
nor U879 (N_879,In_222,In_20);
and U880 (N_880,In_945,In_136);
nor U881 (N_881,In_806,In_674);
or U882 (N_882,In_55,In_311);
nor U883 (N_883,In_394,In_813);
nand U884 (N_884,In_188,In_473);
and U885 (N_885,In_159,In_630);
and U886 (N_886,In_111,In_443);
or U887 (N_887,In_932,In_155);
nand U888 (N_888,In_491,In_834);
or U889 (N_889,In_813,In_748);
or U890 (N_890,In_440,In_338);
and U891 (N_891,In_184,In_707);
nand U892 (N_892,In_887,In_658);
nor U893 (N_893,In_111,In_65);
nor U894 (N_894,In_782,In_121);
nand U895 (N_895,In_818,In_865);
nand U896 (N_896,In_189,In_79);
or U897 (N_897,In_355,In_748);
nor U898 (N_898,In_64,In_668);
nand U899 (N_899,In_877,In_609);
and U900 (N_900,In_967,In_551);
nand U901 (N_901,In_754,In_365);
nand U902 (N_902,In_20,In_649);
nand U903 (N_903,In_784,In_273);
and U904 (N_904,In_7,In_174);
or U905 (N_905,In_715,In_550);
nor U906 (N_906,In_396,In_427);
nor U907 (N_907,In_510,In_718);
nand U908 (N_908,In_266,In_48);
and U909 (N_909,In_113,In_454);
and U910 (N_910,In_341,In_986);
nand U911 (N_911,In_99,In_480);
xnor U912 (N_912,In_652,In_194);
and U913 (N_913,In_719,In_1);
nand U914 (N_914,In_77,In_43);
nand U915 (N_915,In_591,In_715);
nor U916 (N_916,In_711,In_728);
or U917 (N_917,In_24,In_745);
nor U918 (N_918,In_175,In_351);
or U919 (N_919,In_305,In_91);
nor U920 (N_920,In_855,In_429);
nand U921 (N_921,In_541,In_878);
and U922 (N_922,In_499,In_310);
nand U923 (N_923,In_171,In_250);
or U924 (N_924,In_972,In_986);
nor U925 (N_925,In_259,In_633);
nand U926 (N_926,In_254,In_799);
and U927 (N_927,In_986,In_707);
and U928 (N_928,In_852,In_925);
nor U929 (N_929,In_453,In_276);
or U930 (N_930,In_342,In_467);
nand U931 (N_931,In_957,In_393);
and U932 (N_932,In_37,In_964);
and U933 (N_933,In_562,In_110);
and U934 (N_934,In_803,In_445);
nor U935 (N_935,In_747,In_456);
nand U936 (N_936,In_749,In_335);
nand U937 (N_937,In_282,In_854);
or U938 (N_938,In_503,In_162);
nor U939 (N_939,In_104,In_142);
or U940 (N_940,In_160,In_502);
or U941 (N_941,In_912,In_9);
and U942 (N_942,In_590,In_223);
or U943 (N_943,In_638,In_959);
nand U944 (N_944,In_786,In_922);
and U945 (N_945,In_851,In_234);
or U946 (N_946,In_363,In_990);
or U947 (N_947,In_521,In_211);
nand U948 (N_948,In_781,In_605);
or U949 (N_949,In_781,In_933);
nand U950 (N_950,In_393,In_80);
nand U951 (N_951,In_87,In_155);
or U952 (N_952,In_223,In_999);
xor U953 (N_953,In_504,In_880);
or U954 (N_954,In_49,In_246);
and U955 (N_955,In_583,In_334);
and U956 (N_956,In_709,In_534);
and U957 (N_957,In_597,In_871);
or U958 (N_958,In_433,In_350);
and U959 (N_959,In_363,In_993);
or U960 (N_960,In_187,In_700);
nand U961 (N_961,In_999,In_29);
or U962 (N_962,In_620,In_114);
nor U963 (N_963,In_140,In_356);
and U964 (N_964,In_833,In_698);
nor U965 (N_965,In_409,In_330);
nand U966 (N_966,In_74,In_872);
and U967 (N_967,In_490,In_220);
nand U968 (N_968,In_899,In_461);
nor U969 (N_969,In_976,In_83);
and U970 (N_970,In_116,In_709);
nor U971 (N_971,In_78,In_987);
and U972 (N_972,In_879,In_460);
or U973 (N_973,In_885,In_142);
nand U974 (N_974,In_243,In_247);
xnor U975 (N_975,In_837,In_850);
and U976 (N_976,In_509,In_0);
nand U977 (N_977,In_42,In_658);
nand U978 (N_978,In_219,In_705);
or U979 (N_979,In_691,In_675);
or U980 (N_980,In_562,In_501);
nor U981 (N_981,In_299,In_838);
or U982 (N_982,In_620,In_524);
or U983 (N_983,In_479,In_180);
nor U984 (N_984,In_155,In_767);
nand U985 (N_985,In_778,In_78);
or U986 (N_986,In_769,In_890);
nand U987 (N_987,In_804,In_550);
nand U988 (N_988,In_670,In_76);
or U989 (N_989,In_459,In_298);
and U990 (N_990,In_632,In_146);
or U991 (N_991,In_618,In_71);
and U992 (N_992,In_264,In_593);
or U993 (N_993,In_490,In_217);
and U994 (N_994,In_182,In_614);
and U995 (N_995,In_149,In_503);
or U996 (N_996,In_530,In_93);
nand U997 (N_997,In_272,In_163);
and U998 (N_998,In_458,In_262);
nor U999 (N_999,In_662,In_19);
nor U1000 (N_1000,N_133,N_818);
nor U1001 (N_1001,N_468,N_250);
nand U1002 (N_1002,N_561,N_348);
or U1003 (N_1003,N_841,N_827);
or U1004 (N_1004,N_56,N_402);
nand U1005 (N_1005,N_738,N_330);
xnor U1006 (N_1006,N_607,N_766);
or U1007 (N_1007,N_62,N_492);
nand U1008 (N_1008,N_374,N_596);
nor U1009 (N_1009,N_150,N_604);
nor U1010 (N_1010,N_430,N_166);
or U1011 (N_1011,N_793,N_942);
or U1012 (N_1012,N_429,N_158);
and U1013 (N_1013,N_851,N_884);
and U1014 (N_1014,N_312,N_603);
or U1015 (N_1015,N_275,N_232);
nand U1016 (N_1016,N_500,N_893);
nand U1017 (N_1017,N_987,N_777);
nor U1018 (N_1018,N_134,N_277);
nand U1019 (N_1019,N_662,N_999);
or U1020 (N_1020,N_555,N_235);
nor U1021 (N_1021,N_170,N_316);
nor U1022 (N_1022,N_979,N_392);
nand U1023 (N_1023,N_257,N_146);
or U1024 (N_1024,N_417,N_87);
and U1025 (N_1025,N_249,N_605);
or U1026 (N_1026,N_618,N_422);
or U1027 (N_1027,N_716,N_84);
nor U1028 (N_1028,N_178,N_912);
nand U1029 (N_1029,N_475,N_85);
nor U1030 (N_1030,N_447,N_209);
and U1031 (N_1031,N_273,N_126);
xor U1032 (N_1032,N_467,N_240);
and U1033 (N_1033,N_742,N_761);
and U1034 (N_1034,N_169,N_537);
and U1035 (N_1035,N_488,N_381);
nor U1036 (N_1036,N_589,N_573);
or U1037 (N_1037,N_53,N_720);
nand U1038 (N_1038,N_687,N_326);
or U1039 (N_1039,N_113,N_509);
and U1040 (N_1040,N_246,N_760);
and U1041 (N_1041,N_152,N_47);
or U1042 (N_1042,N_67,N_175);
and U1043 (N_1043,N_365,N_837);
nand U1044 (N_1044,N_506,N_242);
nand U1045 (N_1045,N_584,N_586);
nor U1046 (N_1046,N_620,N_754);
and U1047 (N_1047,N_413,N_737);
nor U1048 (N_1048,N_254,N_878);
nor U1049 (N_1049,N_951,N_991);
nor U1050 (N_1050,N_495,N_251);
or U1051 (N_1051,N_937,N_272);
or U1052 (N_1052,N_141,N_773);
and U1053 (N_1053,N_703,N_86);
nor U1054 (N_1054,N_576,N_787);
nor U1055 (N_1055,N_947,N_915);
nand U1056 (N_1056,N_568,N_310);
or U1057 (N_1057,N_428,N_439);
or U1058 (N_1058,N_921,N_805);
nand U1059 (N_1059,N_803,N_354);
and U1060 (N_1060,N_271,N_23);
nor U1061 (N_1061,N_698,N_383);
nand U1062 (N_1062,N_798,N_627);
nor U1063 (N_1063,N_828,N_99);
nor U1064 (N_1064,N_465,N_398);
nor U1065 (N_1065,N_955,N_905);
or U1066 (N_1066,N_518,N_785);
or U1067 (N_1067,N_40,N_83);
nor U1068 (N_1068,N_78,N_347);
and U1069 (N_1069,N_297,N_213);
and U1070 (N_1070,N_815,N_558);
nor U1071 (N_1071,N_744,N_385);
nand U1072 (N_1072,N_957,N_714);
and U1073 (N_1073,N_180,N_515);
or U1074 (N_1074,N_30,N_567);
or U1075 (N_1075,N_974,N_850);
nor U1076 (N_1076,N_194,N_711);
or U1077 (N_1077,N_438,N_16);
nand U1078 (N_1078,N_239,N_635);
or U1079 (N_1079,N_994,N_17);
nand U1080 (N_1080,N_253,N_114);
or U1081 (N_1081,N_0,N_42);
nor U1082 (N_1082,N_2,N_368);
and U1083 (N_1083,N_886,N_221);
nand U1084 (N_1084,N_733,N_412);
nand U1085 (N_1085,N_591,N_410);
nand U1086 (N_1086,N_625,N_795);
and U1087 (N_1087,N_369,N_963);
and U1088 (N_1088,N_58,N_964);
nand U1089 (N_1089,N_968,N_334);
and U1090 (N_1090,N_525,N_517);
or U1091 (N_1091,N_357,N_936);
or U1092 (N_1092,N_167,N_661);
and U1093 (N_1093,N_772,N_634);
or U1094 (N_1094,N_395,N_732);
nand U1095 (N_1095,N_228,N_643);
and U1096 (N_1096,N_177,N_13);
and U1097 (N_1097,N_918,N_204);
and U1098 (N_1098,N_457,N_350);
xnor U1099 (N_1099,N_888,N_751);
or U1100 (N_1100,N_973,N_847);
nand U1101 (N_1101,N_340,N_959);
and U1102 (N_1102,N_9,N_355);
and U1103 (N_1103,N_444,N_94);
nand U1104 (N_1104,N_538,N_63);
or U1105 (N_1105,N_230,N_51);
or U1106 (N_1106,N_692,N_375);
and U1107 (N_1107,N_341,N_107);
xor U1108 (N_1108,N_343,N_989);
and U1109 (N_1109,N_535,N_472);
and U1110 (N_1110,N_44,N_702);
nor U1111 (N_1111,N_466,N_932);
and U1112 (N_1112,N_753,N_746);
nor U1113 (N_1113,N_922,N_728);
nor U1114 (N_1114,N_299,N_524);
or U1115 (N_1115,N_840,N_206);
nor U1116 (N_1116,N_119,N_481);
and U1117 (N_1117,N_45,N_967);
nand U1118 (N_1118,N_432,N_657);
or U1119 (N_1119,N_41,N_770);
nor U1120 (N_1120,N_889,N_322);
and U1121 (N_1121,N_306,N_266);
nor U1122 (N_1122,N_755,N_757);
nand U1123 (N_1123,N_1,N_91);
or U1124 (N_1124,N_387,N_880);
or U1125 (N_1125,N_482,N_715);
or U1126 (N_1126,N_844,N_890);
nand U1127 (N_1127,N_258,N_445);
and U1128 (N_1128,N_806,N_476);
and U1129 (N_1129,N_871,N_335);
and U1130 (N_1130,N_210,N_164);
xor U1131 (N_1131,N_54,N_581);
and U1132 (N_1132,N_900,N_110);
and U1133 (N_1133,N_799,N_867);
and U1134 (N_1134,N_223,N_224);
nand U1135 (N_1135,N_642,N_252);
nand U1136 (N_1136,N_440,N_424);
nor U1137 (N_1137,N_135,N_193);
or U1138 (N_1138,N_965,N_65);
nand U1139 (N_1139,N_647,N_870);
nor U1140 (N_1140,N_786,N_508);
nor U1141 (N_1141,N_609,N_804);
xnor U1142 (N_1142,N_590,N_699);
nor U1143 (N_1143,N_529,N_353);
nor U1144 (N_1144,N_924,N_856);
and U1145 (N_1145,N_628,N_283);
or U1146 (N_1146,N_174,N_961);
and U1147 (N_1147,N_400,N_911);
nand U1148 (N_1148,N_274,N_520);
nor U1149 (N_1149,N_366,N_825);
xor U1150 (N_1150,N_521,N_512);
nand U1151 (N_1151,N_676,N_27);
nand U1152 (N_1152,N_291,N_280);
nand U1153 (N_1153,N_588,N_667);
or U1154 (N_1154,N_4,N_903);
nand U1155 (N_1155,N_248,N_490);
nand U1156 (N_1156,N_995,N_983);
and U1157 (N_1157,N_90,N_115);
xor U1158 (N_1158,N_877,N_547);
nand U1159 (N_1159,N_39,N_990);
and U1160 (N_1160,N_68,N_172);
and U1161 (N_1161,N_247,N_441);
nor U1162 (N_1162,N_314,N_927);
and U1163 (N_1163,N_631,N_191);
and U1164 (N_1164,N_727,N_833);
and U1165 (N_1165,N_632,N_677);
nand U1166 (N_1166,N_653,N_626);
and U1167 (N_1167,N_846,N_323);
nand U1168 (N_1168,N_153,N_22);
nor U1169 (N_1169,N_516,N_189);
and U1170 (N_1170,N_938,N_843);
or U1171 (N_1171,N_98,N_443);
nor U1172 (N_1172,N_104,N_35);
or U1173 (N_1173,N_928,N_759);
and U1174 (N_1174,N_415,N_469);
and U1175 (N_1175,N_984,N_553);
nor U1176 (N_1176,N_199,N_906);
nand U1177 (N_1177,N_33,N_278);
xnor U1178 (N_1178,N_982,N_648);
nand U1179 (N_1179,N_97,N_225);
and U1180 (N_1180,N_95,N_775);
and U1181 (N_1181,N_998,N_971);
and U1182 (N_1182,N_265,N_736);
nand U1183 (N_1183,N_981,N_872);
or U1184 (N_1184,N_459,N_564);
and U1185 (N_1185,N_543,N_941);
and U1186 (N_1186,N_860,N_378);
nor U1187 (N_1187,N_931,N_790);
nand U1188 (N_1188,N_92,N_705);
nor U1189 (N_1189,N_8,N_857);
nand U1190 (N_1190,N_619,N_691);
nand U1191 (N_1191,N_969,N_106);
or U1192 (N_1192,N_132,N_282);
and U1193 (N_1193,N_60,N_245);
nand U1194 (N_1194,N_414,N_32);
nor U1195 (N_1195,N_531,N_497);
and U1196 (N_1196,N_261,N_52);
or U1197 (N_1197,N_863,N_997);
or U1198 (N_1198,N_909,N_136);
nand U1199 (N_1199,N_286,N_303);
nand U1200 (N_1200,N_845,N_934);
xnor U1201 (N_1201,N_658,N_156);
xor U1202 (N_1202,N_259,N_784);
or U1203 (N_1203,N_236,N_608);
or U1204 (N_1204,N_861,N_168);
or U1205 (N_1205,N_907,N_663);
and U1206 (N_1206,N_190,N_587);
or U1207 (N_1207,N_382,N_655);
nor U1208 (N_1208,N_401,N_202);
and U1209 (N_1209,N_866,N_621);
and U1210 (N_1210,N_570,N_701);
nor U1211 (N_1211,N_741,N_752);
or U1212 (N_1212,N_454,N_717);
nand U1213 (N_1213,N_853,N_838);
and U1214 (N_1214,N_214,N_317);
nand U1215 (N_1215,N_73,N_530);
and U1216 (N_1216,N_583,N_883);
and U1217 (N_1217,N_142,N_36);
nor U1218 (N_1218,N_11,N_796);
nor U1219 (N_1219,N_187,N_565);
nand U1220 (N_1220,N_666,N_638);
nor U1221 (N_1221,N_37,N_954);
nor U1222 (N_1222,N_739,N_260);
or U1223 (N_1223,N_645,N_49);
or U1224 (N_1224,N_380,N_532);
or U1225 (N_1225,N_735,N_217);
nor U1226 (N_1226,N_898,N_894);
or U1227 (N_1227,N_933,N_449);
nand U1228 (N_1228,N_143,N_970);
nor U1229 (N_1229,N_534,N_270);
nand U1230 (N_1230,N_814,N_307);
nor U1231 (N_1231,N_745,N_925);
nor U1232 (N_1232,N_498,N_820);
and U1233 (N_1233,N_528,N_293);
nand U1234 (N_1234,N_656,N_822);
nor U1235 (N_1235,N_102,N_862);
and U1236 (N_1236,N_5,N_539);
or U1237 (N_1237,N_423,N_18);
and U1238 (N_1238,N_526,N_302);
or U1239 (N_1239,N_418,N_899);
nand U1240 (N_1240,N_816,N_391);
and U1241 (N_1241,N_962,N_285);
and U1242 (N_1242,N_124,N_131);
nand U1243 (N_1243,N_318,N_208);
nand U1244 (N_1244,N_671,N_494);
and U1245 (N_1245,N_29,N_810);
or U1246 (N_1246,N_471,N_145);
or U1247 (N_1247,N_578,N_780);
nand U1248 (N_1248,N_926,N_950);
nor U1249 (N_1249,N_743,N_876);
nand U1250 (N_1250,N_849,N_923);
nor U1251 (N_1251,N_783,N_352);
nand U1252 (N_1252,N_858,N_376);
and U1253 (N_1253,N_304,N_309);
nor U1254 (N_1254,N_24,N_522);
nor U1255 (N_1255,N_96,N_461);
nand U1256 (N_1256,N_680,N_144);
nor U1257 (N_1257,N_519,N_707);
nand U1258 (N_1258,N_292,N_460);
nor U1259 (N_1259,N_329,N_474);
nand U1260 (N_1260,N_479,N_154);
or U1261 (N_1261,N_389,N_864);
nor U1262 (N_1262,N_345,N_137);
nand U1263 (N_1263,N_678,N_268);
nor U1264 (N_1264,N_89,N_483);
and U1265 (N_1265,N_823,N_569);
and U1266 (N_1266,N_593,N_425);
and U1267 (N_1267,N_713,N_74);
or U1268 (N_1268,N_956,N_197);
nor U1269 (N_1269,N_697,N_473);
and U1270 (N_1270,N_219,N_176);
nand U1271 (N_1271,N_70,N_262);
or U1272 (N_1272,N_895,N_364);
nand U1273 (N_1273,N_882,N_544);
nand U1274 (N_1274,N_767,N_750);
and U1275 (N_1275,N_386,N_377);
or U1276 (N_1276,N_267,N_493);
or U1277 (N_1277,N_649,N_551);
and U1278 (N_1278,N_416,N_88);
or U1279 (N_1279,N_173,N_76);
or U1280 (N_1280,N_712,N_298);
and U1281 (N_1281,N_477,N_399);
or U1282 (N_1282,N_611,N_81);
or U1283 (N_1283,N_276,N_462);
nand U1284 (N_1284,N_161,N_367);
or U1285 (N_1285,N_617,N_978);
and U1286 (N_1286,N_865,N_287);
or U1287 (N_1287,N_346,N_875);
nand U1288 (N_1288,N_43,N_220);
nand U1289 (N_1289,N_129,N_216);
nor U1290 (N_1290,N_103,N_935);
or U1291 (N_1291,N_710,N_301);
nand U1292 (N_1292,N_433,N_66);
nor U1293 (N_1293,N_940,N_264);
or U1294 (N_1294,N_646,N_390);
or U1295 (N_1295,N_533,N_25);
nor U1296 (N_1296,N_300,N_308);
or U1297 (N_1297,N_830,N_571);
or U1298 (N_1298,N_130,N_237);
and U1299 (N_1299,N_859,N_993);
or U1300 (N_1300,N_123,N_327);
and U1301 (N_1301,N_211,N_238);
and U1302 (N_1302,N_665,N_71);
nor U1303 (N_1303,N_781,N_10);
nand U1304 (N_1304,N_910,N_975);
nor U1305 (N_1305,N_188,N_797);
or U1306 (N_1306,N_652,N_641);
or U1307 (N_1307,N_511,N_908);
nor U1308 (N_1308,N_769,N_171);
and U1309 (N_1309,N_536,N_949);
nor U1310 (N_1310,N_779,N_855);
nand U1311 (N_1311,N_791,N_675);
or U1312 (N_1312,N_801,N_336);
nand U1313 (N_1313,N_580,N_943);
and U1314 (N_1314,N_195,N_852);
or U1315 (N_1315,N_747,N_332);
nor U1316 (N_1316,N_572,N_320);
or U1317 (N_1317,N_879,N_255);
xnor U1318 (N_1318,N_28,N_198);
or U1319 (N_1319,N_234,N_765);
nand U1320 (N_1320,N_405,N_944);
nand U1321 (N_1321,N_478,N_985);
and U1322 (N_1322,N_694,N_157);
nor U1323 (N_1323,N_231,N_61);
nand U1324 (N_1324,N_953,N_284);
nor U1325 (N_1325,N_807,N_901);
nand U1326 (N_1326,N_723,N_696);
nand U1327 (N_1327,N_939,N_59);
nand U1328 (N_1328,N_470,N_598);
or U1329 (N_1329,N_541,N_919);
nor U1330 (N_1330,N_6,N_281);
nand U1331 (N_1331,N_328,N_196);
or U1332 (N_1332,N_624,N_279);
nand U1333 (N_1333,N_361,N_480);
nor U1334 (N_1334,N_486,N_319);
nor U1335 (N_1335,N_453,N_514);
and U1336 (N_1336,N_562,N_162);
and U1337 (N_1337,N_792,N_930);
or U1338 (N_1338,N_778,N_200);
or U1339 (N_1339,N_668,N_585);
nand U1340 (N_1340,N_77,N_148);
xnor U1341 (N_1341,N_874,N_574);
and U1342 (N_1342,N_724,N_689);
nand U1343 (N_1343,N_325,N_730);
or U1344 (N_1344,N_673,N_637);
nand U1345 (N_1345,N_913,N_105);
nor U1346 (N_1346,N_125,N_693);
or U1347 (N_1347,N_324,N_813);
and U1348 (N_1348,N_505,N_669);
or U1349 (N_1349,N_679,N_660);
nor U1350 (N_1350,N_409,N_542);
nor U1351 (N_1351,N_149,N_550);
or U1352 (N_1352,N_873,N_700);
and U1353 (N_1353,N_996,N_456);
and U1354 (N_1354,N_575,N_545);
and U1355 (N_1355,N_892,N_321);
xor U1356 (N_1356,N_331,N_116);
nand U1357 (N_1357,N_19,N_159);
or U1358 (N_1358,N_640,N_359);
nor U1359 (N_1359,N_826,N_370);
or U1360 (N_1360,N_834,N_458);
nor U1361 (N_1361,N_758,N_311);
and U1362 (N_1362,N_427,N_147);
and U1363 (N_1363,N_295,N_421);
nor U1364 (N_1364,N_362,N_450);
and U1365 (N_1365,N_501,N_948);
or U1366 (N_1366,N_21,N_333);
or U1367 (N_1367,N_904,N_832);
and U1368 (N_1368,N_269,N_546);
nor U1369 (N_1369,N_139,N_920);
nand U1370 (N_1370,N_182,N_442);
and U1371 (N_1371,N_384,N_437);
nand U1372 (N_1372,N_681,N_127);
and U1373 (N_1373,N_756,N_50);
nand U1374 (N_1374,N_774,N_672);
nand U1375 (N_1375,N_848,N_740);
and U1376 (N_1376,N_379,N_557);
and U1377 (N_1377,N_579,N_674);
or U1378 (N_1378,N_592,N_902);
nand U1379 (N_1379,N_686,N_819);
nor U1380 (N_1380,N_824,N_577);
or U1381 (N_1381,N_722,N_601);
and U1382 (N_1382,N_349,N_946);
nor U1383 (N_1383,N_205,N_109);
nand U1384 (N_1384,N_695,N_891);
nand U1385 (N_1385,N_363,N_455);
and U1386 (N_1386,N_184,N_929);
or U1387 (N_1387,N_771,N_633);
and U1388 (N_1388,N_831,N_48);
and U1389 (N_1389,N_484,N_725);
nor U1390 (N_1390,N_683,N_463);
nand U1391 (N_1391,N_315,N_600);
nand U1392 (N_1392,N_836,N_881);
nand U1393 (N_1393,N_226,N_958);
xnor U1394 (N_1394,N_227,N_811);
or U1395 (N_1395,N_407,N_839);
nand U1396 (N_1396,N_977,N_80);
nand U1397 (N_1397,N_185,N_101);
xor U1398 (N_1398,N_305,N_966);
and U1399 (N_1399,N_339,N_290);
nor U1400 (N_1400,N_615,N_491);
xor U1401 (N_1401,N_393,N_606);
and U1402 (N_1402,N_972,N_748);
nor U1403 (N_1403,N_639,N_731);
or U1404 (N_1404,N_289,N_594);
nor U1405 (N_1405,N_782,N_64);
nor U1406 (N_1406,N_201,N_842);
or U1407 (N_1407,N_706,N_342);
nor U1408 (N_1408,N_485,N_802);
nor U1409 (N_1409,N_595,N_708);
or U1410 (N_1410,N_897,N_749);
nand U1411 (N_1411,N_75,N_582);
and U1412 (N_1412,N_622,N_344);
nand U1413 (N_1413,N_854,N_294);
and U1414 (N_1414,N_34,N_718);
and U1415 (N_1415,N_3,N_829);
nor U1416 (N_1416,N_82,N_207);
nor U1417 (N_1417,N_690,N_659);
or U1418 (N_1418,N_436,N_613);
or U1419 (N_1419,N_650,N_644);
nor U1420 (N_1420,N_869,N_121);
nand U1421 (N_1421,N_719,N_118);
and U1422 (N_1422,N_729,N_396);
nor U1423 (N_1423,N_15,N_599);
nand U1424 (N_1424,N_682,N_945);
nand U1425 (N_1425,N_808,N_434);
or U1426 (N_1426,N_452,N_373);
nand U1427 (N_1427,N_358,N_835);
or U1428 (N_1428,N_215,N_431);
nor U1429 (N_1429,N_885,N_241);
and U1430 (N_1430,N_426,N_112);
nand U1431 (N_1431,N_14,N_549);
nand U1432 (N_1432,N_868,N_630);
or U1433 (N_1433,N_79,N_420);
nand U1434 (N_1434,N_563,N_20);
or U1435 (N_1435,N_155,N_952);
nor U1436 (N_1436,N_411,N_548);
or U1437 (N_1437,N_288,N_685);
and U1438 (N_1438,N_654,N_165);
nand U1439 (N_1439,N_111,N_183);
and U1440 (N_1440,N_72,N_108);
xor U1441 (N_1441,N_960,N_916);
or U1442 (N_1442,N_489,N_917);
nand U1443 (N_1443,N_616,N_222);
nand U1444 (N_1444,N_100,N_93);
nor U1445 (N_1445,N_122,N_554);
and U1446 (N_1446,N_404,N_408);
or U1447 (N_1447,N_186,N_38);
nand U1448 (N_1448,N_734,N_179);
nand U1449 (N_1449,N_496,N_448);
and U1450 (N_1450,N_992,N_513);
or U1451 (N_1451,N_768,N_233);
nor U1452 (N_1452,N_800,N_614);
nor U1453 (N_1453,N_629,N_120);
or U1454 (N_1454,N_762,N_986);
nor U1455 (N_1455,N_651,N_523);
xnor U1456 (N_1456,N_503,N_789);
nor U1457 (N_1457,N_403,N_709);
or U1458 (N_1458,N_721,N_419);
and U1459 (N_1459,N_487,N_360);
or U1460 (N_1460,N_504,N_559);
nand U1461 (N_1461,N_540,N_151);
nand U1462 (N_1462,N_812,N_57);
or U1463 (N_1463,N_502,N_988);
or U1464 (N_1464,N_636,N_464);
nand U1465 (N_1465,N_338,N_809);
and U1466 (N_1466,N_212,N_181);
and U1467 (N_1467,N_764,N_46);
nor U1468 (N_1468,N_263,N_31);
and U1469 (N_1469,N_69,N_821);
nor U1470 (N_1470,N_296,N_976);
nor U1471 (N_1471,N_356,N_527);
nor U1472 (N_1472,N_612,N_435);
and U1473 (N_1473,N_566,N_664);
nor U1474 (N_1474,N_794,N_26);
nor U1475 (N_1475,N_704,N_788);
or U1476 (N_1476,N_160,N_218);
or U1477 (N_1477,N_117,N_914);
or U1478 (N_1478,N_256,N_371);
and U1479 (N_1479,N_388,N_980);
or U1480 (N_1480,N_372,N_337);
and U1481 (N_1481,N_140,N_394);
and U1482 (N_1482,N_244,N_510);
and U1483 (N_1483,N_556,N_406);
and U1484 (N_1484,N_688,N_763);
nand U1485 (N_1485,N_229,N_776);
or U1486 (N_1486,N_12,N_313);
or U1487 (N_1487,N_610,N_446);
nor U1488 (N_1488,N_684,N_602);
nor U1489 (N_1489,N_560,N_507);
nand U1490 (N_1490,N_397,N_351);
nor U1491 (N_1491,N_163,N_243);
and U1492 (N_1492,N_203,N_138);
or U1493 (N_1493,N_192,N_128);
nor U1494 (N_1494,N_499,N_670);
and U1495 (N_1495,N_7,N_817);
and U1496 (N_1496,N_726,N_597);
and U1497 (N_1497,N_552,N_623);
or U1498 (N_1498,N_451,N_887);
or U1499 (N_1499,N_55,N_896);
nor U1500 (N_1500,N_90,N_677);
and U1501 (N_1501,N_118,N_508);
nor U1502 (N_1502,N_939,N_723);
nor U1503 (N_1503,N_334,N_759);
nand U1504 (N_1504,N_140,N_360);
or U1505 (N_1505,N_806,N_609);
nor U1506 (N_1506,N_920,N_8);
nor U1507 (N_1507,N_214,N_375);
nand U1508 (N_1508,N_618,N_606);
or U1509 (N_1509,N_809,N_578);
nand U1510 (N_1510,N_484,N_73);
nor U1511 (N_1511,N_580,N_565);
or U1512 (N_1512,N_306,N_238);
or U1513 (N_1513,N_87,N_400);
or U1514 (N_1514,N_602,N_78);
nand U1515 (N_1515,N_74,N_362);
nor U1516 (N_1516,N_857,N_880);
and U1517 (N_1517,N_679,N_326);
nand U1518 (N_1518,N_382,N_127);
nand U1519 (N_1519,N_620,N_962);
and U1520 (N_1520,N_597,N_263);
or U1521 (N_1521,N_516,N_300);
and U1522 (N_1522,N_91,N_652);
and U1523 (N_1523,N_380,N_467);
nor U1524 (N_1524,N_156,N_487);
nor U1525 (N_1525,N_703,N_722);
nor U1526 (N_1526,N_868,N_826);
or U1527 (N_1527,N_162,N_680);
and U1528 (N_1528,N_542,N_344);
nor U1529 (N_1529,N_96,N_365);
xnor U1530 (N_1530,N_621,N_130);
and U1531 (N_1531,N_852,N_358);
nand U1532 (N_1532,N_621,N_920);
and U1533 (N_1533,N_929,N_810);
or U1534 (N_1534,N_552,N_512);
and U1535 (N_1535,N_197,N_320);
or U1536 (N_1536,N_487,N_466);
nand U1537 (N_1537,N_719,N_917);
and U1538 (N_1538,N_115,N_33);
and U1539 (N_1539,N_227,N_551);
xor U1540 (N_1540,N_381,N_584);
nand U1541 (N_1541,N_950,N_994);
or U1542 (N_1542,N_921,N_675);
or U1543 (N_1543,N_622,N_476);
or U1544 (N_1544,N_973,N_611);
nand U1545 (N_1545,N_848,N_522);
and U1546 (N_1546,N_17,N_196);
and U1547 (N_1547,N_404,N_799);
xnor U1548 (N_1548,N_662,N_393);
or U1549 (N_1549,N_578,N_115);
or U1550 (N_1550,N_821,N_944);
and U1551 (N_1551,N_508,N_954);
or U1552 (N_1552,N_50,N_426);
or U1553 (N_1553,N_239,N_971);
nor U1554 (N_1554,N_749,N_685);
nand U1555 (N_1555,N_340,N_963);
nand U1556 (N_1556,N_503,N_924);
or U1557 (N_1557,N_939,N_42);
or U1558 (N_1558,N_30,N_63);
nand U1559 (N_1559,N_702,N_253);
or U1560 (N_1560,N_617,N_648);
nand U1561 (N_1561,N_935,N_634);
or U1562 (N_1562,N_741,N_414);
nand U1563 (N_1563,N_603,N_255);
or U1564 (N_1564,N_9,N_80);
and U1565 (N_1565,N_370,N_973);
and U1566 (N_1566,N_158,N_241);
nand U1567 (N_1567,N_493,N_544);
and U1568 (N_1568,N_863,N_662);
nor U1569 (N_1569,N_395,N_510);
nor U1570 (N_1570,N_277,N_438);
nand U1571 (N_1571,N_493,N_903);
and U1572 (N_1572,N_230,N_346);
nor U1573 (N_1573,N_493,N_758);
and U1574 (N_1574,N_859,N_989);
nor U1575 (N_1575,N_304,N_950);
nor U1576 (N_1576,N_581,N_418);
or U1577 (N_1577,N_762,N_22);
or U1578 (N_1578,N_423,N_5);
nor U1579 (N_1579,N_71,N_868);
or U1580 (N_1580,N_6,N_785);
and U1581 (N_1581,N_379,N_922);
nor U1582 (N_1582,N_558,N_415);
nand U1583 (N_1583,N_504,N_85);
nand U1584 (N_1584,N_627,N_497);
nand U1585 (N_1585,N_970,N_888);
or U1586 (N_1586,N_356,N_395);
nand U1587 (N_1587,N_910,N_713);
nand U1588 (N_1588,N_387,N_423);
nand U1589 (N_1589,N_405,N_628);
nor U1590 (N_1590,N_138,N_713);
nor U1591 (N_1591,N_647,N_284);
xnor U1592 (N_1592,N_519,N_534);
xor U1593 (N_1593,N_64,N_67);
or U1594 (N_1594,N_91,N_339);
nor U1595 (N_1595,N_480,N_685);
nand U1596 (N_1596,N_381,N_679);
or U1597 (N_1597,N_346,N_195);
nor U1598 (N_1598,N_380,N_119);
and U1599 (N_1599,N_915,N_772);
nor U1600 (N_1600,N_661,N_859);
nor U1601 (N_1601,N_851,N_137);
and U1602 (N_1602,N_808,N_402);
or U1603 (N_1603,N_627,N_843);
or U1604 (N_1604,N_494,N_32);
nand U1605 (N_1605,N_791,N_659);
and U1606 (N_1606,N_769,N_651);
and U1607 (N_1607,N_493,N_800);
or U1608 (N_1608,N_883,N_498);
nor U1609 (N_1609,N_322,N_885);
or U1610 (N_1610,N_151,N_291);
nor U1611 (N_1611,N_306,N_466);
and U1612 (N_1612,N_404,N_776);
or U1613 (N_1613,N_633,N_902);
nand U1614 (N_1614,N_2,N_538);
and U1615 (N_1615,N_492,N_29);
nand U1616 (N_1616,N_192,N_50);
xnor U1617 (N_1617,N_10,N_397);
nand U1618 (N_1618,N_725,N_338);
nand U1619 (N_1619,N_372,N_507);
and U1620 (N_1620,N_805,N_584);
or U1621 (N_1621,N_237,N_663);
or U1622 (N_1622,N_316,N_972);
nand U1623 (N_1623,N_241,N_682);
or U1624 (N_1624,N_727,N_989);
and U1625 (N_1625,N_555,N_200);
xnor U1626 (N_1626,N_11,N_745);
or U1627 (N_1627,N_127,N_983);
and U1628 (N_1628,N_62,N_522);
and U1629 (N_1629,N_825,N_940);
nor U1630 (N_1630,N_521,N_767);
nand U1631 (N_1631,N_465,N_275);
nor U1632 (N_1632,N_358,N_108);
nand U1633 (N_1633,N_208,N_275);
or U1634 (N_1634,N_582,N_951);
nor U1635 (N_1635,N_897,N_177);
nor U1636 (N_1636,N_614,N_730);
and U1637 (N_1637,N_174,N_936);
nor U1638 (N_1638,N_279,N_746);
or U1639 (N_1639,N_249,N_16);
nand U1640 (N_1640,N_107,N_786);
nor U1641 (N_1641,N_773,N_695);
nor U1642 (N_1642,N_979,N_884);
nand U1643 (N_1643,N_830,N_695);
nand U1644 (N_1644,N_252,N_888);
or U1645 (N_1645,N_536,N_543);
or U1646 (N_1646,N_198,N_101);
or U1647 (N_1647,N_575,N_620);
nand U1648 (N_1648,N_877,N_842);
or U1649 (N_1649,N_614,N_138);
and U1650 (N_1650,N_501,N_982);
and U1651 (N_1651,N_837,N_333);
nand U1652 (N_1652,N_527,N_177);
and U1653 (N_1653,N_401,N_217);
or U1654 (N_1654,N_582,N_720);
and U1655 (N_1655,N_82,N_876);
nor U1656 (N_1656,N_734,N_89);
and U1657 (N_1657,N_733,N_627);
nand U1658 (N_1658,N_108,N_883);
nand U1659 (N_1659,N_618,N_95);
nand U1660 (N_1660,N_231,N_506);
nand U1661 (N_1661,N_722,N_810);
nor U1662 (N_1662,N_713,N_826);
nor U1663 (N_1663,N_430,N_758);
and U1664 (N_1664,N_333,N_565);
xnor U1665 (N_1665,N_312,N_182);
nor U1666 (N_1666,N_534,N_377);
or U1667 (N_1667,N_216,N_839);
nand U1668 (N_1668,N_240,N_935);
nor U1669 (N_1669,N_74,N_992);
nor U1670 (N_1670,N_581,N_328);
nor U1671 (N_1671,N_415,N_308);
nor U1672 (N_1672,N_459,N_117);
and U1673 (N_1673,N_137,N_455);
nand U1674 (N_1674,N_854,N_554);
nand U1675 (N_1675,N_10,N_472);
or U1676 (N_1676,N_247,N_418);
nor U1677 (N_1677,N_919,N_743);
nand U1678 (N_1678,N_863,N_515);
or U1679 (N_1679,N_928,N_413);
nor U1680 (N_1680,N_327,N_263);
xor U1681 (N_1681,N_462,N_54);
or U1682 (N_1682,N_939,N_726);
nand U1683 (N_1683,N_657,N_590);
and U1684 (N_1684,N_619,N_588);
or U1685 (N_1685,N_23,N_528);
nor U1686 (N_1686,N_657,N_566);
nor U1687 (N_1687,N_141,N_845);
or U1688 (N_1688,N_85,N_193);
and U1689 (N_1689,N_133,N_618);
nor U1690 (N_1690,N_189,N_96);
nor U1691 (N_1691,N_548,N_362);
and U1692 (N_1692,N_702,N_146);
nand U1693 (N_1693,N_262,N_659);
nand U1694 (N_1694,N_413,N_736);
nand U1695 (N_1695,N_818,N_270);
nand U1696 (N_1696,N_874,N_98);
nor U1697 (N_1697,N_353,N_156);
nor U1698 (N_1698,N_257,N_625);
nor U1699 (N_1699,N_232,N_612);
and U1700 (N_1700,N_345,N_19);
nand U1701 (N_1701,N_510,N_594);
and U1702 (N_1702,N_332,N_310);
or U1703 (N_1703,N_240,N_548);
or U1704 (N_1704,N_965,N_856);
nor U1705 (N_1705,N_758,N_390);
nor U1706 (N_1706,N_651,N_211);
nor U1707 (N_1707,N_582,N_959);
nand U1708 (N_1708,N_993,N_775);
nor U1709 (N_1709,N_202,N_351);
or U1710 (N_1710,N_863,N_89);
nor U1711 (N_1711,N_962,N_766);
nand U1712 (N_1712,N_821,N_225);
or U1713 (N_1713,N_9,N_372);
or U1714 (N_1714,N_793,N_796);
nand U1715 (N_1715,N_23,N_994);
nor U1716 (N_1716,N_255,N_89);
nor U1717 (N_1717,N_964,N_498);
nand U1718 (N_1718,N_721,N_994);
or U1719 (N_1719,N_66,N_631);
and U1720 (N_1720,N_862,N_400);
or U1721 (N_1721,N_12,N_138);
or U1722 (N_1722,N_67,N_194);
nand U1723 (N_1723,N_822,N_632);
or U1724 (N_1724,N_942,N_822);
and U1725 (N_1725,N_664,N_412);
or U1726 (N_1726,N_13,N_298);
and U1727 (N_1727,N_430,N_94);
and U1728 (N_1728,N_940,N_855);
or U1729 (N_1729,N_731,N_313);
nand U1730 (N_1730,N_997,N_856);
or U1731 (N_1731,N_406,N_916);
nand U1732 (N_1732,N_526,N_428);
and U1733 (N_1733,N_246,N_104);
or U1734 (N_1734,N_782,N_489);
xnor U1735 (N_1735,N_997,N_734);
nand U1736 (N_1736,N_926,N_970);
nand U1737 (N_1737,N_837,N_118);
or U1738 (N_1738,N_952,N_781);
nor U1739 (N_1739,N_266,N_852);
nand U1740 (N_1740,N_210,N_239);
and U1741 (N_1741,N_181,N_407);
or U1742 (N_1742,N_647,N_918);
nand U1743 (N_1743,N_853,N_979);
nor U1744 (N_1744,N_145,N_870);
or U1745 (N_1745,N_137,N_638);
nor U1746 (N_1746,N_545,N_258);
nand U1747 (N_1747,N_593,N_900);
and U1748 (N_1748,N_270,N_662);
or U1749 (N_1749,N_258,N_896);
nand U1750 (N_1750,N_220,N_775);
or U1751 (N_1751,N_543,N_294);
nor U1752 (N_1752,N_256,N_511);
nand U1753 (N_1753,N_522,N_667);
nand U1754 (N_1754,N_149,N_474);
and U1755 (N_1755,N_584,N_473);
and U1756 (N_1756,N_391,N_637);
xnor U1757 (N_1757,N_241,N_863);
nor U1758 (N_1758,N_155,N_135);
xor U1759 (N_1759,N_616,N_225);
or U1760 (N_1760,N_200,N_195);
or U1761 (N_1761,N_497,N_899);
and U1762 (N_1762,N_834,N_537);
nor U1763 (N_1763,N_57,N_535);
and U1764 (N_1764,N_511,N_512);
nor U1765 (N_1765,N_940,N_886);
nor U1766 (N_1766,N_646,N_589);
nor U1767 (N_1767,N_532,N_159);
and U1768 (N_1768,N_870,N_577);
nand U1769 (N_1769,N_753,N_137);
nand U1770 (N_1770,N_348,N_773);
or U1771 (N_1771,N_431,N_766);
nor U1772 (N_1772,N_54,N_193);
or U1773 (N_1773,N_253,N_179);
or U1774 (N_1774,N_967,N_947);
or U1775 (N_1775,N_591,N_555);
nand U1776 (N_1776,N_246,N_466);
or U1777 (N_1777,N_233,N_860);
and U1778 (N_1778,N_750,N_552);
or U1779 (N_1779,N_300,N_28);
nor U1780 (N_1780,N_276,N_55);
nor U1781 (N_1781,N_952,N_605);
nand U1782 (N_1782,N_44,N_244);
nor U1783 (N_1783,N_200,N_992);
nand U1784 (N_1784,N_821,N_951);
or U1785 (N_1785,N_685,N_303);
or U1786 (N_1786,N_487,N_320);
nand U1787 (N_1787,N_299,N_975);
or U1788 (N_1788,N_981,N_381);
or U1789 (N_1789,N_103,N_891);
nand U1790 (N_1790,N_674,N_97);
nand U1791 (N_1791,N_335,N_141);
nand U1792 (N_1792,N_201,N_831);
nor U1793 (N_1793,N_880,N_303);
nor U1794 (N_1794,N_655,N_844);
nor U1795 (N_1795,N_765,N_209);
nand U1796 (N_1796,N_377,N_100);
or U1797 (N_1797,N_523,N_787);
nor U1798 (N_1798,N_282,N_883);
or U1799 (N_1799,N_468,N_276);
and U1800 (N_1800,N_167,N_529);
and U1801 (N_1801,N_645,N_246);
and U1802 (N_1802,N_367,N_528);
xnor U1803 (N_1803,N_229,N_87);
and U1804 (N_1804,N_811,N_941);
and U1805 (N_1805,N_137,N_967);
nor U1806 (N_1806,N_61,N_502);
and U1807 (N_1807,N_972,N_513);
xnor U1808 (N_1808,N_702,N_741);
nand U1809 (N_1809,N_172,N_296);
nand U1810 (N_1810,N_592,N_711);
and U1811 (N_1811,N_123,N_221);
nand U1812 (N_1812,N_450,N_736);
or U1813 (N_1813,N_693,N_565);
or U1814 (N_1814,N_500,N_888);
nand U1815 (N_1815,N_419,N_907);
nor U1816 (N_1816,N_216,N_188);
nand U1817 (N_1817,N_208,N_7);
nand U1818 (N_1818,N_368,N_621);
nor U1819 (N_1819,N_32,N_287);
nand U1820 (N_1820,N_25,N_78);
nor U1821 (N_1821,N_618,N_398);
and U1822 (N_1822,N_641,N_947);
nand U1823 (N_1823,N_702,N_96);
nor U1824 (N_1824,N_224,N_354);
nor U1825 (N_1825,N_79,N_73);
and U1826 (N_1826,N_322,N_684);
nor U1827 (N_1827,N_351,N_460);
and U1828 (N_1828,N_421,N_422);
nor U1829 (N_1829,N_600,N_613);
nor U1830 (N_1830,N_379,N_609);
nand U1831 (N_1831,N_601,N_735);
nand U1832 (N_1832,N_338,N_284);
or U1833 (N_1833,N_691,N_364);
nor U1834 (N_1834,N_137,N_289);
nor U1835 (N_1835,N_378,N_577);
or U1836 (N_1836,N_970,N_916);
and U1837 (N_1837,N_20,N_351);
nor U1838 (N_1838,N_739,N_191);
nor U1839 (N_1839,N_617,N_191);
nor U1840 (N_1840,N_423,N_701);
nand U1841 (N_1841,N_968,N_911);
nand U1842 (N_1842,N_428,N_892);
nor U1843 (N_1843,N_44,N_397);
and U1844 (N_1844,N_590,N_340);
and U1845 (N_1845,N_582,N_48);
and U1846 (N_1846,N_820,N_612);
nor U1847 (N_1847,N_962,N_335);
and U1848 (N_1848,N_930,N_63);
nor U1849 (N_1849,N_265,N_581);
nand U1850 (N_1850,N_833,N_457);
or U1851 (N_1851,N_120,N_756);
nand U1852 (N_1852,N_627,N_309);
and U1853 (N_1853,N_284,N_738);
nand U1854 (N_1854,N_864,N_210);
or U1855 (N_1855,N_76,N_457);
or U1856 (N_1856,N_610,N_769);
nand U1857 (N_1857,N_861,N_853);
nand U1858 (N_1858,N_967,N_451);
nand U1859 (N_1859,N_880,N_960);
xor U1860 (N_1860,N_59,N_787);
xnor U1861 (N_1861,N_862,N_106);
nor U1862 (N_1862,N_478,N_817);
and U1863 (N_1863,N_447,N_825);
nor U1864 (N_1864,N_12,N_845);
nand U1865 (N_1865,N_909,N_789);
nor U1866 (N_1866,N_995,N_128);
nand U1867 (N_1867,N_196,N_48);
or U1868 (N_1868,N_960,N_664);
and U1869 (N_1869,N_603,N_887);
xnor U1870 (N_1870,N_824,N_895);
nor U1871 (N_1871,N_496,N_907);
and U1872 (N_1872,N_338,N_577);
or U1873 (N_1873,N_594,N_966);
and U1874 (N_1874,N_850,N_852);
and U1875 (N_1875,N_281,N_662);
or U1876 (N_1876,N_329,N_800);
and U1877 (N_1877,N_317,N_980);
nor U1878 (N_1878,N_848,N_793);
nand U1879 (N_1879,N_478,N_147);
or U1880 (N_1880,N_913,N_655);
or U1881 (N_1881,N_458,N_574);
and U1882 (N_1882,N_766,N_236);
nor U1883 (N_1883,N_57,N_600);
or U1884 (N_1884,N_396,N_401);
nor U1885 (N_1885,N_926,N_421);
xor U1886 (N_1886,N_270,N_748);
nor U1887 (N_1887,N_179,N_475);
nand U1888 (N_1888,N_319,N_553);
or U1889 (N_1889,N_412,N_305);
and U1890 (N_1890,N_988,N_745);
or U1891 (N_1891,N_165,N_429);
nor U1892 (N_1892,N_623,N_103);
nand U1893 (N_1893,N_889,N_278);
nor U1894 (N_1894,N_499,N_377);
nand U1895 (N_1895,N_593,N_789);
and U1896 (N_1896,N_477,N_743);
nor U1897 (N_1897,N_720,N_704);
nand U1898 (N_1898,N_459,N_44);
xor U1899 (N_1899,N_960,N_89);
nand U1900 (N_1900,N_761,N_180);
and U1901 (N_1901,N_878,N_59);
and U1902 (N_1902,N_592,N_954);
or U1903 (N_1903,N_679,N_525);
and U1904 (N_1904,N_0,N_460);
nor U1905 (N_1905,N_131,N_71);
and U1906 (N_1906,N_523,N_865);
nor U1907 (N_1907,N_606,N_793);
nand U1908 (N_1908,N_931,N_921);
nor U1909 (N_1909,N_735,N_553);
and U1910 (N_1910,N_583,N_385);
or U1911 (N_1911,N_453,N_230);
nor U1912 (N_1912,N_128,N_248);
or U1913 (N_1913,N_403,N_203);
and U1914 (N_1914,N_412,N_171);
nor U1915 (N_1915,N_719,N_727);
and U1916 (N_1916,N_454,N_119);
or U1917 (N_1917,N_910,N_247);
and U1918 (N_1918,N_428,N_571);
nor U1919 (N_1919,N_971,N_67);
nand U1920 (N_1920,N_758,N_1);
nand U1921 (N_1921,N_970,N_774);
or U1922 (N_1922,N_369,N_848);
nor U1923 (N_1923,N_876,N_621);
nand U1924 (N_1924,N_726,N_46);
or U1925 (N_1925,N_628,N_943);
nand U1926 (N_1926,N_898,N_798);
nand U1927 (N_1927,N_896,N_557);
nand U1928 (N_1928,N_902,N_188);
or U1929 (N_1929,N_232,N_741);
or U1930 (N_1930,N_741,N_78);
nand U1931 (N_1931,N_316,N_835);
nor U1932 (N_1932,N_752,N_220);
or U1933 (N_1933,N_993,N_632);
nand U1934 (N_1934,N_421,N_562);
or U1935 (N_1935,N_232,N_370);
nand U1936 (N_1936,N_602,N_619);
and U1937 (N_1937,N_484,N_974);
or U1938 (N_1938,N_123,N_728);
and U1939 (N_1939,N_183,N_843);
and U1940 (N_1940,N_55,N_935);
nor U1941 (N_1941,N_902,N_737);
nor U1942 (N_1942,N_179,N_642);
nor U1943 (N_1943,N_562,N_336);
nand U1944 (N_1944,N_111,N_859);
nor U1945 (N_1945,N_529,N_737);
nor U1946 (N_1946,N_933,N_831);
nor U1947 (N_1947,N_914,N_39);
and U1948 (N_1948,N_330,N_4);
nand U1949 (N_1949,N_326,N_104);
and U1950 (N_1950,N_790,N_734);
nor U1951 (N_1951,N_159,N_781);
or U1952 (N_1952,N_105,N_41);
and U1953 (N_1953,N_900,N_17);
nand U1954 (N_1954,N_474,N_89);
and U1955 (N_1955,N_707,N_64);
and U1956 (N_1956,N_533,N_771);
and U1957 (N_1957,N_829,N_187);
and U1958 (N_1958,N_404,N_305);
nor U1959 (N_1959,N_297,N_813);
nand U1960 (N_1960,N_792,N_858);
and U1961 (N_1961,N_574,N_611);
nor U1962 (N_1962,N_624,N_844);
nand U1963 (N_1963,N_85,N_666);
and U1964 (N_1964,N_710,N_233);
and U1965 (N_1965,N_513,N_535);
and U1966 (N_1966,N_964,N_339);
nor U1967 (N_1967,N_962,N_893);
and U1968 (N_1968,N_592,N_377);
nor U1969 (N_1969,N_168,N_493);
nor U1970 (N_1970,N_844,N_648);
or U1971 (N_1971,N_995,N_239);
xnor U1972 (N_1972,N_172,N_159);
nand U1973 (N_1973,N_938,N_584);
nor U1974 (N_1974,N_310,N_384);
and U1975 (N_1975,N_795,N_95);
nand U1976 (N_1976,N_996,N_88);
or U1977 (N_1977,N_932,N_208);
nand U1978 (N_1978,N_96,N_257);
or U1979 (N_1979,N_674,N_506);
and U1980 (N_1980,N_583,N_225);
nor U1981 (N_1981,N_654,N_308);
or U1982 (N_1982,N_572,N_892);
nand U1983 (N_1983,N_9,N_308);
or U1984 (N_1984,N_964,N_697);
or U1985 (N_1985,N_577,N_235);
nor U1986 (N_1986,N_731,N_49);
or U1987 (N_1987,N_247,N_930);
nor U1988 (N_1988,N_930,N_203);
nor U1989 (N_1989,N_298,N_374);
nand U1990 (N_1990,N_683,N_55);
or U1991 (N_1991,N_786,N_427);
nand U1992 (N_1992,N_899,N_433);
nor U1993 (N_1993,N_200,N_167);
or U1994 (N_1994,N_652,N_426);
or U1995 (N_1995,N_897,N_920);
nor U1996 (N_1996,N_376,N_432);
nand U1997 (N_1997,N_660,N_142);
and U1998 (N_1998,N_750,N_512);
nor U1999 (N_1999,N_858,N_266);
and U2000 (N_2000,N_1939,N_1078);
nor U2001 (N_2001,N_1179,N_1795);
and U2002 (N_2002,N_1706,N_1432);
nand U2003 (N_2003,N_1354,N_1808);
nor U2004 (N_2004,N_1680,N_1736);
nor U2005 (N_2005,N_1880,N_1642);
nor U2006 (N_2006,N_1957,N_1198);
nand U2007 (N_2007,N_1782,N_1127);
nor U2008 (N_2008,N_1761,N_1787);
and U2009 (N_2009,N_1257,N_1550);
or U2010 (N_2010,N_1340,N_1687);
and U2011 (N_2011,N_1435,N_1363);
nand U2012 (N_2012,N_1730,N_1241);
or U2013 (N_2013,N_1572,N_1816);
nand U2014 (N_2014,N_1597,N_1935);
nor U2015 (N_2015,N_1608,N_1181);
or U2016 (N_2016,N_1359,N_1999);
and U2017 (N_2017,N_1470,N_1058);
nor U2018 (N_2018,N_1892,N_1203);
or U2019 (N_2019,N_1882,N_1881);
and U2020 (N_2020,N_1139,N_1667);
nand U2021 (N_2021,N_1543,N_1475);
nor U2022 (N_2022,N_1765,N_1162);
nor U2023 (N_2023,N_1638,N_1512);
xor U2024 (N_2024,N_1751,N_1073);
or U2025 (N_2025,N_1451,N_1873);
or U2026 (N_2026,N_1352,N_1106);
nand U2027 (N_2027,N_1871,N_1517);
nand U2028 (N_2028,N_1626,N_1226);
xor U2029 (N_2029,N_1801,N_1605);
xor U2030 (N_2030,N_1250,N_1938);
nand U2031 (N_2031,N_1306,N_1773);
nand U2032 (N_2032,N_1911,N_1169);
and U2033 (N_2033,N_1212,N_1615);
xor U2034 (N_2034,N_1423,N_1130);
and U2035 (N_2035,N_1324,N_1217);
nand U2036 (N_2036,N_1546,N_1102);
or U2037 (N_2037,N_1369,N_1184);
or U2038 (N_2038,N_1152,N_1399);
nand U2039 (N_2039,N_1180,N_1850);
and U2040 (N_2040,N_1558,N_1442);
and U2041 (N_2041,N_1658,N_1937);
nand U2042 (N_2042,N_1804,N_1504);
and U2043 (N_2043,N_1523,N_1815);
or U2044 (N_2044,N_1049,N_1720);
nand U2045 (N_2045,N_1270,N_1421);
or U2046 (N_2046,N_1814,N_1068);
or U2047 (N_2047,N_1409,N_1280);
nand U2048 (N_2048,N_1439,N_1383);
or U2049 (N_2049,N_1516,N_1308);
and U2050 (N_2050,N_1894,N_1243);
nand U2051 (N_2051,N_1040,N_1681);
or U2052 (N_2052,N_1271,N_1618);
nand U2053 (N_2053,N_1222,N_1121);
nand U2054 (N_2054,N_1659,N_1066);
nor U2055 (N_2055,N_1603,N_1725);
and U2056 (N_2056,N_1839,N_1144);
nor U2057 (N_2057,N_1494,N_1551);
nand U2058 (N_2058,N_1819,N_1582);
nor U2059 (N_2059,N_1416,N_1207);
nor U2060 (N_2060,N_1900,N_1348);
nor U2061 (N_2061,N_1678,N_1899);
nand U2062 (N_2062,N_1138,N_1006);
and U2063 (N_2063,N_1171,N_1797);
nor U2064 (N_2064,N_1168,N_1836);
or U2065 (N_2065,N_1488,N_1807);
nor U2066 (N_2066,N_1395,N_1933);
and U2067 (N_2067,N_1278,N_1921);
nand U2068 (N_2068,N_1110,N_1499);
nand U2069 (N_2069,N_1994,N_1763);
nand U2070 (N_2070,N_1230,N_1483);
nand U2071 (N_2071,N_1234,N_1617);
and U2072 (N_2072,N_1444,N_1592);
nand U2073 (N_2073,N_1097,N_1657);
nor U2074 (N_2074,N_1347,N_1455);
and U2075 (N_2075,N_1844,N_1920);
xnor U2076 (N_2076,N_1949,N_1780);
and U2077 (N_2077,N_1770,N_1950);
xor U2078 (N_2078,N_1313,N_1150);
and U2079 (N_2079,N_1898,N_1244);
or U2080 (N_2080,N_1232,N_1620);
or U2081 (N_2081,N_1792,N_1785);
nand U2082 (N_2082,N_1974,N_1178);
and U2083 (N_2083,N_1126,N_1426);
or U2084 (N_2084,N_1120,N_1033);
nand U2085 (N_2085,N_1878,N_1365);
and U2086 (N_2086,N_1041,N_1074);
nand U2087 (N_2087,N_1979,N_1134);
nand U2088 (N_2088,N_1132,N_1916);
nand U2089 (N_2089,N_1349,N_1598);
or U2090 (N_2090,N_1298,N_1918);
nand U2091 (N_2091,N_1641,N_1701);
nor U2092 (N_2092,N_1789,N_1849);
nand U2093 (N_2093,N_1374,N_1166);
nand U2094 (N_2094,N_1440,N_1133);
or U2095 (N_2095,N_1404,N_1759);
and U2096 (N_2096,N_1087,N_1955);
or U2097 (N_2097,N_1284,N_1204);
nor U2098 (N_2098,N_1290,N_1755);
nor U2099 (N_2099,N_1427,N_1491);
or U2100 (N_2100,N_1568,N_1584);
and U2101 (N_2101,N_1889,N_1958);
and U2102 (N_2102,N_1748,N_1077);
and U2103 (N_2103,N_1036,N_1414);
or U2104 (N_2104,N_1852,N_1874);
nor U2105 (N_2105,N_1972,N_1535);
or U2106 (N_2106,N_1745,N_1824);
nand U2107 (N_2107,N_1500,N_1925);
or U2108 (N_2108,N_1205,N_1960);
and U2109 (N_2109,N_1868,N_1161);
and U2110 (N_2110,N_1739,N_1345);
and U2111 (N_2111,N_1070,N_1710);
or U2112 (N_2112,N_1406,N_1276);
nor U2113 (N_2113,N_1309,N_1017);
nor U2114 (N_2114,N_1214,N_1413);
nor U2115 (N_2115,N_1740,N_1282);
xnor U2116 (N_2116,N_1614,N_1688);
and U2117 (N_2117,N_1445,N_1832);
or U2118 (N_2118,N_1101,N_1553);
nand U2119 (N_2119,N_1586,N_1624);
or U2120 (N_2120,N_1301,N_1071);
nand U2121 (N_2121,N_1945,N_1754);
nand U2122 (N_2122,N_1197,N_1337);
and U2123 (N_2123,N_1025,N_1677);
or U2124 (N_2124,N_1090,N_1741);
or U2125 (N_2125,N_1587,N_1631);
or U2126 (N_2126,N_1718,N_1987);
nand U2127 (N_2127,N_1990,N_1112);
or U2128 (N_2128,N_1652,N_1331);
and U2129 (N_2129,N_1952,N_1190);
and U2130 (N_2130,N_1764,N_1621);
and U2131 (N_2131,N_1733,N_1788);
nand U2132 (N_2132,N_1569,N_1965);
or U2133 (N_2133,N_1387,N_1928);
xor U2134 (N_2134,N_1859,N_1148);
and U2135 (N_2135,N_1534,N_1183);
or U2136 (N_2136,N_1502,N_1011);
or U2137 (N_2137,N_1325,N_1408);
or U2138 (N_2138,N_1573,N_1342);
and U2139 (N_2139,N_1547,N_1647);
and U2140 (N_2140,N_1526,N_1224);
nand U2141 (N_2141,N_1154,N_1583);
and U2142 (N_2142,N_1842,N_1089);
nor U2143 (N_2143,N_1403,N_1355);
and U2144 (N_2144,N_1312,N_1047);
nand U2145 (N_2145,N_1200,N_1279);
nand U2146 (N_2146,N_1827,N_1570);
and U2147 (N_2147,N_1109,N_1428);
nor U2148 (N_2148,N_1735,N_1307);
or U2149 (N_2149,N_1683,N_1386);
nand U2150 (N_2150,N_1216,N_1564);
nand U2151 (N_2151,N_1825,N_1042);
or U2152 (N_2152,N_1039,N_1784);
or U2153 (N_2153,N_1746,N_1919);
nand U2154 (N_2154,N_1622,N_1732);
nor U2155 (N_2155,N_1867,N_1277);
nor U2156 (N_2156,N_1287,N_1269);
or U2157 (N_2157,N_1895,N_1799);
or U2158 (N_2158,N_1501,N_1668);
nor U2159 (N_2159,N_1100,N_1971);
or U2160 (N_2160,N_1713,N_1976);
or U2161 (N_2161,N_1639,N_1076);
and U2162 (N_2162,N_1989,N_1548);
and U2163 (N_2163,N_1790,N_1015);
nand U2164 (N_2164,N_1385,N_1590);
and U2165 (N_2165,N_1465,N_1258);
and U2166 (N_2166,N_1601,N_1019);
nand U2167 (N_2167,N_1092,N_1061);
xnor U2168 (N_2168,N_1968,N_1973);
nand U2169 (N_2169,N_1752,N_1956);
nor U2170 (N_2170,N_1360,N_1637);
nand U2171 (N_2171,N_1443,N_1646);
or U2172 (N_2172,N_1314,N_1196);
or U2173 (N_2173,N_1020,N_1136);
nand U2174 (N_2174,N_1460,N_1378);
nand U2175 (N_2175,N_1219,N_1125);
nand U2176 (N_2176,N_1487,N_1779);
and U2177 (N_2177,N_1063,N_1757);
nor U2178 (N_2178,N_1293,N_1259);
nor U2179 (N_2179,N_1915,N_1192);
nor U2180 (N_2180,N_1820,N_1239);
or U2181 (N_2181,N_1091,N_1660);
nor U2182 (N_2182,N_1388,N_1265);
nor U2183 (N_2183,N_1519,N_1604);
or U2184 (N_2184,N_1158,N_1209);
or U2185 (N_2185,N_1887,N_1630);
nand U2186 (N_2186,N_1533,N_1984);
and U2187 (N_2187,N_1571,N_1907);
nor U2188 (N_2188,N_1142,N_1817);
nor U2189 (N_2189,N_1610,N_1013);
nor U2190 (N_2190,N_1247,N_1344);
nor U2191 (N_2191,N_1128,N_1469);
nor U2192 (N_2192,N_1145,N_1322);
nor U2193 (N_2193,N_1069,N_1855);
or U2194 (N_2194,N_1143,N_1872);
nand U2195 (N_2195,N_1157,N_1402);
nand U2196 (N_2196,N_1124,N_1530);
nand U2197 (N_2197,N_1320,N_1875);
nand U2198 (N_2198,N_1316,N_1518);
nor U2199 (N_2199,N_1609,N_1381);
and U2200 (N_2200,N_1228,N_1291);
xor U2201 (N_2201,N_1371,N_1458);
nand U2202 (N_2202,N_1245,N_1167);
or U2203 (N_2203,N_1947,N_1311);
and U2204 (N_2204,N_1299,N_1031);
or U2205 (N_2205,N_1351,N_1653);
nor U2206 (N_2206,N_1929,N_1305);
nand U2207 (N_2207,N_1507,N_1537);
nor U2208 (N_2208,N_1461,N_1140);
nand U2209 (N_2209,N_1991,N_1043);
and U2210 (N_2210,N_1430,N_1264);
or U2211 (N_2211,N_1625,N_1865);
or U2212 (N_2212,N_1922,N_1176);
nand U2213 (N_2213,N_1260,N_1699);
and U2214 (N_2214,N_1397,N_1497);
nand U2215 (N_2215,N_1449,N_1159);
and U2216 (N_2216,N_1803,N_1393);
nand U2217 (N_2217,N_1318,N_1317);
nand U2218 (N_2218,N_1493,N_1188);
and U2219 (N_2219,N_1137,N_1229);
nand U2220 (N_2220,N_1712,N_1093);
nand U2221 (N_2221,N_1303,N_1923);
nand U2222 (N_2222,N_1951,N_1786);
nor U2223 (N_2223,N_1525,N_1566);
and U2224 (N_2224,N_1946,N_1187);
or U2225 (N_2225,N_1064,N_1372);
nor U2226 (N_2226,N_1108,N_1080);
nand U2227 (N_2227,N_1753,N_1731);
nand U2228 (N_2228,N_1062,N_1542);
nand U2229 (N_2229,N_1904,N_1422);
or U2230 (N_2230,N_1716,N_1391);
or U2231 (N_2231,N_1116,N_1117);
or U2232 (N_2232,N_1253,N_1705);
or U2233 (N_2233,N_1028,N_1329);
and U2234 (N_2234,N_1480,N_1319);
nor U2235 (N_2235,N_1942,N_1485);
nand U2236 (N_2236,N_1707,N_1001);
nand U2237 (N_2237,N_1811,N_1562);
nor U2238 (N_2238,N_1988,N_1085);
or U2239 (N_2239,N_1629,N_1812);
nand U2240 (N_2240,N_1223,N_1924);
nand U2241 (N_2241,N_1323,N_1632);
nand U2242 (N_2242,N_1088,N_1577);
or U2243 (N_2243,N_1729,N_1709);
and U2244 (N_2244,N_1237,N_1056);
or U2245 (N_2245,N_1723,N_1356);
and U2246 (N_2246,N_1377,N_1415);
and U2247 (N_2247,N_1281,N_1310);
or U2248 (N_2248,N_1823,N_1978);
nand U2249 (N_2249,N_1420,N_1035);
or U2250 (N_2250,N_1453,N_1560);
and U2251 (N_2251,N_1454,N_1541);
nand U2252 (N_2252,N_1338,N_1644);
nand U2253 (N_2253,N_1514,N_1805);
and U2254 (N_2254,N_1103,N_1302);
nand U2255 (N_2255,N_1255,N_1396);
nor U2256 (N_2256,N_1419,N_1696);
nor U2257 (N_2257,N_1682,N_1489);
or U2258 (N_2258,N_1822,N_1877);
and U2259 (N_2259,N_1524,N_1589);
nor U2260 (N_2260,N_1697,N_1781);
nor U2261 (N_2261,N_1131,N_1715);
nand U2262 (N_2262,N_1446,N_1431);
nand U2263 (N_2263,N_1515,N_1595);
nor U2264 (N_2264,N_1633,N_1858);
nand U2265 (N_2265,N_1806,N_1864);
or U2266 (N_2266,N_1686,N_1235);
nor U2267 (N_2267,N_1195,N_1249);
nand U2268 (N_2268,N_1242,N_1719);
nand U2269 (N_2269,N_1208,N_1008);
nor U2270 (N_2270,N_1679,N_1457);
and U2271 (N_2271,N_1540,N_1272);
or U2272 (N_2272,N_1775,N_1410);
nand U2273 (N_2273,N_1472,N_1665);
or U2274 (N_2274,N_1450,N_1151);
and U2275 (N_2275,N_1700,N_1417);
and U2276 (N_2276,N_1045,N_1016);
nor U2277 (N_2277,N_1671,N_1050);
and U2278 (N_2278,N_1390,N_1285);
and U2279 (N_2279,N_1802,N_1173);
or U2280 (N_2280,N_1048,N_1254);
and U2281 (N_2281,N_1766,N_1111);
nor U2282 (N_2282,N_1970,N_1906);
or U2283 (N_2283,N_1714,N_1052);
nor U2284 (N_2284,N_1998,N_1172);
nand U2285 (N_2285,N_1539,N_1645);
and U2286 (N_2286,N_1908,N_1940);
nor U2287 (N_2287,N_1580,N_1901);
nor U2288 (N_2288,N_1495,N_1612);
or U2289 (N_2289,N_1983,N_1010);
nor U2290 (N_2290,N_1896,N_1596);
or U2291 (N_2291,N_1776,N_1563);
nand U2292 (N_2292,N_1777,N_1405);
nand U2293 (N_2293,N_1623,N_1591);
or U2294 (N_2294,N_1655,N_1910);
nand U2295 (N_2295,N_1466,N_1905);
nand U2296 (N_2296,N_1934,N_1611);
nor U2297 (N_2297,N_1220,N_1708);
and U2298 (N_2298,N_1704,N_1012);
nor U2299 (N_2299,N_1467,N_1651);
or U2300 (N_2300,N_1856,N_1155);
nand U2301 (N_2301,N_1462,N_1005);
nor U2302 (N_2302,N_1527,N_1189);
or U2303 (N_2303,N_1554,N_1174);
nor U2304 (N_2304,N_1436,N_1099);
nand U2305 (N_2305,N_1559,N_1857);
nand U2306 (N_2306,N_1756,N_1879);
or U2307 (N_2307,N_1160,N_1883);
nor U2308 (N_2308,N_1376,N_1536);
or U2309 (N_2309,N_1600,N_1456);
or U2310 (N_2310,N_1474,N_1791);
nor U2311 (N_2311,N_1927,N_1296);
and U2312 (N_2312,N_1826,N_1574);
or U2313 (N_2313,N_1818,N_1231);
nand U2314 (N_2314,N_1175,N_1747);
nand U2315 (N_2315,N_1476,N_1698);
nor U2316 (N_2316,N_1201,N_1084);
and U2317 (N_2317,N_1643,N_1486);
nor U2318 (N_2318,N_1967,N_1141);
and U2319 (N_2319,N_1024,N_1441);
nand U2320 (N_2320,N_1105,N_1496);
or U2321 (N_2321,N_1774,N_1424);
nor U2322 (N_2322,N_1521,N_1743);
and U2323 (N_2323,N_1726,N_1627);
nor U2324 (N_2324,N_1002,N_1581);
nor U2325 (N_2325,N_1392,N_1398);
nand U2326 (N_2326,N_1619,N_1966);
nand U2327 (N_2327,N_1297,N_1914);
nand U2328 (N_2328,N_1032,N_1186);
and U2329 (N_2329,N_1863,N_1944);
nor U2330 (N_2330,N_1164,N_1202);
nor U2331 (N_2331,N_1022,N_1588);
and U2332 (N_2332,N_1636,N_1663);
or U2333 (N_2333,N_1593,N_1156);
nor U2334 (N_2334,N_1327,N_1382);
nor U2335 (N_2335,N_1552,N_1594);
and U2336 (N_2336,N_1054,N_1809);
nand U2337 (N_2337,N_1362,N_1350);
or U2338 (N_2338,N_1628,N_1503);
and U2339 (N_2339,N_1650,N_1266);
or U2340 (N_2340,N_1727,N_1007);
and U2341 (N_2341,N_1030,N_1607);
nor U2342 (N_2342,N_1575,N_1407);
and U2343 (N_2343,N_1119,N_1848);
xor U2344 (N_2344,N_1545,N_1912);
nand U2345 (N_2345,N_1676,N_1268);
nand U2346 (N_2346,N_1821,N_1694);
and U2347 (N_2347,N_1263,N_1640);
nor U2348 (N_2348,N_1096,N_1506);
or U2349 (N_2349,N_1165,N_1691);
nor U2350 (N_2350,N_1834,N_1982);
or U2351 (N_2351,N_1029,N_1051);
nor U2352 (N_2352,N_1926,N_1860);
nor U2353 (N_2353,N_1225,N_1885);
nor U2354 (N_2354,N_1578,N_1375);
nand U2355 (N_2355,N_1490,N_1059);
and U2356 (N_2356,N_1634,N_1869);
nand U2357 (N_2357,N_1557,N_1336);
and U2358 (N_2358,N_1902,N_1954);
and U2359 (N_2359,N_1662,N_1693);
and U2360 (N_2360,N_1330,N_1847);
or U2361 (N_2361,N_1086,N_1664);
nor U2362 (N_2362,N_1484,N_1602);
nor U2363 (N_2363,N_1044,N_1962);
and U2364 (N_2364,N_1616,N_1528);
nor U2365 (N_2365,N_1034,N_1037);
and U2366 (N_2366,N_1995,N_1418);
nor U2367 (N_2367,N_1884,N_1018);
and U2368 (N_2368,N_1251,N_1373);
and U2369 (N_2369,N_1288,N_1026);
nand U2370 (N_2370,N_1561,N_1749);
nand U2371 (N_2371,N_1837,N_1447);
nand U2372 (N_2372,N_1931,N_1300);
or U2373 (N_2373,N_1964,N_1959);
or U2374 (N_2374,N_1233,N_1104);
nand U2375 (N_2375,N_1835,N_1193);
or U2376 (N_2376,N_1674,N_1082);
or U2377 (N_2377,N_1843,N_1332);
nor U2378 (N_2378,N_1492,N_1221);
or U2379 (N_2379,N_1380,N_1838);
nand U2380 (N_2380,N_1948,N_1256);
nor U2381 (N_2381,N_1685,N_1742);
nand U2382 (N_2382,N_1509,N_1115);
nand U2383 (N_2383,N_1913,N_1648);
or U2384 (N_2384,N_1851,N_1210);
or U2385 (N_2385,N_1544,N_1997);
and U2386 (N_2386,N_1796,N_1023);
nand U2387 (N_2387,N_1315,N_1464);
and U2388 (N_2388,N_1163,N_1118);
and U2389 (N_2389,N_1936,N_1890);
and U2390 (N_2390,N_1370,N_1334);
nand U2391 (N_2391,N_1072,N_1961);
nand U2392 (N_2392,N_1888,N_1829);
or U2393 (N_2393,N_1767,N_1149);
xnor U2394 (N_2394,N_1567,N_1861);
or U2395 (N_2395,N_1830,N_1692);
nand U2396 (N_2396,N_1075,N_1576);
and U2397 (N_2397,N_1146,N_1666);
nand U2398 (N_2398,N_1341,N_1909);
nor U2399 (N_2399,N_1262,N_1695);
nand U2400 (N_2400,N_1147,N_1452);
nor U2401 (N_2401,N_1425,N_1943);
or U2402 (N_2402,N_1672,N_1194);
or U2403 (N_2403,N_1981,N_1122);
and U2404 (N_2404,N_1903,N_1252);
xor U2405 (N_2405,N_1434,N_1177);
nor U2406 (N_2406,N_1478,N_1283);
or U2407 (N_2407,N_1538,N_1286);
and U2408 (N_2408,N_1346,N_1364);
or U2409 (N_2409,N_1661,N_1236);
and U2410 (N_2410,N_1227,N_1366);
nand U2411 (N_2411,N_1841,N_1482);
and U2412 (N_2412,N_1673,N_1459);
and U2413 (N_2413,N_1379,N_1897);
and U2414 (N_2414,N_1793,N_1060);
nor U2415 (N_2415,N_1339,N_1170);
and U2416 (N_2416,N_1734,N_1840);
and U2417 (N_2417,N_1513,N_1199);
or U2418 (N_2418,N_1750,N_1702);
nor U2419 (N_2419,N_1599,N_1772);
nor U2420 (N_2420,N_1046,N_1508);
and U2421 (N_2421,N_1684,N_1182);
or U2422 (N_2422,N_1003,N_1505);
xor U2423 (N_2423,N_1274,N_1289);
nor U2424 (N_2424,N_1367,N_1891);
or U2425 (N_2425,N_1304,N_1738);
nor U2426 (N_2426,N_1246,N_1649);
nand U2427 (N_2427,N_1448,N_1328);
and U2428 (N_2428,N_1930,N_1401);
nor U2429 (N_2429,N_1992,N_1703);
or U2430 (N_2430,N_1481,N_1326);
and U2431 (N_2431,N_1980,N_1565);
nand U2432 (N_2432,N_1275,N_1079);
nor U2433 (N_2433,N_1211,N_1768);
nand U2434 (N_2434,N_1067,N_1009);
or U2435 (N_2435,N_1675,N_1218);
or U2436 (N_2436,N_1065,N_1267);
or U2437 (N_2437,N_1261,N_1057);
nor U2438 (N_2438,N_1853,N_1654);
nor U2439 (N_2439,N_1081,N_1532);
nor U2440 (N_2440,N_1000,N_1555);
nand U2441 (N_2441,N_1027,N_1737);
nor U2442 (N_2442,N_1511,N_1353);
nor U2443 (N_2443,N_1917,N_1129);
nor U2444 (N_2444,N_1831,N_1095);
or U2445 (N_2445,N_1969,N_1021);
nor U2446 (N_2446,N_1473,N_1744);
nand U2447 (N_2447,N_1690,N_1014);
and U2448 (N_2448,N_1986,N_1670);
and U2449 (N_2449,N_1114,N_1977);
and U2450 (N_2450,N_1728,N_1669);
and U2451 (N_2451,N_1498,N_1556);
xor U2452 (N_2452,N_1606,N_1724);
nor U2453 (N_2453,N_1053,N_1238);
nor U2454 (N_2454,N_1522,N_1479);
and U2455 (N_2455,N_1993,N_1721);
nand U2456 (N_2456,N_1876,N_1463);
or U2457 (N_2457,N_1361,N_1711);
nand U2458 (N_2458,N_1866,N_1384);
and U2459 (N_2459,N_1333,N_1813);
and U2460 (N_2460,N_1429,N_1004);
nor U2461 (N_2461,N_1794,N_1240);
nand U2462 (N_2462,N_1038,N_1579);
nor U2463 (N_2463,N_1335,N_1689);
and U2464 (N_2464,N_1098,N_1531);
or U2465 (N_2465,N_1549,N_1292);
nand U2466 (N_2466,N_1758,N_1358);
or U2467 (N_2467,N_1438,N_1113);
nand U2468 (N_2468,N_1471,N_1294);
and U2469 (N_2469,N_1191,N_1389);
nor U2470 (N_2470,N_1778,N_1783);
nand U2471 (N_2471,N_1394,N_1055);
and U2472 (N_2472,N_1932,N_1833);
nand U2473 (N_2473,N_1762,N_1321);
nor U2474 (N_2474,N_1343,N_1635);
nor U2475 (N_2475,N_1963,N_1510);
nor U2476 (N_2476,N_1529,N_1094);
and U2477 (N_2477,N_1845,N_1717);
nand U2478 (N_2478,N_1135,N_1886);
and U2479 (N_2479,N_1828,N_1862);
and U2480 (N_2480,N_1411,N_1760);
or U2481 (N_2481,N_1585,N_1215);
or U2482 (N_2482,N_1722,N_1941);
or U2483 (N_2483,N_1975,N_1213);
or U2484 (N_2484,N_1412,N_1870);
nand U2485 (N_2485,N_1893,N_1357);
and U2486 (N_2486,N_1185,N_1769);
nand U2487 (N_2487,N_1810,N_1368);
nor U2488 (N_2488,N_1206,N_1153);
or U2489 (N_2489,N_1433,N_1854);
and U2490 (N_2490,N_1437,N_1985);
nor U2491 (N_2491,N_1468,N_1477);
or U2492 (N_2492,N_1123,N_1295);
nand U2493 (N_2493,N_1771,N_1846);
and U2494 (N_2494,N_1083,N_1656);
and U2495 (N_2495,N_1107,N_1613);
and U2496 (N_2496,N_1996,N_1953);
and U2497 (N_2497,N_1273,N_1800);
and U2498 (N_2498,N_1248,N_1520);
and U2499 (N_2499,N_1798,N_1400);
nand U2500 (N_2500,N_1211,N_1654);
and U2501 (N_2501,N_1341,N_1759);
and U2502 (N_2502,N_1624,N_1858);
and U2503 (N_2503,N_1164,N_1852);
nand U2504 (N_2504,N_1758,N_1849);
and U2505 (N_2505,N_1219,N_1332);
or U2506 (N_2506,N_1002,N_1795);
and U2507 (N_2507,N_1151,N_1193);
or U2508 (N_2508,N_1746,N_1819);
and U2509 (N_2509,N_1415,N_1080);
nand U2510 (N_2510,N_1439,N_1014);
nor U2511 (N_2511,N_1764,N_1898);
nor U2512 (N_2512,N_1814,N_1470);
and U2513 (N_2513,N_1672,N_1205);
or U2514 (N_2514,N_1067,N_1991);
or U2515 (N_2515,N_1224,N_1290);
nor U2516 (N_2516,N_1440,N_1575);
or U2517 (N_2517,N_1440,N_1979);
nor U2518 (N_2518,N_1990,N_1713);
and U2519 (N_2519,N_1681,N_1462);
and U2520 (N_2520,N_1039,N_1131);
nand U2521 (N_2521,N_1516,N_1525);
xor U2522 (N_2522,N_1434,N_1429);
or U2523 (N_2523,N_1844,N_1751);
or U2524 (N_2524,N_1483,N_1226);
nor U2525 (N_2525,N_1777,N_1657);
and U2526 (N_2526,N_1192,N_1725);
nand U2527 (N_2527,N_1670,N_1460);
and U2528 (N_2528,N_1049,N_1482);
nor U2529 (N_2529,N_1018,N_1065);
or U2530 (N_2530,N_1921,N_1458);
nand U2531 (N_2531,N_1739,N_1053);
nor U2532 (N_2532,N_1637,N_1757);
nand U2533 (N_2533,N_1880,N_1211);
and U2534 (N_2534,N_1247,N_1048);
and U2535 (N_2535,N_1487,N_1142);
nand U2536 (N_2536,N_1460,N_1270);
or U2537 (N_2537,N_1869,N_1312);
nor U2538 (N_2538,N_1151,N_1582);
nor U2539 (N_2539,N_1894,N_1039);
and U2540 (N_2540,N_1994,N_1636);
or U2541 (N_2541,N_1383,N_1380);
or U2542 (N_2542,N_1371,N_1924);
nand U2543 (N_2543,N_1810,N_1265);
and U2544 (N_2544,N_1036,N_1889);
or U2545 (N_2545,N_1138,N_1451);
or U2546 (N_2546,N_1113,N_1772);
nand U2547 (N_2547,N_1682,N_1828);
and U2548 (N_2548,N_1909,N_1580);
and U2549 (N_2549,N_1530,N_1203);
nor U2550 (N_2550,N_1861,N_1489);
nor U2551 (N_2551,N_1516,N_1094);
nand U2552 (N_2552,N_1654,N_1206);
nor U2553 (N_2553,N_1431,N_1945);
or U2554 (N_2554,N_1941,N_1466);
and U2555 (N_2555,N_1927,N_1668);
or U2556 (N_2556,N_1525,N_1405);
or U2557 (N_2557,N_1614,N_1547);
and U2558 (N_2558,N_1696,N_1431);
nand U2559 (N_2559,N_1637,N_1058);
and U2560 (N_2560,N_1723,N_1320);
nand U2561 (N_2561,N_1073,N_1695);
nand U2562 (N_2562,N_1336,N_1038);
nand U2563 (N_2563,N_1221,N_1507);
and U2564 (N_2564,N_1494,N_1071);
nor U2565 (N_2565,N_1459,N_1550);
and U2566 (N_2566,N_1646,N_1685);
or U2567 (N_2567,N_1354,N_1710);
nor U2568 (N_2568,N_1089,N_1426);
or U2569 (N_2569,N_1022,N_1728);
or U2570 (N_2570,N_1140,N_1296);
nand U2571 (N_2571,N_1919,N_1467);
xor U2572 (N_2572,N_1773,N_1354);
nand U2573 (N_2573,N_1303,N_1059);
and U2574 (N_2574,N_1393,N_1415);
nand U2575 (N_2575,N_1235,N_1140);
nand U2576 (N_2576,N_1306,N_1438);
or U2577 (N_2577,N_1370,N_1181);
nand U2578 (N_2578,N_1090,N_1635);
and U2579 (N_2579,N_1695,N_1367);
and U2580 (N_2580,N_1119,N_1545);
or U2581 (N_2581,N_1441,N_1019);
and U2582 (N_2582,N_1737,N_1720);
nor U2583 (N_2583,N_1792,N_1182);
and U2584 (N_2584,N_1127,N_1349);
nor U2585 (N_2585,N_1518,N_1046);
or U2586 (N_2586,N_1795,N_1604);
nand U2587 (N_2587,N_1376,N_1117);
or U2588 (N_2588,N_1970,N_1524);
and U2589 (N_2589,N_1215,N_1764);
or U2590 (N_2590,N_1833,N_1903);
or U2591 (N_2591,N_1499,N_1736);
nor U2592 (N_2592,N_1840,N_1169);
nand U2593 (N_2593,N_1553,N_1869);
or U2594 (N_2594,N_1318,N_1658);
nor U2595 (N_2595,N_1264,N_1305);
or U2596 (N_2596,N_1037,N_1430);
nor U2597 (N_2597,N_1949,N_1948);
nor U2598 (N_2598,N_1410,N_1425);
or U2599 (N_2599,N_1969,N_1803);
nor U2600 (N_2600,N_1712,N_1708);
nand U2601 (N_2601,N_1207,N_1656);
nor U2602 (N_2602,N_1226,N_1996);
nor U2603 (N_2603,N_1066,N_1838);
nand U2604 (N_2604,N_1925,N_1744);
nand U2605 (N_2605,N_1906,N_1844);
nand U2606 (N_2606,N_1652,N_1866);
nand U2607 (N_2607,N_1341,N_1331);
nand U2608 (N_2608,N_1546,N_1357);
nand U2609 (N_2609,N_1342,N_1698);
xnor U2610 (N_2610,N_1719,N_1627);
or U2611 (N_2611,N_1408,N_1128);
nand U2612 (N_2612,N_1592,N_1668);
nand U2613 (N_2613,N_1495,N_1276);
and U2614 (N_2614,N_1061,N_1197);
nor U2615 (N_2615,N_1568,N_1487);
nor U2616 (N_2616,N_1512,N_1618);
and U2617 (N_2617,N_1250,N_1077);
or U2618 (N_2618,N_1213,N_1019);
and U2619 (N_2619,N_1509,N_1202);
nand U2620 (N_2620,N_1921,N_1636);
nor U2621 (N_2621,N_1755,N_1702);
or U2622 (N_2622,N_1857,N_1475);
nand U2623 (N_2623,N_1728,N_1122);
nand U2624 (N_2624,N_1659,N_1504);
and U2625 (N_2625,N_1641,N_1891);
nand U2626 (N_2626,N_1977,N_1683);
nand U2627 (N_2627,N_1431,N_1565);
and U2628 (N_2628,N_1079,N_1226);
and U2629 (N_2629,N_1205,N_1339);
and U2630 (N_2630,N_1252,N_1676);
nor U2631 (N_2631,N_1063,N_1337);
and U2632 (N_2632,N_1119,N_1444);
and U2633 (N_2633,N_1725,N_1904);
nor U2634 (N_2634,N_1739,N_1789);
nor U2635 (N_2635,N_1998,N_1766);
or U2636 (N_2636,N_1762,N_1388);
nand U2637 (N_2637,N_1081,N_1070);
nor U2638 (N_2638,N_1297,N_1764);
or U2639 (N_2639,N_1699,N_1248);
nand U2640 (N_2640,N_1974,N_1233);
or U2641 (N_2641,N_1315,N_1137);
or U2642 (N_2642,N_1626,N_1135);
and U2643 (N_2643,N_1045,N_1155);
and U2644 (N_2644,N_1758,N_1088);
nand U2645 (N_2645,N_1567,N_1943);
or U2646 (N_2646,N_1133,N_1515);
or U2647 (N_2647,N_1765,N_1560);
xor U2648 (N_2648,N_1573,N_1692);
nand U2649 (N_2649,N_1905,N_1026);
and U2650 (N_2650,N_1479,N_1893);
or U2651 (N_2651,N_1844,N_1694);
nor U2652 (N_2652,N_1762,N_1047);
or U2653 (N_2653,N_1752,N_1078);
nor U2654 (N_2654,N_1424,N_1422);
nor U2655 (N_2655,N_1026,N_1996);
and U2656 (N_2656,N_1520,N_1435);
or U2657 (N_2657,N_1061,N_1193);
nand U2658 (N_2658,N_1545,N_1403);
nand U2659 (N_2659,N_1658,N_1675);
and U2660 (N_2660,N_1341,N_1023);
nor U2661 (N_2661,N_1190,N_1878);
and U2662 (N_2662,N_1415,N_1322);
nand U2663 (N_2663,N_1065,N_1617);
nand U2664 (N_2664,N_1479,N_1664);
nor U2665 (N_2665,N_1704,N_1811);
and U2666 (N_2666,N_1031,N_1138);
or U2667 (N_2667,N_1491,N_1908);
or U2668 (N_2668,N_1310,N_1219);
nand U2669 (N_2669,N_1107,N_1791);
and U2670 (N_2670,N_1390,N_1666);
nor U2671 (N_2671,N_1476,N_1200);
and U2672 (N_2672,N_1366,N_1744);
nand U2673 (N_2673,N_1707,N_1187);
and U2674 (N_2674,N_1279,N_1280);
nor U2675 (N_2675,N_1054,N_1343);
xor U2676 (N_2676,N_1870,N_1760);
or U2677 (N_2677,N_1384,N_1578);
xnor U2678 (N_2678,N_1673,N_1597);
and U2679 (N_2679,N_1301,N_1436);
nand U2680 (N_2680,N_1897,N_1087);
nor U2681 (N_2681,N_1204,N_1902);
or U2682 (N_2682,N_1736,N_1221);
or U2683 (N_2683,N_1545,N_1612);
and U2684 (N_2684,N_1496,N_1860);
nand U2685 (N_2685,N_1730,N_1268);
or U2686 (N_2686,N_1831,N_1903);
nand U2687 (N_2687,N_1507,N_1268);
nor U2688 (N_2688,N_1073,N_1450);
or U2689 (N_2689,N_1474,N_1812);
nand U2690 (N_2690,N_1048,N_1320);
nand U2691 (N_2691,N_1025,N_1880);
and U2692 (N_2692,N_1069,N_1071);
or U2693 (N_2693,N_1568,N_1199);
nor U2694 (N_2694,N_1002,N_1872);
or U2695 (N_2695,N_1917,N_1480);
nor U2696 (N_2696,N_1331,N_1649);
nand U2697 (N_2697,N_1297,N_1776);
nor U2698 (N_2698,N_1335,N_1251);
nand U2699 (N_2699,N_1367,N_1485);
or U2700 (N_2700,N_1886,N_1805);
nand U2701 (N_2701,N_1966,N_1000);
nand U2702 (N_2702,N_1374,N_1217);
or U2703 (N_2703,N_1464,N_1185);
and U2704 (N_2704,N_1006,N_1508);
nand U2705 (N_2705,N_1045,N_1463);
and U2706 (N_2706,N_1689,N_1723);
nand U2707 (N_2707,N_1482,N_1490);
or U2708 (N_2708,N_1614,N_1523);
or U2709 (N_2709,N_1092,N_1563);
nand U2710 (N_2710,N_1021,N_1515);
and U2711 (N_2711,N_1948,N_1691);
nor U2712 (N_2712,N_1425,N_1558);
nor U2713 (N_2713,N_1514,N_1192);
and U2714 (N_2714,N_1094,N_1258);
nand U2715 (N_2715,N_1642,N_1092);
nand U2716 (N_2716,N_1882,N_1931);
nand U2717 (N_2717,N_1590,N_1011);
and U2718 (N_2718,N_1375,N_1376);
and U2719 (N_2719,N_1668,N_1060);
and U2720 (N_2720,N_1350,N_1919);
or U2721 (N_2721,N_1102,N_1780);
nor U2722 (N_2722,N_1302,N_1479);
and U2723 (N_2723,N_1319,N_1726);
nor U2724 (N_2724,N_1110,N_1848);
nand U2725 (N_2725,N_1775,N_1794);
xor U2726 (N_2726,N_1835,N_1041);
nor U2727 (N_2727,N_1553,N_1843);
nor U2728 (N_2728,N_1677,N_1089);
nand U2729 (N_2729,N_1235,N_1906);
or U2730 (N_2730,N_1069,N_1546);
nor U2731 (N_2731,N_1406,N_1792);
and U2732 (N_2732,N_1932,N_1023);
nor U2733 (N_2733,N_1402,N_1785);
nor U2734 (N_2734,N_1531,N_1104);
nand U2735 (N_2735,N_1265,N_1831);
or U2736 (N_2736,N_1529,N_1421);
nor U2737 (N_2737,N_1046,N_1276);
or U2738 (N_2738,N_1787,N_1407);
and U2739 (N_2739,N_1764,N_1697);
nand U2740 (N_2740,N_1740,N_1051);
nand U2741 (N_2741,N_1395,N_1799);
or U2742 (N_2742,N_1794,N_1515);
or U2743 (N_2743,N_1564,N_1764);
or U2744 (N_2744,N_1214,N_1583);
nor U2745 (N_2745,N_1311,N_1993);
nor U2746 (N_2746,N_1724,N_1401);
nand U2747 (N_2747,N_1550,N_1227);
nor U2748 (N_2748,N_1130,N_1560);
nand U2749 (N_2749,N_1507,N_1041);
nor U2750 (N_2750,N_1155,N_1698);
or U2751 (N_2751,N_1192,N_1461);
and U2752 (N_2752,N_1555,N_1660);
nand U2753 (N_2753,N_1421,N_1111);
nor U2754 (N_2754,N_1392,N_1722);
and U2755 (N_2755,N_1884,N_1720);
nand U2756 (N_2756,N_1634,N_1098);
nor U2757 (N_2757,N_1509,N_1634);
nor U2758 (N_2758,N_1052,N_1802);
nor U2759 (N_2759,N_1907,N_1769);
or U2760 (N_2760,N_1060,N_1495);
or U2761 (N_2761,N_1611,N_1727);
or U2762 (N_2762,N_1823,N_1986);
nor U2763 (N_2763,N_1419,N_1603);
nor U2764 (N_2764,N_1156,N_1068);
nor U2765 (N_2765,N_1704,N_1534);
nor U2766 (N_2766,N_1401,N_1919);
or U2767 (N_2767,N_1715,N_1868);
nand U2768 (N_2768,N_1693,N_1940);
nand U2769 (N_2769,N_1620,N_1446);
or U2770 (N_2770,N_1637,N_1735);
or U2771 (N_2771,N_1008,N_1163);
nor U2772 (N_2772,N_1630,N_1645);
and U2773 (N_2773,N_1568,N_1620);
nand U2774 (N_2774,N_1947,N_1405);
or U2775 (N_2775,N_1755,N_1639);
xor U2776 (N_2776,N_1286,N_1577);
nor U2777 (N_2777,N_1865,N_1383);
or U2778 (N_2778,N_1769,N_1058);
nand U2779 (N_2779,N_1557,N_1966);
nor U2780 (N_2780,N_1591,N_1989);
and U2781 (N_2781,N_1135,N_1903);
nand U2782 (N_2782,N_1283,N_1078);
nand U2783 (N_2783,N_1398,N_1725);
nand U2784 (N_2784,N_1139,N_1527);
nand U2785 (N_2785,N_1871,N_1605);
nand U2786 (N_2786,N_1356,N_1043);
or U2787 (N_2787,N_1018,N_1496);
nor U2788 (N_2788,N_1480,N_1048);
and U2789 (N_2789,N_1238,N_1493);
nor U2790 (N_2790,N_1423,N_1903);
nor U2791 (N_2791,N_1653,N_1178);
nand U2792 (N_2792,N_1776,N_1030);
nand U2793 (N_2793,N_1195,N_1395);
nand U2794 (N_2794,N_1570,N_1528);
or U2795 (N_2795,N_1913,N_1224);
or U2796 (N_2796,N_1147,N_1278);
and U2797 (N_2797,N_1559,N_1218);
and U2798 (N_2798,N_1576,N_1906);
nor U2799 (N_2799,N_1464,N_1118);
and U2800 (N_2800,N_1896,N_1122);
or U2801 (N_2801,N_1521,N_1784);
and U2802 (N_2802,N_1505,N_1814);
and U2803 (N_2803,N_1590,N_1580);
and U2804 (N_2804,N_1483,N_1332);
nand U2805 (N_2805,N_1525,N_1981);
nand U2806 (N_2806,N_1859,N_1558);
and U2807 (N_2807,N_1476,N_1187);
nand U2808 (N_2808,N_1536,N_1750);
nand U2809 (N_2809,N_1536,N_1322);
or U2810 (N_2810,N_1342,N_1251);
nand U2811 (N_2811,N_1970,N_1170);
or U2812 (N_2812,N_1210,N_1695);
nand U2813 (N_2813,N_1405,N_1866);
and U2814 (N_2814,N_1818,N_1718);
nor U2815 (N_2815,N_1933,N_1251);
or U2816 (N_2816,N_1545,N_1017);
xor U2817 (N_2817,N_1046,N_1215);
or U2818 (N_2818,N_1750,N_1759);
nor U2819 (N_2819,N_1727,N_1819);
nor U2820 (N_2820,N_1000,N_1314);
or U2821 (N_2821,N_1754,N_1328);
or U2822 (N_2822,N_1145,N_1649);
and U2823 (N_2823,N_1335,N_1494);
and U2824 (N_2824,N_1735,N_1708);
and U2825 (N_2825,N_1449,N_1440);
nor U2826 (N_2826,N_1811,N_1646);
nand U2827 (N_2827,N_1648,N_1458);
or U2828 (N_2828,N_1630,N_1141);
nor U2829 (N_2829,N_1727,N_1989);
and U2830 (N_2830,N_1237,N_1890);
and U2831 (N_2831,N_1710,N_1157);
nand U2832 (N_2832,N_1732,N_1825);
nor U2833 (N_2833,N_1466,N_1841);
and U2834 (N_2834,N_1510,N_1297);
and U2835 (N_2835,N_1972,N_1492);
or U2836 (N_2836,N_1903,N_1065);
and U2837 (N_2837,N_1159,N_1174);
and U2838 (N_2838,N_1253,N_1446);
and U2839 (N_2839,N_1682,N_1583);
and U2840 (N_2840,N_1492,N_1794);
nor U2841 (N_2841,N_1257,N_1562);
or U2842 (N_2842,N_1055,N_1106);
or U2843 (N_2843,N_1952,N_1734);
nor U2844 (N_2844,N_1010,N_1163);
nand U2845 (N_2845,N_1692,N_1448);
or U2846 (N_2846,N_1288,N_1220);
or U2847 (N_2847,N_1799,N_1726);
nand U2848 (N_2848,N_1734,N_1077);
and U2849 (N_2849,N_1729,N_1465);
and U2850 (N_2850,N_1170,N_1487);
nor U2851 (N_2851,N_1212,N_1994);
nand U2852 (N_2852,N_1698,N_1206);
nand U2853 (N_2853,N_1810,N_1914);
nand U2854 (N_2854,N_1421,N_1452);
nand U2855 (N_2855,N_1760,N_1315);
or U2856 (N_2856,N_1162,N_1883);
nor U2857 (N_2857,N_1762,N_1203);
or U2858 (N_2858,N_1109,N_1090);
nor U2859 (N_2859,N_1311,N_1874);
xnor U2860 (N_2860,N_1714,N_1285);
nor U2861 (N_2861,N_1432,N_1714);
nor U2862 (N_2862,N_1988,N_1195);
nand U2863 (N_2863,N_1490,N_1045);
nor U2864 (N_2864,N_1059,N_1697);
nor U2865 (N_2865,N_1287,N_1082);
or U2866 (N_2866,N_1960,N_1620);
or U2867 (N_2867,N_1926,N_1012);
or U2868 (N_2868,N_1924,N_1673);
nand U2869 (N_2869,N_1580,N_1822);
nor U2870 (N_2870,N_1027,N_1408);
and U2871 (N_2871,N_1483,N_1661);
and U2872 (N_2872,N_1560,N_1864);
nor U2873 (N_2873,N_1683,N_1627);
and U2874 (N_2874,N_1159,N_1413);
nor U2875 (N_2875,N_1791,N_1441);
nor U2876 (N_2876,N_1519,N_1695);
and U2877 (N_2877,N_1571,N_1769);
and U2878 (N_2878,N_1381,N_1895);
nor U2879 (N_2879,N_1010,N_1443);
xor U2880 (N_2880,N_1089,N_1273);
and U2881 (N_2881,N_1407,N_1863);
and U2882 (N_2882,N_1767,N_1439);
nor U2883 (N_2883,N_1264,N_1401);
nand U2884 (N_2884,N_1628,N_1529);
nor U2885 (N_2885,N_1938,N_1162);
and U2886 (N_2886,N_1060,N_1776);
or U2887 (N_2887,N_1108,N_1572);
nor U2888 (N_2888,N_1927,N_1297);
nor U2889 (N_2889,N_1324,N_1479);
nand U2890 (N_2890,N_1853,N_1841);
and U2891 (N_2891,N_1831,N_1192);
or U2892 (N_2892,N_1502,N_1110);
nand U2893 (N_2893,N_1720,N_1847);
or U2894 (N_2894,N_1549,N_1784);
xor U2895 (N_2895,N_1578,N_1936);
or U2896 (N_2896,N_1624,N_1275);
nand U2897 (N_2897,N_1948,N_1828);
nor U2898 (N_2898,N_1106,N_1514);
xor U2899 (N_2899,N_1169,N_1588);
nor U2900 (N_2900,N_1287,N_1185);
or U2901 (N_2901,N_1040,N_1212);
nor U2902 (N_2902,N_1764,N_1531);
and U2903 (N_2903,N_1861,N_1867);
nor U2904 (N_2904,N_1935,N_1458);
and U2905 (N_2905,N_1737,N_1552);
and U2906 (N_2906,N_1757,N_1542);
or U2907 (N_2907,N_1020,N_1110);
and U2908 (N_2908,N_1019,N_1183);
and U2909 (N_2909,N_1121,N_1710);
nor U2910 (N_2910,N_1987,N_1595);
nor U2911 (N_2911,N_1951,N_1443);
nand U2912 (N_2912,N_1536,N_1957);
xnor U2913 (N_2913,N_1843,N_1718);
nor U2914 (N_2914,N_1823,N_1458);
nand U2915 (N_2915,N_1943,N_1162);
and U2916 (N_2916,N_1528,N_1858);
or U2917 (N_2917,N_1363,N_1911);
or U2918 (N_2918,N_1634,N_1870);
nand U2919 (N_2919,N_1742,N_1848);
or U2920 (N_2920,N_1264,N_1382);
nor U2921 (N_2921,N_1790,N_1056);
or U2922 (N_2922,N_1131,N_1763);
nor U2923 (N_2923,N_1025,N_1834);
and U2924 (N_2924,N_1287,N_1995);
nor U2925 (N_2925,N_1357,N_1655);
nand U2926 (N_2926,N_1498,N_1382);
or U2927 (N_2927,N_1248,N_1640);
nand U2928 (N_2928,N_1198,N_1707);
and U2929 (N_2929,N_1190,N_1855);
or U2930 (N_2930,N_1351,N_1066);
nand U2931 (N_2931,N_1334,N_1349);
or U2932 (N_2932,N_1942,N_1795);
nor U2933 (N_2933,N_1853,N_1295);
or U2934 (N_2934,N_1594,N_1880);
and U2935 (N_2935,N_1119,N_1443);
nand U2936 (N_2936,N_1669,N_1696);
or U2937 (N_2937,N_1842,N_1232);
xnor U2938 (N_2938,N_1542,N_1416);
nor U2939 (N_2939,N_1875,N_1922);
and U2940 (N_2940,N_1766,N_1570);
or U2941 (N_2941,N_1165,N_1823);
and U2942 (N_2942,N_1231,N_1183);
and U2943 (N_2943,N_1062,N_1633);
or U2944 (N_2944,N_1527,N_1740);
nor U2945 (N_2945,N_1013,N_1615);
nand U2946 (N_2946,N_1834,N_1026);
nand U2947 (N_2947,N_1716,N_1539);
xor U2948 (N_2948,N_1758,N_1061);
nand U2949 (N_2949,N_1615,N_1873);
nor U2950 (N_2950,N_1770,N_1608);
or U2951 (N_2951,N_1566,N_1325);
and U2952 (N_2952,N_1948,N_1951);
and U2953 (N_2953,N_1656,N_1116);
or U2954 (N_2954,N_1067,N_1907);
nor U2955 (N_2955,N_1295,N_1260);
and U2956 (N_2956,N_1992,N_1705);
or U2957 (N_2957,N_1518,N_1274);
nor U2958 (N_2958,N_1777,N_1528);
xnor U2959 (N_2959,N_1398,N_1643);
or U2960 (N_2960,N_1524,N_1460);
nor U2961 (N_2961,N_1808,N_1302);
nor U2962 (N_2962,N_1664,N_1061);
nor U2963 (N_2963,N_1484,N_1808);
nor U2964 (N_2964,N_1257,N_1402);
and U2965 (N_2965,N_1629,N_1576);
nor U2966 (N_2966,N_1414,N_1584);
or U2967 (N_2967,N_1157,N_1859);
or U2968 (N_2968,N_1760,N_1003);
or U2969 (N_2969,N_1643,N_1640);
and U2970 (N_2970,N_1259,N_1694);
and U2971 (N_2971,N_1437,N_1138);
nand U2972 (N_2972,N_1349,N_1980);
and U2973 (N_2973,N_1192,N_1651);
nand U2974 (N_2974,N_1343,N_1986);
or U2975 (N_2975,N_1568,N_1052);
and U2976 (N_2976,N_1969,N_1089);
and U2977 (N_2977,N_1896,N_1228);
and U2978 (N_2978,N_1353,N_1865);
or U2979 (N_2979,N_1099,N_1964);
nor U2980 (N_2980,N_1807,N_1402);
nand U2981 (N_2981,N_1943,N_1627);
nand U2982 (N_2982,N_1107,N_1740);
nor U2983 (N_2983,N_1399,N_1506);
or U2984 (N_2984,N_1541,N_1321);
or U2985 (N_2985,N_1235,N_1479);
and U2986 (N_2986,N_1764,N_1061);
nand U2987 (N_2987,N_1856,N_1551);
nand U2988 (N_2988,N_1182,N_1977);
nand U2989 (N_2989,N_1785,N_1218);
nor U2990 (N_2990,N_1033,N_1495);
nor U2991 (N_2991,N_1099,N_1810);
nor U2992 (N_2992,N_1120,N_1046);
and U2993 (N_2993,N_1237,N_1004);
or U2994 (N_2994,N_1704,N_1105);
nand U2995 (N_2995,N_1878,N_1313);
and U2996 (N_2996,N_1353,N_1482);
or U2997 (N_2997,N_1677,N_1223);
nand U2998 (N_2998,N_1583,N_1055);
nor U2999 (N_2999,N_1815,N_1754);
nand U3000 (N_3000,N_2652,N_2536);
or U3001 (N_3001,N_2722,N_2811);
nor U3002 (N_3002,N_2119,N_2593);
nand U3003 (N_3003,N_2233,N_2420);
and U3004 (N_3004,N_2134,N_2918);
and U3005 (N_3005,N_2560,N_2237);
and U3006 (N_3006,N_2923,N_2479);
and U3007 (N_3007,N_2699,N_2188);
or U3008 (N_3008,N_2276,N_2186);
nor U3009 (N_3009,N_2824,N_2809);
nand U3010 (N_3010,N_2498,N_2093);
nor U3011 (N_3011,N_2489,N_2300);
or U3012 (N_3012,N_2054,N_2143);
nand U3013 (N_3013,N_2278,N_2499);
and U3014 (N_3014,N_2465,N_2749);
nor U3015 (N_3015,N_2603,N_2960);
xor U3016 (N_3016,N_2883,N_2306);
nor U3017 (N_3017,N_2669,N_2955);
or U3018 (N_3018,N_2321,N_2155);
nand U3019 (N_3019,N_2708,N_2302);
or U3020 (N_3020,N_2452,N_2158);
nand U3021 (N_3021,N_2059,N_2950);
and U3022 (N_3022,N_2545,N_2151);
nand U3023 (N_3023,N_2087,N_2152);
nor U3024 (N_3024,N_2739,N_2798);
and U3025 (N_3025,N_2348,N_2915);
nor U3026 (N_3026,N_2174,N_2873);
and U3027 (N_3027,N_2964,N_2185);
and U3028 (N_3028,N_2380,N_2965);
nand U3029 (N_3029,N_2289,N_2642);
or U3030 (N_3030,N_2308,N_2694);
or U3031 (N_3031,N_2561,N_2311);
nor U3032 (N_3032,N_2013,N_2100);
nand U3033 (N_3033,N_2983,N_2564);
nand U3034 (N_3034,N_2880,N_2274);
and U3035 (N_3035,N_2901,N_2931);
or U3036 (N_3036,N_2800,N_2926);
nor U3037 (N_3037,N_2412,N_2558);
and U3038 (N_3038,N_2025,N_2191);
nor U3039 (N_3039,N_2695,N_2241);
nor U3040 (N_3040,N_2862,N_2655);
nand U3041 (N_3041,N_2644,N_2555);
nand U3042 (N_3042,N_2074,N_2261);
or U3043 (N_3043,N_2223,N_2127);
nand U3044 (N_3044,N_2539,N_2106);
and U3045 (N_3045,N_2653,N_2864);
nor U3046 (N_3046,N_2852,N_2036);
xor U3047 (N_3047,N_2411,N_2734);
and U3048 (N_3048,N_2598,N_2641);
and U3049 (N_3049,N_2827,N_2362);
or U3050 (N_3050,N_2688,N_2126);
nand U3051 (N_3051,N_2386,N_2647);
nor U3052 (N_3052,N_2872,N_2586);
nand U3053 (N_3053,N_2906,N_2407);
nand U3054 (N_3054,N_2635,N_2557);
nor U3055 (N_3055,N_2510,N_2092);
or U3056 (N_3056,N_2843,N_2091);
nor U3057 (N_3057,N_2360,N_2773);
nor U3058 (N_3058,N_2267,N_2890);
nand U3059 (N_3059,N_2513,N_2951);
nor U3060 (N_3060,N_2627,N_2972);
xor U3061 (N_3061,N_2636,N_2044);
nor U3062 (N_3062,N_2405,N_2661);
or U3063 (N_3063,N_2710,N_2194);
xor U3064 (N_3064,N_2264,N_2856);
or U3065 (N_3065,N_2995,N_2372);
and U3066 (N_3066,N_2830,N_2347);
and U3067 (N_3067,N_2161,N_2008);
and U3068 (N_3068,N_2527,N_2224);
and U3069 (N_3069,N_2822,N_2375);
or U3070 (N_3070,N_2902,N_2582);
nand U3071 (N_3071,N_2860,N_2885);
and U3072 (N_3072,N_2572,N_2802);
xor U3073 (N_3073,N_2107,N_2521);
nor U3074 (N_3074,N_2390,N_2720);
nand U3075 (N_3075,N_2497,N_2870);
and U3076 (N_3076,N_2385,N_2529);
nor U3077 (N_3077,N_2729,N_2989);
or U3078 (N_3078,N_2445,N_2110);
xor U3079 (N_3079,N_2469,N_2842);
or U3080 (N_3080,N_2226,N_2674);
nand U3081 (N_3081,N_2975,N_2559);
nand U3082 (N_3082,N_2028,N_2114);
or U3083 (N_3083,N_2022,N_2982);
nor U3084 (N_3084,N_2630,N_2506);
or U3085 (N_3085,N_2696,N_2150);
or U3086 (N_3086,N_2820,N_2512);
and U3087 (N_3087,N_2903,N_2904);
and U3088 (N_3088,N_2429,N_2767);
and U3089 (N_3089,N_2941,N_2602);
nor U3090 (N_3090,N_2382,N_2604);
or U3091 (N_3091,N_2379,N_2128);
nand U3092 (N_3092,N_2569,N_2549);
nand U3093 (N_3093,N_2966,N_2631);
nand U3094 (N_3094,N_2578,N_2509);
and U3095 (N_3095,N_2922,N_2164);
or U3096 (N_3096,N_2472,N_2252);
and U3097 (N_3097,N_2098,N_2553);
or U3098 (N_3098,N_2763,N_2285);
or U3099 (N_3099,N_2944,N_2011);
nand U3100 (N_3100,N_2473,N_2755);
and U3101 (N_3101,N_2242,N_2425);
nor U3102 (N_3102,N_2159,N_2665);
nand U3103 (N_3103,N_2646,N_2096);
or U3104 (N_3104,N_2577,N_2184);
nand U3105 (N_3105,N_2166,N_2954);
and U3106 (N_3106,N_2381,N_2033);
nand U3107 (N_3107,N_2222,N_2131);
nand U3108 (N_3108,N_2774,N_2209);
and U3109 (N_3109,N_2490,N_2094);
nor U3110 (N_3110,N_2384,N_2788);
nand U3111 (N_3111,N_2515,N_2592);
nor U3112 (N_3112,N_2866,N_2459);
and U3113 (N_3113,N_2446,N_2973);
nor U3114 (N_3114,N_2725,N_2912);
nand U3115 (N_3115,N_2762,N_2244);
and U3116 (N_3116,N_2340,N_2879);
or U3117 (N_3117,N_2370,N_2449);
or U3118 (N_3118,N_2895,N_2238);
nor U3119 (N_3119,N_2142,N_2974);
and U3120 (N_3120,N_2045,N_2507);
nor U3121 (N_3121,N_2551,N_2139);
nor U3122 (N_3122,N_2178,N_2393);
and U3123 (N_3123,N_2021,N_2248);
nand U3124 (N_3124,N_2190,N_2101);
nor U3125 (N_3125,N_2826,N_2475);
xnor U3126 (N_3126,N_2138,N_2171);
nand U3127 (N_3127,N_2132,N_2791);
or U3128 (N_3128,N_2388,N_2316);
and U3129 (N_3129,N_2858,N_2849);
xnor U3130 (N_3130,N_2286,N_2476);
nor U3131 (N_3131,N_2658,N_2697);
xor U3132 (N_3132,N_2109,N_2061);
nand U3133 (N_3133,N_2819,N_2454);
nand U3134 (N_3134,N_2525,N_2060);
nand U3135 (N_3135,N_2344,N_2993);
nor U3136 (N_3136,N_2992,N_2976);
or U3137 (N_3137,N_2085,N_2324);
nand U3138 (N_3138,N_2361,N_2605);
nand U3139 (N_3139,N_2530,N_2784);
or U3140 (N_3140,N_2543,N_2905);
and U3141 (N_3141,N_2260,N_2103);
or U3142 (N_3142,N_2900,N_2594);
nand U3143 (N_3143,N_2235,N_2312);
nor U3144 (N_3144,N_2197,N_2778);
nand U3145 (N_3145,N_2769,N_2421);
nor U3146 (N_3146,N_2201,N_2043);
or U3147 (N_3147,N_2398,N_2567);
and U3148 (N_3148,N_2258,N_2181);
nand U3149 (N_3149,N_2154,N_2437);
nand U3150 (N_3150,N_2496,N_2032);
nand U3151 (N_3151,N_2548,N_2313);
or U3152 (N_3152,N_2735,N_2083);
and U3153 (N_3153,N_2969,N_2997);
nand U3154 (N_3154,N_2643,N_2392);
and U3155 (N_3155,N_2123,N_2840);
or U3156 (N_3156,N_2246,N_2520);
nand U3157 (N_3157,N_2511,N_2700);
and U3158 (N_3158,N_2550,N_2262);
and U3159 (N_3159,N_2371,N_2568);
or U3160 (N_3160,N_2495,N_2713);
nand U3161 (N_3161,N_2257,N_2337);
or U3162 (N_3162,N_2066,N_2198);
and U3163 (N_3163,N_2364,N_2399);
xor U3164 (N_3164,N_2205,N_2829);
or U3165 (N_3165,N_2366,N_2216);
nand U3166 (N_3166,N_2322,N_2422);
nor U3167 (N_3167,N_2744,N_2136);
and U3168 (N_3168,N_2081,N_2948);
nand U3169 (N_3169,N_2812,N_2051);
nand U3170 (N_3170,N_2048,N_2491);
or U3171 (N_3171,N_2396,N_2967);
and U3172 (N_3172,N_2149,N_2365);
and U3173 (N_3173,N_2637,N_2374);
or U3174 (N_3174,N_2428,N_2005);
nand U3175 (N_3175,N_2911,N_2323);
nor U3176 (N_3176,N_2419,N_2522);
nand U3177 (N_3177,N_2508,N_2991);
nand U3178 (N_3178,N_2438,N_2494);
nor U3179 (N_3179,N_2227,N_2884);
or U3180 (N_3180,N_2736,N_2664);
or U3181 (N_3181,N_2462,N_2591);
and U3182 (N_3182,N_2971,N_2432);
xor U3183 (N_3183,N_2783,N_2657);
nand U3184 (N_3184,N_2433,N_2474);
or U3185 (N_3185,N_2724,N_2280);
nand U3186 (N_3186,N_2533,N_2733);
nand U3187 (N_3187,N_2439,N_2231);
or U3188 (N_3188,N_2301,N_2999);
xnor U3189 (N_3189,N_2305,N_2893);
nor U3190 (N_3190,N_2546,N_2263);
and U3191 (N_3191,N_2481,N_2024);
nor U3192 (N_3192,N_2482,N_2140);
or U3193 (N_3193,N_2804,N_2668);
and U3194 (N_3194,N_2701,N_2335);
or U3195 (N_3195,N_2875,N_2757);
nor U3196 (N_3196,N_2981,N_2493);
nor U3197 (N_3197,N_2534,N_2979);
and U3198 (N_3198,N_2987,N_2213);
and U3199 (N_3199,N_2619,N_2790);
or U3200 (N_3200,N_2590,N_2857);
nand U3201 (N_3201,N_2125,N_2503);
nor U3202 (N_3202,N_2120,N_2104);
or U3203 (N_3203,N_2986,N_2633);
and U3204 (N_3204,N_2715,N_2610);
or U3205 (N_3205,N_2055,N_2097);
and U3206 (N_3206,N_2684,N_2281);
nand U3207 (N_3207,N_2378,N_2679);
and U3208 (N_3208,N_2464,N_2618);
nand U3209 (N_3209,N_2326,N_2881);
nand U3210 (N_3210,N_2389,N_2929);
nor U3211 (N_3211,N_2741,N_2220);
nand U3212 (N_3212,N_2841,N_2761);
nor U3213 (N_3213,N_2676,N_2654);
nand U3214 (N_3214,N_2189,N_2214);
and U3215 (N_3215,N_2062,N_2265);
or U3216 (N_3216,N_2453,N_2990);
nor U3217 (N_3217,N_2620,N_2805);
or U3218 (N_3218,N_2565,N_2383);
or U3219 (N_3219,N_2772,N_2484);
or U3220 (N_3220,N_2949,N_2770);
and U3221 (N_3221,N_2271,N_2523);
or U3222 (N_3222,N_2693,N_2208);
or U3223 (N_3223,N_2651,N_2318);
nand U3224 (N_3224,N_2759,N_2165);
and U3225 (N_3225,N_2451,N_2650);
nand U3226 (N_3226,N_2573,N_2579);
nor U3227 (N_3227,N_2207,N_2272);
nor U3228 (N_3228,N_2299,N_2455);
and U3229 (N_3229,N_2984,N_2834);
nand U3230 (N_3230,N_2049,N_2738);
nand U3231 (N_3231,N_2065,N_2962);
nor U3232 (N_3232,N_2638,N_2850);
and U3233 (N_3233,N_2718,N_2239);
xnor U3234 (N_3234,N_2339,N_2556);
nand U3235 (N_3235,N_2698,N_2273);
or U3236 (N_3236,N_2745,N_2814);
and U3237 (N_3237,N_2341,N_2501);
nand U3238 (N_3238,N_2293,N_2566);
nand U3239 (N_3239,N_2825,N_2443);
nand U3240 (N_3240,N_2765,N_2963);
nand U3241 (N_3241,N_2562,N_2907);
nor U3242 (N_3242,N_2373,N_2867);
and U3243 (N_3243,N_2342,N_2423);
nor U3244 (N_3244,N_2920,N_2253);
or U3245 (N_3245,N_2703,N_2606);
nand U3246 (N_3246,N_2358,N_2531);
and U3247 (N_3247,N_2355,N_2625);
and U3248 (N_3248,N_2859,N_2417);
nor U3249 (N_3249,N_2839,N_2019);
nand U3250 (N_3250,N_2404,N_2041);
nand U3251 (N_3251,N_2892,N_2775);
nand U3252 (N_3252,N_2387,N_2518);
and U3253 (N_3253,N_2175,N_2897);
and U3254 (N_3254,N_2996,N_2416);
or U3255 (N_3255,N_2219,N_2928);
or U3256 (N_3256,N_2970,N_2868);
and U3257 (N_3257,N_2243,N_2467);
and U3258 (N_3258,N_2538,N_2946);
nor U3259 (N_3259,N_2781,N_2147);
nor U3260 (N_3260,N_2570,N_2616);
nand U3261 (N_3261,N_2052,N_2779);
and U3262 (N_3262,N_2563,N_2847);
nor U3263 (N_3263,N_2848,N_2346);
and U3264 (N_3264,N_2532,N_2672);
and U3265 (N_3265,N_2933,N_2292);
nand U3266 (N_3266,N_2742,N_2303);
nand U3267 (N_3267,N_2111,N_2082);
nand U3268 (N_3268,N_2448,N_2815);
nor U3269 (N_3269,N_2296,N_2776);
nor U3270 (N_3270,N_2617,N_2891);
or U3271 (N_3271,N_2117,N_2345);
and U3272 (N_3272,N_2528,N_2349);
or U3273 (N_3273,N_2719,N_2206);
nand U3274 (N_3274,N_2599,N_2634);
xor U3275 (N_3275,N_2232,N_2705);
and U3276 (N_3276,N_2029,N_2471);
nand U3277 (N_3277,N_2410,N_2747);
or U3278 (N_3278,N_2351,N_2689);
and U3279 (N_3279,N_2327,N_2415);
and U3280 (N_3280,N_2331,N_2200);
or U3281 (N_3281,N_2752,N_2486);
nand U3282 (N_3282,N_2608,N_2943);
nor U3283 (N_3283,N_2363,N_2600);
or U3284 (N_3284,N_2913,N_2137);
or U3285 (N_3285,N_2196,N_2047);
nor U3286 (N_3286,N_2660,N_2766);
or U3287 (N_3287,N_2728,N_2040);
or U3288 (N_3288,N_2487,N_2806);
or U3289 (N_3289,N_2921,N_2210);
and U3290 (N_3290,N_2488,N_2894);
nand U3291 (N_3291,N_2332,N_2927);
and U3292 (N_3292,N_2105,N_2282);
nor U3293 (N_3293,N_2640,N_2027);
nor U3294 (N_3294,N_2576,N_2042);
and U3295 (N_3295,N_2869,N_2748);
or U3296 (N_3296,N_2707,N_2945);
or U3297 (N_3297,N_2932,N_2780);
or U3298 (N_3298,N_2026,N_2124);
or U3299 (N_3299,N_2334,N_2317);
and U3300 (N_3300,N_2162,N_2799);
nand U3301 (N_3301,N_2397,N_2070);
nor U3302 (N_3302,N_2882,N_2418);
or U3303 (N_3303,N_2878,N_2596);
nor U3304 (N_3304,N_2255,N_2067);
nand U3305 (N_3305,N_2069,N_2977);
and U3306 (N_3306,N_2998,N_2807);
or U3307 (N_3307,N_2259,N_2009);
nand U3308 (N_3308,N_2007,N_2477);
or U3309 (N_3309,N_2702,N_2785);
xor U3310 (N_3310,N_2073,N_2659);
or U3311 (N_3311,N_2671,N_2730);
and U3312 (N_3312,N_2771,N_2035);
or U3313 (N_3313,N_2519,N_2450);
nor U3314 (N_3314,N_2202,N_2217);
nor U3315 (N_3315,N_2251,N_2304);
and U3316 (N_3316,N_2645,N_2835);
nor U3317 (N_3317,N_2172,N_2298);
nand U3318 (N_3318,N_2275,N_2517);
nand U3319 (N_3319,N_2086,N_2402);
nor U3320 (N_3320,N_2177,N_2743);
xnor U3321 (N_3321,N_2006,N_2924);
or U3322 (N_3322,N_2670,N_2176);
nand U3323 (N_3323,N_2144,N_2084);
or U3324 (N_3324,N_2795,N_2199);
and U3325 (N_3325,N_2575,N_2367);
and U3326 (N_3326,N_2621,N_2376);
nor U3327 (N_3327,N_2667,N_2692);
or U3328 (N_3328,N_2723,N_2677);
or U3329 (N_3329,N_2683,N_2108);
nor U3330 (N_3330,N_2803,N_2942);
nor U3331 (N_3331,N_2102,N_2716);
nand U3332 (N_3332,N_2797,N_2832);
nand U3333 (N_3333,N_2288,N_2838);
nor U3334 (N_3334,N_2810,N_2956);
and U3335 (N_3335,N_2754,N_2876);
or U3336 (N_3336,N_2121,N_2204);
nand U3337 (N_3337,N_2156,N_2940);
nand U3338 (N_3338,N_2034,N_2247);
nand U3339 (N_3339,N_2666,N_2195);
or U3340 (N_3340,N_2173,N_2690);
nor U3341 (N_3341,N_2187,N_2325);
nor U3342 (N_3342,N_2330,N_2662);
and U3343 (N_3343,N_2003,N_2406);
nand U3344 (N_3344,N_2268,N_2169);
nor U3345 (N_3345,N_2607,N_2221);
nand U3346 (N_3346,N_2240,N_2413);
or U3347 (N_3347,N_2629,N_2552);
nor U3348 (N_3348,N_2249,N_2831);
nand U3349 (N_3349,N_2250,N_2823);
nor U3350 (N_3350,N_2010,N_2711);
nor U3351 (N_3351,N_2935,N_2076);
nand U3352 (N_3352,N_2183,N_2369);
or U3353 (N_3353,N_2504,N_2612);
nand U3354 (N_3354,N_2535,N_2444);
or U3355 (N_3355,N_2581,N_2595);
and U3356 (N_3356,N_2297,N_2153);
nor U3357 (N_3357,N_2587,N_2391);
and U3358 (N_3358,N_2801,N_2714);
nor U3359 (N_3359,N_2789,N_2192);
nand U3360 (N_3360,N_2320,N_2203);
or U3361 (N_3361,N_2343,N_2333);
nand U3362 (N_3362,N_2018,N_2046);
nor U3363 (N_3363,N_2908,N_2266);
nand U3364 (N_3364,N_2886,N_2000);
and U3365 (N_3365,N_2492,N_2833);
or U3366 (N_3366,N_2540,N_2329);
or U3367 (N_3367,N_2685,N_2245);
or U3368 (N_3368,N_2211,N_2115);
xnor U3369 (N_3369,N_2768,N_2163);
or U3370 (N_3370,N_2394,N_2717);
and U3371 (N_3371,N_2628,N_2632);
nor U3372 (N_3372,N_2461,N_2130);
nand U3373 (N_3373,N_2064,N_2314);
or U3374 (N_3374,N_2792,N_2352);
or U3375 (N_3375,N_2914,N_2080);
nand U3376 (N_3376,N_2936,N_2157);
or U3377 (N_3377,N_2704,N_2377);
and U3378 (N_3378,N_2088,N_2182);
and U3379 (N_3379,N_2571,N_2338);
nand U3380 (N_3380,N_2502,N_2639);
nor U3381 (N_3381,N_2017,N_2403);
or U3382 (N_3382,N_2440,N_2648);
nor U3383 (N_3383,N_2930,N_2853);
or U3384 (N_3384,N_2855,N_2112);
and U3385 (N_3385,N_2786,N_2751);
or U3386 (N_3386,N_2544,N_2816);
and U3387 (N_3387,N_2818,N_2691);
or U3388 (N_3388,N_2952,N_2782);
nor U3389 (N_3389,N_2170,N_2284);
nor U3390 (N_3390,N_2328,N_2959);
or U3391 (N_3391,N_2270,N_2218);
or U3392 (N_3392,N_2611,N_2077);
nand U3393 (N_3393,N_2712,N_2427);
nor U3394 (N_3394,N_2113,N_2898);
nand U3395 (N_3395,N_2758,N_2500);
nand U3396 (N_3396,N_2409,N_2436);
nor U3397 (N_3397,N_2938,N_2874);
or U3398 (N_3398,N_2597,N_2828);
and U3399 (N_3399,N_2680,N_2071);
and U3400 (N_3400,N_2023,N_2589);
and U3401 (N_3401,N_2309,N_2287);
nand U3402 (N_3402,N_2649,N_2424);
or U3403 (N_3403,N_2953,N_2505);
nand U3404 (N_3404,N_2031,N_2686);
nand U3405 (N_3405,N_2229,N_2146);
nand U3406 (N_3406,N_2078,N_2687);
nand U3407 (N_3407,N_2468,N_2957);
and U3408 (N_3408,N_2584,N_2994);
or U3409 (N_3409,N_2609,N_2793);
and U3410 (N_3410,N_2678,N_2601);
nor U3411 (N_3411,N_2269,N_2463);
or U3412 (N_3412,N_2063,N_2526);
and U3413 (N_3413,N_2291,N_2148);
nor U3414 (N_3414,N_2871,N_2746);
nand U3415 (N_3415,N_2614,N_2541);
and U3416 (N_3416,N_2050,N_2777);
and U3417 (N_3417,N_2845,N_2426);
nor U3418 (N_3418,N_2256,N_2731);
and U3419 (N_3419,N_2414,N_2079);
or U3420 (N_3420,N_2038,N_2431);
or U3421 (N_3421,N_2588,N_2726);
nor U3422 (N_3422,N_2160,N_2447);
nor U3423 (N_3423,N_2727,N_2057);
nor U3424 (N_3424,N_2435,N_2613);
or U3425 (N_3425,N_2909,N_2012);
nand U3426 (N_3426,N_2167,N_2179);
or U3427 (N_3427,N_2889,N_2910);
and U3428 (N_3428,N_2095,N_2899);
nand U3429 (N_3429,N_2622,N_2837);
nor U3430 (N_3430,N_2919,N_2014);
or U3431 (N_3431,N_2626,N_2836);
nor U3432 (N_3432,N_2787,N_2254);
or U3433 (N_3433,N_2934,N_2075);
or U3434 (N_3434,N_2978,N_2395);
nand U3435 (N_3435,N_2234,N_2813);
nor U3436 (N_3436,N_2817,N_2656);
nand U3437 (N_3437,N_2861,N_2039);
nor U3438 (N_3438,N_2037,N_2053);
nor U3439 (N_3439,N_2917,N_2236);
and U3440 (N_3440,N_2673,N_2133);
nand U3441 (N_3441,N_2277,N_2480);
nor U3442 (N_3442,N_2958,N_2542);
nor U3443 (N_3443,N_2980,N_2030);
or U3444 (N_3444,N_2888,N_2135);
or U3445 (N_3445,N_2740,N_2916);
nor U3446 (N_3446,N_2460,N_2709);
nor U3447 (N_3447,N_2336,N_2004);
or U3448 (N_3448,N_2225,N_2015);
nor U3449 (N_3449,N_2089,N_2681);
nor U3450 (N_3450,N_2001,N_2441);
nor U3451 (N_3451,N_2821,N_2400);
and U3452 (N_3452,N_2808,N_2228);
nor U3453 (N_3453,N_2887,N_2430);
nor U3454 (N_3454,N_2547,N_2583);
or U3455 (N_3455,N_2353,N_2099);
nor U3456 (N_3456,N_2068,N_2230);
or U3457 (N_3457,N_2968,N_2356);
or U3458 (N_3458,N_2756,N_2129);
nand U3459 (N_3459,N_2947,N_2796);
nor U3460 (N_3460,N_2675,N_2794);
and U3461 (N_3461,N_2307,N_2753);
nand U3462 (N_3462,N_2401,N_2846);
and U3463 (N_3463,N_2457,N_2434);
nand U3464 (N_3464,N_2863,N_2721);
and U3465 (N_3465,N_2706,N_2554);
nor U3466 (N_3466,N_2058,N_2310);
nor U3467 (N_3467,N_2002,N_2574);
nand U3468 (N_3468,N_2016,N_2865);
nor U3469 (N_3469,N_2283,N_2485);
and U3470 (N_3470,N_2319,N_2524);
and U3471 (N_3471,N_2116,N_2764);
nand U3472 (N_3472,N_2939,N_2478);
nand U3473 (N_3473,N_2985,N_2193);
and U3474 (N_3474,N_2877,N_2056);
nor U3475 (N_3475,N_2357,N_2470);
and U3476 (N_3476,N_2122,N_2896);
or U3477 (N_3477,N_2854,N_2458);
nor U3478 (N_3478,N_2483,N_2514);
or U3479 (N_3479,N_2760,N_2682);
nor U3480 (N_3480,N_2844,N_2295);
nor U3481 (N_3481,N_2580,N_2212);
nor U3482 (N_3482,N_2279,N_2615);
nor U3483 (N_3483,N_2315,N_2294);
or U3484 (N_3484,N_2118,N_2516);
or U3485 (N_3485,N_2145,N_2988);
nand U3486 (N_3486,N_2585,N_2851);
and U3487 (N_3487,N_2180,N_2072);
and U3488 (N_3488,N_2624,N_2750);
nor U3489 (N_3489,N_2290,N_2354);
or U3490 (N_3490,N_2408,N_2350);
or U3491 (N_3491,N_2663,N_2456);
nor U3492 (N_3492,N_2925,N_2141);
or U3493 (N_3493,N_2623,N_2215);
nand U3494 (N_3494,N_2732,N_2466);
nor U3495 (N_3495,N_2090,N_2168);
or U3496 (N_3496,N_2961,N_2442);
or U3497 (N_3497,N_2359,N_2368);
nor U3498 (N_3498,N_2537,N_2937);
and U3499 (N_3499,N_2020,N_2737);
xor U3500 (N_3500,N_2221,N_2878);
and U3501 (N_3501,N_2774,N_2843);
nand U3502 (N_3502,N_2942,N_2274);
and U3503 (N_3503,N_2346,N_2972);
and U3504 (N_3504,N_2899,N_2371);
nor U3505 (N_3505,N_2575,N_2269);
and U3506 (N_3506,N_2756,N_2070);
or U3507 (N_3507,N_2634,N_2152);
nand U3508 (N_3508,N_2759,N_2662);
or U3509 (N_3509,N_2601,N_2165);
and U3510 (N_3510,N_2950,N_2207);
nand U3511 (N_3511,N_2282,N_2011);
or U3512 (N_3512,N_2912,N_2630);
and U3513 (N_3513,N_2544,N_2836);
or U3514 (N_3514,N_2215,N_2161);
or U3515 (N_3515,N_2975,N_2749);
and U3516 (N_3516,N_2186,N_2188);
or U3517 (N_3517,N_2417,N_2867);
nor U3518 (N_3518,N_2762,N_2604);
and U3519 (N_3519,N_2041,N_2336);
and U3520 (N_3520,N_2181,N_2519);
or U3521 (N_3521,N_2366,N_2889);
nand U3522 (N_3522,N_2078,N_2521);
or U3523 (N_3523,N_2530,N_2246);
and U3524 (N_3524,N_2126,N_2807);
xor U3525 (N_3525,N_2955,N_2274);
nand U3526 (N_3526,N_2667,N_2691);
nand U3527 (N_3527,N_2339,N_2366);
nand U3528 (N_3528,N_2845,N_2207);
or U3529 (N_3529,N_2652,N_2169);
nand U3530 (N_3530,N_2795,N_2776);
or U3531 (N_3531,N_2641,N_2078);
nor U3532 (N_3532,N_2166,N_2070);
nand U3533 (N_3533,N_2979,N_2548);
nand U3534 (N_3534,N_2667,N_2718);
nand U3535 (N_3535,N_2425,N_2297);
nor U3536 (N_3536,N_2055,N_2018);
or U3537 (N_3537,N_2546,N_2222);
and U3538 (N_3538,N_2141,N_2195);
and U3539 (N_3539,N_2862,N_2899);
nor U3540 (N_3540,N_2234,N_2467);
and U3541 (N_3541,N_2735,N_2657);
and U3542 (N_3542,N_2345,N_2682);
nor U3543 (N_3543,N_2413,N_2941);
or U3544 (N_3544,N_2400,N_2463);
and U3545 (N_3545,N_2394,N_2578);
or U3546 (N_3546,N_2193,N_2475);
or U3547 (N_3547,N_2222,N_2197);
or U3548 (N_3548,N_2085,N_2364);
nand U3549 (N_3549,N_2457,N_2530);
nand U3550 (N_3550,N_2929,N_2932);
nor U3551 (N_3551,N_2834,N_2844);
nor U3552 (N_3552,N_2664,N_2574);
nand U3553 (N_3553,N_2397,N_2616);
nor U3554 (N_3554,N_2543,N_2691);
or U3555 (N_3555,N_2142,N_2672);
nand U3556 (N_3556,N_2977,N_2641);
nor U3557 (N_3557,N_2032,N_2903);
nand U3558 (N_3558,N_2184,N_2692);
nand U3559 (N_3559,N_2367,N_2824);
nand U3560 (N_3560,N_2246,N_2663);
and U3561 (N_3561,N_2939,N_2615);
and U3562 (N_3562,N_2305,N_2356);
xor U3563 (N_3563,N_2252,N_2801);
nand U3564 (N_3564,N_2490,N_2541);
or U3565 (N_3565,N_2646,N_2374);
nor U3566 (N_3566,N_2517,N_2046);
and U3567 (N_3567,N_2886,N_2644);
nor U3568 (N_3568,N_2083,N_2202);
and U3569 (N_3569,N_2605,N_2471);
or U3570 (N_3570,N_2061,N_2052);
or U3571 (N_3571,N_2261,N_2742);
or U3572 (N_3572,N_2282,N_2593);
and U3573 (N_3573,N_2960,N_2851);
or U3574 (N_3574,N_2861,N_2991);
nand U3575 (N_3575,N_2952,N_2232);
or U3576 (N_3576,N_2883,N_2311);
nand U3577 (N_3577,N_2973,N_2561);
and U3578 (N_3578,N_2530,N_2934);
nor U3579 (N_3579,N_2560,N_2787);
nor U3580 (N_3580,N_2857,N_2943);
nand U3581 (N_3581,N_2389,N_2995);
or U3582 (N_3582,N_2756,N_2520);
or U3583 (N_3583,N_2695,N_2214);
and U3584 (N_3584,N_2482,N_2479);
nor U3585 (N_3585,N_2907,N_2659);
nor U3586 (N_3586,N_2039,N_2385);
and U3587 (N_3587,N_2648,N_2214);
or U3588 (N_3588,N_2880,N_2258);
nor U3589 (N_3589,N_2641,N_2493);
or U3590 (N_3590,N_2797,N_2667);
xor U3591 (N_3591,N_2243,N_2395);
or U3592 (N_3592,N_2996,N_2594);
nand U3593 (N_3593,N_2404,N_2375);
or U3594 (N_3594,N_2678,N_2312);
and U3595 (N_3595,N_2550,N_2436);
nand U3596 (N_3596,N_2898,N_2725);
and U3597 (N_3597,N_2944,N_2720);
nor U3598 (N_3598,N_2167,N_2557);
nor U3599 (N_3599,N_2986,N_2005);
nand U3600 (N_3600,N_2799,N_2122);
nand U3601 (N_3601,N_2494,N_2680);
or U3602 (N_3602,N_2358,N_2525);
xnor U3603 (N_3603,N_2958,N_2977);
and U3604 (N_3604,N_2424,N_2220);
nor U3605 (N_3605,N_2978,N_2030);
nor U3606 (N_3606,N_2852,N_2660);
and U3607 (N_3607,N_2093,N_2820);
or U3608 (N_3608,N_2029,N_2441);
and U3609 (N_3609,N_2234,N_2025);
or U3610 (N_3610,N_2429,N_2921);
xor U3611 (N_3611,N_2845,N_2464);
nand U3612 (N_3612,N_2791,N_2415);
and U3613 (N_3613,N_2809,N_2362);
or U3614 (N_3614,N_2979,N_2408);
and U3615 (N_3615,N_2126,N_2712);
or U3616 (N_3616,N_2747,N_2670);
nor U3617 (N_3617,N_2278,N_2589);
nor U3618 (N_3618,N_2993,N_2941);
nand U3619 (N_3619,N_2002,N_2153);
xor U3620 (N_3620,N_2057,N_2048);
nand U3621 (N_3621,N_2309,N_2606);
and U3622 (N_3622,N_2511,N_2153);
nor U3623 (N_3623,N_2236,N_2803);
nor U3624 (N_3624,N_2057,N_2863);
xnor U3625 (N_3625,N_2645,N_2531);
and U3626 (N_3626,N_2838,N_2990);
and U3627 (N_3627,N_2466,N_2672);
xnor U3628 (N_3628,N_2167,N_2894);
or U3629 (N_3629,N_2178,N_2201);
nand U3630 (N_3630,N_2497,N_2321);
or U3631 (N_3631,N_2301,N_2277);
or U3632 (N_3632,N_2202,N_2771);
nand U3633 (N_3633,N_2359,N_2384);
nand U3634 (N_3634,N_2076,N_2442);
nand U3635 (N_3635,N_2428,N_2561);
and U3636 (N_3636,N_2068,N_2185);
or U3637 (N_3637,N_2195,N_2138);
nand U3638 (N_3638,N_2157,N_2254);
or U3639 (N_3639,N_2468,N_2372);
nor U3640 (N_3640,N_2401,N_2736);
nand U3641 (N_3641,N_2927,N_2548);
nand U3642 (N_3642,N_2869,N_2886);
nor U3643 (N_3643,N_2940,N_2661);
nor U3644 (N_3644,N_2620,N_2804);
nor U3645 (N_3645,N_2374,N_2946);
nor U3646 (N_3646,N_2299,N_2324);
nand U3647 (N_3647,N_2968,N_2413);
or U3648 (N_3648,N_2725,N_2360);
and U3649 (N_3649,N_2450,N_2336);
nor U3650 (N_3650,N_2727,N_2247);
and U3651 (N_3651,N_2594,N_2640);
and U3652 (N_3652,N_2095,N_2162);
nand U3653 (N_3653,N_2899,N_2146);
and U3654 (N_3654,N_2341,N_2374);
or U3655 (N_3655,N_2582,N_2953);
nand U3656 (N_3656,N_2466,N_2778);
nor U3657 (N_3657,N_2419,N_2820);
nand U3658 (N_3658,N_2023,N_2070);
or U3659 (N_3659,N_2927,N_2568);
nand U3660 (N_3660,N_2197,N_2491);
nor U3661 (N_3661,N_2882,N_2054);
or U3662 (N_3662,N_2947,N_2830);
or U3663 (N_3663,N_2605,N_2730);
xor U3664 (N_3664,N_2341,N_2352);
nor U3665 (N_3665,N_2625,N_2975);
or U3666 (N_3666,N_2340,N_2017);
nor U3667 (N_3667,N_2755,N_2588);
nor U3668 (N_3668,N_2147,N_2374);
nor U3669 (N_3669,N_2873,N_2025);
nand U3670 (N_3670,N_2588,N_2514);
nor U3671 (N_3671,N_2407,N_2709);
nand U3672 (N_3672,N_2891,N_2803);
and U3673 (N_3673,N_2170,N_2580);
or U3674 (N_3674,N_2971,N_2045);
or U3675 (N_3675,N_2878,N_2446);
or U3676 (N_3676,N_2005,N_2313);
or U3677 (N_3677,N_2262,N_2661);
nand U3678 (N_3678,N_2085,N_2094);
xor U3679 (N_3679,N_2555,N_2753);
or U3680 (N_3680,N_2648,N_2339);
nand U3681 (N_3681,N_2506,N_2172);
or U3682 (N_3682,N_2143,N_2290);
and U3683 (N_3683,N_2909,N_2861);
nor U3684 (N_3684,N_2765,N_2855);
and U3685 (N_3685,N_2586,N_2584);
or U3686 (N_3686,N_2461,N_2631);
xor U3687 (N_3687,N_2874,N_2450);
and U3688 (N_3688,N_2143,N_2959);
or U3689 (N_3689,N_2916,N_2269);
nand U3690 (N_3690,N_2030,N_2855);
nor U3691 (N_3691,N_2932,N_2927);
or U3692 (N_3692,N_2274,N_2019);
and U3693 (N_3693,N_2648,N_2608);
nor U3694 (N_3694,N_2068,N_2595);
and U3695 (N_3695,N_2665,N_2731);
or U3696 (N_3696,N_2826,N_2657);
xor U3697 (N_3697,N_2442,N_2680);
or U3698 (N_3698,N_2955,N_2762);
or U3699 (N_3699,N_2879,N_2007);
nor U3700 (N_3700,N_2337,N_2571);
nor U3701 (N_3701,N_2468,N_2576);
nand U3702 (N_3702,N_2837,N_2685);
nor U3703 (N_3703,N_2086,N_2917);
or U3704 (N_3704,N_2990,N_2669);
nand U3705 (N_3705,N_2752,N_2912);
and U3706 (N_3706,N_2324,N_2633);
or U3707 (N_3707,N_2667,N_2319);
nor U3708 (N_3708,N_2291,N_2561);
nor U3709 (N_3709,N_2171,N_2611);
nand U3710 (N_3710,N_2166,N_2862);
or U3711 (N_3711,N_2825,N_2690);
or U3712 (N_3712,N_2844,N_2342);
or U3713 (N_3713,N_2782,N_2001);
and U3714 (N_3714,N_2155,N_2594);
nand U3715 (N_3715,N_2070,N_2031);
or U3716 (N_3716,N_2668,N_2488);
xnor U3717 (N_3717,N_2542,N_2963);
xor U3718 (N_3718,N_2521,N_2942);
nand U3719 (N_3719,N_2571,N_2124);
nor U3720 (N_3720,N_2463,N_2881);
nand U3721 (N_3721,N_2314,N_2310);
or U3722 (N_3722,N_2106,N_2406);
xnor U3723 (N_3723,N_2071,N_2220);
nor U3724 (N_3724,N_2471,N_2130);
or U3725 (N_3725,N_2866,N_2884);
nand U3726 (N_3726,N_2420,N_2056);
nand U3727 (N_3727,N_2738,N_2141);
xnor U3728 (N_3728,N_2058,N_2725);
nor U3729 (N_3729,N_2805,N_2077);
nor U3730 (N_3730,N_2276,N_2077);
nor U3731 (N_3731,N_2446,N_2668);
or U3732 (N_3732,N_2387,N_2144);
and U3733 (N_3733,N_2090,N_2154);
and U3734 (N_3734,N_2289,N_2814);
and U3735 (N_3735,N_2809,N_2399);
nand U3736 (N_3736,N_2030,N_2900);
nor U3737 (N_3737,N_2796,N_2741);
nand U3738 (N_3738,N_2510,N_2263);
or U3739 (N_3739,N_2174,N_2834);
nand U3740 (N_3740,N_2042,N_2503);
nand U3741 (N_3741,N_2801,N_2737);
nand U3742 (N_3742,N_2908,N_2936);
nand U3743 (N_3743,N_2189,N_2622);
nand U3744 (N_3744,N_2585,N_2328);
nand U3745 (N_3745,N_2357,N_2278);
and U3746 (N_3746,N_2308,N_2040);
and U3747 (N_3747,N_2896,N_2224);
or U3748 (N_3748,N_2773,N_2925);
nor U3749 (N_3749,N_2356,N_2596);
and U3750 (N_3750,N_2915,N_2736);
xnor U3751 (N_3751,N_2615,N_2716);
and U3752 (N_3752,N_2664,N_2841);
nor U3753 (N_3753,N_2891,N_2036);
or U3754 (N_3754,N_2261,N_2510);
and U3755 (N_3755,N_2538,N_2761);
and U3756 (N_3756,N_2606,N_2469);
nor U3757 (N_3757,N_2102,N_2417);
xor U3758 (N_3758,N_2254,N_2497);
xor U3759 (N_3759,N_2331,N_2994);
nand U3760 (N_3760,N_2350,N_2954);
or U3761 (N_3761,N_2834,N_2114);
nor U3762 (N_3762,N_2703,N_2900);
nor U3763 (N_3763,N_2364,N_2091);
nor U3764 (N_3764,N_2549,N_2233);
nand U3765 (N_3765,N_2305,N_2852);
or U3766 (N_3766,N_2236,N_2001);
and U3767 (N_3767,N_2472,N_2204);
or U3768 (N_3768,N_2780,N_2528);
or U3769 (N_3769,N_2028,N_2275);
nand U3770 (N_3770,N_2041,N_2330);
and U3771 (N_3771,N_2930,N_2957);
and U3772 (N_3772,N_2882,N_2767);
nor U3773 (N_3773,N_2581,N_2366);
and U3774 (N_3774,N_2525,N_2464);
nor U3775 (N_3775,N_2831,N_2932);
nor U3776 (N_3776,N_2879,N_2947);
and U3777 (N_3777,N_2807,N_2249);
and U3778 (N_3778,N_2755,N_2893);
nor U3779 (N_3779,N_2348,N_2865);
xor U3780 (N_3780,N_2591,N_2404);
nor U3781 (N_3781,N_2062,N_2040);
nor U3782 (N_3782,N_2622,N_2008);
or U3783 (N_3783,N_2265,N_2389);
and U3784 (N_3784,N_2167,N_2755);
nand U3785 (N_3785,N_2744,N_2627);
nand U3786 (N_3786,N_2814,N_2914);
nor U3787 (N_3787,N_2676,N_2095);
or U3788 (N_3788,N_2596,N_2191);
and U3789 (N_3789,N_2239,N_2038);
or U3790 (N_3790,N_2383,N_2347);
nand U3791 (N_3791,N_2681,N_2704);
and U3792 (N_3792,N_2441,N_2859);
or U3793 (N_3793,N_2168,N_2748);
nand U3794 (N_3794,N_2842,N_2718);
and U3795 (N_3795,N_2219,N_2073);
nor U3796 (N_3796,N_2098,N_2361);
nor U3797 (N_3797,N_2407,N_2302);
or U3798 (N_3798,N_2651,N_2461);
nand U3799 (N_3799,N_2684,N_2022);
nand U3800 (N_3800,N_2829,N_2164);
and U3801 (N_3801,N_2562,N_2908);
nor U3802 (N_3802,N_2154,N_2585);
or U3803 (N_3803,N_2898,N_2154);
nand U3804 (N_3804,N_2878,N_2603);
nor U3805 (N_3805,N_2784,N_2495);
nor U3806 (N_3806,N_2317,N_2542);
or U3807 (N_3807,N_2950,N_2360);
nor U3808 (N_3808,N_2276,N_2152);
and U3809 (N_3809,N_2811,N_2255);
or U3810 (N_3810,N_2087,N_2218);
nor U3811 (N_3811,N_2437,N_2877);
and U3812 (N_3812,N_2757,N_2388);
or U3813 (N_3813,N_2426,N_2453);
nand U3814 (N_3814,N_2797,N_2956);
and U3815 (N_3815,N_2991,N_2742);
and U3816 (N_3816,N_2933,N_2016);
and U3817 (N_3817,N_2184,N_2081);
nand U3818 (N_3818,N_2893,N_2815);
and U3819 (N_3819,N_2139,N_2972);
and U3820 (N_3820,N_2016,N_2445);
nor U3821 (N_3821,N_2155,N_2577);
and U3822 (N_3822,N_2828,N_2177);
or U3823 (N_3823,N_2539,N_2640);
and U3824 (N_3824,N_2477,N_2870);
and U3825 (N_3825,N_2741,N_2815);
or U3826 (N_3826,N_2615,N_2609);
nand U3827 (N_3827,N_2851,N_2532);
or U3828 (N_3828,N_2238,N_2156);
nor U3829 (N_3829,N_2186,N_2306);
nand U3830 (N_3830,N_2562,N_2983);
nor U3831 (N_3831,N_2402,N_2469);
nor U3832 (N_3832,N_2009,N_2157);
nor U3833 (N_3833,N_2220,N_2761);
and U3834 (N_3834,N_2968,N_2602);
nand U3835 (N_3835,N_2061,N_2021);
and U3836 (N_3836,N_2892,N_2063);
or U3837 (N_3837,N_2857,N_2065);
nand U3838 (N_3838,N_2144,N_2491);
nor U3839 (N_3839,N_2402,N_2014);
nand U3840 (N_3840,N_2069,N_2200);
or U3841 (N_3841,N_2604,N_2480);
nand U3842 (N_3842,N_2261,N_2730);
nand U3843 (N_3843,N_2875,N_2453);
or U3844 (N_3844,N_2548,N_2945);
nand U3845 (N_3845,N_2967,N_2183);
or U3846 (N_3846,N_2103,N_2742);
or U3847 (N_3847,N_2053,N_2059);
nand U3848 (N_3848,N_2184,N_2987);
nor U3849 (N_3849,N_2782,N_2293);
nor U3850 (N_3850,N_2799,N_2369);
nor U3851 (N_3851,N_2281,N_2136);
and U3852 (N_3852,N_2275,N_2754);
nor U3853 (N_3853,N_2789,N_2371);
nand U3854 (N_3854,N_2674,N_2269);
nor U3855 (N_3855,N_2003,N_2390);
nor U3856 (N_3856,N_2458,N_2701);
or U3857 (N_3857,N_2539,N_2919);
nor U3858 (N_3858,N_2210,N_2218);
and U3859 (N_3859,N_2733,N_2436);
xor U3860 (N_3860,N_2917,N_2527);
nand U3861 (N_3861,N_2465,N_2256);
or U3862 (N_3862,N_2129,N_2357);
nor U3863 (N_3863,N_2874,N_2347);
or U3864 (N_3864,N_2491,N_2314);
and U3865 (N_3865,N_2960,N_2363);
nand U3866 (N_3866,N_2198,N_2985);
or U3867 (N_3867,N_2443,N_2719);
or U3868 (N_3868,N_2869,N_2994);
nand U3869 (N_3869,N_2669,N_2577);
xnor U3870 (N_3870,N_2919,N_2197);
or U3871 (N_3871,N_2950,N_2998);
nor U3872 (N_3872,N_2062,N_2678);
nand U3873 (N_3873,N_2947,N_2717);
or U3874 (N_3874,N_2071,N_2863);
or U3875 (N_3875,N_2708,N_2651);
and U3876 (N_3876,N_2597,N_2842);
nor U3877 (N_3877,N_2245,N_2993);
and U3878 (N_3878,N_2610,N_2657);
nand U3879 (N_3879,N_2511,N_2543);
and U3880 (N_3880,N_2269,N_2173);
and U3881 (N_3881,N_2486,N_2961);
or U3882 (N_3882,N_2786,N_2602);
and U3883 (N_3883,N_2070,N_2018);
nor U3884 (N_3884,N_2459,N_2325);
nor U3885 (N_3885,N_2302,N_2676);
nand U3886 (N_3886,N_2773,N_2278);
nor U3887 (N_3887,N_2551,N_2496);
xor U3888 (N_3888,N_2934,N_2250);
xnor U3889 (N_3889,N_2324,N_2896);
nor U3890 (N_3890,N_2250,N_2821);
and U3891 (N_3891,N_2656,N_2854);
nand U3892 (N_3892,N_2224,N_2577);
or U3893 (N_3893,N_2584,N_2429);
or U3894 (N_3894,N_2182,N_2757);
and U3895 (N_3895,N_2238,N_2291);
nand U3896 (N_3896,N_2029,N_2458);
nor U3897 (N_3897,N_2199,N_2723);
nor U3898 (N_3898,N_2072,N_2422);
nand U3899 (N_3899,N_2289,N_2878);
nand U3900 (N_3900,N_2082,N_2051);
and U3901 (N_3901,N_2327,N_2796);
nand U3902 (N_3902,N_2269,N_2059);
nand U3903 (N_3903,N_2638,N_2932);
nor U3904 (N_3904,N_2201,N_2698);
nand U3905 (N_3905,N_2684,N_2527);
nand U3906 (N_3906,N_2730,N_2039);
nand U3907 (N_3907,N_2763,N_2761);
and U3908 (N_3908,N_2181,N_2930);
and U3909 (N_3909,N_2547,N_2217);
or U3910 (N_3910,N_2088,N_2468);
nor U3911 (N_3911,N_2538,N_2573);
or U3912 (N_3912,N_2014,N_2171);
nor U3913 (N_3913,N_2932,N_2548);
or U3914 (N_3914,N_2708,N_2240);
nand U3915 (N_3915,N_2306,N_2876);
nand U3916 (N_3916,N_2426,N_2248);
nor U3917 (N_3917,N_2071,N_2074);
xnor U3918 (N_3918,N_2704,N_2128);
or U3919 (N_3919,N_2644,N_2460);
nor U3920 (N_3920,N_2374,N_2360);
or U3921 (N_3921,N_2216,N_2629);
and U3922 (N_3922,N_2681,N_2646);
nor U3923 (N_3923,N_2604,N_2242);
or U3924 (N_3924,N_2625,N_2889);
or U3925 (N_3925,N_2108,N_2048);
nor U3926 (N_3926,N_2491,N_2202);
or U3927 (N_3927,N_2252,N_2290);
and U3928 (N_3928,N_2877,N_2120);
nor U3929 (N_3929,N_2602,N_2734);
nor U3930 (N_3930,N_2822,N_2775);
or U3931 (N_3931,N_2015,N_2690);
and U3932 (N_3932,N_2486,N_2034);
and U3933 (N_3933,N_2922,N_2085);
nor U3934 (N_3934,N_2644,N_2182);
nand U3935 (N_3935,N_2762,N_2353);
nor U3936 (N_3936,N_2496,N_2066);
nand U3937 (N_3937,N_2182,N_2699);
nor U3938 (N_3938,N_2443,N_2348);
and U3939 (N_3939,N_2667,N_2081);
nand U3940 (N_3940,N_2476,N_2530);
or U3941 (N_3941,N_2824,N_2236);
and U3942 (N_3942,N_2466,N_2758);
or U3943 (N_3943,N_2866,N_2557);
and U3944 (N_3944,N_2074,N_2667);
or U3945 (N_3945,N_2189,N_2678);
nor U3946 (N_3946,N_2895,N_2987);
and U3947 (N_3947,N_2037,N_2477);
or U3948 (N_3948,N_2972,N_2130);
and U3949 (N_3949,N_2568,N_2258);
and U3950 (N_3950,N_2296,N_2350);
nand U3951 (N_3951,N_2537,N_2223);
nor U3952 (N_3952,N_2759,N_2259);
nor U3953 (N_3953,N_2538,N_2146);
or U3954 (N_3954,N_2538,N_2364);
or U3955 (N_3955,N_2618,N_2834);
nand U3956 (N_3956,N_2318,N_2539);
nand U3957 (N_3957,N_2049,N_2566);
nor U3958 (N_3958,N_2894,N_2726);
or U3959 (N_3959,N_2254,N_2810);
nand U3960 (N_3960,N_2811,N_2123);
and U3961 (N_3961,N_2794,N_2477);
nor U3962 (N_3962,N_2623,N_2861);
nand U3963 (N_3963,N_2953,N_2868);
nand U3964 (N_3964,N_2742,N_2975);
nand U3965 (N_3965,N_2949,N_2290);
or U3966 (N_3966,N_2979,N_2371);
and U3967 (N_3967,N_2063,N_2392);
nor U3968 (N_3968,N_2363,N_2040);
or U3969 (N_3969,N_2859,N_2505);
and U3970 (N_3970,N_2302,N_2328);
or U3971 (N_3971,N_2853,N_2024);
or U3972 (N_3972,N_2891,N_2409);
nor U3973 (N_3973,N_2042,N_2618);
nand U3974 (N_3974,N_2687,N_2518);
nor U3975 (N_3975,N_2365,N_2524);
nand U3976 (N_3976,N_2494,N_2575);
and U3977 (N_3977,N_2439,N_2641);
nor U3978 (N_3978,N_2287,N_2185);
and U3979 (N_3979,N_2085,N_2759);
nor U3980 (N_3980,N_2537,N_2675);
xnor U3981 (N_3981,N_2286,N_2691);
and U3982 (N_3982,N_2983,N_2859);
and U3983 (N_3983,N_2969,N_2961);
or U3984 (N_3984,N_2977,N_2623);
nand U3985 (N_3985,N_2751,N_2418);
nand U3986 (N_3986,N_2868,N_2085);
nand U3987 (N_3987,N_2077,N_2802);
and U3988 (N_3988,N_2707,N_2502);
and U3989 (N_3989,N_2509,N_2169);
and U3990 (N_3990,N_2349,N_2843);
or U3991 (N_3991,N_2998,N_2194);
or U3992 (N_3992,N_2976,N_2894);
nor U3993 (N_3993,N_2707,N_2383);
and U3994 (N_3994,N_2725,N_2373);
and U3995 (N_3995,N_2472,N_2275);
and U3996 (N_3996,N_2006,N_2407);
and U3997 (N_3997,N_2167,N_2525);
nand U3998 (N_3998,N_2323,N_2857);
xor U3999 (N_3999,N_2155,N_2785);
xnor U4000 (N_4000,N_3270,N_3027);
and U4001 (N_4001,N_3300,N_3405);
or U4002 (N_4002,N_3559,N_3040);
nor U4003 (N_4003,N_3606,N_3190);
nand U4004 (N_4004,N_3883,N_3809);
xor U4005 (N_4005,N_3851,N_3562);
nand U4006 (N_4006,N_3867,N_3574);
or U4007 (N_4007,N_3039,N_3436);
nand U4008 (N_4008,N_3875,N_3331);
nand U4009 (N_4009,N_3191,N_3912);
and U4010 (N_4010,N_3825,N_3857);
or U4011 (N_4011,N_3662,N_3595);
nor U4012 (N_4012,N_3048,N_3236);
and U4013 (N_4013,N_3090,N_3541);
and U4014 (N_4014,N_3426,N_3406);
nor U4015 (N_4015,N_3959,N_3932);
nand U4016 (N_4016,N_3686,N_3837);
nor U4017 (N_4017,N_3336,N_3395);
or U4018 (N_4018,N_3946,N_3636);
nand U4019 (N_4019,N_3930,N_3112);
nor U4020 (N_4020,N_3613,N_3435);
or U4021 (N_4021,N_3420,N_3326);
and U4022 (N_4022,N_3088,N_3251);
nand U4023 (N_4023,N_3836,N_3294);
nand U4024 (N_4024,N_3681,N_3460);
nor U4025 (N_4025,N_3927,N_3659);
nand U4026 (N_4026,N_3956,N_3709);
and U4027 (N_4027,N_3219,N_3340);
nand U4028 (N_4028,N_3753,N_3441);
nor U4029 (N_4029,N_3532,N_3856);
and U4030 (N_4030,N_3063,N_3355);
nor U4031 (N_4031,N_3119,N_3175);
nand U4032 (N_4032,N_3644,N_3120);
nand U4033 (N_4033,N_3128,N_3020);
xor U4034 (N_4034,N_3747,N_3834);
and U4035 (N_4035,N_3670,N_3873);
or U4036 (N_4036,N_3654,N_3743);
nor U4037 (N_4037,N_3168,N_3019);
nand U4038 (N_4038,N_3131,N_3201);
nor U4039 (N_4039,N_3230,N_3638);
xnor U4040 (N_4040,N_3003,N_3671);
nor U4041 (N_4041,N_3576,N_3879);
nand U4042 (N_4042,N_3023,N_3471);
nand U4043 (N_4043,N_3192,N_3101);
nand U4044 (N_4044,N_3596,N_3727);
and U4045 (N_4045,N_3194,N_3418);
and U4046 (N_4046,N_3521,N_3216);
and U4047 (N_4047,N_3695,N_3828);
or U4048 (N_4048,N_3928,N_3892);
and U4049 (N_4049,N_3459,N_3153);
or U4050 (N_4050,N_3220,N_3782);
nand U4051 (N_4051,N_3433,N_3047);
nand U4052 (N_4052,N_3007,N_3379);
nand U4053 (N_4053,N_3292,N_3324);
and U4054 (N_4054,N_3165,N_3132);
nor U4055 (N_4055,N_3762,N_3456);
and U4056 (N_4056,N_3731,N_3372);
nand U4057 (N_4057,N_3184,N_3622);
nor U4058 (N_4058,N_3462,N_3213);
nor U4059 (N_4059,N_3854,N_3560);
or U4060 (N_4060,N_3965,N_3181);
and U4061 (N_4061,N_3581,N_3949);
or U4062 (N_4062,N_3641,N_3899);
nand U4063 (N_4063,N_3672,N_3885);
or U4064 (N_4064,N_3751,N_3086);
nor U4065 (N_4065,N_3350,N_3640);
and U4066 (N_4066,N_3908,N_3818);
nor U4067 (N_4067,N_3226,N_3035);
and U4068 (N_4068,N_3732,N_3455);
nand U4069 (N_4069,N_3780,N_3994);
xor U4070 (N_4070,N_3208,N_3593);
nor U4071 (N_4071,N_3682,N_3363);
nor U4072 (N_4072,N_3673,N_3282);
nand U4073 (N_4073,N_3787,N_3133);
nand U4074 (N_4074,N_3152,N_3764);
and U4075 (N_4075,N_3164,N_3888);
nor U4076 (N_4076,N_3900,N_3674);
or U4077 (N_4077,N_3632,N_3617);
or U4078 (N_4078,N_3947,N_3159);
and U4079 (N_4079,N_3445,N_3345);
nor U4080 (N_4080,N_3820,N_3609);
nand U4081 (N_4081,N_3136,N_3468);
nand U4082 (N_4082,N_3470,N_3806);
nand U4083 (N_4083,N_3333,N_3493);
and U4084 (N_4084,N_3943,N_3006);
nor U4085 (N_4085,N_3678,N_3683);
or U4086 (N_4086,N_3388,N_3091);
nor U4087 (N_4087,N_3948,N_3146);
and U4088 (N_4088,N_3733,N_3328);
and U4089 (N_4089,N_3171,N_3921);
or U4090 (N_4090,N_3688,N_3805);
or U4091 (N_4091,N_3620,N_3938);
nand U4092 (N_4092,N_3740,N_3111);
nor U4093 (N_4093,N_3001,N_3509);
or U4094 (N_4094,N_3123,N_3544);
nand U4095 (N_4095,N_3660,N_3561);
or U4096 (N_4096,N_3630,N_3701);
nand U4097 (N_4097,N_3500,N_3793);
xor U4098 (N_4098,N_3507,N_3629);
and U4099 (N_4099,N_3718,N_3481);
or U4100 (N_4100,N_3483,N_3295);
or U4101 (N_4101,N_3502,N_3030);
nor U4102 (N_4102,N_3619,N_3266);
nand U4103 (N_4103,N_3401,N_3341);
nor U4104 (N_4104,N_3317,N_3477);
or U4105 (N_4105,N_3204,N_3827);
nor U4106 (N_4106,N_3163,N_3774);
or U4107 (N_4107,N_3643,N_3071);
nor U4108 (N_4108,N_3278,N_3982);
or U4109 (N_4109,N_3752,N_3992);
nand U4110 (N_4110,N_3253,N_3303);
and U4111 (N_4111,N_3375,N_3017);
nand U4112 (N_4112,N_3097,N_3922);
nand U4113 (N_4113,N_3438,N_3987);
nor U4114 (N_4114,N_3423,N_3575);
and U4115 (N_4115,N_3931,N_3816);
nand U4116 (N_4116,N_3657,N_3222);
and U4117 (N_4117,N_3891,N_3840);
nor U4118 (N_4118,N_3627,N_3392);
nor U4119 (N_4119,N_3158,N_3316);
and U4120 (N_4120,N_3410,N_3556);
nor U4121 (N_4121,N_3980,N_3868);
and U4122 (N_4122,N_3140,N_3663);
nand U4123 (N_4123,N_3099,N_3797);
or U4124 (N_4124,N_3170,N_3103);
nor U4125 (N_4125,N_3991,N_3371);
and U4126 (N_4126,N_3461,N_3916);
nand U4127 (N_4127,N_3605,N_3722);
nor U4128 (N_4128,N_3070,N_3193);
nand U4129 (N_4129,N_3254,N_3188);
nor U4130 (N_4130,N_3092,N_3325);
and U4131 (N_4131,N_3452,N_3697);
nor U4132 (N_4132,N_3304,N_3963);
and U4133 (N_4133,N_3690,N_3053);
nand U4134 (N_4134,N_3506,N_3069);
or U4135 (N_4135,N_3463,N_3050);
or U4136 (N_4136,N_3218,N_3798);
nor U4137 (N_4137,N_3894,N_3967);
and U4138 (N_4138,N_3385,N_3079);
nand U4139 (N_4139,N_3961,N_3234);
nand U4140 (N_4140,N_3784,N_3275);
nand U4141 (N_4141,N_3167,N_3373);
nand U4142 (N_4142,N_3364,N_3056);
or U4143 (N_4143,N_3450,N_3298);
nand U4144 (N_4144,N_3589,N_3439);
or U4145 (N_4145,N_3978,N_3497);
nor U4146 (N_4146,N_3166,N_3279);
and U4147 (N_4147,N_3878,N_3807);
and U4148 (N_4148,N_3511,N_3425);
nand U4149 (N_4149,N_3923,N_3842);
nor U4150 (N_4150,N_3647,N_3615);
or U4151 (N_4151,N_3874,N_3272);
xor U4152 (N_4152,N_3705,N_3361);
nand U4153 (N_4153,N_3434,N_3687);
nand U4154 (N_4154,N_3501,N_3046);
and U4155 (N_4155,N_3065,N_3513);
and U4156 (N_4156,N_3107,N_3238);
and U4157 (N_4157,N_3149,N_3397);
or U4158 (N_4158,N_3999,N_3646);
nand U4159 (N_4159,N_3198,N_3905);
xnor U4160 (N_4160,N_3320,N_3739);
nor U4161 (N_4161,N_3877,N_3958);
nand U4162 (N_4162,N_3799,N_3221);
nand U4163 (N_4163,N_3383,N_3839);
or U4164 (N_4164,N_3485,N_3239);
nor U4165 (N_4165,N_3349,N_3206);
nand U4166 (N_4166,N_3637,N_3977);
nand U4167 (N_4167,N_3259,N_3391);
and U4168 (N_4168,N_3849,N_3016);
and U4169 (N_4169,N_3095,N_3384);
or U4170 (N_4170,N_3172,N_3941);
nand U4171 (N_4171,N_3680,N_3366);
nor U4172 (N_4172,N_3360,N_3548);
and U4173 (N_4173,N_3811,N_3783);
nor U4174 (N_4174,N_3995,N_3726);
or U4175 (N_4175,N_3015,N_3712);
and U4176 (N_4176,N_3389,N_3742);
or U4177 (N_4177,N_3962,N_3285);
nor U4178 (N_4178,N_3792,N_3309);
and U4179 (N_4179,N_3546,N_3321);
nand U4180 (N_4180,N_3018,N_3185);
nand U4181 (N_4181,N_3415,N_3318);
or U4182 (N_4182,N_3555,N_3414);
or U4183 (N_4183,N_3058,N_3177);
nor U4184 (N_4184,N_3422,N_3872);
nor U4185 (N_4185,N_3429,N_3665);
or U4186 (N_4186,N_3209,N_3494);
xor U4187 (N_4187,N_3145,N_3076);
nor U4188 (N_4188,N_3247,N_3297);
nand U4189 (N_4189,N_3844,N_3186);
and U4190 (N_4190,N_3344,N_3700);
nand U4191 (N_4191,N_3979,N_3808);
nand U4192 (N_4192,N_3248,N_3728);
nor U4193 (N_4193,N_3668,N_3903);
or U4194 (N_4194,N_3975,N_3684);
and U4195 (N_4195,N_3520,N_3597);
nand U4196 (N_4196,N_3458,N_3582);
or U4197 (N_4197,N_3108,N_3926);
nand U4198 (N_4198,N_3523,N_3486);
nor U4199 (N_4199,N_3710,N_3760);
or U4200 (N_4200,N_3072,N_3860);
nor U4201 (N_4201,N_3954,N_3729);
or U4202 (N_4202,N_3081,N_3639);
nand U4203 (N_4203,N_3524,N_3538);
nor U4204 (N_4204,N_3587,N_3886);
and U4205 (N_4205,N_3085,N_3504);
and U4206 (N_4206,N_3199,N_3910);
nor U4207 (N_4207,N_3604,N_3887);
nand U4208 (N_4208,N_3557,N_3082);
xor U4209 (N_4209,N_3531,N_3658);
and U4210 (N_4210,N_3351,N_3386);
nor U4211 (N_4211,N_3368,N_3855);
nor U4212 (N_4212,N_3770,N_3256);
nor U4213 (N_4213,N_3565,N_3723);
nor U4214 (N_4214,N_3346,N_3583);
nand U4215 (N_4215,N_3358,N_3735);
nor U4216 (N_4216,N_3096,N_3314);
nand U4217 (N_4217,N_3424,N_3319);
nand U4218 (N_4218,N_3154,N_3713);
nor U4219 (N_4219,N_3568,N_3696);
or U4220 (N_4220,N_3578,N_3871);
or U4221 (N_4221,N_3968,N_3866);
and U4222 (N_4222,N_3276,N_3600);
xor U4223 (N_4223,N_3518,N_3214);
nor U4224 (N_4224,N_3525,N_3540);
or U4225 (N_4225,N_3655,N_3161);
nand U4226 (N_4226,N_3196,N_3308);
nor U4227 (N_4227,N_3530,N_3858);
nand U4228 (N_4228,N_3109,N_3042);
xnor U4229 (N_4229,N_3289,N_3265);
nor U4230 (N_4230,N_3974,N_3902);
nor U4231 (N_4231,N_3178,N_3964);
nor U4232 (N_4232,N_3411,N_3933);
or U4233 (N_4233,N_3400,N_3261);
and U4234 (N_4234,N_3950,N_3551);
or U4235 (N_4235,N_3488,N_3353);
nand U4236 (N_4236,N_3648,N_3362);
nor U4237 (N_4237,N_3431,N_3491);
or U4238 (N_4238,N_3078,N_3898);
nor U4239 (N_4239,N_3651,N_3692);
and U4240 (N_4240,N_3614,N_3989);
or U4241 (N_4241,N_3129,N_3267);
nor U4242 (N_4242,N_3527,N_3352);
nor U4243 (N_4243,N_3759,N_3232);
nand U4244 (N_4244,N_3610,N_3881);
and U4245 (N_4245,N_3066,N_3327);
nand U4246 (N_4246,N_3124,N_3484);
xnor U4247 (N_4247,N_3847,N_3767);
and U4248 (N_4248,N_3835,N_3707);
and U4249 (N_4249,N_3077,N_3197);
nand U4250 (N_4250,N_3374,N_3517);
nand U4251 (N_4251,N_3955,N_3832);
nor U4252 (N_4252,N_3758,N_3051);
nor U4253 (N_4253,N_3734,N_3339);
nor U4254 (N_4254,N_3675,N_3183);
nor U4255 (N_4255,N_3624,N_3939);
nor U4256 (N_4256,N_3252,N_3679);
nor U4257 (N_4257,N_3510,N_3880);
nor U4258 (N_4258,N_3157,N_3570);
or U4259 (N_4259,N_3473,N_3223);
nand U4260 (N_4260,N_3785,N_3026);
and U4261 (N_4261,N_3380,N_3716);
nor U4262 (N_4262,N_3169,N_3296);
nor U4263 (N_4263,N_3915,N_3031);
or U4264 (N_4264,N_3233,N_3376);
nand U4265 (N_4265,N_3093,N_3976);
nor U4266 (N_4266,N_3616,N_3599);
nand U4267 (N_4267,N_3160,N_3853);
nand U4268 (N_4268,N_3117,N_3087);
or U4269 (N_4269,N_3717,N_3571);
nor U4270 (N_4270,N_3281,N_3393);
nor U4271 (N_4271,N_3846,N_3579);
nand U4272 (N_4272,N_3904,N_3761);
and U4273 (N_4273,N_3156,N_3572);
or U4274 (N_4274,N_3075,N_3567);
and U4275 (N_4275,N_3588,N_3553);
or U4276 (N_4276,N_3408,N_3356);
or U4277 (N_4277,N_3952,N_3508);
or U4278 (N_4278,N_3529,N_3498);
nand U4279 (N_4279,N_3496,N_3914);
nor U4280 (N_4280,N_3741,N_3286);
and U4281 (N_4281,N_3765,N_3049);
and U4282 (N_4282,N_3135,N_3273);
nor U4283 (N_4283,N_3147,N_3310);
and U4284 (N_4284,N_3134,N_3307);
and U4285 (N_4285,N_3795,N_3611);
xor U4286 (N_4286,N_3843,N_3480);
and U4287 (N_4287,N_3306,N_3812);
xor U4288 (N_4288,N_3487,N_3449);
nand U4289 (N_4289,N_3357,N_3021);
or U4290 (N_4290,N_3004,N_3791);
nor U4291 (N_4291,N_3736,N_3802);
nor U4292 (N_4292,N_3427,N_3882);
nand U4293 (N_4293,N_3769,N_3519);
and U4294 (N_4294,N_3211,N_3584);
nand U4295 (N_4295,N_3257,N_3499);
nor U4296 (N_4296,N_3522,N_3864);
xnor U4297 (N_4297,N_3210,N_3036);
nor U4298 (N_4298,N_3466,N_3002);
nand U4299 (N_4299,N_3789,N_3585);
or U4300 (N_4300,N_3944,N_3264);
nand U4301 (N_4301,N_3008,N_3876);
nor U4302 (N_4302,N_3246,N_3777);
xor U4303 (N_4303,N_3815,N_3187);
and U4304 (N_4304,N_3010,N_3550);
nand U4305 (N_4305,N_3746,N_3446);
xor U4306 (N_4306,N_3890,N_3012);
nor U4307 (N_4307,N_3800,N_3444);
nand U4308 (N_4308,N_3953,N_3786);
nand U4309 (N_4309,N_3258,N_3838);
or U4310 (N_4310,N_3334,N_3503);
or U4311 (N_4311,N_3116,N_3301);
or U4312 (N_4312,N_3409,N_3073);
and U4313 (N_4313,N_3542,N_3896);
or U4314 (N_4314,N_3775,N_3173);
and U4315 (N_4315,N_3055,N_3598);
or U4316 (N_4316,N_3533,N_3635);
nor U4317 (N_4317,N_3537,N_3033);
nor U4318 (N_4318,N_3271,N_3906);
nor U4319 (N_4319,N_3057,N_3863);
or U4320 (N_4320,N_3750,N_3212);
nor U4321 (N_4321,N_3677,N_3725);
and U4322 (N_4322,N_3241,N_3195);
nand U4323 (N_4323,N_3889,N_3378);
nor U4324 (N_4324,N_3794,N_3676);
or U4325 (N_4325,N_3407,N_3179);
nand U4326 (N_4326,N_3607,N_3623);
and U4327 (N_4327,N_3102,N_3702);
and U4328 (N_4328,N_3884,N_3390);
nor U4329 (N_4329,N_3972,N_3924);
or U4330 (N_4330,N_3283,N_3831);
and U4331 (N_4331,N_3404,N_3901);
nand U4332 (N_4332,N_3951,N_3650);
or U4333 (N_4333,N_3329,N_3826);
nor U4334 (N_4334,N_3694,N_3105);
and U4335 (N_4335,N_3564,N_3810);
or U4336 (N_4336,N_3457,N_3067);
nor U4337 (N_4337,N_3098,N_3859);
nor U4338 (N_4338,N_3437,N_3022);
or U4339 (N_4339,N_3269,N_3768);
nand U4340 (N_4340,N_3203,N_3115);
nand U4341 (N_4341,N_3689,N_3287);
nand U4342 (N_4342,N_3505,N_3412);
nor U4343 (N_4343,N_3652,N_3416);
or U4344 (N_4344,N_3074,N_3645);
nor U4345 (N_4345,N_3060,N_3014);
xnor U4346 (N_4346,N_3649,N_3748);
nand U4347 (N_4347,N_3447,N_3998);
or U4348 (N_4348,N_3249,N_3453);
and U4349 (N_4349,N_3005,N_3824);
nor U4350 (N_4350,N_3763,N_3284);
or U4351 (N_4351,N_3817,N_3207);
or U4352 (N_4352,N_3240,N_3162);
nor U4353 (N_4353,N_3515,N_3969);
nand U4354 (N_4354,N_3291,N_3813);
or U4355 (N_4355,N_3413,N_3942);
nand U4356 (N_4356,N_3142,N_3322);
nand U4357 (N_4357,N_3382,N_3029);
nand U4358 (N_4358,N_3569,N_3492);
nor U4359 (N_4359,N_3299,N_3981);
nand U4360 (N_4360,N_3714,N_3244);
nand U4361 (N_4361,N_3189,N_3653);
xor U4362 (N_4362,N_3268,N_3469);
and U4363 (N_4363,N_3845,N_3667);
and U4364 (N_4364,N_3454,N_3305);
nor U4365 (N_4365,N_3034,N_3394);
or U4366 (N_4366,N_3430,N_3642);
and U4367 (N_4367,N_3144,N_3052);
or U4368 (N_4368,N_3313,N_3343);
xor U4369 (N_4369,N_3428,N_3476);
nand U4370 (N_4370,N_3474,N_3054);
nand U4371 (N_4371,N_3536,N_3061);
nor U4372 (N_4372,N_3543,N_3495);
or U4373 (N_4373,N_3862,N_3591);
or U4374 (N_4374,N_3822,N_3586);
or U4375 (N_4375,N_3790,N_3526);
nor U4376 (N_4376,N_3365,N_3801);
or U4377 (N_4377,N_3242,N_3841);
nor U4378 (N_4378,N_3971,N_3829);
nand U4379 (N_4379,N_3897,N_3370);
nand U4380 (N_4380,N_3895,N_3068);
nand U4381 (N_4381,N_3089,N_3465);
nand U4382 (N_4382,N_3479,N_3960);
or U4383 (N_4383,N_3514,N_3985);
and U4384 (N_4384,N_3997,N_3122);
or U4385 (N_4385,N_3293,N_3094);
nor U4386 (N_4386,N_3766,N_3781);
or U4387 (N_4387,N_3118,N_3626);
nor U4388 (N_4388,N_3592,N_3545);
or U4389 (N_4389,N_3633,N_3940);
and U4390 (N_4390,N_3000,N_3909);
or U4391 (N_4391,N_3125,N_3262);
nor U4392 (N_4392,N_3130,N_3970);
nand U4393 (N_4393,N_3552,N_3715);
nor U4394 (N_4394,N_3139,N_3621);
or U4395 (N_4395,N_3549,N_3554);
or U4396 (N_4396,N_3243,N_3440);
and U4397 (N_4397,N_3011,N_3573);
or U4398 (N_4398,N_3749,N_3467);
or U4399 (N_4399,N_3983,N_3711);
or U4400 (N_4400,N_3217,N_3302);
nor U4401 (N_4401,N_3323,N_3402);
nand U4402 (N_4402,N_3369,N_3064);
and U4403 (N_4403,N_3566,N_3698);
or U4404 (N_4404,N_3730,N_3148);
or U4405 (N_4405,N_3347,N_3041);
nor U4406 (N_4406,N_3850,N_3594);
nor U4407 (N_4407,N_3993,N_3009);
nor U4408 (N_4408,N_3603,N_3126);
or U4409 (N_4409,N_3110,N_3337);
xnor U4410 (N_4410,N_3925,N_3451);
nor U4411 (N_4411,N_3539,N_3945);
xnor U4412 (N_4412,N_3990,N_3803);
or U4413 (N_4413,N_3547,N_3235);
nor U4414 (N_4414,N_3100,N_3315);
and U4415 (N_4415,N_3848,N_3771);
nor U4416 (N_4416,N_3907,N_3691);
and U4417 (N_4417,N_3776,N_3202);
xnor U4418 (N_4418,N_3038,N_3044);
or U4419 (N_4419,N_3720,N_3478);
xnor U4420 (N_4420,N_3744,N_3708);
nor U4421 (N_4421,N_3819,N_3280);
nor U4422 (N_4422,N_3988,N_3754);
nor U4423 (N_4423,N_3490,N_3399);
nor U4424 (N_4424,N_3666,N_3704);
xor U4425 (N_4425,N_3934,N_3417);
and U4426 (N_4426,N_3516,N_3475);
xnor U4427 (N_4427,N_3288,N_3260);
nor U4428 (N_4428,N_3277,N_3229);
nor U4429 (N_4429,N_3037,N_3200);
nand U4430 (N_4430,N_3535,N_3917);
nand U4431 (N_4431,N_3861,N_3150);
nor U4432 (N_4432,N_3755,N_3918);
nand U4433 (N_4433,N_3104,N_3330);
nor U4434 (N_4434,N_3772,N_3121);
nor U4435 (N_4435,N_3577,N_3359);
or U4436 (N_4436,N_3865,N_3778);
nor U4437 (N_4437,N_3719,N_3332);
nor U4438 (N_4438,N_3724,N_3274);
nand U4439 (N_4439,N_3984,N_3669);
or U4440 (N_4440,N_3664,N_3127);
nand U4441 (N_4441,N_3174,N_3608);
nor U4442 (N_4442,N_3788,N_3448);
nor U4443 (N_4443,N_3986,N_3348);
nand U4444 (N_4444,N_3237,N_3432);
nand U4445 (N_4445,N_3113,N_3245);
nor U4446 (N_4446,N_3354,N_3141);
nor U4447 (N_4447,N_3738,N_3137);
and U4448 (N_4448,N_3312,N_3601);
and U4449 (N_4449,N_3143,N_3263);
and U4450 (N_4450,N_3464,N_3106);
nor U4451 (N_4451,N_3602,N_3224);
or U4452 (N_4452,N_3737,N_3396);
nand U4453 (N_4453,N_3893,N_3114);
or U4454 (N_4454,N_3180,N_3138);
and U4455 (N_4455,N_3699,N_3580);
or U4456 (N_4456,N_3290,N_3756);
nor U4457 (N_4457,N_3387,N_3852);
nand U4458 (N_4458,N_3796,N_3913);
or U4459 (N_4459,N_3830,N_3869);
nand U4460 (N_4460,N_3013,N_3528);
nand U4461 (N_4461,N_3176,N_3773);
nor U4462 (N_4462,N_3335,N_3215);
nor U4463 (N_4463,N_3024,N_3377);
nand U4464 (N_4464,N_3062,N_3661);
or U4465 (N_4465,N_3182,N_3966);
nand U4466 (N_4466,N_3957,N_3472);
nand U4467 (N_4467,N_3757,N_3618);
nor U4468 (N_4468,N_3631,N_3398);
nor U4469 (N_4469,N_3421,N_3703);
xnor U4470 (N_4470,N_3804,N_3628);
or U4471 (N_4471,N_3227,N_3381);
and U4472 (N_4472,N_3032,N_3059);
nor U4473 (N_4473,N_3255,N_3419);
nor U4474 (N_4474,N_3693,N_3721);
or U4475 (N_4475,N_3814,N_3045);
nand U4476 (N_4476,N_3656,N_3084);
and U4477 (N_4477,N_3973,N_3534);
or U4478 (N_4478,N_3342,N_3779);
nor U4479 (N_4479,N_3745,N_3920);
nand U4480 (N_4480,N_3911,N_3833);
or U4481 (N_4481,N_3311,N_3706);
and U4482 (N_4482,N_3612,N_3367);
nand U4483 (N_4483,N_3028,N_3443);
and U4484 (N_4484,N_3205,N_3870);
nand U4485 (N_4485,N_3442,N_3935);
nand U4486 (N_4486,N_3338,N_3043);
xnor U4487 (N_4487,N_3625,N_3403);
or U4488 (N_4488,N_3228,N_3634);
nand U4489 (N_4489,N_3025,N_3155);
or U4490 (N_4490,N_3231,N_3083);
or U4491 (N_4491,N_3919,N_3558);
nand U4492 (N_4492,N_3225,N_3590);
and U4493 (N_4493,N_3512,N_3929);
or U4494 (N_4494,N_3936,N_3685);
nand U4495 (N_4495,N_3482,N_3151);
or U4496 (N_4496,N_3823,N_3563);
nor U4497 (N_4497,N_3250,N_3489);
or U4498 (N_4498,N_3821,N_3996);
nor U4499 (N_4499,N_3080,N_3937);
and U4500 (N_4500,N_3987,N_3318);
or U4501 (N_4501,N_3879,N_3555);
nor U4502 (N_4502,N_3144,N_3494);
nor U4503 (N_4503,N_3807,N_3161);
and U4504 (N_4504,N_3591,N_3970);
nand U4505 (N_4505,N_3471,N_3539);
nand U4506 (N_4506,N_3070,N_3805);
nor U4507 (N_4507,N_3552,N_3081);
or U4508 (N_4508,N_3809,N_3924);
nand U4509 (N_4509,N_3461,N_3413);
nor U4510 (N_4510,N_3690,N_3399);
nor U4511 (N_4511,N_3938,N_3195);
or U4512 (N_4512,N_3814,N_3616);
nand U4513 (N_4513,N_3491,N_3471);
or U4514 (N_4514,N_3562,N_3346);
nor U4515 (N_4515,N_3921,N_3451);
nand U4516 (N_4516,N_3381,N_3625);
or U4517 (N_4517,N_3539,N_3894);
nor U4518 (N_4518,N_3939,N_3746);
nand U4519 (N_4519,N_3307,N_3924);
and U4520 (N_4520,N_3639,N_3296);
nand U4521 (N_4521,N_3865,N_3565);
and U4522 (N_4522,N_3694,N_3755);
nor U4523 (N_4523,N_3265,N_3946);
nand U4524 (N_4524,N_3143,N_3210);
nor U4525 (N_4525,N_3717,N_3257);
nand U4526 (N_4526,N_3923,N_3629);
and U4527 (N_4527,N_3821,N_3524);
or U4528 (N_4528,N_3161,N_3346);
nand U4529 (N_4529,N_3316,N_3105);
and U4530 (N_4530,N_3616,N_3239);
and U4531 (N_4531,N_3148,N_3538);
and U4532 (N_4532,N_3087,N_3886);
and U4533 (N_4533,N_3995,N_3266);
and U4534 (N_4534,N_3596,N_3346);
nand U4535 (N_4535,N_3593,N_3561);
and U4536 (N_4536,N_3014,N_3618);
nor U4537 (N_4537,N_3528,N_3116);
or U4538 (N_4538,N_3324,N_3061);
nor U4539 (N_4539,N_3493,N_3453);
or U4540 (N_4540,N_3607,N_3104);
nor U4541 (N_4541,N_3298,N_3664);
and U4542 (N_4542,N_3267,N_3768);
nand U4543 (N_4543,N_3947,N_3943);
or U4544 (N_4544,N_3681,N_3769);
nand U4545 (N_4545,N_3579,N_3334);
nand U4546 (N_4546,N_3397,N_3116);
or U4547 (N_4547,N_3073,N_3413);
nand U4548 (N_4548,N_3678,N_3045);
or U4549 (N_4549,N_3082,N_3766);
or U4550 (N_4550,N_3154,N_3551);
and U4551 (N_4551,N_3601,N_3798);
nand U4552 (N_4552,N_3906,N_3377);
nand U4553 (N_4553,N_3233,N_3203);
nor U4554 (N_4554,N_3766,N_3381);
or U4555 (N_4555,N_3652,N_3196);
or U4556 (N_4556,N_3857,N_3672);
or U4557 (N_4557,N_3596,N_3352);
xnor U4558 (N_4558,N_3689,N_3552);
nand U4559 (N_4559,N_3150,N_3380);
or U4560 (N_4560,N_3540,N_3799);
nand U4561 (N_4561,N_3380,N_3963);
and U4562 (N_4562,N_3209,N_3554);
nor U4563 (N_4563,N_3260,N_3373);
and U4564 (N_4564,N_3410,N_3458);
or U4565 (N_4565,N_3375,N_3317);
nand U4566 (N_4566,N_3950,N_3158);
xnor U4567 (N_4567,N_3719,N_3455);
or U4568 (N_4568,N_3985,N_3510);
nor U4569 (N_4569,N_3819,N_3586);
or U4570 (N_4570,N_3818,N_3389);
or U4571 (N_4571,N_3223,N_3721);
or U4572 (N_4572,N_3871,N_3604);
or U4573 (N_4573,N_3932,N_3641);
and U4574 (N_4574,N_3268,N_3409);
or U4575 (N_4575,N_3720,N_3179);
nor U4576 (N_4576,N_3252,N_3263);
or U4577 (N_4577,N_3310,N_3604);
nor U4578 (N_4578,N_3555,N_3823);
or U4579 (N_4579,N_3833,N_3347);
nand U4580 (N_4580,N_3896,N_3252);
nand U4581 (N_4581,N_3338,N_3921);
and U4582 (N_4582,N_3354,N_3967);
or U4583 (N_4583,N_3181,N_3631);
or U4584 (N_4584,N_3130,N_3500);
nor U4585 (N_4585,N_3299,N_3263);
or U4586 (N_4586,N_3097,N_3356);
or U4587 (N_4587,N_3937,N_3007);
or U4588 (N_4588,N_3636,N_3589);
nor U4589 (N_4589,N_3989,N_3687);
or U4590 (N_4590,N_3732,N_3704);
and U4591 (N_4591,N_3062,N_3023);
nor U4592 (N_4592,N_3254,N_3187);
nor U4593 (N_4593,N_3323,N_3723);
or U4594 (N_4594,N_3551,N_3662);
or U4595 (N_4595,N_3859,N_3515);
or U4596 (N_4596,N_3690,N_3586);
nor U4597 (N_4597,N_3286,N_3884);
nor U4598 (N_4598,N_3974,N_3511);
or U4599 (N_4599,N_3829,N_3979);
nand U4600 (N_4600,N_3759,N_3913);
or U4601 (N_4601,N_3037,N_3693);
nand U4602 (N_4602,N_3991,N_3662);
and U4603 (N_4603,N_3148,N_3135);
and U4604 (N_4604,N_3537,N_3475);
nor U4605 (N_4605,N_3107,N_3034);
or U4606 (N_4606,N_3420,N_3026);
nand U4607 (N_4607,N_3657,N_3655);
nand U4608 (N_4608,N_3160,N_3099);
nand U4609 (N_4609,N_3761,N_3396);
nand U4610 (N_4610,N_3179,N_3317);
nor U4611 (N_4611,N_3833,N_3251);
nand U4612 (N_4612,N_3021,N_3489);
and U4613 (N_4613,N_3683,N_3345);
nand U4614 (N_4614,N_3573,N_3313);
nand U4615 (N_4615,N_3293,N_3412);
nand U4616 (N_4616,N_3269,N_3529);
xor U4617 (N_4617,N_3433,N_3210);
or U4618 (N_4618,N_3567,N_3159);
nor U4619 (N_4619,N_3686,N_3745);
nor U4620 (N_4620,N_3155,N_3298);
nor U4621 (N_4621,N_3394,N_3585);
or U4622 (N_4622,N_3214,N_3684);
nor U4623 (N_4623,N_3967,N_3277);
nand U4624 (N_4624,N_3428,N_3949);
or U4625 (N_4625,N_3069,N_3454);
nor U4626 (N_4626,N_3629,N_3409);
or U4627 (N_4627,N_3581,N_3328);
or U4628 (N_4628,N_3287,N_3447);
nand U4629 (N_4629,N_3859,N_3342);
nor U4630 (N_4630,N_3198,N_3897);
and U4631 (N_4631,N_3594,N_3671);
nand U4632 (N_4632,N_3063,N_3020);
xor U4633 (N_4633,N_3088,N_3389);
and U4634 (N_4634,N_3694,N_3451);
or U4635 (N_4635,N_3889,N_3569);
and U4636 (N_4636,N_3021,N_3110);
nor U4637 (N_4637,N_3889,N_3160);
or U4638 (N_4638,N_3339,N_3428);
and U4639 (N_4639,N_3690,N_3305);
and U4640 (N_4640,N_3259,N_3875);
and U4641 (N_4641,N_3058,N_3424);
or U4642 (N_4642,N_3202,N_3279);
or U4643 (N_4643,N_3393,N_3585);
nor U4644 (N_4644,N_3420,N_3084);
or U4645 (N_4645,N_3564,N_3449);
nor U4646 (N_4646,N_3469,N_3102);
and U4647 (N_4647,N_3691,N_3069);
or U4648 (N_4648,N_3186,N_3129);
or U4649 (N_4649,N_3171,N_3007);
and U4650 (N_4650,N_3385,N_3145);
nand U4651 (N_4651,N_3557,N_3850);
nand U4652 (N_4652,N_3961,N_3211);
nor U4653 (N_4653,N_3184,N_3343);
and U4654 (N_4654,N_3917,N_3739);
or U4655 (N_4655,N_3308,N_3908);
and U4656 (N_4656,N_3235,N_3705);
and U4657 (N_4657,N_3204,N_3298);
nor U4658 (N_4658,N_3523,N_3715);
nor U4659 (N_4659,N_3957,N_3385);
xnor U4660 (N_4660,N_3692,N_3123);
nand U4661 (N_4661,N_3806,N_3375);
or U4662 (N_4662,N_3394,N_3254);
or U4663 (N_4663,N_3875,N_3743);
nor U4664 (N_4664,N_3719,N_3498);
nor U4665 (N_4665,N_3290,N_3842);
or U4666 (N_4666,N_3729,N_3657);
and U4667 (N_4667,N_3676,N_3514);
nand U4668 (N_4668,N_3988,N_3690);
and U4669 (N_4669,N_3603,N_3493);
and U4670 (N_4670,N_3584,N_3989);
nor U4671 (N_4671,N_3213,N_3841);
nor U4672 (N_4672,N_3196,N_3942);
nor U4673 (N_4673,N_3922,N_3850);
and U4674 (N_4674,N_3878,N_3279);
nor U4675 (N_4675,N_3871,N_3942);
nor U4676 (N_4676,N_3989,N_3718);
and U4677 (N_4677,N_3182,N_3991);
nand U4678 (N_4678,N_3414,N_3998);
nand U4679 (N_4679,N_3624,N_3963);
or U4680 (N_4680,N_3005,N_3871);
or U4681 (N_4681,N_3293,N_3926);
and U4682 (N_4682,N_3855,N_3259);
xnor U4683 (N_4683,N_3935,N_3233);
nand U4684 (N_4684,N_3735,N_3309);
nand U4685 (N_4685,N_3500,N_3806);
nand U4686 (N_4686,N_3866,N_3391);
nand U4687 (N_4687,N_3777,N_3775);
or U4688 (N_4688,N_3050,N_3669);
nand U4689 (N_4689,N_3765,N_3386);
nand U4690 (N_4690,N_3095,N_3308);
nand U4691 (N_4691,N_3651,N_3419);
or U4692 (N_4692,N_3798,N_3888);
and U4693 (N_4693,N_3934,N_3878);
and U4694 (N_4694,N_3426,N_3312);
and U4695 (N_4695,N_3029,N_3410);
nor U4696 (N_4696,N_3904,N_3773);
nand U4697 (N_4697,N_3540,N_3223);
nor U4698 (N_4698,N_3110,N_3460);
nor U4699 (N_4699,N_3545,N_3896);
or U4700 (N_4700,N_3348,N_3800);
nor U4701 (N_4701,N_3802,N_3903);
nor U4702 (N_4702,N_3488,N_3920);
or U4703 (N_4703,N_3438,N_3576);
and U4704 (N_4704,N_3907,N_3873);
nand U4705 (N_4705,N_3546,N_3289);
nand U4706 (N_4706,N_3240,N_3785);
nand U4707 (N_4707,N_3717,N_3703);
nand U4708 (N_4708,N_3372,N_3440);
nor U4709 (N_4709,N_3985,N_3818);
nand U4710 (N_4710,N_3206,N_3319);
and U4711 (N_4711,N_3707,N_3223);
and U4712 (N_4712,N_3837,N_3597);
or U4713 (N_4713,N_3155,N_3858);
nor U4714 (N_4714,N_3493,N_3313);
and U4715 (N_4715,N_3881,N_3168);
or U4716 (N_4716,N_3964,N_3705);
or U4717 (N_4717,N_3040,N_3488);
nand U4718 (N_4718,N_3966,N_3011);
and U4719 (N_4719,N_3161,N_3132);
nor U4720 (N_4720,N_3924,N_3439);
nand U4721 (N_4721,N_3054,N_3592);
and U4722 (N_4722,N_3556,N_3777);
nor U4723 (N_4723,N_3448,N_3413);
and U4724 (N_4724,N_3168,N_3166);
nor U4725 (N_4725,N_3442,N_3407);
nor U4726 (N_4726,N_3322,N_3160);
and U4727 (N_4727,N_3917,N_3153);
or U4728 (N_4728,N_3484,N_3794);
xor U4729 (N_4729,N_3509,N_3454);
nand U4730 (N_4730,N_3383,N_3160);
and U4731 (N_4731,N_3192,N_3493);
xnor U4732 (N_4732,N_3458,N_3273);
nand U4733 (N_4733,N_3166,N_3392);
and U4734 (N_4734,N_3302,N_3371);
or U4735 (N_4735,N_3816,N_3079);
and U4736 (N_4736,N_3277,N_3139);
nor U4737 (N_4737,N_3876,N_3202);
and U4738 (N_4738,N_3981,N_3048);
or U4739 (N_4739,N_3438,N_3693);
and U4740 (N_4740,N_3508,N_3592);
or U4741 (N_4741,N_3849,N_3568);
or U4742 (N_4742,N_3231,N_3518);
nand U4743 (N_4743,N_3499,N_3909);
or U4744 (N_4744,N_3903,N_3159);
nor U4745 (N_4745,N_3885,N_3040);
and U4746 (N_4746,N_3386,N_3380);
nor U4747 (N_4747,N_3975,N_3284);
and U4748 (N_4748,N_3453,N_3475);
and U4749 (N_4749,N_3596,N_3282);
nand U4750 (N_4750,N_3516,N_3453);
nand U4751 (N_4751,N_3121,N_3443);
or U4752 (N_4752,N_3049,N_3716);
nor U4753 (N_4753,N_3258,N_3151);
or U4754 (N_4754,N_3453,N_3206);
nand U4755 (N_4755,N_3654,N_3314);
nand U4756 (N_4756,N_3171,N_3216);
or U4757 (N_4757,N_3074,N_3988);
and U4758 (N_4758,N_3788,N_3610);
and U4759 (N_4759,N_3315,N_3711);
nand U4760 (N_4760,N_3671,N_3288);
xnor U4761 (N_4761,N_3922,N_3690);
xnor U4762 (N_4762,N_3189,N_3615);
nand U4763 (N_4763,N_3515,N_3268);
xnor U4764 (N_4764,N_3900,N_3010);
nor U4765 (N_4765,N_3542,N_3016);
or U4766 (N_4766,N_3996,N_3982);
and U4767 (N_4767,N_3633,N_3271);
nor U4768 (N_4768,N_3526,N_3043);
nand U4769 (N_4769,N_3573,N_3228);
and U4770 (N_4770,N_3461,N_3165);
nor U4771 (N_4771,N_3708,N_3049);
nand U4772 (N_4772,N_3733,N_3852);
nor U4773 (N_4773,N_3571,N_3104);
or U4774 (N_4774,N_3455,N_3024);
and U4775 (N_4775,N_3121,N_3643);
nor U4776 (N_4776,N_3945,N_3814);
and U4777 (N_4777,N_3539,N_3801);
nand U4778 (N_4778,N_3007,N_3197);
nor U4779 (N_4779,N_3984,N_3524);
nand U4780 (N_4780,N_3804,N_3605);
nand U4781 (N_4781,N_3273,N_3650);
nand U4782 (N_4782,N_3154,N_3307);
or U4783 (N_4783,N_3015,N_3156);
and U4784 (N_4784,N_3394,N_3774);
xor U4785 (N_4785,N_3217,N_3379);
and U4786 (N_4786,N_3931,N_3777);
or U4787 (N_4787,N_3488,N_3498);
nand U4788 (N_4788,N_3112,N_3582);
nand U4789 (N_4789,N_3187,N_3452);
and U4790 (N_4790,N_3410,N_3156);
or U4791 (N_4791,N_3474,N_3102);
or U4792 (N_4792,N_3670,N_3329);
and U4793 (N_4793,N_3709,N_3683);
or U4794 (N_4794,N_3443,N_3805);
nor U4795 (N_4795,N_3262,N_3950);
and U4796 (N_4796,N_3665,N_3195);
or U4797 (N_4797,N_3590,N_3467);
nor U4798 (N_4798,N_3778,N_3438);
and U4799 (N_4799,N_3439,N_3693);
and U4800 (N_4800,N_3206,N_3248);
nor U4801 (N_4801,N_3077,N_3035);
or U4802 (N_4802,N_3392,N_3282);
nor U4803 (N_4803,N_3592,N_3632);
nand U4804 (N_4804,N_3762,N_3422);
or U4805 (N_4805,N_3933,N_3985);
nand U4806 (N_4806,N_3858,N_3476);
or U4807 (N_4807,N_3832,N_3321);
or U4808 (N_4808,N_3699,N_3639);
nand U4809 (N_4809,N_3976,N_3542);
nor U4810 (N_4810,N_3976,N_3331);
nor U4811 (N_4811,N_3953,N_3857);
nor U4812 (N_4812,N_3409,N_3324);
or U4813 (N_4813,N_3603,N_3907);
and U4814 (N_4814,N_3159,N_3616);
and U4815 (N_4815,N_3510,N_3485);
and U4816 (N_4816,N_3032,N_3697);
nand U4817 (N_4817,N_3276,N_3098);
nand U4818 (N_4818,N_3983,N_3065);
nand U4819 (N_4819,N_3055,N_3804);
or U4820 (N_4820,N_3520,N_3627);
nor U4821 (N_4821,N_3884,N_3085);
nor U4822 (N_4822,N_3541,N_3655);
or U4823 (N_4823,N_3601,N_3487);
and U4824 (N_4824,N_3632,N_3506);
and U4825 (N_4825,N_3549,N_3978);
nor U4826 (N_4826,N_3841,N_3478);
nand U4827 (N_4827,N_3967,N_3283);
or U4828 (N_4828,N_3301,N_3907);
and U4829 (N_4829,N_3524,N_3619);
nand U4830 (N_4830,N_3394,N_3540);
nand U4831 (N_4831,N_3710,N_3122);
nor U4832 (N_4832,N_3178,N_3014);
or U4833 (N_4833,N_3711,N_3919);
nand U4834 (N_4834,N_3758,N_3228);
or U4835 (N_4835,N_3297,N_3640);
nor U4836 (N_4836,N_3373,N_3996);
and U4837 (N_4837,N_3377,N_3665);
and U4838 (N_4838,N_3414,N_3880);
or U4839 (N_4839,N_3773,N_3630);
nand U4840 (N_4840,N_3186,N_3806);
or U4841 (N_4841,N_3575,N_3641);
and U4842 (N_4842,N_3796,N_3760);
nand U4843 (N_4843,N_3934,N_3382);
nand U4844 (N_4844,N_3178,N_3445);
or U4845 (N_4845,N_3783,N_3387);
nand U4846 (N_4846,N_3729,N_3765);
nand U4847 (N_4847,N_3699,N_3676);
or U4848 (N_4848,N_3246,N_3308);
nand U4849 (N_4849,N_3715,N_3054);
or U4850 (N_4850,N_3086,N_3657);
and U4851 (N_4851,N_3260,N_3412);
nand U4852 (N_4852,N_3533,N_3438);
and U4853 (N_4853,N_3570,N_3228);
nor U4854 (N_4854,N_3047,N_3223);
or U4855 (N_4855,N_3319,N_3904);
and U4856 (N_4856,N_3926,N_3775);
or U4857 (N_4857,N_3246,N_3662);
and U4858 (N_4858,N_3649,N_3404);
and U4859 (N_4859,N_3789,N_3365);
nand U4860 (N_4860,N_3679,N_3104);
nand U4861 (N_4861,N_3831,N_3015);
or U4862 (N_4862,N_3691,N_3405);
or U4863 (N_4863,N_3939,N_3604);
nor U4864 (N_4864,N_3948,N_3080);
xnor U4865 (N_4865,N_3248,N_3319);
or U4866 (N_4866,N_3937,N_3071);
and U4867 (N_4867,N_3788,N_3152);
nor U4868 (N_4868,N_3740,N_3670);
and U4869 (N_4869,N_3060,N_3735);
and U4870 (N_4870,N_3693,N_3797);
nor U4871 (N_4871,N_3278,N_3488);
nor U4872 (N_4872,N_3605,N_3450);
and U4873 (N_4873,N_3002,N_3884);
nand U4874 (N_4874,N_3324,N_3545);
and U4875 (N_4875,N_3638,N_3060);
and U4876 (N_4876,N_3510,N_3906);
nand U4877 (N_4877,N_3661,N_3547);
nor U4878 (N_4878,N_3552,N_3534);
nor U4879 (N_4879,N_3989,N_3542);
and U4880 (N_4880,N_3612,N_3723);
nand U4881 (N_4881,N_3029,N_3629);
and U4882 (N_4882,N_3907,N_3218);
or U4883 (N_4883,N_3360,N_3353);
and U4884 (N_4884,N_3438,N_3017);
nor U4885 (N_4885,N_3326,N_3530);
and U4886 (N_4886,N_3761,N_3303);
xnor U4887 (N_4887,N_3111,N_3726);
nor U4888 (N_4888,N_3750,N_3379);
and U4889 (N_4889,N_3407,N_3213);
nor U4890 (N_4890,N_3707,N_3394);
nor U4891 (N_4891,N_3917,N_3979);
and U4892 (N_4892,N_3505,N_3330);
and U4893 (N_4893,N_3818,N_3331);
nor U4894 (N_4894,N_3967,N_3003);
and U4895 (N_4895,N_3805,N_3866);
and U4896 (N_4896,N_3953,N_3171);
nand U4897 (N_4897,N_3798,N_3603);
nor U4898 (N_4898,N_3731,N_3753);
xnor U4899 (N_4899,N_3184,N_3769);
or U4900 (N_4900,N_3865,N_3494);
nor U4901 (N_4901,N_3822,N_3548);
nand U4902 (N_4902,N_3076,N_3771);
nand U4903 (N_4903,N_3373,N_3464);
and U4904 (N_4904,N_3991,N_3007);
or U4905 (N_4905,N_3116,N_3351);
and U4906 (N_4906,N_3958,N_3597);
nor U4907 (N_4907,N_3037,N_3338);
nand U4908 (N_4908,N_3874,N_3240);
and U4909 (N_4909,N_3753,N_3715);
nor U4910 (N_4910,N_3996,N_3238);
and U4911 (N_4911,N_3387,N_3219);
or U4912 (N_4912,N_3370,N_3371);
nor U4913 (N_4913,N_3391,N_3710);
nand U4914 (N_4914,N_3413,N_3170);
or U4915 (N_4915,N_3402,N_3125);
nand U4916 (N_4916,N_3881,N_3210);
nand U4917 (N_4917,N_3556,N_3814);
and U4918 (N_4918,N_3896,N_3920);
nand U4919 (N_4919,N_3847,N_3672);
nor U4920 (N_4920,N_3297,N_3509);
and U4921 (N_4921,N_3876,N_3841);
nand U4922 (N_4922,N_3471,N_3680);
and U4923 (N_4923,N_3232,N_3864);
or U4924 (N_4924,N_3570,N_3387);
nor U4925 (N_4925,N_3908,N_3413);
nand U4926 (N_4926,N_3796,N_3143);
or U4927 (N_4927,N_3059,N_3051);
and U4928 (N_4928,N_3617,N_3525);
nand U4929 (N_4929,N_3754,N_3195);
and U4930 (N_4930,N_3576,N_3433);
nor U4931 (N_4931,N_3937,N_3974);
or U4932 (N_4932,N_3499,N_3067);
nand U4933 (N_4933,N_3529,N_3223);
nor U4934 (N_4934,N_3169,N_3858);
and U4935 (N_4935,N_3028,N_3011);
nand U4936 (N_4936,N_3543,N_3778);
nor U4937 (N_4937,N_3726,N_3729);
nand U4938 (N_4938,N_3656,N_3249);
nor U4939 (N_4939,N_3489,N_3383);
nand U4940 (N_4940,N_3720,N_3413);
xnor U4941 (N_4941,N_3793,N_3944);
nor U4942 (N_4942,N_3716,N_3698);
nor U4943 (N_4943,N_3719,N_3442);
nand U4944 (N_4944,N_3600,N_3856);
or U4945 (N_4945,N_3267,N_3536);
and U4946 (N_4946,N_3700,N_3880);
nand U4947 (N_4947,N_3487,N_3026);
or U4948 (N_4948,N_3882,N_3311);
or U4949 (N_4949,N_3848,N_3537);
and U4950 (N_4950,N_3822,N_3630);
and U4951 (N_4951,N_3842,N_3859);
nand U4952 (N_4952,N_3115,N_3747);
nand U4953 (N_4953,N_3272,N_3633);
or U4954 (N_4954,N_3314,N_3441);
nand U4955 (N_4955,N_3643,N_3252);
nor U4956 (N_4956,N_3453,N_3707);
nand U4957 (N_4957,N_3120,N_3083);
xor U4958 (N_4958,N_3010,N_3450);
or U4959 (N_4959,N_3442,N_3267);
nand U4960 (N_4960,N_3477,N_3842);
and U4961 (N_4961,N_3170,N_3709);
or U4962 (N_4962,N_3496,N_3684);
nand U4963 (N_4963,N_3075,N_3530);
nand U4964 (N_4964,N_3242,N_3386);
nor U4965 (N_4965,N_3811,N_3700);
or U4966 (N_4966,N_3892,N_3255);
and U4967 (N_4967,N_3067,N_3335);
and U4968 (N_4968,N_3893,N_3417);
nand U4969 (N_4969,N_3611,N_3024);
nor U4970 (N_4970,N_3297,N_3148);
or U4971 (N_4971,N_3033,N_3739);
and U4972 (N_4972,N_3360,N_3318);
nor U4973 (N_4973,N_3170,N_3951);
nor U4974 (N_4974,N_3253,N_3912);
or U4975 (N_4975,N_3053,N_3747);
or U4976 (N_4976,N_3962,N_3223);
or U4977 (N_4977,N_3972,N_3286);
or U4978 (N_4978,N_3019,N_3271);
nand U4979 (N_4979,N_3039,N_3298);
or U4980 (N_4980,N_3577,N_3568);
and U4981 (N_4981,N_3128,N_3952);
nor U4982 (N_4982,N_3176,N_3249);
nor U4983 (N_4983,N_3589,N_3509);
and U4984 (N_4984,N_3994,N_3991);
nor U4985 (N_4985,N_3034,N_3555);
or U4986 (N_4986,N_3457,N_3542);
or U4987 (N_4987,N_3942,N_3248);
nor U4988 (N_4988,N_3708,N_3611);
nand U4989 (N_4989,N_3711,N_3726);
nor U4990 (N_4990,N_3811,N_3967);
and U4991 (N_4991,N_3235,N_3909);
and U4992 (N_4992,N_3626,N_3821);
and U4993 (N_4993,N_3499,N_3595);
and U4994 (N_4994,N_3306,N_3626);
and U4995 (N_4995,N_3699,N_3169);
or U4996 (N_4996,N_3890,N_3029);
and U4997 (N_4997,N_3823,N_3020);
or U4998 (N_4998,N_3502,N_3768);
nand U4999 (N_4999,N_3006,N_3909);
and U5000 (N_5000,N_4192,N_4838);
nand U5001 (N_5001,N_4482,N_4212);
nand U5002 (N_5002,N_4275,N_4501);
and U5003 (N_5003,N_4557,N_4395);
nor U5004 (N_5004,N_4590,N_4336);
and U5005 (N_5005,N_4668,N_4868);
nor U5006 (N_5006,N_4848,N_4358);
or U5007 (N_5007,N_4393,N_4337);
or U5008 (N_5008,N_4761,N_4435);
or U5009 (N_5009,N_4574,N_4602);
nand U5010 (N_5010,N_4624,N_4439);
nor U5011 (N_5011,N_4216,N_4985);
and U5012 (N_5012,N_4186,N_4208);
or U5013 (N_5013,N_4823,N_4324);
nand U5014 (N_5014,N_4375,N_4901);
and U5015 (N_5015,N_4132,N_4203);
nor U5016 (N_5016,N_4524,N_4314);
or U5017 (N_5017,N_4717,N_4535);
nand U5018 (N_5018,N_4019,N_4799);
nor U5019 (N_5019,N_4096,N_4757);
or U5020 (N_5020,N_4503,N_4102);
nand U5021 (N_5021,N_4413,N_4093);
and U5022 (N_5022,N_4549,N_4999);
or U5023 (N_5023,N_4671,N_4774);
or U5024 (N_5024,N_4633,N_4729);
and U5025 (N_5025,N_4384,N_4014);
nor U5026 (N_5026,N_4425,N_4458);
or U5027 (N_5027,N_4230,N_4837);
or U5028 (N_5028,N_4855,N_4719);
nor U5029 (N_5029,N_4742,N_4510);
or U5030 (N_5030,N_4608,N_4890);
nor U5031 (N_5031,N_4387,N_4781);
nor U5032 (N_5032,N_4021,N_4410);
and U5033 (N_5033,N_4233,N_4052);
nand U5034 (N_5034,N_4639,N_4184);
and U5035 (N_5035,N_4533,N_4892);
and U5036 (N_5036,N_4397,N_4017);
nand U5037 (N_5037,N_4190,N_4516);
nor U5038 (N_5038,N_4552,N_4048);
nand U5039 (N_5039,N_4694,N_4264);
and U5040 (N_5040,N_4810,N_4910);
and U5041 (N_5041,N_4344,N_4955);
and U5042 (N_5042,N_4127,N_4968);
or U5043 (N_5043,N_4762,N_4972);
and U5044 (N_5044,N_4860,N_4942);
and U5045 (N_5045,N_4200,N_4281);
or U5046 (N_5046,N_4297,N_4016);
and U5047 (N_5047,N_4683,N_4941);
xnor U5048 (N_5048,N_4261,N_4670);
and U5049 (N_5049,N_4565,N_4229);
xor U5050 (N_5050,N_4666,N_4060);
and U5051 (N_5051,N_4152,N_4912);
nor U5052 (N_5052,N_4622,N_4389);
or U5053 (N_5053,N_4915,N_4926);
nand U5054 (N_5054,N_4921,N_4707);
or U5055 (N_5055,N_4328,N_4592);
and U5056 (N_5056,N_4073,N_4824);
or U5057 (N_5057,N_4778,N_4436);
or U5058 (N_5058,N_4422,N_4561);
or U5059 (N_5059,N_4087,N_4718);
or U5060 (N_5060,N_4852,N_4064);
nand U5061 (N_5061,N_4569,N_4366);
and U5062 (N_5062,N_4791,N_4356);
nand U5063 (N_5063,N_4593,N_4946);
and U5064 (N_5064,N_4245,N_4692);
or U5065 (N_5065,N_4898,N_4759);
or U5066 (N_5066,N_4933,N_4071);
and U5067 (N_5067,N_4571,N_4169);
and U5068 (N_5068,N_4417,N_4431);
and U5069 (N_5069,N_4513,N_4251);
nor U5070 (N_5070,N_4749,N_4051);
nand U5071 (N_5071,N_4079,N_4721);
and U5072 (N_5072,N_4638,N_4495);
nor U5073 (N_5073,N_4564,N_4256);
nand U5074 (N_5074,N_4101,N_4609);
nand U5075 (N_5075,N_4173,N_4641);
nor U5076 (N_5076,N_4025,N_4411);
nor U5077 (N_5077,N_4630,N_4441);
nor U5078 (N_5078,N_4235,N_4359);
nand U5079 (N_5079,N_4874,N_4620);
and U5080 (N_5080,N_4760,N_4685);
nand U5081 (N_5081,N_4548,N_4714);
nor U5082 (N_5082,N_4003,N_4164);
and U5083 (N_5083,N_4489,N_4792);
and U5084 (N_5084,N_4734,N_4930);
nor U5085 (N_5085,N_4637,N_4134);
nor U5086 (N_5086,N_4790,N_4427);
nand U5087 (N_5087,N_4372,N_4407);
or U5088 (N_5088,N_4330,N_4944);
nor U5089 (N_5089,N_4811,N_4089);
or U5090 (N_5090,N_4857,N_4065);
or U5091 (N_5091,N_4405,N_4464);
nor U5092 (N_5092,N_4131,N_4211);
and U5093 (N_5093,N_4383,N_4900);
or U5094 (N_5094,N_4300,N_4704);
nand U5095 (N_5095,N_4376,N_4711);
nor U5096 (N_5096,N_4394,N_4047);
or U5097 (N_5097,N_4399,N_4904);
or U5098 (N_5098,N_4023,N_4554);
nand U5099 (N_5099,N_4306,N_4728);
or U5100 (N_5100,N_4409,N_4515);
or U5101 (N_5101,N_4743,N_4614);
nand U5102 (N_5102,N_4716,N_4696);
or U5103 (N_5103,N_4882,N_4911);
and U5104 (N_5104,N_4176,N_4750);
nand U5105 (N_5105,N_4850,N_4339);
xnor U5106 (N_5106,N_4978,N_4856);
or U5107 (N_5107,N_4688,N_4830);
nor U5108 (N_5108,N_4794,N_4136);
nand U5109 (N_5109,N_4701,N_4672);
and U5110 (N_5110,N_4543,N_4568);
or U5111 (N_5111,N_4445,N_4053);
or U5112 (N_5112,N_4806,N_4475);
and U5113 (N_5113,N_4899,N_4844);
and U5114 (N_5114,N_4954,N_4936);
and U5115 (N_5115,N_4018,N_4326);
nor U5116 (N_5116,N_4284,N_4305);
nand U5117 (N_5117,N_4545,N_4125);
or U5118 (N_5118,N_4962,N_4459);
nand U5119 (N_5119,N_4538,N_4576);
and U5120 (N_5120,N_4536,N_4527);
and U5121 (N_5121,N_4897,N_4272);
and U5122 (N_5122,N_4476,N_4656);
or U5123 (N_5123,N_4865,N_4138);
nor U5124 (N_5124,N_4010,N_4128);
nand U5125 (N_5125,N_4710,N_4075);
and U5126 (N_5126,N_4600,N_4834);
or U5127 (N_5127,N_4595,N_4509);
nor U5128 (N_5128,N_4634,N_4908);
and U5129 (N_5129,N_4000,N_4274);
nor U5130 (N_5130,N_4814,N_4673);
nand U5131 (N_5131,N_4323,N_4241);
or U5132 (N_5132,N_4345,N_4078);
or U5133 (N_5133,N_4380,N_4960);
nand U5134 (N_5134,N_4088,N_4555);
nor U5135 (N_5135,N_4661,N_4290);
and U5136 (N_5136,N_4286,N_4130);
or U5137 (N_5137,N_4821,N_4097);
nor U5138 (N_5138,N_4460,N_4179);
and U5139 (N_5139,N_4041,N_4686);
or U5140 (N_5140,N_4948,N_4334);
and U5141 (N_5141,N_4950,N_4866);
nor U5142 (N_5142,N_4709,N_4123);
nor U5143 (N_5143,N_4304,N_4497);
or U5144 (N_5144,N_4829,N_4582);
nand U5145 (N_5145,N_4373,N_4815);
nand U5146 (N_5146,N_4362,N_4107);
nand U5147 (N_5147,N_4193,N_4804);
nor U5148 (N_5148,N_4544,N_4008);
and U5149 (N_5149,N_4808,N_4349);
or U5150 (N_5150,N_4428,N_4414);
nand U5151 (N_5151,N_4061,N_4687);
nand U5152 (N_5152,N_4020,N_4378);
nor U5153 (N_5153,N_4415,N_4802);
nand U5154 (N_5154,N_4207,N_4454);
and U5155 (N_5155,N_4753,N_4421);
nand U5156 (N_5156,N_4880,N_4221);
nand U5157 (N_5157,N_4492,N_4888);
or U5158 (N_5158,N_4733,N_4213);
nor U5159 (N_5159,N_4452,N_4963);
or U5160 (N_5160,N_4652,N_4189);
nand U5161 (N_5161,N_4843,N_4177);
and U5162 (N_5162,N_4283,N_4572);
nand U5163 (N_5163,N_4045,N_4801);
nand U5164 (N_5164,N_4063,N_4196);
nand U5165 (N_5165,N_4905,N_4773);
and U5166 (N_5166,N_4679,N_4684);
or U5167 (N_5167,N_4234,N_4562);
or U5168 (N_5168,N_4606,N_4118);
or U5169 (N_5169,N_4805,N_4462);
or U5170 (N_5170,N_4917,N_4981);
nand U5171 (N_5171,N_4271,N_4161);
nor U5172 (N_5172,N_4891,N_4315);
nor U5173 (N_5173,N_4222,N_4440);
nand U5174 (N_5174,N_4114,N_4491);
nor U5175 (N_5175,N_4085,N_4004);
or U5176 (N_5176,N_4741,N_4346);
and U5177 (N_5177,N_4626,N_4259);
nor U5178 (N_5178,N_4043,N_4112);
or U5179 (N_5179,N_4282,N_4156);
nor U5180 (N_5180,N_4227,N_4586);
or U5181 (N_5181,N_4158,N_4969);
nor U5182 (N_5182,N_4708,N_4443);
or U5183 (N_5183,N_4232,N_4833);
or U5184 (N_5184,N_4612,N_4160);
or U5185 (N_5185,N_4007,N_4472);
or U5186 (N_5186,N_4166,N_4976);
nor U5187 (N_5187,N_4444,N_4325);
and U5188 (N_5188,N_4034,N_4520);
nor U5189 (N_5189,N_4991,N_4214);
nand U5190 (N_5190,N_4285,N_4889);
or U5191 (N_5191,N_4257,N_4418);
nand U5192 (N_5192,N_4858,N_4191);
nand U5193 (N_5193,N_4647,N_4426);
nand U5194 (N_5194,N_4803,N_4605);
and U5195 (N_5195,N_4374,N_4363);
nand U5196 (N_5196,N_4697,N_4455);
nand U5197 (N_5197,N_4722,N_4157);
or U5198 (N_5198,N_4594,N_4862);
and U5199 (N_5199,N_4506,N_4108);
nor U5200 (N_5200,N_4507,N_4525);
or U5201 (N_5201,N_4360,N_4481);
and U5202 (N_5202,N_4278,N_4066);
or U5203 (N_5203,N_4247,N_4086);
or U5204 (N_5204,N_4110,N_4840);
nor U5205 (N_5205,N_4649,N_4474);
nand U5206 (N_5206,N_4989,N_4252);
or U5207 (N_5207,N_4117,N_4797);
and U5208 (N_5208,N_4578,N_4416);
nand U5209 (N_5209,N_4433,N_4607);
or U5210 (N_5210,N_4279,N_4404);
nand U5211 (N_5211,N_4547,N_4224);
nor U5212 (N_5212,N_4062,N_4635);
nand U5213 (N_5213,N_4785,N_4570);
nor U5214 (N_5214,N_4896,N_4269);
nor U5215 (N_5215,N_4437,N_4154);
or U5216 (N_5216,N_4277,N_4250);
xor U5217 (N_5217,N_4703,N_4738);
nand U5218 (N_5218,N_4825,N_4292);
nor U5219 (N_5219,N_4456,N_4260);
xor U5220 (N_5220,N_4386,N_4432);
nor U5221 (N_5221,N_4243,N_4116);
or U5222 (N_5222,N_4313,N_4654);
nand U5223 (N_5223,N_4690,N_4477);
or U5224 (N_5224,N_4957,N_4522);
nand U5225 (N_5225,N_4723,N_4341);
or U5226 (N_5226,N_4922,N_4529);
nor U5227 (N_5227,N_4457,N_4309);
and U5228 (N_5228,N_4450,N_4057);
nand U5229 (N_5229,N_4970,N_4975);
nor U5230 (N_5230,N_4747,N_4756);
nor U5231 (N_5231,N_4831,N_4371);
and U5232 (N_5232,N_4669,N_4887);
or U5233 (N_5233,N_4597,N_4903);
or U5234 (N_5234,N_4228,N_4782);
nand U5235 (N_5235,N_4849,N_4388);
and U5236 (N_5236,N_4493,N_4551);
or U5237 (N_5237,N_4348,N_4682);
and U5238 (N_5238,N_4170,N_4141);
nand U5239 (N_5239,N_4965,N_4643);
and U5240 (N_5240,N_4220,N_4906);
or U5241 (N_5241,N_4142,N_4751);
nor U5242 (N_5242,N_4406,N_4488);
or U5243 (N_5243,N_4937,N_4009);
and U5244 (N_5244,N_4081,N_4657);
nor U5245 (N_5245,N_4333,N_4712);
nand U5246 (N_5246,N_4699,N_4943);
nor U5247 (N_5247,N_4006,N_4604);
and U5248 (N_5248,N_4319,N_4391);
nor U5249 (N_5249,N_4320,N_4530);
nand U5250 (N_5250,N_4775,N_4736);
or U5251 (N_5251,N_4822,N_4812);
or U5252 (N_5252,N_4788,N_4990);
nand U5253 (N_5253,N_4466,N_4240);
and U5254 (N_5254,N_4449,N_4178);
nand U5255 (N_5255,N_4998,N_4013);
or U5256 (N_5256,N_4869,N_4321);
nand U5257 (N_5257,N_4180,N_4451);
nor U5258 (N_5258,N_4223,N_4039);
nand U5259 (N_5259,N_4162,N_4758);
nand U5260 (N_5260,N_4650,N_4980);
nor U5261 (N_5261,N_4959,N_4129);
and U5262 (N_5262,N_4542,N_4206);
and U5263 (N_5263,N_4469,N_4769);
and U5264 (N_5264,N_4603,N_4423);
or U5265 (N_5265,N_4238,N_4343);
nor U5266 (N_5266,N_4977,N_4149);
and U5267 (N_5267,N_4667,N_4816);
or U5268 (N_5268,N_4902,N_4379);
or U5269 (N_5269,N_4645,N_4453);
nor U5270 (N_5270,N_4988,N_4702);
nor U5271 (N_5271,N_4070,N_4541);
xnor U5272 (N_5272,N_4106,N_4266);
and U5273 (N_5273,N_4771,N_4776);
nand U5274 (N_5274,N_4148,N_4745);
and U5275 (N_5275,N_4573,N_4658);
or U5276 (N_5276,N_4448,N_4677);
nand U5277 (N_5277,N_4155,N_4528);
and U5278 (N_5278,N_4273,N_4642);
and U5279 (N_5279,N_4183,N_4767);
nor U5280 (N_5280,N_4119,N_4952);
xnor U5281 (N_5281,N_4144,N_4310);
nand U5282 (N_5282,N_4828,N_4953);
and U5283 (N_5283,N_4011,N_4361);
and U5284 (N_5284,N_4648,N_4210);
or U5285 (N_5285,N_4610,N_4322);
or U5286 (N_5286,N_4982,N_4150);
nand U5287 (N_5287,N_4966,N_4122);
xor U5288 (N_5288,N_4487,N_4581);
nor U5289 (N_5289,N_4770,N_4293);
or U5290 (N_5290,N_4651,N_4298);
and U5291 (N_5291,N_4611,N_4698);
nor U5292 (N_5292,N_4486,N_4974);
and U5293 (N_5293,N_4591,N_4598);
or U5294 (N_5294,N_4146,N_4546);
or U5295 (N_5295,N_4997,N_4032);
nor U5296 (N_5296,N_4059,N_4517);
nor U5297 (N_5297,N_4498,N_4438);
and U5298 (N_5298,N_4468,N_4248);
nand U5299 (N_5299,N_4201,N_4935);
or U5300 (N_5300,N_4700,N_4430);
nand U5301 (N_5301,N_4764,N_4042);
nand U5302 (N_5302,N_4172,N_4907);
nor U5303 (N_5303,N_4140,N_4861);
nand U5304 (N_5304,N_4022,N_4137);
nand U5305 (N_5305,N_4332,N_4680);
and U5306 (N_5306,N_4766,N_4030);
or U5307 (N_5307,N_4185,N_4931);
or U5308 (N_5308,N_4015,N_4135);
or U5309 (N_5309,N_4473,N_4928);
and U5310 (N_5310,N_4705,N_4884);
nand U5311 (N_5311,N_4396,N_4217);
nor U5312 (N_5312,N_4925,N_4263);
nor U5313 (N_5313,N_4398,N_4923);
nand U5314 (N_5314,N_4002,N_4082);
xnor U5315 (N_5315,N_4105,N_4353);
nand U5316 (N_5316,N_4402,N_4827);
and U5317 (N_5317,N_4244,N_4873);
nand U5318 (N_5318,N_4636,N_4553);
or U5319 (N_5319,N_4947,N_4851);
and U5320 (N_5320,N_4613,N_4099);
and U5321 (N_5321,N_4480,N_4909);
and U5322 (N_5322,N_4335,N_4817);
or U5323 (N_5323,N_4746,N_4199);
or U5324 (N_5324,N_4956,N_4986);
nor U5325 (N_5325,N_4979,N_4385);
nand U5326 (N_5326,N_4104,N_4893);
or U5327 (N_5327,N_4895,N_4663);
or U5328 (N_5328,N_4329,N_4069);
or U5329 (N_5329,N_4567,N_4854);
or U5330 (N_5330,N_4268,N_4054);
and U5331 (N_5331,N_4331,N_4713);
nand U5332 (N_5332,N_4442,N_4876);
nor U5333 (N_5333,N_4674,N_4072);
and U5334 (N_5334,N_4539,N_4288);
and U5335 (N_5335,N_4165,N_4505);
nand U5336 (N_5336,N_4617,N_4067);
nor U5337 (N_5337,N_4735,N_4001);
and U5338 (N_5338,N_4342,N_4845);
nor U5339 (N_5339,N_4504,N_4074);
and U5340 (N_5340,N_4198,N_4951);
nand U5341 (N_5341,N_4035,N_4847);
nand U5342 (N_5342,N_4878,N_4737);
or U5343 (N_5343,N_4945,N_4618);
or U5344 (N_5344,N_4644,N_4560);
nand U5345 (N_5345,N_4147,N_4126);
nor U5346 (N_5346,N_4133,N_4381);
or U5347 (N_5347,N_4752,N_4471);
and U5348 (N_5348,N_4163,N_4296);
and U5349 (N_5349,N_4579,N_4226);
nor U5350 (N_5350,N_4689,N_4971);
or U5351 (N_5351,N_4789,N_4357);
and U5352 (N_5352,N_4625,N_4258);
and U5353 (N_5353,N_4090,N_4446);
nand U5354 (N_5354,N_4168,N_4660);
and U5355 (N_5355,N_4365,N_4276);
or U5356 (N_5356,N_4103,N_4655);
xnor U5357 (N_5357,N_4139,N_4691);
or U5358 (N_5358,N_4094,N_4676);
nor U5359 (N_5359,N_4559,N_4080);
nor U5360 (N_5360,N_4351,N_4370);
and U5361 (N_5361,N_4631,N_4294);
and U5362 (N_5362,N_4403,N_4031);
nand U5363 (N_5363,N_4932,N_4632);
and U5364 (N_5364,N_4367,N_4540);
and U5365 (N_5365,N_4076,N_4870);
nand U5366 (N_5366,N_4352,N_4779);
nor U5367 (N_5367,N_4091,N_4744);
or U5368 (N_5368,N_4115,N_4312);
and U5369 (N_5369,N_4280,N_4470);
xnor U5370 (N_5370,N_4532,N_4665);
nand U5371 (N_5371,N_4871,N_4036);
nand U5372 (N_5372,N_4739,N_4826);
xor U5373 (N_5373,N_4024,N_4596);
nand U5374 (N_5374,N_4188,N_4846);
nor U5375 (N_5375,N_4585,N_4005);
and U5376 (N_5376,N_4627,N_4502);
nand U5377 (N_5377,N_4724,N_4434);
nor U5378 (N_5378,N_4589,N_4143);
nand U5379 (N_5379,N_4863,N_4040);
or U5380 (N_5380,N_4958,N_4120);
or U5381 (N_5381,N_4084,N_4623);
nor U5382 (N_5382,N_4732,N_4886);
or U5383 (N_5383,N_4029,N_4796);
nand U5384 (N_5384,N_4317,N_4167);
nand U5385 (N_5385,N_4995,N_4299);
and U5386 (N_5386,N_4187,N_4237);
nor U5387 (N_5387,N_4026,N_4795);
nor U5388 (N_5388,N_4316,N_4046);
and U5389 (N_5389,N_4174,N_4270);
nor U5390 (N_5390,N_4056,N_4973);
nor U5391 (N_5391,N_4994,N_4558);
and U5392 (N_5392,N_4731,N_4772);
nor U5393 (N_5393,N_4408,N_4302);
or U5394 (N_5394,N_4483,N_4249);
or U5395 (N_5395,N_4727,N_4835);
nor U5396 (N_5396,N_4621,N_4253);
or U5397 (N_5397,N_4798,N_4355);
nand U5398 (N_5398,N_4748,N_4028);
nand U5399 (N_5399,N_4267,N_4151);
nand U5400 (N_5400,N_4100,N_4659);
nor U5401 (N_5401,N_4725,N_4095);
or U5402 (N_5402,N_4204,N_4307);
and U5403 (N_5403,N_4098,N_4914);
or U5404 (N_5404,N_4526,N_4254);
or U5405 (N_5405,N_4996,N_4836);
nand U5406 (N_5406,N_4420,N_4777);
and U5407 (N_5407,N_4083,N_4494);
and U5408 (N_5408,N_4784,N_4246);
or U5409 (N_5409,N_4153,N_4340);
and U5410 (N_5410,N_4308,N_4881);
nor U5411 (N_5411,N_4949,N_4938);
or U5412 (N_5412,N_4490,N_4171);
or U5413 (N_5413,N_4992,N_4720);
nor U5414 (N_5414,N_4050,N_4311);
nor U5415 (N_5415,N_4629,N_4390);
nor U5416 (N_5416,N_4077,N_4755);
or U5417 (N_5417,N_4033,N_4514);
or U5418 (N_5418,N_4049,N_4807);
and U5419 (N_5419,N_4215,N_4419);
nor U5420 (N_5420,N_4412,N_4392);
or U5421 (N_5421,N_4820,N_4236);
nand U5422 (N_5422,N_4231,N_4940);
nor U5423 (N_5423,N_4500,N_4809);
or U5424 (N_5424,N_4800,N_4841);
and U5425 (N_5425,N_4653,N_4984);
nor U5426 (N_5426,N_4550,N_4175);
nand U5427 (N_5427,N_4429,N_4287);
and U5428 (N_5428,N_4463,N_4038);
and U5429 (N_5429,N_4338,N_4853);
and U5430 (N_5430,N_4145,N_4793);
xor U5431 (N_5431,N_4675,N_4424);
and U5432 (N_5432,N_4646,N_4864);
and U5433 (N_5433,N_4218,N_4584);
or U5434 (N_5434,N_4839,N_4382);
nand U5435 (N_5435,N_4113,N_4111);
nand U5436 (N_5436,N_4364,N_4347);
or U5437 (N_5437,N_4983,N_4918);
nand U5438 (N_5438,N_4109,N_4012);
nor U5439 (N_5439,N_4939,N_4588);
and U5440 (N_5440,N_4523,N_4681);
and U5441 (N_5441,N_4879,N_4695);
nand U5442 (N_5442,N_4662,N_4478);
nand U5443 (N_5443,N_4883,N_4255);
nor U5444 (N_5444,N_4465,N_4508);
and U5445 (N_5445,N_4401,N_4730);
nor U5446 (N_5446,N_4819,N_4616);
nor U5447 (N_5447,N_4842,N_4859);
nor U5448 (N_5448,N_4205,N_4563);
and U5449 (N_5449,N_4182,N_4885);
and U5450 (N_5450,N_4239,N_4499);
nor U5451 (N_5451,N_4219,N_4531);
and U5452 (N_5452,N_4587,N_4262);
nor U5453 (N_5453,N_4194,N_4664);
xnor U5454 (N_5454,N_4044,N_4303);
or U5455 (N_5455,N_4534,N_4875);
or U5456 (N_5456,N_4181,N_4818);
nor U5457 (N_5457,N_4461,N_4058);
or U5458 (N_5458,N_4092,N_4615);
nor U5459 (N_5459,N_4877,N_4159);
and U5460 (N_5460,N_4027,N_4715);
nor U5461 (N_5461,N_4195,N_4291);
nand U5462 (N_5462,N_4872,N_4518);
nor U5463 (N_5463,N_4927,N_4961);
and U5464 (N_5464,N_4786,N_4678);
and U5465 (N_5465,N_4354,N_4566);
nand U5466 (N_5466,N_4295,N_4783);
nor U5467 (N_5467,N_4916,N_4377);
and U5468 (N_5468,N_4934,N_4068);
nand U5469 (N_5469,N_4121,N_4467);
nor U5470 (N_5470,N_4301,N_4209);
nor U5471 (N_5471,N_4599,N_4740);
or U5472 (N_5472,N_4583,N_4037);
or U5473 (N_5473,N_4512,N_4318);
nand U5474 (N_5474,N_4628,N_4787);
nor U5475 (N_5475,N_4619,N_4580);
and U5476 (N_5476,N_4265,N_4726);
or U5477 (N_5477,N_4919,N_4400);
nand U5478 (N_5478,N_4369,N_4496);
or U5479 (N_5479,N_4350,N_4055);
or U5480 (N_5480,N_4521,N_4754);
nand U5481 (N_5481,N_4556,N_4601);
nor U5482 (N_5482,N_4484,N_4894);
nand U5483 (N_5483,N_4706,N_4327);
and U5484 (N_5484,N_4813,N_4537);
nand U5485 (N_5485,N_4640,N_4832);
or U5486 (N_5486,N_4967,N_4242);
nor U5487 (N_5487,N_4289,N_4867);
nand U5488 (N_5488,N_4763,N_4964);
nand U5489 (N_5489,N_4913,N_4225);
and U5490 (N_5490,N_4768,N_4987);
nor U5491 (N_5491,N_4197,N_4575);
nand U5492 (N_5492,N_4693,N_4765);
nand U5493 (N_5493,N_4124,N_4368);
nor U5494 (N_5494,N_4511,N_4202);
and U5495 (N_5495,N_4447,N_4993);
and U5496 (N_5496,N_4780,N_4920);
and U5497 (N_5497,N_4929,N_4485);
nand U5498 (N_5498,N_4479,N_4519);
or U5499 (N_5499,N_4577,N_4924);
and U5500 (N_5500,N_4157,N_4220);
nand U5501 (N_5501,N_4499,N_4684);
and U5502 (N_5502,N_4218,N_4574);
nor U5503 (N_5503,N_4525,N_4072);
or U5504 (N_5504,N_4947,N_4113);
or U5505 (N_5505,N_4839,N_4573);
nand U5506 (N_5506,N_4318,N_4906);
nand U5507 (N_5507,N_4926,N_4596);
nand U5508 (N_5508,N_4290,N_4014);
or U5509 (N_5509,N_4770,N_4732);
nor U5510 (N_5510,N_4317,N_4354);
or U5511 (N_5511,N_4330,N_4569);
nand U5512 (N_5512,N_4111,N_4126);
nor U5513 (N_5513,N_4553,N_4743);
or U5514 (N_5514,N_4092,N_4567);
or U5515 (N_5515,N_4710,N_4476);
nor U5516 (N_5516,N_4967,N_4871);
nor U5517 (N_5517,N_4540,N_4115);
and U5518 (N_5518,N_4923,N_4445);
and U5519 (N_5519,N_4313,N_4418);
nand U5520 (N_5520,N_4697,N_4579);
or U5521 (N_5521,N_4854,N_4164);
nand U5522 (N_5522,N_4280,N_4981);
nor U5523 (N_5523,N_4983,N_4598);
or U5524 (N_5524,N_4932,N_4199);
nand U5525 (N_5525,N_4958,N_4069);
and U5526 (N_5526,N_4278,N_4161);
nand U5527 (N_5527,N_4650,N_4552);
nand U5528 (N_5528,N_4295,N_4822);
and U5529 (N_5529,N_4491,N_4962);
and U5530 (N_5530,N_4078,N_4756);
nor U5531 (N_5531,N_4541,N_4815);
or U5532 (N_5532,N_4261,N_4799);
xor U5533 (N_5533,N_4229,N_4477);
or U5534 (N_5534,N_4560,N_4539);
nor U5535 (N_5535,N_4235,N_4953);
or U5536 (N_5536,N_4317,N_4707);
and U5537 (N_5537,N_4467,N_4577);
nor U5538 (N_5538,N_4543,N_4757);
nor U5539 (N_5539,N_4983,N_4022);
or U5540 (N_5540,N_4353,N_4571);
and U5541 (N_5541,N_4698,N_4574);
nor U5542 (N_5542,N_4794,N_4793);
nand U5543 (N_5543,N_4242,N_4623);
or U5544 (N_5544,N_4527,N_4011);
or U5545 (N_5545,N_4632,N_4063);
or U5546 (N_5546,N_4702,N_4422);
nand U5547 (N_5547,N_4109,N_4928);
and U5548 (N_5548,N_4923,N_4391);
and U5549 (N_5549,N_4437,N_4747);
and U5550 (N_5550,N_4699,N_4127);
nand U5551 (N_5551,N_4021,N_4303);
and U5552 (N_5552,N_4327,N_4540);
nor U5553 (N_5553,N_4871,N_4161);
xor U5554 (N_5554,N_4309,N_4813);
nor U5555 (N_5555,N_4619,N_4284);
nand U5556 (N_5556,N_4489,N_4177);
nand U5557 (N_5557,N_4068,N_4879);
and U5558 (N_5558,N_4830,N_4443);
nand U5559 (N_5559,N_4089,N_4341);
nand U5560 (N_5560,N_4922,N_4366);
or U5561 (N_5561,N_4477,N_4990);
or U5562 (N_5562,N_4682,N_4245);
nor U5563 (N_5563,N_4889,N_4934);
or U5564 (N_5564,N_4409,N_4737);
and U5565 (N_5565,N_4404,N_4176);
nand U5566 (N_5566,N_4647,N_4165);
and U5567 (N_5567,N_4938,N_4144);
and U5568 (N_5568,N_4523,N_4691);
nor U5569 (N_5569,N_4109,N_4241);
or U5570 (N_5570,N_4244,N_4022);
and U5571 (N_5571,N_4383,N_4439);
and U5572 (N_5572,N_4858,N_4088);
nand U5573 (N_5573,N_4839,N_4212);
and U5574 (N_5574,N_4874,N_4033);
and U5575 (N_5575,N_4105,N_4058);
nor U5576 (N_5576,N_4663,N_4799);
nand U5577 (N_5577,N_4657,N_4028);
nand U5578 (N_5578,N_4772,N_4086);
nand U5579 (N_5579,N_4743,N_4719);
and U5580 (N_5580,N_4149,N_4899);
or U5581 (N_5581,N_4894,N_4275);
or U5582 (N_5582,N_4884,N_4596);
and U5583 (N_5583,N_4018,N_4363);
or U5584 (N_5584,N_4691,N_4562);
nand U5585 (N_5585,N_4011,N_4229);
and U5586 (N_5586,N_4884,N_4433);
xnor U5587 (N_5587,N_4328,N_4695);
and U5588 (N_5588,N_4162,N_4324);
nand U5589 (N_5589,N_4161,N_4078);
and U5590 (N_5590,N_4722,N_4518);
or U5591 (N_5591,N_4510,N_4206);
and U5592 (N_5592,N_4175,N_4874);
nor U5593 (N_5593,N_4035,N_4755);
nor U5594 (N_5594,N_4667,N_4121);
or U5595 (N_5595,N_4442,N_4170);
or U5596 (N_5596,N_4765,N_4964);
and U5597 (N_5597,N_4117,N_4684);
nor U5598 (N_5598,N_4842,N_4836);
nor U5599 (N_5599,N_4220,N_4874);
and U5600 (N_5600,N_4337,N_4934);
or U5601 (N_5601,N_4377,N_4570);
nor U5602 (N_5602,N_4881,N_4995);
or U5603 (N_5603,N_4089,N_4006);
nor U5604 (N_5604,N_4556,N_4664);
nand U5605 (N_5605,N_4689,N_4968);
and U5606 (N_5606,N_4864,N_4687);
nor U5607 (N_5607,N_4542,N_4955);
nand U5608 (N_5608,N_4414,N_4769);
or U5609 (N_5609,N_4364,N_4384);
or U5610 (N_5610,N_4078,N_4483);
and U5611 (N_5611,N_4128,N_4415);
and U5612 (N_5612,N_4343,N_4015);
nand U5613 (N_5613,N_4321,N_4134);
and U5614 (N_5614,N_4039,N_4344);
or U5615 (N_5615,N_4209,N_4923);
nand U5616 (N_5616,N_4236,N_4758);
nand U5617 (N_5617,N_4472,N_4454);
or U5618 (N_5618,N_4025,N_4079);
nand U5619 (N_5619,N_4917,N_4234);
and U5620 (N_5620,N_4542,N_4815);
or U5621 (N_5621,N_4242,N_4688);
nand U5622 (N_5622,N_4618,N_4233);
nand U5623 (N_5623,N_4644,N_4866);
and U5624 (N_5624,N_4839,N_4300);
or U5625 (N_5625,N_4366,N_4706);
or U5626 (N_5626,N_4164,N_4381);
and U5627 (N_5627,N_4531,N_4917);
nor U5628 (N_5628,N_4449,N_4707);
nand U5629 (N_5629,N_4841,N_4596);
and U5630 (N_5630,N_4293,N_4851);
and U5631 (N_5631,N_4974,N_4903);
nor U5632 (N_5632,N_4393,N_4999);
and U5633 (N_5633,N_4841,N_4243);
or U5634 (N_5634,N_4651,N_4542);
or U5635 (N_5635,N_4605,N_4298);
and U5636 (N_5636,N_4521,N_4562);
nand U5637 (N_5637,N_4326,N_4826);
nor U5638 (N_5638,N_4930,N_4631);
or U5639 (N_5639,N_4568,N_4826);
nand U5640 (N_5640,N_4851,N_4506);
nor U5641 (N_5641,N_4380,N_4464);
or U5642 (N_5642,N_4678,N_4975);
and U5643 (N_5643,N_4698,N_4822);
or U5644 (N_5644,N_4189,N_4882);
and U5645 (N_5645,N_4502,N_4724);
and U5646 (N_5646,N_4035,N_4711);
nor U5647 (N_5647,N_4214,N_4976);
and U5648 (N_5648,N_4937,N_4076);
nand U5649 (N_5649,N_4979,N_4478);
nand U5650 (N_5650,N_4410,N_4941);
or U5651 (N_5651,N_4240,N_4781);
nand U5652 (N_5652,N_4881,N_4169);
and U5653 (N_5653,N_4288,N_4876);
and U5654 (N_5654,N_4318,N_4120);
or U5655 (N_5655,N_4805,N_4770);
and U5656 (N_5656,N_4232,N_4891);
or U5657 (N_5657,N_4029,N_4113);
nor U5658 (N_5658,N_4483,N_4114);
nor U5659 (N_5659,N_4541,N_4214);
nor U5660 (N_5660,N_4268,N_4406);
and U5661 (N_5661,N_4918,N_4296);
nor U5662 (N_5662,N_4145,N_4925);
and U5663 (N_5663,N_4696,N_4954);
nor U5664 (N_5664,N_4377,N_4198);
or U5665 (N_5665,N_4775,N_4007);
nand U5666 (N_5666,N_4781,N_4748);
nand U5667 (N_5667,N_4266,N_4912);
nor U5668 (N_5668,N_4633,N_4710);
nor U5669 (N_5669,N_4019,N_4043);
and U5670 (N_5670,N_4302,N_4007);
nand U5671 (N_5671,N_4253,N_4481);
nand U5672 (N_5672,N_4157,N_4790);
nor U5673 (N_5673,N_4180,N_4574);
nor U5674 (N_5674,N_4485,N_4648);
or U5675 (N_5675,N_4569,N_4794);
nand U5676 (N_5676,N_4844,N_4656);
nand U5677 (N_5677,N_4795,N_4627);
and U5678 (N_5678,N_4741,N_4798);
nor U5679 (N_5679,N_4409,N_4796);
nand U5680 (N_5680,N_4151,N_4686);
and U5681 (N_5681,N_4619,N_4212);
or U5682 (N_5682,N_4692,N_4893);
and U5683 (N_5683,N_4770,N_4580);
nor U5684 (N_5684,N_4693,N_4929);
or U5685 (N_5685,N_4554,N_4557);
nor U5686 (N_5686,N_4548,N_4336);
or U5687 (N_5687,N_4932,N_4960);
or U5688 (N_5688,N_4235,N_4002);
nand U5689 (N_5689,N_4213,N_4770);
nor U5690 (N_5690,N_4536,N_4058);
nor U5691 (N_5691,N_4533,N_4240);
nor U5692 (N_5692,N_4440,N_4523);
nor U5693 (N_5693,N_4701,N_4197);
or U5694 (N_5694,N_4028,N_4241);
and U5695 (N_5695,N_4156,N_4947);
nor U5696 (N_5696,N_4767,N_4740);
or U5697 (N_5697,N_4351,N_4131);
nor U5698 (N_5698,N_4458,N_4172);
nor U5699 (N_5699,N_4247,N_4273);
nor U5700 (N_5700,N_4447,N_4180);
and U5701 (N_5701,N_4672,N_4236);
or U5702 (N_5702,N_4827,N_4369);
and U5703 (N_5703,N_4427,N_4103);
nor U5704 (N_5704,N_4637,N_4710);
and U5705 (N_5705,N_4071,N_4301);
and U5706 (N_5706,N_4113,N_4202);
and U5707 (N_5707,N_4534,N_4052);
nor U5708 (N_5708,N_4174,N_4874);
nand U5709 (N_5709,N_4650,N_4690);
or U5710 (N_5710,N_4339,N_4245);
nor U5711 (N_5711,N_4256,N_4175);
or U5712 (N_5712,N_4617,N_4112);
or U5713 (N_5713,N_4113,N_4888);
or U5714 (N_5714,N_4987,N_4609);
nand U5715 (N_5715,N_4423,N_4599);
nor U5716 (N_5716,N_4711,N_4263);
nand U5717 (N_5717,N_4745,N_4582);
nand U5718 (N_5718,N_4015,N_4120);
nor U5719 (N_5719,N_4904,N_4322);
nor U5720 (N_5720,N_4280,N_4333);
xnor U5721 (N_5721,N_4104,N_4054);
nor U5722 (N_5722,N_4734,N_4736);
nor U5723 (N_5723,N_4577,N_4785);
nor U5724 (N_5724,N_4657,N_4178);
nand U5725 (N_5725,N_4899,N_4425);
nor U5726 (N_5726,N_4816,N_4290);
and U5727 (N_5727,N_4295,N_4776);
nand U5728 (N_5728,N_4155,N_4612);
nor U5729 (N_5729,N_4463,N_4325);
nor U5730 (N_5730,N_4460,N_4165);
xor U5731 (N_5731,N_4412,N_4075);
nor U5732 (N_5732,N_4928,N_4309);
nor U5733 (N_5733,N_4209,N_4362);
nor U5734 (N_5734,N_4785,N_4083);
and U5735 (N_5735,N_4575,N_4110);
nand U5736 (N_5736,N_4718,N_4991);
or U5737 (N_5737,N_4551,N_4824);
or U5738 (N_5738,N_4412,N_4167);
nand U5739 (N_5739,N_4053,N_4167);
and U5740 (N_5740,N_4327,N_4610);
nor U5741 (N_5741,N_4384,N_4374);
nand U5742 (N_5742,N_4857,N_4332);
nor U5743 (N_5743,N_4727,N_4618);
nand U5744 (N_5744,N_4226,N_4496);
nand U5745 (N_5745,N_4451,N_4852);
nand U5746 (N_5746,N_4469,N_4868);
or U5747 (N_5747,N_4649,N_4553);
xor U5748 (N_5748,N_4705,N_4350);
or U5749 (N_5749,N_4671,N_4698);
or U5750 (N_5750,N_4232,N_4861);
nand U5751 (N_5751,N_4520,N_4636);
nor U5752 (N_5752,N_4664,N_4935);
nor U5753 (N_5753,N_4340,N_4070);
nand U5754 (N_5754,N_4088,N_4112);
nor U5755 (N_5755,N_4230,N_4854);
nor U5756 (N_5756,N_4450,N_4244);
nand U5757 (N_5757,N_4592,N_4794);
nor U5758 (N_5758,N_4542,N_4809);
xor U5759 (N_5759,N_4084,N_4262);
nand U5760 (N_5760,N_4722,N_4929);
and U5761 (N_5761,N_4694,N_4760);
nor U5762 (N_5762,N_4675,N_4965);
or U5763 (N_5763,N_4595,N_4326);
or U5764 (N_5764,N_4384,N_4081);
nand U5765 (N_5765,N_4171,N_4127);
nor U5766 (N_5766,N_4984,N_4330);
xnor U5767 (N_5767,N_4401,N_4290);
nand U5768 (N_5768,N_4262,N_4616);
nor U5769 (N_5769,N_4228,N_4438);
nor U5770 (N_5770,N_4957,N_4152);
nand U5771 (N_5771,N_4542,N_4276);
nor U5772 (N_5772,N_4507,N_4853);
nand U5773 (N_5773,N_4849,N_4493);
nor U5774 (N_5774,N_4261,N_4628);
nand U5775 (N_5775,N_4558,N_4991);
nor U5776 (N_5776,N_4152,N_4250);
nand U5777 (N_5777,N_4309,N_4700);
nand U5778 (N_5778,N_4856,N_4108);
or U5779 (N_5779,N_4476,N_4005);
or U5780 (N_5780,N_4969,N_4676);
nor U5781 (N_5781,N_4409,N_4206);
and U5782 (N_5782,N_4523,N_4469);
and U5783 (N_5783,N_4650,N_4410);
xnor U5784 (N_5784,N_4150,N_4598);
xnor U5785 (N_5785,N_4094,N_4316);
nor U5786 (N_5786,N_4001,N_4804);
nor U5787 (N_5787,N_4421,N_4936);
nand U5788 (N_5788,N_4023,N_4031);
and U5789 (N_5789,N_4105,N_4699);
or U5790 (N_5790,N_4862,N_4599);
xnor U5791 (N_5791,N_4869,N_4152);
nor U5792 (N_5792,N_4974,N_4056);
nand U5793 (N_5793,N_4166,N_4230);
nor U5794 (N_5794,N_4775,N_4847);
nand U5795 (N_5795,N_4971,N_4275);
and U5796 (N_5796,N_4444,N_4788);
and U5797 (N_5797,N_4255,N_4257);
or U5798 (N_5798,N_4246,N_4513);
nand U5799 (N_5799,N_4312,N_4382);
nor U5800 (N_5800,N_4282,N_4046);
and U5801 (N_5801,N_4487,N_4526);
or U5802 (N_5802,N_4898,N_4956);
nand U5803 (N_5803,N_4956,N_4034);
or U5804 (N_5804,N_4756,N_4394);
or U5805 (N_5805,N_4863,N_4117);
nor U5806 (N_5806,N_4631,N_4194);
nor U5807 (N_5807,N_4022,N_4017);
nand U5808 (N_5808,N_4718,N_4933);
and U5809 (N_5809,N_4726,N_4003);
nand U5810 (N_5810,N_4429,N_4004);
or U5811 (N_5811,N_4698,N_4106);
nor U5812 (N_5812,N_4051,N_4086);
nand U5813 (N_5813,N_4520,N_4362);
and U5814 (N_5814,N_4525,N_4750);
nor U5815 (N_5815,N_4920,N_4060);
nor U5816 (N_5816,N_4377,N_4013);
or U5817 (N_5817,N_4394,N_4143);
nand U5818 (N_5818,N_4282,N_4841);
and U5819 (N_5819,N_4628,N_4509);
or U5820 (N_5820,N_4206,N_4148);
nor U5821 (N_5821,N_4913,N_4096);
nand U5822 (N_5822,N_4039,N_4728);
nor U5823 (N_5823,N_4251,N_4272);
or U5824 (N_5824,N_4489,N_4807);
and U5825 (N_5825,N_4540,N_4791);
xor U5826 (N_5826,N_4679,N_4394);
nand U5827 (N_5827,N_4527,N_4698);
nand U5828 (N_5828,N_4498,N_4534);
nand U5829 (N_5829,N_4957,N_4482);
nor U5830 (N_5830,N_4381,N_4765);
and U5831 (N_5831,N_4123,N_4256);
nor U5832 (N_5832,N_4123,N_4097);
xnor U5833 (N_5833,N_4356,N_4098);
or U5834 (N_5834,N_4455,N_4803);
or U5835 (N_5835,N_4819,N_4955);
and U5836 (N_5836,N_4464,N_4155);
nand U5837 (N_5837,N_4806,N_4742);
and U5838 (N_5838,N_4933,N_4078);
nand U5839 (N_5839,N_4644,N_4535);
and U5840 (N_5840,N_4620,N_4355);
nor U5841 (N_5841,N_4809,N_4748);
nor U5842 (N_5842,N_4295,N_4657);
nor U5843 (N_5843,N_4003,N_4391);
or U5844 (N_5844,N_4348,N_4409);
nor U5845 (N_5845,N_4571,N_4982);
and U5846 (N_5846,N_4070,N_4203);
nor U5847 (N_5847,N_4270,N_4999);
and U5848 (N_5848,N_4422,N_4487);
or U5849 (N_5849,N_4605,N_4020);
and U5850 (N_5850,N_4238,N_4148);
and U5851 (N_5851,N_4779,N_4386);
or U5852 (N_5852,N_4980,N_4371);
or U5853 (N_5853,N_4399,N_4673);
or U5854 (N_5854,N_4297,N_4926);
and U5855 (N_5855,N_4077,N_4195);
nor U5856 (N_5856,N_4786,N_4801);
nand U5857 (N_5857,N_4644,N_4986);
nor U5858 (N_5858,N_4297,N_4425);
xor U5859 (N_5859,N_4446,N_4900);
and U5860 (N_5860,N_4494,N_4928);
nand U5861 (N_5861,N_4300,N_4618);
nand U5862 (N_5862,N_4486,N_4659);
nand U5863 (N_5863,N_4855,N_4495);
or U5864 (N_5864,N_4008,N_4408);
or U5865 (N_5865,N_4324,N_4934);
and U5866 (N_5866,N_4200,N_4919);
and U5867 (N_5867,N_4109,N_4593);
or U5868 (N_5868,N_4312,N_4940);
or U5869 (N_5869,N_4135,N_4430);
nor U5870 (N_5870,N_4804,N_4831);
or U5871 (N_5871,N_4341,N_4395);
nor U5872 (N_5872,N_4832,N_4900);
and U5873 (N_5873,N_4398,N_4726);
nand U5874 (N_5874,N_4503,N_4363);
and U5875 (N_5875,N_4622,N_4400);
or U5876 (N_5876,N_4241,N_4467);
nor U5877 (N_5877,N_4645,N_4158);
nor U5878 (N_5878,N_4157,N_4586);
xnor U5879 (N_5879,N_4343,N_4751);
or U5880 (N_5880,N_4162,N_4826);
or U5881 (N_5881,N_4347,N_4542);
and U5882 (N_5882,N_4489,N_4479);
nor U5883 (N_5883,N_4757,N_4885);
nor U5884 (N_5884,N_4665,N_4840);
or U5885 (N_5885,N_4702,N_4853);
and U5886 (N_5886,N_4269,N_4608);
and U5887 (N_5887,N_4430,N_4660);
nand U5888 (N_5888,N_4629,N_4908);
xor U5889 (N_5889,N_4733,N_4677);
or U5890 (N_5890,N_4297,N_4298);
or U5891 (N_5891,N_4130,N_4793);
or U5892 (N_5892,N_4212,N_4435);
xor U5893 (N_5893,N_4220,N_4467);
or U5894 (N_5894,N_4046,N_4949);
and U5895 (N_5895,N_4584,N_4453);
or U5896 (N_5896,N_4358,N_4925);
and U5897 (N_5897,N_4609,N_4785);
nand U5898 (N_5898,N_4215,N_4988);
and U5899 (N_5899,N_4160,N_4254);
nand U5900 (N_5900,N_4186,N_4277);
and U5901 (N_5901,N_4989,N_4280);
nor U5902 (N_5902,N_4067,N_4460);
nor U5903 (N_5903,N_4927,N_4807);
nand U5904 (N_5904,N_4949,N_4549);
nor U5905 (N_5905,N_4435,N_4792);
or U5906 (N_5906,N_4242,N_4912);
nand U5907 (N_5907,N_4237,N_4585);
nand U5908 (N_5908,N_4763,N_4995);
nand U5909 (N_5909,N_4812,N_4305);
or U5910 (N_5910,N_4086,N_4105);
nand U5911 (N_5911,N_4543,N_4501);
nor U5912 (N_5912,N_4981,N_4228);
or U5913 (N_5913,N_4001,N_4741);
or U5914 (N_5914,N_4274,N_4441);
xnor U5915 (N_5915,N_4618,N_4483);
or U5916 (N_5916,N_4041,N_4666);
and U5917 (N_5917,N_4089,N_4951);
or U5918 (N_5918,N_4167,N_4014);
nor U5919 (N_5919,N_4731,N_4926);
nand U5920 (N_5920,N_4408,N_4669);
nand U5921 (N_5921,N_4195,N_4386);
nor U5922 (N_5922,N_4948,N_4812);
or U5923 (N_5923,N_4327,N_4237);
nor U5924 (N_5924,N_4532,N_4748);
nand U5925 (N_5925,N_4308,N_4843);
nand U5926 (N_5926,N_4405,N_4570);
and U5927 (N_5927,N_4310,N_4266);
or U5928 (N_5928,N_4923,N_4878);
nand U5929 (N_5929,N_4461,N_4705);
or U5930 (N_5930,N_4629,N_4688);
nand U5931 (N_5931,N_4901,N_4502);
or U5932 (N_5932,N_4229,N_4006);
and U5933 (N_5933,N_4361,N_4303);
nor U5934 (N_5934,N_4587,N_4139);
nand U5935 (N_5935,N_4972,N_4188);
or U5936 (N_5936,N_4092,N_4135);
and U5937 (N_5937,N_4621,N_4635);
or U5938 (N_5938,N_4485,N_4203);
and U5939 (N_5939,N_4219,N_4053);
and U5940 (N_5940,N_4722,N_4630);
or U5941 (N_5941,N_4863,N_4710);
and U5942 (N_5942,N_4155,N_4076);
nand U5943 (N_5943,N_4950,N_4819);
and U5944 (N_5944,N_4495,N_4553);
nand U5945 (N_5945,N_4539,N_4428);
or U5946 (N_5946,N_4042,N_4428);
or U5947 (N_5947,N_4364,N_4918);
nor U5948 (N_5948,N_4698,N_4746);
nor U5949 (N_5949,N_4377,N_4378);
and U5950 (N_5950,N_4835,N_4015);
nor U5951 (N_5951,N_4167,N_4798);
or U5952 (N_5952,N_4239,N_4354);
or U5953 (N_5953,N_4983,N_4781);
nand U5954 (N_5954,N_4411,N_4991);
nand U5955 (N_5955,N_4724,N_4031);
or U5956 (N_5956,N_4941,N_4797);
nand U5957 (N_5957,N_4907,N_4804);
nor U5958 (N_5958,N_4422,N_4948);
and U5959 (N_5959,N_4541,N_4692);
and U5960 (N_5960,N_4780,N_4071);
nand U5961 (N_5961,N_4952,N_4065);
or U5962 (N_5962,N_4398,N_4560);
or U5963 (N_5963,N_4087,N_4090);
nand U5964 (N_5964,N_4306,N_4051);
or U5965 (N_5965,N_4344,N_4459);
nand U5966 (N_5966,N_4416,N_4039);
nand U5967 (N_5967,N_4426,N_4148);
or U5968 (N_5968,N_4653,N_4127);
and U5969 (N_5969,N_4951,N_4456);
nor U5970 (N_5970,N_4579,N_4875);
nor U5971 (N_5971,N_4496,N_4331);
nand U5972 (N_5972,N_4950,N_4923);
nor U5973 (N_5973,N_4700,N_4570);
and U5974 (N_5974,N_4194,N_4884);
nand U5975 (N_5975,N_4496,N_4261);
or U5976 (N_5976,N_4957,N_4491);
nor U5977 (N_5977,N_4251,N_4738);
nor U5978 (N_5978,N_4644,N_4750);
nand U5979 (N_5979,N_4472,N_4311);
nor U5980 (N_5980,N_4658,N_4924);
nand U5981 (N_5981,N_4173,N_4795);
and U5982 (N_5982,N_4551,N_4369);
and U5983 (N_5983,N_4972,N_4420);
and U5984 (N_5984,N_4575,N_4180);
and U5985 (N_5985,N_4694,N_4332);
or U5986 (N_5986,N_4596,N_4743);
nand U5987 (N_5987,N_4223,N_4322);
or U5988 (N_5988,N_4232,N_4566);
or U5989 (N_5989,N_4476,N_4249);
nand U5990 (N_5990,N_4544,N_4191);
and U5991 (N_5991,N_4714,N_4902);
nand U5992 (N_5992,N_4158,N_4777);
nor U5993 (N_5993,N_4107,N_4047);
nor U5994 (N_5994,N_4457,N_4746);
or U5995 (N_5995,N_4145,N_4640);
nand U5996 (N_5996,N_4908,N_4571);
or U5997 (N_5997,N_4808,N_4897);
or U5998 (N_5998,N_4274,N_4233);
nand U5999 (N_5999,N_4652,N_4906);
nand U6000 (N_6000,N_5328,N_5163);
nor U6001 (N_6001,N_5860,N_5824);
nand U6002 (N_6002,N_5287,N_5435);
nand U6003 (N_6003,N_5588,N_5696);
and U6004 (N_6004,N_5181,N_5322);
and U6005 (N_6005,N_5316,N_5686);
nand U6006 (N_6006,N_5647,N_5036);
nand U6007 (N_6007,N_5775,N_5285);
xor U6008 (N_6008,N_5528,N_5858);
nand U6009 (N_6009,N_5545,N_5275);
or U6010 (N_6010,N_5204,N_5025);
or U6011 (N_6011,N_5792,N_5683);
nor U6012 (N_6012,N_5185,N_5042);
nand U6013 (N_6013,N_5644,N_5561);
or U6014 (N_6014,N_5235,N_5305);
nand U6015 (N_6015,N_5665,N_5315);
nor U6016 (N_6016,N_5299,N_5355);
nor U6017 (N_6017,N_5820,N_5425);
nor U6018 (N_6018,N_5700,N_5623);
and U6019 (N_6019,N_5766,N_5648);
and U6020 (N_6020,N_5241,N_5890);
or U6021 (N_6021,N_5747,N_5332);
and U6022 (N_6022,N_5104,N_5074);
nor U6023 (N_6023,N_5082,N_5256);
nand U6024 (N_6024,N_5539,N_5306);
nor U6025 (N_6025,N_5385,N_5353);
nand U6026 (N_6026,N_5952,N_5313);
nor U6027 (N_6027,N_5897,N_5230);
or U6028 (N_6028,N_5610,N_5872);
nor U6029 (N_6029,N_5857,N_5838);
or U6030 (N_6030,N_5251,N_5409);
or U6031 (N_6031,N_5173,N_5264);
nor U6032 (N_6032,N_5200,N_5221);
nand U6033 (N_6033,N_5721,N_5568);
nor U6034 (N_6034,N_5601,N_5517);
or U6035 (N_6035,N_5366,N_5718);
and U6036 (N_6036,N_5951,N_5995);
xnor U6037 (N_6037,N_5945,N_5319);
nand U6038 (N_6038,N_5189,N_5988);
nand U6039 (N_6039,N_5598,N_5302);
nor U6040 (N_6040,N_5000,N_5632);
and U6041 (N_6041,N_5252,N_5667);
nand U6042 (N_6042,N_5845,N_5158);
nand U6043 (N_6043,N_5039,N_5006);
or U6044 (N_6044,N_5183,N_5453);
nor U6045 (N_6045,N_5541,N_5512);
nand U6046 (N_6046,N_5909,N_5882);
or U6047 (N_6047,N_5819,N_5320);
or U6048 (N_6048,N_5123,N_5680);
and U6049 (N_6049,N_5823,N_5768);
nor U6050 (N_6050,N_5154,N_5867);
or U6051 (N_6051,N_5645,N_5776);
nor U6052 (N_6052,N_5078,N_5854);
and U6053 (N_6053,N_5965,N_5091);
nand U6054 (N_6054,N_5238,N_5046);
nand U6055 (N_6055,N_5658,N_5779);
nand U6056 (N_6056,N_5757,N_5628);
or U6057 (N_6057,N_5467,N_5578);
or U6058 (N_6058,N_5605,N_5651);
nor U6059 (N_6059,N_5919,N_5770);
nand U6060 (N_6060,N_5953,N_5184);
xnor U6061 (N_6061,N_5224,N_5276);
or U6062 (N_6062,N_5745,N_5210);
and U6063 (N_6063,N_5755,N_5912);
nand U6064 (N_6064,N_5109,N_5612);
nor U6065 (N_6065,N_5841,N_5936);
and U6066 (N_6066,N_5688,N_5192);
or U6067 (N_6067,N_5582,N_5636);
or U6068 (N_6068,N_5484,N_5555);
nand U6069 (N_6069,N_5284,N_5124);
or U6070 (N_6070,N_5174,N_5629);
and U6071 (N_6071,N_5321,N_5834);
nor U6072 (N_6072,N_5412,N_5070);
nor U6073 (N_6073,N_5434,N_5053);
nand U6074 (N_6074,N_5452,N_5408);
and U6075 (N_6075,N_5771,N_5971);
nor U6076 (N_6076,N_5538,N_5175);
xor U6077 (N_6077,N_5339,N_5195);
nor U6078 (N_6078,N_5169,N_5215);
or U6079 (N_6079,N_5875,N_5527);
xor U6080 (N_6080,N_5933,N_5944);
nand U6081 (N_6081,N_5607,N_5630);
or U6082 (N_6082,N_5915,N_5788);
nor U6083 (N_6083,N_5448,N_5551);
xnor U6084 (N_6084,N_5116,N_5827);
nor U6085 (N_6085,N_5344,N_5120);
or U6086 (N_6086,N_5507,N_5115);
and U6087 (N_6087,N_5994,N_5444);
xor U6088 (N_6088,N_5013,N_5048);
xor U6089 (N_6089,N_5996,N_5007);
or U6090 (N_6090,N_5505,N_5217);
nor U6091 (N_6091,N_5659,N_5061);
and U6092 (N_6092,N_5278,N_5341);
nand U6093 (N_6093,N_5022,N_5863);
nand U6094 (N_6094,N_5375,N_5575);
or U6095 (N_6095,N_5808,N_5938);
and U6096 (N_6096,N_5350,N_5990);
nor U6097 (N_6097,N_5619,N_5734);
or U6098 (N_6098,N_5811,N_5018);
and U6099 (N_6099,N_5564,N_5725);
or U6100 (N_6100,N_5798,N_5684);
and U6101 (N_6101,N_5262,N_5443);
and U6102 (N_6102,N_5088,N_5511);
nor U6103 (N_6103,N_5325,N_5806);
nor U6104 (N_6104,N_5168,N_5327);
and U6105 (N_6105,N_5099,N_5454);
xnor U6106 (N_6106,N_5514,N_5490);
nand U6107 (N_6107,N_5597,N_5232);
nand U6108 (N_6108,N_5144,N_5420);
or U6109 (N_6109,N_5159,N_5386);
and U6110 (N_6110,N_5577,N_5281);
and U6111 (N_6111,N_5843,N_5624);
or U6112 (N_6112,N_5874,N_5141);
and U6113 (N_6113,N_5803,N_5787);
nor U6114 (N_6114,N_5001,N_5333);
nand U6115 (N_6115,N_5250,N_5016);
xnor U6116 (N_6116,N_5428,N_5298);
xnor U6117 (N_6117,N_5859,N_5615);
nand U6118 (N_6118,N_5201,N_5323);
and U6119 (N_6119,N_5458,N_5566);
and U6120 (N_6120,N_5913,N_5495);
nor U6121 (N_6121,N_5966,N_5712);
nand U6122 (N_6122,N_5924,N_5969);
and U6123 (N_6123,N_5796,N_5460);
or U6124 (N_6124,N_5893,N_5621);
nand U6125 (N_6125,N_5393,N_5655);
nand U6126 (N_6126,N_5160,N_5885);
nor U6127 (N_6127,N_5617,N_5149);
nor U6128 (N_6128,N_5678,N_5589);
nand U6129 (N_6129,N_5852,N_5613);
or U6130 (N_6130,N_5590,N_5892);
nor U6131 (N_6131,N_5973,N_5842);
and U6132 (N_6132,N_5161,N_5482);
nand U6133 (N_6133,N_5401,N_5832);
nor U6134 (N_6134,N_5244,N_5957);
or U6135 (N_6135,N_5382,N_5853);
or U6136 (N_6136,N_5245,N_5100);
and U6137 (N_6137,N_5999,N_5439);
or U6138 (N_6138,N_5081,N_5270);
or U6139 (N_6139,N_5818,N_5113);
and U6140 (N_6140,N_5553,N_5704);
or U6141 (N_6141,N_5743,N_5034);
nor U6142 (N_6142,N_5493,N_5504);
nor U6143 (N_6143,N_5812,N_5560);
nand U6144 (N_6144,N_5054,N_5030);
or U6145 (N_6145,N_5438,N_5941);
nand U6146 (N_6146,N_5170,N_5019);
or U6147 (N_6147,N_5431,N_5653);
and U6148 (N_6148,N_5228,N_5259);
nand U6149 (N_6149,N_5660,N_5419);
nor U6150 (N_6150,N_5058,N_5057);
nand U6151 (N_6151,N_5426,N_5318);
nor U6152 (N_6152,N_5172,N_5643);
nand U6153 (N_6153,N_5027,N_5413);
and U6154 (N_6154,N_5571,N_5646);
or U6155 (N_6155,N_5668,N_5871);
xnor U6156 (N_6156,N_5804,N_5047);
nor U6157 (N_6157,N_5411,N_5637);
nand U6158 (N_6158,N_5618,N_5675);
or U6159 (N_6159,N_5503,N_5279);
xnor U6160 (N_6160,N_5772,N_5155);
nand U6161 (N_6161,N_5334,N_5194);
nor U6162 (N_6162,N_5178,N_5023);
and U6163 (N_6163,N_5106,N_5947);
nand U6164 (N_6164,N_5979,N_5083);
nand U6165 (N_6165,N_5710,N_5707);
or U6166 (N_6166,N_5657,N_5906);
nand U6167 (N_6167,N_5763,N_5379);
nand U6168 (N_6168,N_5098,N_5166);
nand U6169 (N_6169,N_5246,N_5716);
nor U6170 (N_6170,N_5369,N_5076);
nand U6171 (N_6171,N_5356,N_5608);
or U6172 (N_6172,N_5662,N_5028);
or U6173 (N_6173,N_5015,N_5186);
and U6174 (N_6174,N_5390,N_5446);
or U6175 (N_6175,N_5067,N_5071);
and U6176 (N_6176,N_5072,N_5457);
nor U6177 (N_6177,N_5301,N_5469);
and U6178 (N_6178,N_5380,N_5694);
and U6179 (N_6179,N_5233,N_5652);
and U6180 (N_6180,N_5993,N_5666);
or U6181 (N_6181,N_5922,N_5569);
and U6182 (N_6182,N_5593,N_5984);
and U6183 (N_6183,N_5263,N_5759);
nand U6184 (N_6184,N_5724,N_5423);
nand U6185 (N_6185,N_5220,N_5849);
or U6186 (N_6186,N_5889,N_5229);
or U6187 (N_6187,N_5272,N_5536);
or U6188 (N_6188,N_5387,N_5131);
or U6189 (N_6189,N_5405,N_5987);
and U6190 (N_6190,N_5801,N_5862);
nand U6191 (N_6191,N_5157,N_5701);
and U6192 (N_6192,N_5898,N_5357);
nor U6193 (N_6193,N_5733,N_5376);
or U6194 (N_6194,N_5231,N_5142);
xor U6195 (N_6195,N_5362,N_5295);
nand U6196 (N_6196,N_5592,N_5679);
nand U6197 (N_6197,N_5153,N_5625);
and U6198 (N_6198,N_5519,N_5171);
and U6199 (N_6199,N_5523,N_5135);
nand U6200 (N_6200,N_5261,N_5762);
and U6201 (N_6201,N_5465,N_5156);
nand U6202 (N_6202,N_5914,N_5080);
nor U6203 (N_6203,N_5440,N_5833);
or U6204 (N_6204,N_5813,N_5449);
nand U6205 (N_6205,N_5329,N_5300);
or U6206 (N_6206,N_5085,N_5211);
or U6207 (N_6207,N_5414,N_5273);
or U6208 (N_6208,N_5126,N_5222);
nand U6209 (N_6209,N_5927,N_5430);
nor U6210 (N_6210,N_5292,N_5873);
and U6211 (N_6211,N_5525,N_5641);
nand U6212 (N_6212,N_5127,N_5374);
nand U6213 (N_6213,N_5587,N_5308);
and U6214 (N_6214,N_5209,N_5243);
and U6215 (N_6215,N_5744,N_5368);
and U6216 (N_6216,N_5370,N_5537);
and U6217 (N_6217,N_5017,N_5840);
and U6218 (N_6218,N_5518,N_5112);
and U6219 (N_6219,N_5214,N_5959);
or U6220 (N_6220,N_5483,N_5522);
or U6221 (N_6221,N_5090,N_5399);
and U6222 (N_6222,N_5753,N_5227);
xor U6223 (N_6223,N_5826,N_5547);
and U6224 (N_6224,N_5976,N_5778);
or U6225 (N_6225,N_5992,N_5946);
nor U6226 (N_6226,N_5242,N_5111);
nor U6227 (N_6227,N_5021,N_5869);
xnor U6228 (N_6228,N_5199,N_5433);
and U6229 (N_6229,N_5935,N_5807);
and U6230 (N_6230,N_5394,N_5499);
nand U6231 (N_6231,N_5478,N_5672);
nor U6232 (N_6232,N_5005,N_5365);
nand U6233 (N_6233,N_5631,N_5087);
nor U6234 (N_6234,N_5014,N_5740);
and U6235 (N_6235,N_5634,N_5572);
and U6236 (N_6236,N_5622,N_5218);
and U6237 (N_6237,N_5925,N_5958);
nand U6238 (N_6238,N_5736,N_5506);
nor U6239 (N_6239,N_5825,N_5654);
nand U6240 (N_6240,N_5343,N_5765);
nand U6241 (N_6241,N_5586,N_5864);
nand U6242 (N_6242,N_5866,N_5462);
nand U6243 (N_6243,N_5468,N_5761);
or U6244 (N_6244,N_5650,N_5777);
nor U6245 (N_6245,N_5312,N_5474);
nand U6246 (N_6246,N_5486,N_5162);
and U6247 (N_6247,N_5554,N_5949);
and U6248 (N_6248,N_5026,N_5052);
nand U6249 (N_6249,N_5865,N_5349);
and U6250 (N_6250,N_5060,N_5364);
or U6251 (N_6251,N_5237,N_5004);
nand U6252 (N_6252,N_5089,N_5533);
nor U6253 (N_6253,N_5702,N_5129);
nor U6254 (N_6254,N_5219,N_5565);
or U6255 (N_6255,N_5513,N_5697);
and U6256 (N_6256,N_5501,N_5682);
or U6257 (N_6257,N_5029,N_5674);
nand U6258 (N_6258,N_5404,N_5427);
and U6259 (N_6259,N_5132,N_5360);
or U6260 (N_6260,N_5836,N_5714);
xnor U6261 (N_6261,N_5746,N_5397);
nand U6262 (N_6262,N_5363,N_5145);
nand U6263 (N_6263,N_5870,N_5955);
and U6264 (N_6264,N_5455,N_5497);
and U6265 (N_6265,N_5311,N_5165);
and U6266 (N_6266,N_5212,N_5754);
or U6267 (N_6267,N_5176,N_5602);
xnor U6268 (N_6268,N_5481,N_5253);
or U6269 (N_6269,N_5708,N_5715);
nand U6270 (N_6270,N_5516,N_5293);
xor U6271 (N_6271,N_5649,N_5283);
and U6272 (N_6272,N_5929,N_5167);
and U6273 (N_6273,N_5239,N_5225);
or U6274 (N_6274,N_5340,N_5208);
nand U6275 (N_6275,N_5422,N_5905);
nor U6276 (N_6276,N_5456,N_5307);
and U6277 (N_6277,N_5730,N_5473);
and U6278 (N_6278,N_5317,N_5839);
and U6279 (N_6279,N_5614,N_5508);
and U6280 (N_6280,N_5290,N_5760);
nor U6281 (N_6281,N_5774,N_5073);
nand U6282 (N_6282,N_5883,N_5748);
nand U6283 (N_6283,N_5773,N_5930);
and U6284 (N_6284,N_5611,N_5732);
nand U6285 (N_6285,N_5559,N_5795);
and U6286 (N_6286,N_5720,N_5346);
nor U6287 (N_6287,N_5020,N_5557);
or U6288 (N_6288,N_5967,N_5280);
and U6289 (N_6289,N_5418,N_5268);
and U6290 (N_6290,N_5920,N_5471);
or U6291 (N_6291,N_5868,N_5240);
and U6292 (N_6292,N_5972,N_5805);
and U6293 (N_6293,N_5193,N_5681);
nor U6294 (N_6294,N_5782,N_5676);
nand U6295 (N_6295,N_5887,N_5596);
nand U6296 (N_6296,N_5670,N_5485);
or U6297 (N_6297,N_5510,N_5410);
or U6298 (N_6298,N_5814,N_5381);
nand U6299 (N_6299,N_5002,N_5878);
and U6300 (N_6300,N_5549,N_5703);
and U6301 (N_6301,N_5729,N_5529);
nand U6302 (N_6302,N_5406,N_5671);
nor U6303 (N_6303,N_5692,N_5981);
nand U6304 (N_6304,N_5378,N_5330);
nor U6305 (N_6305,N_5271,N_5828);
and U6306 (N_6306,N_5540,N_5881);
xor U6307 (N_6307,N_5041,N_5921);
nand U6308 (N_6308,N_5861,N_5303);
and U6309 (N_6309,N_5846,N_5459);
or U6310 (N_6310,N_5437,N_5147);
or U6311 (N_6311,N_5249,N_5635);
nand U6312 (N_6312,N_5476,N_5573);
nand U6313 (N_6313,N_5255,N_5847);
or U6314 (N_6314,N_5267,N_5962);
and U6315 (N_6315,N_5102,N_5500);
and U6316 (N_6316,N_5886,N_5257);
or U6317 (N_6317,N_5982,N_5741);
nand U6318 (N_6318,N_5960,N_5896);
nand U6319 (N_6319,N_5354,N_5128);
nand U6320 (N_6320,N_5661,N_5558);
and U6321 (N_6321,N_5384,N_5130);
nor U6322 (N_6322,N_5373,N_5463);
and U6323 (N_6323,N_5737,N_5923);
and U6324 (N_6324,N_5574,N_5134);
nor U6325 (N_6325,N_5093,N_5509);
and U6326 (N_6326,N_5790,N_5136);
xor U6327 (N_6327,N_5361,N_5785);
or U6328 (N_6328,N_5639,N_5822);
nand U6329 (N_6329,N_5584,N_5583);
nand U6330 (N_6330,N_5282,N_5050);
xnor U6331 (N_6331,N_5464,N_5851);
or U6332 (N_6332,N_5855,N_5544);
nand U6333 (N_6333,N_5910,N_5799);
nand U6334 (N_6334,N_5726,N_5604);
or U6335 (N_6335,N_5931,N_5656);
and U6336 (N_6336,N_5236,N_5829);
nand U6337 (N_6337,N_5880,N_5442);
or U6338 (N_6338,N_5148,N_5198);
and U6339 (N_6339,N_5024,N_5092);
or U6340 (N_6340,N_5901,N_5108);
and U6341 (N_6341,N_5068,N_5358);
and U6342 (N_6342,N_5391,N_5884);
nand U6343 (N_6343,N_5977,N_5722);
nor U6344 (N_6344,N_5690,N_5043);
or U6345 (N_6345,N_5556,N_5717);
nand U6346 (N_6346,N_5105,N_5943);
nand U6347 (N_6347,N_5942,N_5530);
nor U6348 (N_6348,N_5638,N_5698);
nand U6349 (N_6349,N_5258,N_5663);
nand U6350 (N_6350,N_5664,N_5395);
and U6351 (N_6351,N_5342,N_5040);
nor U6352 (N_6352,N_5207,N_5084);
nor U6353 (N_6353,N_5968,N_5314);
and U6354 (N_6354,N_5196,N_5324);
nand U6355 (N_6355,N_5937,N_5576);
or U6356 (N_6356,N_5064,N_5786);
and U6357 (N_6357,N_5673,N_5907);
and U6358 (N_6358,N_5062,N_5254);
and U6359 (N_6359,N_5352,N_5494);
nand U6360 (N_6360,N_5521,N_5415);
and U6361 (N_6361,N_5269,N_5917);
nor U6362 (N_6362,N_5986,N_5187);
nor U6363 (N_6363,N_5543,N_5642);
xnor U6364 (N_6364,N_5294,N_5107);
and U6365 (N_6365,N_5223,N_5902);
nor U6366 (N_6366,N_5837,N_5095);
nor U6367 (N_6367,N_5580,N_5830);
or U6368 (N_6368,N_5756,N_5336);
and U6369 (N_6369,N_5248,N_5784);
nand U6370 (N_6370,N_5562,N_5003);
nor U6371 (N_6371,N_5570,N_5980);
or U6372 (N_6372,N_5164,N_5532);
and U6373 (N_6373,N_5934,N_5472);
or U6374 (N_6374,N_5809,N_5479);
nor U6375 (N_6375,N_5338,N_5677);
and U6376 (N_6376,N_5203,N_5388);
or U6377 (N_6377,N_5531,N_5975);
nand U6378 (N_6378,N_5009,N_5594);
or U6379 (N_6379,N_5691,N_5769);
or U6380 (N_6380,N_5234,N_5146);
or U6381 (N_6381,N_5407,N_5151);
nand U6382 (N_6382,N_5265,N_5288);
and U6383 (N_6383,N_5140,N_5125);
or U6384 (N_6384,N_5488,N_5010);
nor U6385 (N_6385,N_5063,N_5821);
or U6386 (N_6386,N_5989,N_5429);
nand U6387 (N_6387,N_5626,N_5856);
and U6388 (N_6388,N_5492,N_5310);
or U6389 (N_6389,N_5075,N_5377);
nor U6390 (N_6390,N_5954,N_5143);
nor U6391 (N_6391,N_5094,N_5445);
nand U6392 (N_6392,N_5752,N_5260);
nor U6393 (N_6393,N_5810,N_5693);
nand U6394 (N_6394,N_5119,N_5879);
or U6395 (N_6395,N_5926,N_5542);
and U6396 (N_6396,N_5266,N_5932);
nand U6397 (N_6397,N_5451,N_5424);
nand U6398 (N_6398,N_5964,N_5117);
nand U6399 (N_6399,N_5206,N_5817);
and U6400 (N_6400,N_5188,N_5038);
or U6401 (N_6401,N_5791,N_5491);
nand U6402 (N_6402,N_5190,N_5940);
and U6403 (N_6403,N_5421,N_5398);
xnor U6404 (N_6404,N_5470,N_5502);
xnor U6405 (N_6405,N_5728,N_5903);
and U6406 (N_6406,N_5815,N_5526);
nor U6407 (N_6407,N_5277,N_5051);
or U6408 (N_6408,N_5037,N_5182);
nor U6409 (N_6409,N_5563,N_5738);
or U6410 (N_6410,N_5480,N_5591);
nand U6411 (N_6411,N_5297,N_5191);
nor U6412 (N_6412,N_5794,N_5735);
and U6413 (N_6413,N_5331,N_5848);
and U6414 (N_6414,N_5035,N_5461);
nor U6415 (N_6415,N_5546,N_5477);
and U6416 (N_6416,N_5606,N_5447);
or U6417 (N_6417,N_5974,N_5751);
and U6418 (N_6418,N_5077,N_5894);
or U6419 (N_6419,N_5065,N_5475);
and U6420 (N_6420,N_5534,N_5432);
and U6421 (N_6421,N_5705,N_5150);
nor U6422 (N_6422,N_5750,N_5520);
nand U6423 (N_6423,N_5689,N_5337);
or U6424 (N_6424,N_5059,N_5783);
and U6425 (N_6425,N_5609,N_5417);
and U6426 (N_6426,N_5079,N_5056);
nand U6427 (N_6427,N_5524,N_5086);
nand U6428 (N_6428,N_5709,N_5326);
nand U6429 (N_6429,N_5797,N_5097);
and U6430 (N_6430,N_5548,N_5139);
nand U6431 (N_6431,N_5758,N_5152);
or U6432 (N_6432,N_5603,N_5891);
nor U6433 (N_6433,N_5888,N_5392);
xor U6434 (N_6434,N_5956,N_5550);
and U6435 (N_6435,N_5296,N_5515);
nand U6436 (N_6436,N_5289,N_5970);
or U6437 (N_6437,N_5213,N_5137);
and U6438 (N_6438,N_5997,N_5844);
xnor U6439 (N_6439,N_5402,N_5695);
and U6440 (N_6440,N_5749,N_5101);
nor U6441 (N_6441,N_5118,N_5291);
or U6442 (N_6442,N_5103,N_5226);
or U6443 (N_6443,N_5496,N_5939);
and U6444 (N_6444,N_5396,N_5348);
and U6445 (N_6445,N_5274,N_5595);
or U6446 (N_6446,N_5309,N_5202);
nor U6447 (N_6447,N_5963,N_5835);
nor U6448 (N_6448,N_5371,N_5950);
or U6449 (N_6449,N_5831,N_5133);
nor U6450 (N_6450,N_5916,N_5948);
and U6451 (N_6451,N_5877,N_5535);
and U6452 (N_6452,N_5895,N_5816);
nor U6453 (N_6453,N_5247,N_5961);
nand U6454 (N_6454,N_5908,N_5335);
nand U6455 (N_6455,N_5985,N_5066);
or U6456 (N_6456,N_5489,N_5567);
nor U6457 (N_6457,N_5627,N_5978);
nand U6458 (N_6458,N_5552,N_5400);
or U6459 (N_6459,N_5789,N_5687);
nand U6460 (N_6460,N_5069,N_5055);
xor U6461 (N_6461,N_5585,N_5347);
or U6462 (N_6462,N_5719,N_5177);
nor U6463 (N_6463,N_5739,N_5928);
nand U6464 (N_6464,N_5731,N_5345);
nand U6465 (N_6465,N_5121,N_5012);
or U6466 (N_6466,N_5723,N_5899);
nand U6467 (N_6467,N_5600,N_5383);
nor U6468 (N_6468,N_5767,N_5049);
nor U6469 (N_6469,N_5579,N_5793);
or U6470 (N_6470,N_5033,N_5850);
nor U6471 (N_6471,N_5403,N_5031);
or U6472 (N_6472,N_5487,N_5599);
nand U6473 (N_6473,N_5742,N_5706);
and U6474 (N_6474,N_5122,N_5699);
and U6475 (N_6475,N_5180,N_5179);
nor U6476 (N_6476,N_5764,N_5367);
or U6477 (N_6477,N_5389,N_5138);
or U6478 (N_6478,N_5205,N_5781);
and U6479 (N_6479,N_5616,N_5466);
or U6480 (N_6480,N_5351,N_5216);
nor U6481 (N_6481,N_5727,N_5876);
nand U6482 (N_6482,N_5450,N_5581);
or U6483 (N_6483,N_5436,N_5900);
or U6484 (N_6484,N_5904,N_5633);
nand U6485 (N_6485,N_5110,N_5286);
or U6486 (N_6486,N_5711,N_5197);
and U6487 (N_6487,N_5713,N_5359);
nor U6488 (N_6488,N_5685,N_5096);
and U6489 (N_6489,N_5991,N_5998);
and U6490 (N_6490,N_5416,N_5802);
and U6491 (N_6491,N_5372,N_5441);
and U6492 (N_6492,N_5983,N_5032);
and U6493 (N_6493,N_5669,N_5620);
xor U6494 (N_6494,N_5911,N_5011);
xor U6495 (N_6495,N_5304,N_5918);
nand U6496 (N_6496,N_5800,N_5044);
and U6497 (N_6497,N_5780,N_5045);
nand U6498 (N_6498,N_5498,N_5640);
nor U6499 (N_6499,N_5008,N_5114);
and U6500 (N_6500,N_5060,N_5216);
or U6501 (N_6501,N_5913,N_5672);
nor U6502 (N_6502,N_5418,N_5007);
nand U6503 (N_6503,N_5450,N_5833);
or U6504 (N_6504,N_5377,N_5634);
nor U6505 (N_6505,N_5319,N_5109);
or U6506 (N_6506,N_5103,N_5901);
and U6507 (N_6507,N_5809,N_5648);
and U6508 (N_6508,N_5437,N_5397);
nor U6509 (N_6509,N_5082,N_5121);
nand U6510 (N_6510,N_5097,N_5350);
and U6511 (N_6511,N_5366,N_5148);
nor U6512 (N_6512,N_5487,N_5697);
nand U6513 (N_6513,N_5894,N_5879);
or U6514 (N_6514,N_5544,N_5758);
xnor U6515 (N_6515,N_5501,N_5618);
nor U6516 (N_6516,N_5428,N_5709);
nand U6517 (N_6517,N_5648,N_5817);
nor U6518 (N_6518,N_5426,N_5790);
and U6519 (N_6519,N_5898,N_5128);
nor U6520 (N_6520,N_5396,N_5045);
nand U6521 (N_6521,N_5159,N_5871);
nor U6522 (N_6522,N_5240,N_5752);
and U6523 (N_6523,N_5926,N_5090);
or U6524 (N_6524,N_5394,N_5455);
and U6525 (N_6525,N_5760,N_5489);
nand U6526 (N_6526,N_5084,N_5788);
or U6527 (N_6527,N_5708,N_5176);
or U6528 (N_6528,N_5830,N_5682);
nand U6529 (N_6529,N_5048,N_5757);
and U6530 (N_6530,N_5805,N_5449);
or U6531 (N_6531,N_5303,N_5482);
nand U6532 (N_6532,N_5561,N_5728);
or U6533 (N_6533,N_5326,N_5973);
or U6534 (N_6534,N_5353,N_5095);
nand U6535 (N_6535,N_5286,N_5139);
nor U6536 (N_6536,N_5403,N_5795);
nor U6537 (N_6537,N_5490,N_5060);
nor U6538 (N_6538,N_5830,N_5406);
and U6539 (N_6539,N_5719,N_5392);
and U6540 (N_6540,N_5058,N_5055);
and U6541 (N_6541,N_5947,N_5823);
or U6542 (N_6542,N_5288,N_5655);
nor U6543 (N_6543,N_5678,N_5395);
nand U6544 (N_6544,N_5509,N_5024);
and U6545 (N_6545,N_5008,N_5596);
and U6546 (N_6546,N_5891,N_5152);
xnor U6547 (N_6547,N_5646,N_5804);
and U6548 (N_6548,N_5823,N_5282);
and U6549 (N_6549,N_5135,N_5295);
or U6550 (N_6550,N_5747,N_5937);
nand U6551 (N_6551,N_5667,N_5634);
and U6552 (N_6552,N_5700,N_5672);
nand U6553 (N_6553,N_5658,N_5669);
and U6554 (N_6554,N_5209,N_5437);
or U6555 (N_6555,N_5732,N_5929);
nor U6556 (N_6556,N_5206,N_5738);
and U6557 (N_6557,N_5298,N_5982);
nand U6558 (N_6558,N_5997,N_5074);
and U6559 (N_6559,N_5259,N_5116);
and U6560 (N_6560,N_5947,N_5537);
or U6561 (N_6561,N_5016,N_5211);
nand U6562 (N_6562,N_5964,N_5482);
and U6563 (N_6563,N_5262,N_5991);
and U6564 (N_6564,N_5931,N_5627);
nand U6565 (N_6565,N_5166,N_5296);
nor U6566 (N_6566,N_5526,N_5415);
nor U6567 (N_6567,N_5499,N_5937);
nand U6568 (N_6568,N_5817,N_5287);
nor U6569 (N_6569,N_5518,N_5455);
or U6570 (N_6570,N_5265,N_5559);
nand U6571 (N_6571,N_5996,N_5514);
and U6572 (N_6572,N_5336,N_5749);
nor U6573 (N_6573,N_5909,N_5447);
nor U6574 (N_6574,N_5990,N_5169);
nor U6575 (N_6575,N_5343,N_5408);
nand U6576 (N_6576,N_5166,N_5734);
nor U6577 (N_6577,N_5093,N_5998);
or U6578 (N_6578,N_5235,N_5389);
or U6579 (N_6579,N_5803,N_5035);
or U6580 (N_6580,N_5913,N_5373);
or U6581 (N_6581,N_5415,N_5169);
nor U6582 (N_6582,N_5537,N_5842);
or U6583 (N_6583,N_5480,N_5280);
nand U6584 (N_6584,N_5730,N_5969);
and U6585 (N_6585,N_5082,N_5050);
nand U6586 (N_6586,N_5706,N_5875);
nor U6587 (N_6587,N_5569,N_5171);
nor U6588 (N_6588,N_5555,N_5090);
or U6589 (N_6589,N_5580,N_5685);
and U6590 (N_6590,N_5729,N_5891);
xor U6591 (N_6591,N_5176,N_5357);
or U6592 (N_6592,N_5840,N_5194);
nor U6593 (N_6593,N_5476,N_5042);
nand U6594 (N_6594,N_5176,N_5840);
and U6595 (N_6595,N_5329,N_5737);
xor U6596 (N_6596,N_5014,N_5680);
and U6597 (N_6597,N_5677,N_5495);
xor U6598 (N_6598,N_5905,N_5657);
nor U6599 (N_6599,N_5143,N_5342);
and U6600 (N_6600,N_5488,N_5114);
or U6601 (N_6601,N_5597,N_5983);
and U6602 (N_6602,N_5277,N_5374);
or U6603 (N_6603,N_5248,N_5466);
nor U6604 (N_6604,N_5201,N_5906);
or U6605 (N_6605,N_5102,N_5748);
nand U6606 (N_6606,N_5578,N_5860);
nand U6607 (N_6607,N_5195,N_5390);
and U6608 (N_6608,N_5551,N_5726);
and U6609 (N_6609,N_5113,N_5530);
nand U6610 (N_6610,N_5259,N_5390);
nand U6611 (N_6611,N_5540,N_5268);
or U6612 (N_6612,N_5117,N_5808);
or U6613 (N_6613,N_5277,N_5643);
or U6614 (N_6614,N_5317,N_5172);
nor U6615 (N_6615,N_5456,N_5468);
and U6616 (N_6616,N_5133,N_5883);
and U6617 (N_6617,N_5502,N_5496);
and U6618 (N_6618,N_5101,N_5502);
nand U6619 (N_6619,N_5212,N_5536);
and U6620 (N_6620,N_5039,N_5659);
nor U6621 (N_6621,N_5487,N_5072);
nor U6622 (N_6622,N_5329,N_5134);
or U6623 (N_6623,N_5505,N_5354);
nand U6624 (N_6624,N_5183,N_5390);
nand U6625 (N_6625,N_5761,N_5138);
nor U6626 (N_6626,N_5904,N_5754);
and U6627 (N_6627,N_5255,N_5849);
or U6628 (N_6628,N_5779,N_5635);
nor U6629 (N_6629,N_5628,N_5030);
nor U6630 (N_6630,N_5603,N_5838);
and U6631 (N_6631,N_5062,N_5531);
nand U6632 (N_6632,N_5611,N_5340);
or U6633 (N_6633,N_5524,N_5815);
nand U6634 (N_6634,N_5080,N_5068);
or U6635 (N_6635,N_5058,N_5115);
and U6636 (N_6636,N_5684,N_5460);
and U6637 (N_6637,N_5615,N_5028);
nand U6638 (N_6638,N_5509,N_5596);
nand U6639 (N_6639,N_5564,N_5798);
and U6640 (N_6640,N_5304,N_5294);
nand U6641 (N_6641,N_5862,N_5306);
nor U6642 (N_6642,N_5154,N_5620);
and U6643 (N_6643,N_5299,N_5678);
or U6644 (N_6644,N_5983,N_5933);
nand U6645 (N_6645,N_5985,N_5420);
nand U6646 (N_6646,N_5357,N_5799);
or U6647 (N_6647,N_5034,N_5678);
or U6648 (N_6648,N_5326,N_5225);
and U6649 (N_6649,N_5992,N_5166);
nor U6650 (N_6650,N_5907,N_5826);
nor U6651 (N_6651,N_5687,N_5366);
or U6652 (N_6652,N_5384,N_5347);
or U6653 (N_6653,N_5818,N_5677);
nand U6654 (N_6654,N_5290,N_5425);
nor U6655 (N_6655,N_5914,N_5093);
and U6656 (N_6656,N_5938,N_5025);
and U6657 (N_6657,N_5316,N_5856);
nor U6658 (N_6658,N_5246,N_5500);
nand U6659 (N_6659,N_5502,N_5346);
and U6660 (N_6660,N_5820,N_5506);
nor U6661 (N_6661,N_5977,N_5932);
nand U6662 (N_6662,N_5110,N_5064);
nand U6663 (N_6663,N_5459,N_5408);
or U6664 (N_6664,N_5127,N_5595);
and U6665 (N_6665,N_5931,N_5486);
and U6666 (N_6666,N_5472,N_5105);
nor U6667 (N_6667,N_5636,N_5923);
nor U6668 (N_6668,N_5131,N_5423);
nor U6669 (N_6669,N_5792,N_5380);
or U6670 (N_6670,N_5014,N_5827);
and U6671 (N_6671,N_5561,N_5134);
and U6672 (N_6672,N_5691,N_5383);
and U6673 (N_6673,N_5412,N_5149);
or U6674 (N_6674,N_5527,N_5590);
or U6675 (N_6675,N_5561,N_5763);
nor U6676 (N_6676,N_5202,N_5724);
or U6677 (N_6677,N_5913,N_5831);
nor U6678 (N_6678,N_5106,N_5146);
nand U6679 (N_6679,N_5944,N_5593);
nor U6680 (N_6680,N_5966,N_5751);
and U6681 (N_6681,N_5113,N_5849);
and U6682 (N_6682,N_5031,N_5626);
and U6683 (N_6683,N_5641,N_5792);
and U6684 (N_6684,N_5116,N_5424);
nand U6685 (N_6685,N_5191,N_5189);
or U6686 (N_6686,N_5376,N_5725);
or U6687 (N_6687,N_5251,N_5015);
nor U6688 (N_6688,N_5402,N_5132);
xnor U6689 (N_6689,N_5063,N_5532);
and U6690 (N_6690,N_5694,N_5516);
nand U6691 (N_6691,N_5394,N_5825);
nand U6692 (N_6692,N_5727,N_5155);
or U6693 (N_6693,N_5651,N_5361);
nand U6694 (N_6694,N_5403,N_5425);
and U6695 (N_6695,N_5646,N_5276);
and U6696 (N_6696,N_5208,N_5377);
or U6697 (N_6697,N_5937,N_5726);
xor U6698 (N_6698,N_5903,N_5617);
nor U6699 (N_6699,N_5609,N_5136);
nand U6700 (N_6700,N_5918,N_5979);
nand U6701 (N_6701,N_5253,N_5383);
nand U6702 (N_6702,N_5332,N_5061);
nand U6703 (N_6703,N_5976,N_5886);
nand U6704 (N_6704,N_5374,N_5129);
or U6705 (N_6705,N_5720,N_5367);
or U6706 (N_6706,N_5651,N_5242);
and U6707 (N_6707,N_5532,N_5178);
or U6708 (N_6708,N_5625,N_5783);
nor U6709 (N_6709,N_5517,N_5482);
nand U6710 (N_6710,N_5902,N_5749);
nand U6711 (N_6711,N_5312,N_5706);
nand U6712 (N_6712,N_5201,N_5539);
or U6713 (N_6713,N_5416,N_5801);
nor U6714 (N_6714,N_5055,N_5458);
nand U6715 (N_6715,N_5146,N_5023);
nor U6716 (N_6716,N_5028,N_5449);
and U6717 (N_6717,N_5510,N_5829);
nand U6718 (N_6718,N_5390,N_5150);
nand U6719 (N_6719,N_5794,N_5040);
nor U6720 (N_6720,N_5047,N_5218);
nor U6721 (N_6721,N_5450,N_5123);
and U6722 (N_6722,N_5882,N_5723);
nor U6723 (N_6723,N_5325,N_5706);
nor U6724 (N_6724,N_5159,N_5542);
nor U6725 (N_6725,N_5852,N_5611);
nor U6726 (N_6726,N_5855,N_5044);
or U6727 (N_6727,N_5717,N_5097);
nand U6728 (N_6728,N_5024,N_5649);
or U6729 (N_6729,N_5919,N_5462);
nor U6730 (N_6730,N_5568,N_5203);
nor U6731 (N_6731,N_5664,N_5658);
xor U6732 (N_6732,N_5207,N_5500);
or U6733 (N_6733,N_5802,N_5901);
nor U6734 (N_6734,N_5402,N_5596);
nor U6735 (N_6735,N_5384,N_5313);
or U6736 (N_6736,N_5303,N_5957);
or U6737 (N_6737,N_5160,N_5326);
nand U6738 (N_6738,N_5401,N_5927);
and U6739 (N_6739,N_5684,N_5373);
nor U6740 (N_6740,N_5279,N_5680);
or U6741 (N_6741,N_5939,N_5734);
and U6742 (N_6742,N_5498,N_5574);
and U6743 (N_6743,N_5821,N_5221);
nand U6744 (N_6744,N_5883,N_5828);
or U6745 (N_6745,N_5057,N_5442);
nand U6746 (N_6746,N_5931,N_5414);
or U6747 (N_6747,N_5212,N_5035);
and U6748 (N_6748,N_5647,N_5294);
nand U6749 (N_6749,N_5009,N_5421);
or U6750 (N_6750,N_5498,N_5654);
nor U6751 (N_6751,N_5286,N_5187);
and U6752 (N_6752,N_5805,N_5672);
and U6753 (N_6753,N_5188,N_5690);
nand U6754 (N_6754,N_5790,N_5829);
or U6755 (N_6755,N_5543,N_5137);
and U6756 (N_6756,N_5356,N_5827);
and U6757 (N_6757,N_5758,N_5436);
and U6758 (N_6758,N_5673,N_5501);
nor U6759 (N_6759,N_5442,N_5253);
nand U6760 (N_6760,N_5160,N_5112);
and U6761 (N_6761,N_5915,N_5048);
and U6762 (N_6762,N_5010,N_5134);
and U6763 (N_6763,N_5265,N_5585);
and U6764 (N_6764,N_5776,N_5848);
nand U6765 (N_6765,N_5640,N_5231);
or U6766 (N_6766,N_5744,N_5364);
and U6767 (N_6767,N_5683,N_5488);
nor U6768 (N_6768,N_5189,N_5361);
nand U6769 (N_6769,N_5450,N_5982);
nand U6770 (N_6770,N_5131,N_5251);
xor U6771 (N_6771,N_5338,N_5398);
nor U6772 (N_6772,N_5090,N_5341);
and U6773 (N_6773,N_5479,N_5190);
nand U6774 (N_6774,N_5333,N_5891);
and U6775 (N_6775,N_5861,N_5544);
or U6776 (N_6776,N_5052,N_5938);
nand U6777 (N_6777,N_5077,N_5055);
or U6778 (N_6778,N_5804,N_5119);
and U6779 (N_6779,N_5179,N_5479);
nand U6780 (N_6780,N_5936,N_5020);
and U6781 (N_6781,N_5119,N_5256);
or U6782 (N_6782,N_5958,N_5489);
and U6783 (N_6783,N_5292,N_5386);
nor U6784 (N_6784,N_5341,N_5140);
and U6785 (N_6785,N_5409,N_5954);
or U6786 (N_6786,N_5822,N_5879);
nand U6787 (N_6787,N_5499,N_5065);
and U6788 (N_6788,N_5742,N_5474);
and U6789 (N_6789,N_5277,N_5425);
or U6790 (N_6790,N_5492,N_5249);
nand U6791 (N_6791,N_5161,N_5745);
nand U6792 (N_6792,N_5668,N_5908);
nor U6793 (N_6793,N_5343,N_5623);
or U6794 (N_6794,N_5940,N_5936);
nand U6795 (N_6795,N_5202,N_5111);
nand U6796 (N_6796,N_5842,N_5477);
or U6797 (N_6797,N_5915,N_5466);
or U6798 (N_6798,N_5107,N_5559);
and U6799 (N_6799,N_5638,N_5657);
nor U6800 (N_6800,N_5351,N_5937);
nand U6801 (N_6801,N_5434,N_5404);
nor U6802 (N_6802,N_5107,N_5330);
or U6803 (N_6803,N_5019,N_5415);
nor U6804 (N_6804,N_5592,N_5970);
or U6805 (N_6805,N_5365,N_5256);
or U6806 (N_6806,N_5775,N_5837);
nand U6807 (N_6807,N_5482,N_5809);
and U6808 (N_6808,N_5003,N_5627);
nand U6809 (N_6809,N_5383,N_5528);
nand U6810 (N_6810,N_5250,N_5242);
or U6811 (N_6811,N_5615,N_5714);
or U6812 (N_6812,N_5577,N_5543);
nand U6813 (N_6813,N_5717,N_5314);
or U6814 (N_6814,N_5298,N_5363);
and U6815 (N_6815,N_5516,N_5305);
nand U6816 (N_6816,N_5076,N_5145);
and U6817 (N_6817,N_5260,N_5179);
or U6818 (N_6818,N_5390,N_5969);
nor U6819 (N_6819,N_5116,N_5964);
or U6820 (N_6820,N_5160,N_5866);
and U6821 (N_6821,N_5209,N_5039);
or U6822 (N_6822,N_5656,N_5014);
or U6823 (N_6823,N_5112,N_5550);
nor U6824 (N_6824,N_5610,N_5492);
or U6825 (N_6825,N_5682,N_5575);
or U6826 (N_6826,N_5367,N_5666);
nand U6827 (N_6827,N_5561,N_5319);
xnor U6828 (N_6828,N_5692,N_5143);
and U6829 (N_6829,N_5888,N_5683);
and U6830 (N_6830,N_5970,N_5544);
and U6831 (N_6831,N_5115,N_5372);
nor U6832 (N_6832,N_5035,N_5681);
or U6833 (N_6833,N_5605,N_5587);
or U6834 (N_6834,N_5355,N_5386);
nor U6835 (N_6835,N_5054,N_5809);
or U6836 (N_6836,N_5734,N_5976);
or U6837 (N_6837,N_5848,N_5947);
or U6838 (N_6838,N_5552,N_5284);
or U6839 (N_6839,N_5577,N_5915);
and U6840 (N_6840,N_5250,N_5284);
nor U6841 (N_6841,N_5207,N_5945);
and U6842 (N_6842,N_5429,N_5774);
nand U6843 (N_6843,N_5363,N_5479);
nand U6844 (N_6844,N_5952,N_5609);
nor U6845 (N_6845,N_5582,N_5438);
nand U6846 (N_6846,N_5725,N_5031);
or U6847 (N_6847,N_5275,N_5560);
or U6848 (N_6848,N_5180,N_5471);
nor U6849 (N_6849,N_5076,N_5098);
nor U6850 (N_6850,N_5848,N_5488);
and U6851 (N_6851,N_5056,N_5051);
nor U6852 (N_6852,N_5697,N_5294);
nand U6853 (N_6853,N_5142,N_5541);
or U6854 (N_6854,N_5734,N_5422);
nand U6855 (N_6855,N_5218,N_5157);
and U6856 (N_6856,N_5505,N_5561);
or U6857 (N_6857,N_5566,N_5095);
nand U6858 (N_6858,N_5300,N_5579);
nand U6859 (N_6859,N_5364,N_5370);
nor U6860 (N_6860,N_5493,N_5011);
and U6861 (N_6861,N_5560,N_5315);
or U6862 (N_6862,N_5155,N_5048);
and U6863 (N_6863,N_5395,N_5642);
and U6864 (N_6864,N_5004,N_5236);
or U6865 (N_6865,N_5106,N_5694);
and U6866 (N_6866,N_5067,N_5126);
nand U6867 (N_6867,N_5352,N_5204);
or U6868 (N_6868,N_5756,N_5548);
and U6869 (N_6869,N_5163,N_5144);
or U6870 (N_6870,N_5702,N_5610);
nand U6871 (N_6871,N_5946,N_5999);
nand U6872 (N_6872,N_5914,N_5129);
nor U6873 (N_6873,N_5966,N_5562);
nand U6874 (N_6874,N_5550,N_5191);
nor U6875 (N_6875,N_5306,N_5231);
nand U6876 (N_6876,N_5427,N_5636);
nand U6877 (N_6877,N_5122,N_5337);
nand U6878 (N_6878,N_5195,N_5058);
nor U6879 (N_6879,N_5010,N_5003);
xor U6880 (N_6880,N_5383,N_5004);
nand U6881 (N_6881,N_5911,N_5599);
and U6882 (N_6882,N_5702,N_5220);
and U6883 (N_6883,N_5060,N_5397);
or U6884 (N_6884,N_5326,N_5352);
or U6885 (N_6885,N_5731,N_5918);
nand U6886 (N_6886,N_5987,N_5710);
and U6887 (N_6887,N_5076,N_5215);
xor U6888 (N_6888,N_5826,N_5612);
or U6889 (N_6889,N_5424,N_5111);
nand U6890 (N_6890,N_5915,N_5922);
and U6891 (N_6891,N_5920,N_5889);
xnor U6892 (N_6892,N_5552,N_5873);
or U6893 (N_6893,N_5734,N_5489);
and U6894 (N_6894,N_5948,N_5145);
and U6895 (N_6895,N_5150,N_5197);
or U6896 (N_6896,N_5944,N_5241);
or U6897 (N_6897,N_5065,N_5610);
xnor U6898 (N_6898,N_5857,N_5151);
and U6899 (N_6899,N_5553,N_5740);
or U6900 (N_6900,N_5607,N_5846);
or U6901 (N_6901,N_5459,N_5880);
and U6902 (N_6902,N_5059,N_5775);
or U6903 (N_6903,N_5527,N_5233);
nor U6904 (N_6904,N_5004,N_5039);
or U6905 (N_6905,N_5920,N_5249);
and U6906 (N_6906,N_5534,N_5180);
or U6907 (N_6907,N_5925,N_5604);
nor U6908 (N_6908,N_5067,N_5265);
nand U6909 (N_6909,N_5947,N_5460);
nand U6910 (N_6910,N_5418,N_5189);
nand U6911 (N_6911,N_5569,N_5511);
or U6912 (N_6912,N_5880,N_5801);
and U6913 (N_6913,N_5637,N_5295);
or U6914 (N_6914,N_5750,N_5354);
and U6915 (N_6915,N_5711,N_5743);
xnor U6916 (N_6916,N_5935,N_5242);
or U6917 (N_6917,N_5869,N_5467);
nor U6918 (N_6918,N_5357,N_5186);
nand U6919 (N_6919,N_5339,N_5132);
or U6920 (N_6920,N_5019,N_5098);
or U6921 (N_6921,N_5545,N_5319);
nand U6922 (N_6922,N_5722,N_5365);
nand U6923 (N_6923,N_5957,N_5256);
or U6924 (N_6924,N_5837,N_5752);
and U6925 (N_6925,N_5925,N_5703);
nor U6926 (N_6926,N_5875,N_5594);
nor U6927 (N_6927,N_5661,N_5431);
and U6928 (N_6928,N_5112,N_5819);
or U6929 (N_6929,N_5273,N_5915);
nand U6930 (N_6930,N_5676,N_5078);
nand U6931 (N_6931,N_5848,N_5936);
and U6932 (N_6932,N_5786,N_5105);
or U6933 (N_6933,N_5589,N_5522);
and U6934 (N_6934,N_5936,N_5765);
nor U6935 (N_6935,N_5320,N_5810);
nor U6936 (N_6936,N_5297,N_5165);
nor U6937 (N_6937,N_5328,N_5387);
and U6938 (N_6938,N_5511,N_5782);
xor U6939 (N_6939,N_5381,N_5425);
nor U6940 (N_6940,N_5277,N_5790);
nor U6941 (N_6941,N_5003,N_5374);
and U6942 (N_6942,N_5121,N_5704);
or U6943 (N_6943,N_5497,N_5242);
nand U6944 (N_6944,N_5921,N_5217);
and U6945 (N_6945,N_5150,N_5476);
nand U6946 (N_6946,N_5413,N_5136);
xnor U6947 (N_6947,N_5180,N_5271);
and U6948 (N_6948,N_5957,N_5005);
or U6949 (N_6949,N_5156,N_5800);
xor U6950 (N_6950,N_5586,N_5821);
or U6951 (N_6951,N_5192,N_5437);
nor U6952 (N_6952,N_5444,N_5317);
and U6953 (N_6953,N_5531,N_5065);
nand U6954 (N_6954,N_5115,N_5172);
or U6955 (N_6955,N_5352,N_5809);
nand U6956 (N_6956,N_5252,N_5908);
or U6957 (N_6957,N_5370,N_5913);
or U6958 (N_6958,N_5969,N_5285);
or U6959 (N_6959,N_5282,N_5031);
or U6960 (N_6960,N_5848,N_5633);
nor U6961 (N_6961,N_5460,N_5101);
and U6962 (N_6962,N_5917,N_5197);
nor U6963 (N_6963,N_5234,N_5471);
nand U6964 (N_6964,N_5465,N_5194);
or U6965 (N_6965,N_5842,N_5522);
or U6966 (N_6966,N_5411,N_5421);
or U6967 (N_6967,N_5148,N_5210);
and U6968 (N_6968,N_5816,N_5349);
xor U6969 (N_6969,N_5156,N_5517);
nand U6970 (N_6970,N_5292,N_5381);
nand U6971 (N_6971,N_5468,N_5557);
nor U6972 (N_6972,N_5877,N_5260);
or U6973 (N_6973,N_5728,N_5215);
nor U6974 (N_6974,N_5696,N_5023);
and U6975 (N_6975,N_5088,N_5211);
nor U6976 (N_6976,N_5199,N_5146);
nand U6977 (N_6977,N_5633,N_5974);
or U6978 (N_6978,N_5482,N_5101);
and U6979 (N_6979,N_5072,N_5623);
nand U6980 (N_6980,N_5800,N_5279);
or U6981 (N_6981,N_5629,N_5472);
nor U6982 (N_6982,N_5315,N_5158);
and U6983 (N_6983,N_5397,N_5819);
or U6984 (N_6984,N_5332,N_5062);
nor U6985 (N_6985,N_5621,N_5878);
nand U6986 (N_6986,N_5669,N_5060);
or U6987 (N_6987,N_5730,N_5192);
nor U6988 (N_6988,N_5621,N_5971);
or U6989 (N_6989,N_5253,N_5794);
or U6990 (N_6990,N_5414,N_5881);
or U6991 (N_6991,N_5487,N_5985);
and U6992 (N_6992,N_5172,N_5120);
or U6993 (N_6993,N_5763,N_5009);
or U6994 (N_6994,N_5122,N_5995);
nand U6995 (N_6995,N_5606,N_5751);
nand U6996 (N_6996,N_5543,N_5651);
or U6997 (N_6997,N_5732,N_5962);
and U6998 (N_6998,N_5643,N_5309);
or U6999 (N_6999,N_5648,N_5859);
nand U7000 (N_7000,N_6067,N_6008);
or U7001 (N_7001,N_6517,N_6194);
xor U7002 (N_7002,N_6559,N_6180);
or U7003 (N_7003,N_6524,N_6701);
nand U7004 (N_7004,N_6987,N_6989);
nand U7005 (N_7005,N_6950,N_6567);
or U7006 (N_7006,N_6032,N_6035);
and U7007 (N_7007,N_6676,N_6202);
nor U7008 (N_7008,N_6974,N_6129);
or U7009 (N_7009,N_6266,N_6314);
nor U7010 (N_7010,N_6907,N_6412);
nor U7011 (N_7011,N_6561,N_6729);
nand U7012 (N_7012,N_6673,N_6714);
nand U7013 (N_7013,N_6077,N_6807);
nor U7014 (N_7014,N_6811,N_6769);
or U7015 (N_7015,N_6912,N_6384);
and U7016 (N_7016,N_6571,N_6763);
nor U7017 (N_7017,N_6473,N_6270);
nand U7018 (N_7018,N_6455,N_6066);
and U7019 (N_7019,N_6297,N_6084);
and U7020 (N_7020,N_6102,N_6363);
and U7021 (N_7021,N_6875,N_6700);
nand U7022 (N_7022,N_6954,N_6512);
nor U7023 (N_7023,N_6014,N_6565);
nand U7024 (N_7024,N_6868,N_6450);
xnor U7025 (N_7025,N_6169,N_6490);
nor U7026 (N_7026,N_6147,N_6534);
and U7027 (N_7027,N_6082,N_6728);
and U7028 (N_7028,N_6911,N_6173);
or U7029 (N_7029,N_6337,N_6731);
nor U7030 (N_7030,N_6167,N_6108);
nor U7031 (N_7031,N_6634,N_6681);
and U7032 (N_7032,N_6364,N_6243);
and U7033 (N_7033,N_6680,N_6047);
and U7034 (N_7034,N_6828,N_6674);
and U7035 (N_7035,N_6981,N_6481);
nor U7036 (N_7036,N_6255,N_6426);
nor U7037 (N_7037,N_6837,N_6573);
nor U7038 (N_7038,N_6550,N_6887);
or U7039 (N_7039,N_6103,N_6521);
nor U7040 (N_7040,N_6187,N_6088);
nor U7041 (N_7041,N_6182,N_6253);
nand U7042 (N_7042,N_6119,N_6752);
or U7043 (N_7043,N_6651,N_6663);
and U7044 (N_7044,N_6283,N_6738);
and U7045 (N_7045,N_6223,N_6895);
and U7046 (N_7046,N_6801,N_6668);
or U7047 (N_7047,N_6348,N_6598);
nand U7048 (N_7048,N_6849,N_6296);
and U7049 (N_7049,N_6351,N_6403);
and U7050 (N_7050,N_6593,N_6639);
nor U7051 (N_7051,N_6896,N_6446);
and U7052 (N_7052,N_6536,N_6300);
nor U7053 (N_7053,N_6137,N_6341);
nand U7054 (N_7054,N_6355,N_6252);
or U7055 (N_7055,N_6349,N_6855);
nor U7056 (N_7056,N_6009,N_6975);
nor U7057 (N_7057,N_6196,N_6206);
and U7058 (N_7058,N_6929,N_6482);
or U7059 (N_7059,N_6884,N_6145);
nand U7060 (N_7060,N_6756,N_6284);
nand U7061 (N_7061,N_6707,N_6564);
or U7062 (N_7062,N_6961,N_6873);
nor U7063 (N_7063,N_6537,N_6215);
or U7064 (N_7064,N_6659,N_6815);
nand U7065 (N_7065,N_6516,N_6079);
or U7066 (N_7066,N_6051,N_6140);
and U7067 (N_7067,N_6267,N_6489);
and U7068 (N_7068,N_6002,N_6375);
nand U7069 (N_7069,N_6785,N_6149);
nand U7070 (N_7070,N_6466,N_6594);
nor U7071 (N_7071,N_6148,N_6393);
or U7072 (N_7072,N_6336,N_6136);
or U7073 (N_7073,N_6445,N_6927);
nand U7074 (N_7074,N_6039,N_6957);
and U7075 (N_7075,N_6750,N_6198);
and U7076 (N_7076,N_6685,N_6759);
nor U7077 (N_7077,N_6784,N_6313);
and U7078 (N_7078,N_6236,N_6599);
and U7079 (N_7079,N_6839,N_6498);
and U7080 (N_7080,N_6309,N_6275);
and U7081 (N_7081,N_6487,N_6919);
or U7082 (N_7082,N_6584,N_6076);
nor U7083 (N_7083,N_6922,N_6062);
nor U7084 (N_7084,N_6812,N_6292);
or U7085 (N_7085,N_6749,N_6859);
nand U7086 (N_7086,N_6802,N_6469);
and U7087 (N_7087,N_6143,N_6387);
and U7088 (N_7088,N_6710,N_6709);
nand U7089 (N_7089,N_6626,N_6118);
or U7090 (N_7090,N_6744,N_6353);
nor U7091 (N_7091,N_6247,N_6982);
nand U7092 (N_7092,N_6753,N_6627);
nand U7093 (N_7093,N_6228,N_6451);
nor U7094 (N_7094,N_6692,N_6789);
and U7095 (N_7095,N_6279,N_6117);
nand U7096 (N_7096,N_6290,N_6834);
and U7097 (N_7097,N_6135,N_6937);
and U7098 (N_7098,N_6658,N_6159);
nand U7099 (N_7099,N_6605,N_6382);
and U7100 (N_7100,N_6074,N_6966);
and U7101 (N_7101,N_6230,N_6029);
and U7102 (N_7102,N_6867,N_6238);
xor U7103 (N_7103,N_6747,N_6513);
nand U7104 (N_7104,N_6732,N_6210);
and U7105 (N_7105,N_6531,N_6320);
nand U7106 (N_7106,N_6872,N_6398);
or U7107 (N_7107,N_6505,N_6156);
or U7108 (N_7108,N_6146,N_6501);
nand U7109 (N_7109,N_6056,N_6303);
and U7110 (N_7110,N_6994,N_6086);
nor U7111 (N_7111,N_6261,N_6092);
and U7112 (N_7112,N_6318,N_6894);
nand U7113 (N_7113,N_6617,N_6064);
nand U7114 (N_7114,N_6171,N_6791);
nand U7115 (N_7115,N_6237,N_6461);
or U7116 (N_7116,N_6754,N_6389);
and U7117 (N_7117,N_6556,N_6025);
and U7118 (N_7118,N_6181,N_6995);
or U7119 (N_7119,N_6444,N_6826);
nor U7120 (N_7120,N_6484,N_6037);
nand U7121 (N_7121,N_6905,N_6452);
or U7122 (N_7122,N_6890,N_6190);
or U7123 (N_7123,N_6971,N_6881);
nand U7124 (N_7124,N_6397,N_6773);
xnor U7125 (N_7125,N_6504,N_6502);
and U7126 (N_7126,N_6439,N_6538);
and U7127 (N_7127,N_6845,N_6876);
nand U7128 (N_7128,N_6376,N_6265);
and U7129 (N_7129,N_6115,N_6603);
and U7130 (N_7130,N_6648,N_6525);
nand U7131 (N_7131,N_6581,N_6254);
nand U7132 (N_7132,N_6740,N_6174);
nand U7133 (N_7133,N_6959,N_6160);
nand U7134 (N_7134,N_6511,N_6916);
nand U7135 (N_7135,N_6438,N_6274);
and U7136 (N_7136,N_6128,N_6479);
nor U7137 (N_7137,N_6507,N_6343);
nor U7138 (N_7138,N_6431,N_6360);
nand U7139 (N_7139,N_6219,N_6184);
nand U7140 (N_7140,N_6533,N_6189);
and U7141 (N_7141,N_6977,N_6662);
and U7142 (N_7142,N_6411,N_6690);
nor U7143 (N_7143,N_6151,N_6378);
nor U7144 (N_7144,N_6790,N_6558);
or U7145 (N_7145,N_6483,N_6606);
nand U7146 (N_7146,N_6608,N_6535);
and U7147 (N_7147,N_6316,N_6224);
nor U7148 (N_7148,N_6724,N_6004);
or U7149 (N_7149,N_6854,N_6509);
nor U7150 (N_7150,N_6453,N_6960);
or U7151 (N_7151,N_6518,N_6979);
and U7152 (N_7152,N_6209,N_6545);
nor U7153 (N_7153,N_6930,N_6847);
xor U7154 (N_7154,N_6891,N_6015);
nand U7155 (N_7155,N_6671,N_6780);
nor U7156 (N_7156,N_6688,N_6327);
nand U7157 (N_7157,N_6460,N_6494);
and U7158 (N_7158,N_6613,N_6414);
or U7159 (N_7159,N_6947,N_6138);
or U7160 (N_7160,N_6248,N_6779);
nand U7161 (N_7161,N_6222,N_6689);
nand U7162 (N_7162,N_6618,N_6861);
or U7163 (N_7163,N_6402,N_6809);
and U7164 (N_7164,N_6063,N_6214);
nand U7165 (N_7165,N_6260,N_6249);
or U7166 (N_7166,N_6120,N_6549);
and U7167 (N_7167,N_6114,N_6670);
and U7168 (N_7168,N_6592,N_6131);
or U7169 (N_7169,N_6672,N_6001);
and U7170 (N_7170,N_6139,N_6677);
nor U7171 (N_7171,N_6038,N_6217);
or U7172 (N_7172,N_6739,N_6976);
nor U7173 (N_7173,N_6301,N_6044);
nor U7174 (N_7174,N_6607,N_6711);
nand U7175 (N_7175,N_6906,N_6175);
or U7176 (N_7176,N_6795,N_6078);
and U7177 (N_7177,N_6956,N_6095);
and U7178 (N_7178,N_6955,N_6863);
and U7179 (N_7179,N_6529,N_6027);
and U7180 (N_7180,N_6016,N_6213);
xnor U7181 (N_7181,N_6322,N_6687);
or U7182 (N_7182,N_6883,N_6649);
nor U7183 (N_7183,N_6186,N_6344);
nor U7184 (N_7184,N_6620,N_6013);
or U7185 (N_7185,N_6601,N_6069);
nor U7186 (N_7186,N_6827,N_6177);
nor U7187 (N_7187,N_6144,N_6201);
and U7188 (N_7188,N_6429,N_6176);
nand U7189 (N_7189,N_6087,N_6269);
and U7190 (N_7190,N_6557,N_6624);
or U7191 (N_7191,N_6262,N_6416);
and U7192 (N_7192,N_6050,N_6359);
and U7193 (N_7193,N_6612,N_6715);
nor U7194 (N_7194,N_6686,N_6619);
or U7195 (N_7195,N_6819,N_6242);
and U7196 (N_7196,N_6589,N_6679);
or U7197 (N_7197,N_6031,N_6797);
and U7198 (N_7198,N_6057,N_6985);
nand U7199 (N_7199,N_6727,N_6833);
nand U7200 (N_7200,N_6365,N_6734);
or U7201 (N_7201,N_6474,N_6562);
nand U7202 (N_7202,N_6582,N_6106);
nand U7203 (N_7203,N_6207,N_6596);
nand U7204 (N_7204,N_6992,N_6287);
nand U7205 (N_7205,N_6105,N_6823);
and U7206 (N_7206,N_6602,N_6133);
or U7207 (N_7207,N_6852,N_6900);
nor U7208 (N_7208,N_6808,N_6475);
nand U7209 (N_7209,N_6478,N_6817);
nand U7210 (N_7210,N_6941,N_6913);
and U7211 (N_7211,N_6054,N_6257);
and U7212 (N_7212,N_6901,N_6288);
xor U7213 (N_7213,N_6241,N_6229);
xor U7214 (N_7214,N_6476,N_6585);
xor U7215 (N_7215,N_6408,N_6081);
nor U7216 (N_7216,N_6286,N_6488);
nand U7217 (N_7217,N_6271,N_6616);
or U7218 (N_7218,N_6704,N_6865);
nor U7219 (N_7219,N_6523,N_6570);
and U7220 (N_7220,N_6306,N_6419);
nand U7221 (N_7221,N_6011,N_6141);
nand U7222 (N_7222,N_6633,N_6527);
or U7223 (N_7223,N_6691,N_6331);
or U7224 (N_7224,N_6888,N_6400);
nor U7225 (N_7225,N_6595,N_6864);
nor U7226 (N_7226,N_6024,N_6540);
or U7227 (N_7227,N_6354,N_6324);
or U7228 (N_7228,N_6276,N_6708);
nor U7229 (N_7229,N_6281,N_6574);
and U7230 (N_7230,N_6666,N_6698);
or U7231 (N_7231,N_6065,N_6792);
or U7232 (N_7232,N_6699,N_6153);
xnor U7233 (N_7233,N_6127,N_6178);
and U7234 (N_7234,N_6736,N_6205);
nand U7235 (N_7235,N_6716,N_6990);
nor U7236 (N_7236,N_6718,N_6409);
nor U7237 (N_7237,N_6667,N_6437);
or U7238 (N_7238,N_6816,N_6334);
nor U7239 (N_7239,N_6315,N_6107);
and U7240 (N_7240,N_6208,N_6577);
nor U7241 (N_7241,N_6635,N_6280);
nand U7242 (N_7242,N_6161,N_6273);
nor U7243 (N_7243,N_6939,N_6305);
nor U7244 (N_7244,N_6477,N_6706);
or U7245 (N_7245,N_6183,N_6949);
or U7246 (N_7246,N_6499,N_6289);
xor U7247 (N_7247,N_6796,N_6328);
and U7248 (N_7248,N_6578,N_6435);
nor U7249 (N_7249,N_6326,N_6164);
nand U7250 (N_7250,N_6434,N_6374);
nand U7251 (N_7251,N_6820,N_6218);
and U7252 (N_7252,N_6394,N_6231);
and U7253 (N_7253,N_6436,N_6737);
and U7254 (N_7254,N_6333,N_6329);
or U7255 (N_7255,N_6193,N_6842);
or U7256 (N_7256,N_6017,N_6251);
or U7257 (N_7257,N_6299,N_6415);
nor U7258 (N_7258,N_6642,N_6925);
or U7259 (N_7259,N_6857,N_6526);
and U7260 (N_7260,N_6999,N_6480);
nor U7261 (N_7261,N_6089,N_6496);
nand U7262 (N_7262,N_6630,N_6302);
or U7263 (N_7263,N_6774,N_6405);
and U7264 (N_7264,N_6225,N_6358);
nand U7265 (N_7265,N_6554,N_6310);
and U7266 (N_7266,N_6410,N_6220);
and U7267 (N_7267,N_6390,N_6682);
or U7268 (N_7268,N_6053,N_6342);
and U7269 (N_7269,N_6885,N_6391);
nand U7270 (N_7270,N_6307,N_6669);
and U7271 (N_7271,N_6972,N_6661);
or U7272 (N_7272,N_6503,N_6413);
nor U7273 (N_7273,N_6468,N_6720);
nor U7274 (N_7274,N_6212,N_6368);
and U7275 (N_7275,N_6377,N_6892);
or U7276 (N_7276,N_6258,N_6803);
nor U7277 (N_7277,N_6694,N_6059);
nand U7278 (N_7278,N_6735,N_6386);
nor U7279 (N_7279,N_6551,N_6030);
or U7280 (N_7280,N_6848,N_6235);
or U7281 (N_7281,N_6000,N_6519);
nand U7282 (N_7282,N_6991,N_6998);
nand U7283 (N_7283,N_6404,N_6109);
or U7284 (N_7284,N_6841,N_6430);
or U7285 (N_7285,N_6070,N_6041);
and U7286 (N_7286,N_6495,N_6471);
nand U7287 (N_7287,N_6268,N_6185);
nor U7288 (N_7288,N_6396,N_6340);
nand U7289 (N_7289,N_6965,N_6958);
nand U7290 (N_7290,N_6683,N_6111);
nor U7291 (N_7291,N_6472,N_6788);
nor U7292 (N_7292,N_6319,N_6866);
and U7293 (N_7293,N_6246,N_6170);
nor U7294 (N_7294,N_6625,N_6058);
and U7295 (N_7295,N_6508,N_6110);
nand U7296 (N_7296,N_6968,N_6264);
and U7297 (N_7297,N_6874,N_6576);
nand U7298 (N_7298,N_6610,N_6832);
or U7299 (N_7299,N_6946,N_6433);
and U7300 (N_7300,N_6870,N_6878);
and U7301 (N_7301,N_6760,N_6915);
or U7302 (N_7302,N_6643,N_6463);
nor U7303 (N_7303,N_6200,N_6285);
nor U7304 (N_7304,N_6500,N_6902);
nand U7305 (N_7305,N_6799,N_6940);
nand U7306 (N_7306,N_6068,N_6563);
xnor U7307 (N_7307,N_6356,N_6745);
nand U7308 (N_7308,N_6132,N_6893);
nor U7309 (N_7309,N_6743,N_6628);
nor U7310 (N_7310,N_6221,N_6497);
or U7311 (N_7311,N_6964,N_6591);
and U7312 (N_7312,N_6928,N_6104);
xor U7313 (N_7313,N_6684,N_6843);
and U7314 (N_7314,N_6712,N_6810);
or U7315 (N_7315,N_6934,N_6530);
nand U7316 (N_7316,N_6470,N_6245);
nand U7317 (N_7317,N_6012,N_6637);
or U7318 (N_7318,N_6098,N_6124);
nor U7319 (N_7319,N_6073,N_6840);
and U7320 (N_7320,N_6350,N_6112);
nor U7321 (N_7321,N_6385,N_6997);
nand U7322 (N_7322,N_6036,N_6005);
or U7323 (N_7323,N_6232,N_6721);
nor U7324 (N_7324,N_6751,N_6432);
nor U7325 (N_7325,N_6742,N_6204);
and U7326 (N_7326,N_6575,N_6986);
or U7327 (N_7327,N_6898,N_6652);
or U7328 (N_7328,N_6988,N_6755);
xor U7329 (N_7329,N_6800,N_6304);
nor U7330 (N_7330,N_6456,N_6019);
nand U7331 (N_7331,N_6548,N_6325);
and U7332 (N_7332,N_6963,N_6099);
or U7333 (N_7333,N_6045,N_6862);
and U7334 (N_7334,N_6851,N_6142);
nor U7335 (N_7335,N_6553,N_6910);
nor U7336 (N_7336,N_6380,N_6983);
and U7337 (N_7337,N_6440,N_6846);
nor U7338 (N_7338,N_6783,N_6165);
or U7339 (N_7339,N_6263,N_6100);
nor U7340 (N_7340,N_6226,N_6973);
nor U7341 (N_7341,N_6122,N_6312);
nand U7342 (N_7342,N_6407,N_6675);
nor U7343 (N_7343,N_6332,N_6043);
nand U7344 (N_7344,N_6935,N_6933);
nand U7345 (N_7345,N_6250,N_6822);
and U7346 (N_7346,N_6869,N_6899);
or U7347 (N_7347,N_6805,N_6458);
nand U7348 (N_7348,N_6943,N_6914);
or U7349 (N_7349,N_6980,N_6395);
nand U7350 (N_7350,N_6049,N_6379);
or U7351 (N_7351,N_6696,N_6770);
and U7352 (N_7352,N_6422,N_6392);
nand U7353 (N_7353,N_6028,N_6748);
nor U7354 (N_7354,N_6560,N_6726);
or U7355 (N_7355,N_6654,N_6665);
and U7356 (N_7356,N_6539,N_6007);
or U7357 (N_7357,N_6814,N_6920);
or U7358 (N_7358,N_6631,N_6566);
and U7359 (N_7359,N_6345,N_6609);
or U7360 (N_7360,N_6162,N_6776);
nor U7361 (N_7361,N_6621,N_6794);
nor U7362 (N_7362,N_6993,N_6424);
nor U7363 (N_7363,N_6762,N_6653);
or U7364 (N_7364,N_6629,N_6777);
and U7365 (N_7365,N_6256,N_6042);
or U7366 (N_7366,N_6768,N_6003);
and U7367 (N_7367,N_6234,N_6335);
or U7368 (N_7368,N_6447,N_6542);
or U7369 (N_7369,N_6775,N_6967);
nand U7370 (N_7370,N_6418,N_6615);
xor U7371 (N_7371,N_6725,N_6787);
nand U7372 (N_7372,N_6216,N_6931);
nand U7373 (N_7373,N_6746,N_6824);
and U7374 (N_7374,N_6702,N_6641);
and U7375 (N_7375,N_6188,N_6373);
or U7376 (N_7376,N_6741,N_6462);
xor U7377 (N_7377,N_6083,N_6157);
xor U7378 (N_7378,N_6798,N_6457);
or U7379 (N_7379,N_6932,N_6614);
nand U7380 (N_7380,N_6158,N_6293);
nand U7381 (N_7381,N_6034,N_6623);
nor U7382 (N_7382,N_6442,N_6061);
or U7383 (N_7383,N_6636,N_6579);
nor U7384 (N_7384,N_6544,N_6514);
nand U7385 (N_7385,N_6239,N_6882);
nor U7386 (N_7386,N_6090,N_6656);
nand U7387 (N_7387,N_6717,N_6569);
nor U7388 (N_7388,N_6272,N_6962);
nand U7389 (N_7389,N_6425,N_6448);
nand U7390 (N_7390,N_6818,N_6485);
nor U7391 (N_7391,N_6339,N_6317);
nor U7392 (N_7392,N_6722,N_6705);
and U7393 (N_7393,N_6370,N_6172);
or U7394 (N_7394,N_6660,N_6401);
and U7395 (N_7395,N_6428,N_6825);
and U7396 (N_7396,N_6046,N_6199);
nand U7397 (N_7397,N_6361,N_6733);
nor U7398 (N_7398,N_6113,N_6203);
nand U7399 (N_7399,N_6179,N_6277);
nor U7400 (N_7400,N_6568,N_6121);
nand U7401 (N_7401,N_6730,N_6022);
or U7402 (N_7402,N_6006,N_6420);
or U7403 (N_7403,N_6033,N_6520);
nor U7404 (N_7404,N_6192,N_6926);
nand U7405 (N_7405,N_6765,N_6723);
and U7406 (N_7406,N_6650,N_6657);
nand U7407 (N_7407,N_6018,N_6506);
nor U7408 (N_7408,N_6093,N_6771);
nor U7409 (N_7409,N_6023,N_6294);
and U7410 (N_7410,N_6055,N_6311);
or U7411 (N_7411,N_6942,N_6917);
nor U7412 (N_7412,N_6091,N_6541);
nand U7413 (N_7413,N_6493,N_6330);
nand U7414 (N_7414,N_6948,N_6632);
and U7415 (N_7415,N_6758,N_6152);
nor U7416 (N_7416,N_6622,N_6010);
nand U7417 (N_7417,N_6323,N_6052);
nand U7418 (N_7418,N_6996,N_6858);
or U7419 (N_7419,N_6879,N_6719);
and U7420 (N_7420,N_6532,N_6836);
and U7421 (N_7421,N_6443,N_6590);
nor U7422 (N_7422,N_6640,N_6647);
or U7423 (N_7423,N_6060,N_6821);
nand U7424 (N_7424,N_6697,N_6655);
or U7425 (N_7425,N_6889,N_6381);
nor U7426 (N_7426,N_6969,N_6600);
or U7427 (N_7427,N_6597,N_6587);
or U7428 (N_7428,N_6150,N_6369);
or U7429 (N_7429,N_6543,N_6282);
or U7430 (N_7430,N_6644,N_6693);
and U7431 (N_7431,N_6829,N_6604);
and U7432 (N_7432,N_6786,N_6951);
nor U7433 (N_7433,N_6850,N_6371);
or U7434 (N_7434,N_6772,N_6080);
or U7435 (N_7435,N_6454,N_6778);
or U7436 (N_7436,N_6586,N_6588);
or U7437 (N_7437,N_6130,N_6767);
nand U7438 (N_7438,N_6844,N_6880);
or U7439 (N_7439,N_6338,N_6921);
nand U7440 (N_7440,N_6166,N_6075);
and U7441 (N_7441,N_6026,N_6321);
nand U7442 (N_7442,N_6347,N_6126);
or U7443 (N_7443,N_6191,N_6945);
nand U7444 (N_7444,N_6465,N_6781);
and U7445 (N_7445,N_6555,N_6154);
nand U7446 (N_7446,N_6766,N_6295);
nand U7447 (N_7447,N_6486,N_6804);
nand U7448 (N_7448,N_6464,N_6163);
or U7449 (N_7449,N_6835,N_6871);
or U7450 (N_7450,N_6886,N_6406);
or U7451 (N_7451,N_6831,N_6938);
or U7452 (N_7452,N_6646,N_6853);
or U7453 (N_7453,N_6491,N_6399);
nor U7454 (N_7454,N_6678,N_6291);
or U7455 (N_7455,N_6233,N_6757);
nor U7456 (N_7456,N_6155,N_6388);
and U7457 (N_7457,N_6713,N_6492);
nor U7458 (N_7458,N_6952,N_6924);
and U7459 (N_7459,N_6793,N_6909);
and U7460 (N_7460,N_6197,N_6423);
nor U7461 (N_7461,N_6580,N_6782);
nor U7462 (N_7462,N_6510,N_6528);
and U7463 (N_7463,N_6071,N_6101);
or U7464 (N_7464,N_6427,N_6908);
and U7465 (N_7465,N_6125,N_6904);
and U7466 (N_7466,N_6813,N_6923);
or U7467 (N_7467,N_6020,N_6021);
or U7468 (N_7468,N_6383,N_6944);
and U7469 (N_7469,N_6695,N_6522);
and U7470 (N_7470,N_6278,N_6372);
nor U7471 (N_7471,N_6195,N_6259);
or U7472 (N_7472,N_6352,N_6308);
and U7473 (N_7473,N_6877,N_6638);
and U7474 (N_7474,N_6048,N_6362);
or U7475 (N_7475,N_6227,N_6583);
or U7476 (N_7476,N_6134,N_6123);
or U7477 (N_7477,N_6552,N_6918);
and U7478 (N_7478,N_6547,N_6357);
nand U7479 (N_7479,N_6094,N_6449);
nand U7480 (N_7480,N_6040,N_6703);
nand U7481 (N_7481,N_6645,N_6572);
or U7482 (N_7482,N_6515,N_6467);
nor U7483 (N_7483,N_6085,N_6096);
and U7484 (N_7484,N_6546,N_6459);
nand U7485 (N_7485,N_6970,N_6838);
nand U7486 (N_7486,N_6244,N_6097);
and U7487 (N_7487,N_6168,N_6417);
or U7488 (N_7488,N_6367,N_6953);
or U7489 (N_7489,N_6116,N_6366);
nand U7490 (N_7490,N_6346,N_6240);
nor U7491 (N_7491,N_6441,N_6897);
xor U7492 (N_7492,N_6903,N_6830);
and U7493 (N_7493,N_6421,N_6984);
or U7494 (N_7494,N_6211,N_6856);
and U7495 (N_7495,N_6860,N_6978);
or U7496 (N_7496,N_6664,N_6936);
or U7497 (N_7497,N_6072,N_6764);
and U7498 (N_7498,N_6761,N_6611);
or U7499 (N_7499,N_6806,N_6298);
and U7500 (N_7500,N_6859,N_6033);
or U7501 (N_7501,N_6043,N_6046);
and U7502 (N_7502,N_6878,N_6537);
or U7503 (N_7503,N_6633,N_6224);
and U7504 (N_7504,N_6362,N_6149);
nand U7505 (N_7505,N_6264,N_6985);
xor U7506 (N_7506,N_6351,N_6649);
nand U7507 (N_7507,N_6822,N_6031);
and U7508 (N_7508,N_6245,N_6619);
or U7509 (N_7509,N_6032,N_6199);
or U7510 (N_7510,N_6915,N_6526);
nand U7511 (N_7511,N_6994,N_6325);
nand U7512 (N_7512,N_6779,N_6945);
and U7513 (N_7513,N_6497,N_6760);
nand U7514 (N_7514,N_6242,N_6007);
nor U7515 (N_7515,N_6946,N_6842);
and U7516 (N_7516,N_6732,N_6862);
and U7517 (N_7517,N_6584,N_6857);
xnor U7518 (N_7518,N_6662,N_6669);
xnor U7519 (N_7519,N_6855,N_6433);
nor U7520 (N_7520,N_6247,N_6448);
and U7521 (N_7521,N_6193,N_6074);
or U7522 (N_7522,N_6710,N_6033);
and U7523 (N_7523,N_6006,N_6458);
or U7524 (N_7524,N_6789,N_6729);
and U7525 (N_7525,N_6549,N_6687);
nor U7526 (N_7526,N_6112,N_6577);
or U7527 (N_7527,N_6630,N_6649);
nand U7528 (N_7528,N_6402,N_6593);
nand U7529 (N_7529,N_6961,N_6321);
nand U7530 (N_7530,N_6306,N_6784);
or U7531 (N_7531,N_6570,N_6674);
or U7532 (N_7532,N_6454,N_6590);
or U7533 (N_7533,N_6556,N_6437);
nor U7534 (N_7534,N_6049,N_6796);
or U7535 (N_7535,N_6426,N_6805);
or U7536 (N_7536,N_6383,N_6284);
and U7537 (N_7537,N_6470,N_6272);
nand U7538 (N_7538,N_6936,N_6204);
nor U7539 (N_7539,N_6984,N_6000);
and U7540 (N_7540,N_6717,N_6444);
nor U7541 (N_7541,N_6028,N_6212);
and U7542 (N_7542,N_6430,N_6339);
or U7543 (N_7543,N_6143,N_6471);
nand U7544 (N_7544,N_6773,N_6019);
nand U7545 (N_7545,N_6846,N_6635);
and U7546 (N_7546,N_6422,N_6860);
nor U7547 (N_7547,N_6743,N_6271);
nand U7548 (N_7548,N_6310,N_6285);
or U7549 (N_7549,N_6361,N_6565);
nor U7550 (N_7550,N_6464,N_6525);
nand U7551 (N_7551,N_6786,N_6533);
and U7552 (N_7552,N_6712,N_6374);
nand U7553 (N_7553,N_6407,N_6672);
or U7554 (N_7554,N_6804,N_6659);
nor U7555 (N_7555,N_6465,N_6733);
nand U7556 (N_7556,N_6882,N_6862);
and U7557 (N_7557,N_6625,N_6466);
nand U7558 (N_7558,N_6469,N_6720);
nor U7559 (N_7559,N_6168,N_6904);
nor U7560 (N_7560,N_6137,N_6511);
nand U7561 (N_7561,N_6395,N_6526);
nor U7562 (N_7562,N_6345,N_6451);
or U7563 (N_7563,N_6044,N_6067);
and U7564 (N_7564,N_6172,N_6420);
and U7565 (N_7565,N_6239,N_6987);
nand U7566 (N_7566,N_6209,N_6310);
and U7567 (N_7567,N_6887,N_6060);
nor U7568 (N_7568,N_6617,N_6194);
and U7569 (N_7569,N_6647,N_6420);
nand U7570 (N_7570,N_6682,N_6246);
or U7571 (N_7571,N_6190,N_6543);
and U7572 (N_7572,N_6994,N_6343);
nand U7573 (N_7573,N_6524,N_6811);
or U7574 (N_7574,N_6562,N_6844);
nor U7575 (N_7575,N_6770,N_6860);
and U7576 (N_7576,N_6039,N_6162);
or U7577 (N_7577,N_6748,N_6969);
nor U7578 (N_7578,N_6313,N_6188);
nor U7579 (N_7579,N_6119,N_6376);
or U7580 (N_7580,N_6507,N_6457);
nand U7581 (N_7581,N_6063,N_6458);
and U7582 (N_7582,N_6238,N_6918);
nand U7583 (N_7583,N_6457,N_6499);
nor U7584 (N_7584,N_6804,N_6339);
or U7585 (N_7585,N_6017,N_6342);
or U7586 (N_7586,N_6979,N_6140);
nor U7587 (N_7587,N_6480,N_6621);
and U7588 (N_7588,N_6272,N_6017);
nand U7589 (N_7589,N_6717,N_6740);
nand U7590 (N_7590,N_6173,N_6053);
or U7591 (N_7591,N_6969,N_6060);
or U7592 (N_7592,N_6541,N_6675);
or U7593 (N_7593,N_6401,N_6804);
nor U7594 (N_7594,N_6951,N_6906);
nor U7595 (N_7595,N_6089,N_6769);
nor U7596 (N_7596,N_6031,N_6991);
or U7597 (N_7597,N_6772,N_6765);
nor U7598 (N_7598,N_6485,N_6450);
nor U7599 (N_7599,N_6534,N_6755);
nor U7600 (N_7600,N_6099,N_6555);
nand U7601 (N_7601,N_6157,N_6448);
and U7602 (N_7602,N_6491,N_6245);
nor U7603 (N_7603,N_6891,N_6706);
nand U7604 (N_7604,N_6342,N_6341);
and U7605 (N_7605,N_6180,N_6723);
and U7606 (N_7606,N_6029,N_6207);
and U7607 (N_7607,N_6752,N_6543);
nand U7608 (N_7608,N_6975,N_6389);
or U7609 (N_7609,N_6880,N_6189);
nor U7610 (N_7610,N_6056,N_6349);
or U7611 (N_7611,N_6750,N_6460);
and U7612 (N_7612,N_6057,N_6404);
nand U7613 (N_7613,N_6982,N_6058);
and U7614 (N_7614,N_6024,N_6104);
nor U7615 (N_7615,N_6833,N_6466);
nand U7616 (N_7616,N_6239,N_6251);
and U7617 (N_7617,N_6618,N_6819);
or U7618 (N_7618,N_6150,N_6522);
nand U7619 (N_7619,N_6752,N_6737);
or U7620 (N_7620,N_6235,N_6445);
nor U7621 (N_7621,N_6383,N_6744);
and U7622 (N_7622,N_6990,N_6660);
nor U7623 (N_7623,N_6099,N_6875);
nand U7624 (N_7624,N_6004,N_6809);
xor U7625 (N_7625,N_6054,N_6392);
and U7626 (N_7626,N_6031,N_6033);
xnor U7627 (N_7627,N_6275,N_6990);
nand U7628 (N_7628,N_6911,N_6854);
nor U7629 (N_7629,N_6583,N_6832);
or U7630 (N_7630,N_6724,N_6921);
nor U7631 (N_7631,N_6533,N_6017);
nand U7632 (N_7632,N_6363,N_6544);
or U7633 (N_7633,N_6362,N_6988);
nor U7634 (N_7634,N_6238,N_6630);
nor U7635 (N_7635,N_6053,N_6326);
xnor U7636 (N_7636,N_6106,N_6149);
and U7637 (N_7637,N_6557,N_6443);
xor U7638 (N_7638,N_6279,N_6669);
nor U7639 (N_7639,N_6297,N_6201);
or U7640 (N_7640,N_6003,N_6540);
nor U7641 (N_7641,N_6654,N_6109);
nand U7642 (N_7642,N_6941,N_6374);
or U7643 (N_7643,N_6152,N_6768);
nand U7644 (N_7644,N_6598,N_6724);
or U7645 (N_7645,N_6608,N_6639);
or U7646 (N_7646,N_6614,N_6489);
nand U7647 (N_7647,N_6438,N_6734);
or U7648 (N_7648,N_6320,N_6126);
and U7649 (N_7649,N_6792,N_6918);
nor U7650 (N_7650,N_6613,N_6082);
or U7651 (N_7651,N_6273,N_6048);
nor U7652 (N_7652,N_6526,N_6469);
nand U7653 (N_7653,N_6502,N_6036);
and U7654 (N_7654,N_6533,N_6724);
nand U7655 (N_7655,N_6584,N_6154);
and U7656 (N_7656,N_6535,N_6778);
nand U7657 (N_7657,N_6440,N_6952);
nor U7658 (N_7658,N_6686,N_6156);
nand U7659 (N_7659,N_6177,N_6903);
and U7660 (N_7660,N_6829,N_6570);
and U7661 (N_7661,N_6694,N_6648);
or U7662 (N_7662,N_6201,N_6887);
xor U7663 (N_7663,N_6566,N_6040);
and U7664 (N_7664,N_6215,N_6994);
nor U7665 (N_7665,N_6671,N_6593);
or U7666 (N_7666,N_6634,N_6482);
nor U7667 (N_7667,N_6879,N_6171);
or U7668 (N_7668,N_6221,N_6700);
nand U7669 (N_7669,N_6652,N_6855);
nor U7670 (N_7670,N_6371,N_6737);
or U7671 (N_7671,N_6626,N_6132);
nor U7672 (N_7672,N_6244,N_6127);
and U7673 (N_7673,N_6856,N_6073);
nand U7674 (N_7674,N_6907,N_6532);
and U7675 (N_7675,N_6458,N_6894);
nor U7676 (N_7676,N_6198,N_6394);
nand U7677 (N_7677,N_6586,N_6232);
and U7678 (N_7678,N_6881,N_6406);
nor U7679 (N_7679,N_6000,N_6965);
nand U7680 (N_7680,N_6393,N_6704);
nor U7681 (N_7681,N_6114,N_6613);
and U7682 (N_7682,N_6118,N_6423);
or U7683 (N_7683,N_6923,N_6289);
and U7684 (N_7684,N_6368,N_6028);
and U7685 (N_7685,N_6248,N_6150);
or U7686 (N_7686,N_6098,N_6042);
or U7687 (N_7687,N_6064,N_6533);
and U7688 (N_7688,N_6150,N_6388);
and U7689 (N_7689,N_6240,N_6052);
or U7690 (N_7690,N_6723,N_6727);
and U7691 (N_7691,N_6676,N_6931);
or U7692 (N_7692,N_6778,N_6085);
and U7693 (N_7693,N_6679,N_6432);
and U7694 (N_7694,N_6925,N_6933);
nand U7695 (N_7695,N_6576,N_6955);
and U7696 (N_7696,N_6727,N_6037);
nor U7697 (N_7697,N_6566,N_6872);
nand U7698 (N_7698,N_6873,N_6754);
or U7699 (N_7699,N_6920,N_6078);
or U7700 (N_7700,N_6505,N_6479);
nand U7701 (N_7701,N_6296,N_6401);
nand U7702 (N_7702,N_6081,N_6317);
nor U7703 (N_7703,N_6992,N_6247);
or U7704 (N_7704,N_6375,N_6473);
or U7705 (N_7705,N_6141,N_6712);
and U7706 (N_7706,N_6382,N_6709);
nand U7707 (N_7707,N_6251,N_6421);
nand U7708 (N_7708,N_6172,N_6919);
nand U7709 (N_7709,N_6559,N_6006);
and U7710 (N_7710,N_6518,N_6536);
and U7711 (N_7711,N_6778,N_6138);
or U7712 (N_7712,N_6189,N_6290);
nand U7713 (N_7713,N_6507,N_6295);
or U7714 (N_7714,N_6629,N_6138);
nor U7715 (N_7715,N_6455,N_6462);
nor U7716 (N_7716,N_6861,N_6852);
nand U7717 (N_7717,N_6354,N_6189);
nor U7718 (N_7718,N_6702,N_6675);
and U7719 (N_7719,N_6262,N_6146);
nand U7720 (N_7720,N_6871,N_6886);
nor U7721 (N_7721,N_6704,N_6822);
and U7722 (N_7722,N_6150,N_6046);
or U7723 (N_7723,N_6045,N_6855);
xnor U7724 (N_7724,N_6838,N_6053);
nor U7725 (N_7725,N_6888,N_6891);
and U7726 (N_7726,N_6369,N_6823);
and U7727 (N_7727,N_6888,N_6758);
or U7728 (N_7728,N_6964,N_6565);
nor U7729 (N_7729,N_6170,N_6173);
xnor U7730 (N_7730,N_6758,N_6302);
and U7731 (N_7731,N_6329,N_6064);
nand U7732 (N_7732,N_6169,N_6648);
and U7733 (N_7733,N_6295,N_6485);
nand U7734 (N_7734,N_6338,N_6670);
nand U7735 (N_7735,N_6447,N_6334);
and U7736 (N_7736,N_6845,N_6763);
nand U7737 (N_7737,N_6006,N_6212);
and U7738 (N_7738,N_6761,N_6030);
or U7739 (N_7739,N_6957,N_6329);
and U7740 (N_7740,N_6691,N_6067);
or U7741 (N_7741,N_6496,N_6422);
nand U7742 (N_7742,N_6701,N_6111);
nor U7743 (N_7743,N_6049,N_6469);
nor U7744 (N_7744,N_6292,N_6734);
or U7745 (N_7745,N_6845,N_6585);
nand U7746 (N_7746,N_6394,N_6920);
or U7747 (N_7747,N_6170,N_6422);
nand U7748 (N_7748,N_6026,N_6316);
nand U7749 (N_7749,N_6489,N_6397);
nor U7750 (N_7750,N_6960,N_6947);
nand U7751 (N_7751,N_6676,N_6662);
nand U7752 (N_7752,N_6849,N_6389);
xnor U7753 (N_7753,N_6759,N_6339);
and U7754 (N_7754,N_6071,N_6511);
or U7755 (N_7755,N_6910,N_6903);
and U7756 (N_7756,N_6510,N_6698);
or U7757 (N_7757,N_6880,N_6356);
nand U7758 (N_7758,N_6274,N_6747);
nor U7759 (N_7759,N_6820,N_6169);
or U7760 (N_7760,N_6871,N_6087);
nand U7761 (N_7761,N_6621,N_6890);
nor U7762 (N_7762,N_6522,N_6102);
nand U7763 (N_7763,N_6721,N_6778);
or U7764 (N_7764,N_6649,N_6927);
or U7765 (N_7765,N_6032,N_6216);
nor U7766 (N_7766,N_6967,N_6855);
nor U7767 (N_7767,N_6732,N_6071);
nor U7768 (N_7768,N_6940,N_6753);
nor U7769 (N_7769,N_6344,N_6538);
and U7770 (N_7770,N_6722,N_6258);
or U7771 (N_7771,N_6731,N_6442);
or U7772 (N_7772,N_6876,N_6554);
nand U7773 (N_7773,N_6034,N_6055);
and U7774 (N_7774,N_6732,N_6579);
or U7775 (N_7775,N_6412,N_6511);
nor U7776 (N_7776,N_6020,N_6527);
or U7777 (N_7777,N_6281,N_6480);
nor U7778 (N_7778,N_6008,N_6304);
and U7779 (N_7779,N_6080,N_6334);
nand U7780 (N_7780,N_6891,N_6022);
or U7781 (N_7781,N_6478,N_6709);
and U7782 (N_7782,N_6400,N_6532);
or U7783 (N_7783,N_6021,N_6949);
or U7784 (N_7784,N_6805,N_6320);
nor U7785 (N_7785,N_6848,N_6362);
nor U7786 (N_7786,N_6294,N_6172);
nor U7787 (N_7787,N_6924,N_6235);
nor U7788 (N_7788,N_6074,N_6783);
nand U7789 (N_7789,N_6105,N_6364);
nor U7790 (N_7790,N_6186,N_6138);
and U7791 (N_7791,N_6553,N_6348);
or U7792 (N_7792,N_6813,N_6881);
or U7793 (N_7793,N_6130,N_6654);
nor U7794 (N_7794,N_6144,N_6512);
nor U7795 (N_7795,N_6817,N_6923);
nor U7796 (N_7796,N_6490,N_6009);
nor U7797 (N_7797,N_6171,N_6851);
and U7798 (N_7798,N_6917,N_6228);
nor U7799 (N_7799,N_6481,N_6989);
nand U7800 (N_7800,N_6849,N_6076);
nand U7801 (N_7801,N_6248,N_6557);
and U7802 (N_7802,N_6652,N_6099);
nor U7803 (N_7803,N_6406,N_6199);
nand U7804 (N_7804,N_6510,N_6176);
or U7805 (N_7805,N_6152,N_6194);
nor U7806 (N_7806,N_6535,N_6431);
or U7807 (N_7807,N_6981,N_6476);
or U7808 (N_7808,N_6350,N_6132);
nor U7809 (N_7809,N_6266,N_6571);
or U7810 (N_7810,N_6917,N_6686);
and U7811 (N_7811,N_6892,N_6116);
and U7812 (N_7812,N_6003,N_6762);
and U7813 (N_7813,N_6850,N_6140);
or U7814 (N_7814,N_6810,N_6819);
and U7815 (N_7815,N_6385,N_6645);
nor U7816 (N_7816,N_6211,N_6492);
nor U7817 (N_7817,N_6268,N_6730);
nor U7818 (N_7818,N_6408,N_6768);
nand U7819 (N_7819,N_6677,N_6900);
or U7820 (N_7820,N_6833,N_6735);
or U7821 (N_7821,N_6244,N_6303);
nor U7822 (N_7822,N_6814,N_6474);
nor U7823 (N_7823,N_6820,N_6207);
and U7824 (N_7824,N_6305,N_6585);
xnor U7825 (N_7825,N_6650,N_6449);
or U7826 (N_7826,N_6991,N_6575);
or U7827 (N_7827,N_6761,N_6777);
nand U7828 (N_7828,N_6611,N_6324);
nor U7829 (N_7829,N_6903,N_6686);
nand U7830 (N_7830,N_6797,N_6074);
or U7831 (N_7831,N_6588,N_6497);
nand U7832 (N_7832,N_6499,N_6623);
nand U7833 (N_7833,N_6787,N_6830);
or U7834 (N_7834,N_6192,N_6587);
and U7835 (N_7835,N_6173,N_6282);
nor U7836 (N_7836,N_6578,N_6604);
nor U7837 (N_7837,N_6991,N_6432);
nand U7838 (N_7838,N_6925,N_6758);
nand U7839 (N_7839,N_6983,N_6038);
nor U7840 (N_7840,N_6379,N_6895);
and U7841 (N_7841,N_6419,N_6246);
nand U7842 (N_7842,N_6336,N_6223);
nand U7843 (N_7843,N_6064,N_6017);
nand U7844 (N_7844,N_6585,N_6173);
nor U7845 (N_7845,N_6157,N_6615);
nand U7846 (N_7846,N_6148,N_6612);
nand U7847 (N_7847,N_6862,N_6343);
and U7848 (N_7848,N_6587,N_6862);
nand U7849 (N_7849,N_6613,N_6584);
or U7850 (N_7850,N_6067,N_6672);
or U7851 (N_7851,N_6348,N_6572);
and U7852 (N_7852,N_6801,N_6594);
nor U7853 (N_7853,N_6556,N_6294);
and U7854 (N_7854,N_6866,N_6181);
and U7855 (N_7855,N_6680,N_6674);
and U7856 (N_7856,N_6706,N_6689);
and U7857 (N_7857,N_6709,N_6807);
or U7858 (N_7858,N_6761,N_6297);
nand U7859 (N_7859,N_6064,N_6273);
and U7860 (N_7860,N_6803,N_6604);
or U7861 (N_7861,N_6121,N_6501);
nand U7862 (N_7862,N_6021,N_6909);
nand U7863 (N_7863,N_6951,N_6677);
xnor U7864 (N_7864,N_6846,N_6933);
or U7865 (N_7865,N_6672,N_6416);
nand U7866 (N_7866,N_6386,N_6470);
or U7867 (N_7867,N_6452,N_6902);
and U7868 (N_7868,N_6456,N_6914);
or U7869 (N_7869,N_6342,N_6376);
or U7870 (N_7870,N_6907,N_6332);
or U7871 (N_7871,N_6551,N_6364);
or U7872 (N_7872,N_6142,N_6546);
nor U7873 (N_7873,N_6519,N_6717);
nor U7874 (N_7874,N_6336,N_6580);
nand U7875 (N_7875,N_6224,N_6542);
nor U7876 (N_7876,N_6639,N_6827);
nand U7877 (N_7877,N_6115,N_6367);
or U7878 (N_7878,N_6365,N_6294);
nor U7879 (N_7879,N_6902,N_6015);
nand U7880 (N_7880,N_6776,N_6890);
nand U7881 (N_7881,N_6258,N_6485);
or U7882 (N_7882,N_6225,N_6189);
and U7883 (N_7883,N_6556,N_6844);
or U7884 (N_7884,N_6279,N_6630);
nor U7885 (N_7885,N_6766,N_6886);
nand U7886 (N_7886,N_6676,N_6472);
and U7887 (N_7887,N_6745,N_6449);
and U7888 (N_7888,N_6214,N_6597);
nand U7889 (N_7889,N_6892,N_6222);
or U7890 (N_7890,N_6813,N_6741);
and U7891 (N_7891,N_6128,N_6429);
or U7892 (N_7892,N_6008,N_6933);
or U7893 (N_7893,N_6985,N_6198);
xnor U7894 (N_7894,N_6652,N_6199);
xor U7895 (N_7895,N_6759,N_6857);
nor U7896 (N_7896,N_6497,N_6790);
nor U7897 (N_7897,N_6959,N_6510);
nor U7898 (N_7898,N_6206,N_6159);
nor U7899 (N_7899,N_6536,N_6751);
nand U7900 (N_7900,N_6890,N_6106);
nand U7901 (N_7901,N_6109,N_6104);
nand U7902 (N_7902,N_6607,N_6240);
nand U7903 (N_7903,N_6486,N_6743);
nand U7904 (N_7904,N_6797,N_6399);
and U7905 (N_7905,N_6475,N_6517);
nor U7906 (N_7906,N_6872,N_6638);
nor U7907 (N_7907,N_6937,N_6938);
and U7908 (N_7908,N_6388,N_6636);
nor U7909 (N_7909,N_6096,N_6683);
nor U7910 (N_7910,N_6409,N_6269);
and U7911 (N_7911,N_6638,N_6454);
or U7912 (N_7912,N_6009,N_6589);
nand U7913 (N_7913,N_6730,N_6312);
nor U7914 (N_7914,N_6474,N_6755);
or U7915 (N_7915,N_6795,N_6014);
and U7916 (N_7916,N_6228,N_6937);
and U7917 (N_7917,N_6237,N_6762);
and U7918 (N_7918,N_6731,N_6148);
nand U7919 (N_7919,N_6594,N_6570);
nor U7920 (N_7920,N_6400,N_6742);
or U7921 (N_7921,N_6298,N_6957);
or U7922 (N_7922,N_6716,N_6313);
xnor U7923 (N_7923,N_6754,N_6158);
nand U7924 (N_7924,N_6775,N_6295);
or U7925 (N_7925,N_6814,N_6557);
nor U7926 (N_7926,N_6489,N_6632);
and U7927 (N_7927,N_6294,N_6758);
nor U7928 (N_7928,N_6944,N_6538);
and U7929 (N_7929,N_6411,N_6873);
nand U7930 (N_7930,N_6277,N_6479);
or U7931 (N_7931,N_6672,N_6261);
and U7932 (N_7932,N_6947,N_6139);
or U7933 (N_7933,N_6162,N_6980);
nand U7934 (N_7934,N_6649,N_6036);
nand U7935 (N_7935,N_6757,N_6150);
or U7936 (N_7936,N_6080,N_6138);
nor U7937 (N_7937,N_6815,N_6921);
nand U7938 (N_7938,N_6035,N_6113);
and U7939 (N_7939,N_6179,N_6505);
nor U7940 (N_7940,N_6866,N_6224);
nor U7941 (N_7941,N_6793,N_6292);
and U7942 (N_7942,N_6792,N_6469);
or U7943 (N_7943,N_6972,N_6897);
nor U7944 (N_7944,N_6732,N_6923);
or U7945 (N_7945,N_6504,N_6744);
and U7946 (N_7946,N_6771,N_6039);
nor U7947 (N_7947,N_6620,N_6313);
and U7948 (N_7948,N_6291,N_6809);
nor U7949 (N_7949,N_6346,N_6428);
nor U7950 (N_7950,N_6231,N_6568);
and U7951 (N_7951,N_6728,N_6749);
nand U7952 (N_7952,N_6337,N_6728);
nand U7953 (N_7953,N_6401,N_6861);
nand U7954 (N_7954,N_6191,N_6496);
xnor U7955 (N_7955,N_6197,N_6376);
nor U7956 (N_7956,N_6822,N_6452);
nor U7957 (N_7957,N_6998,N_6659);
nor U7958 (N_7958,N_6048,N_6711);
xnor U7959 (N_7959,N_6923,N_6672);
nand U7960 (N_7960,N_6227,N_6815);
nor U7961 (N_7961,N_6944,N_6652);
or U7962 (N_7962,N_6370,N_6141);
or U7963 (N_7963,N_6622,N_6874);
and U7964 (N_7964,N_6281,N_6900);
xor U7965 (N_7965,N_6952,N_6976);
or U7966 (N_7966,N_6661,N_6939);
and U7967 (N_7967,N_6619,N_6709);
and U7968 (N_7968,N_6860,N_6890);
or U7969 (N_7969,N_6696,N_6550);
nor U7970 (N_7970,N_6254,N_6268);
and U7971 (N_7971,N_6512,N_6028);
and U7972 (N_7972,N_6884,N_6210);
nand U7973 (N_7973,N_6056,N_6216);
or U7974 (N_7974,N_6579,N_6197);
and U7975 (N_7975,N_6513,N_6018);
or U7976 (N_7976,N_6010,N_6503);
nand U7977 (N_7977,N_6243,N_6845);
and U7978 (N_7978,N_6374,N_6226);
xor U7979 (N_7979,N_6558,N_6415);
nor U7980 (N_7980,N_6714,N_6893);
or U7981 (N_7981,N_6577,N_6858);
or U7982 (N_7982,N_6504,N_6186);
nand U7983 (N_7983,N_6627,N_6135);
or U7984 (N_7984,N_6481,N_6337);
nand U7985 (N_7985,N_6647,N_6793);
or U7986 (N_7986,N_6238,N_6651);
and U7987 (N_7987,N_6641,N_6082);
and U7988 (N_7988,N_6299,N_6094);
or U7989 (N_7989,N_6702,N_6764);
nand U7990 (N_7990,N_6497,N_6661);
and U7991 (N_7991,N_6719,N_6097);
and U7992 (N_7992,N_6440,N_6451);
and U7993 (N_7993,N_6178,N_6337);
or U7994 (N_7994,N_6876,N_6351);
nor U7995 (N_7995,N_6734,N_6828);
nand U7996 (N_7996,N_6470,N_6140);
nor U7997 (N_7997,N_6395,N_6563);
xnor U7998 (N_7998,N_6436,N_6094);
nor U7999 (N_7999,N_6638,N_6613);
and U8000 (N_8000,N_7264,N_7033);
nand U8001 (N_8001,N_7096,N_7823);
nand U8002 (N_8002,N_7135,N_7552);
and U8003 (N_8003,N_7628,N_7496);
or U8004 (N_8004,N_7151,N_7962);
and U8005 (N_8005,N_7736,N_7269);
or U8006 (N_8006,N_7539,N_7755);
and U8007 (N_8007,N_7193,N_7906);
nand U8008 (N_8008,N_7716,N_7863);
nand U8009 (N_8009,N_7171,N_7372);
or U8010 (N_8010,N_7396,N_7040);
and U8011 (N_8011,N_7585,N_7146);
nor U8012 (N_8012,N_7510,N_7702);
and U8013 (N_8013,N_7069,N_7262);
and U8014 (N_8014,N_7435,N_7909);
nor U8015 (N_8015,N_7215,N_7361);
or U8016 (N_8016,N_7106,N_7518);
or U8017 (N_8017,N_7908,N_7444);
nand U8018 (N_8018,N_7390,N_7085);
and U8019 (N_8019,N_7242,N_7216);
or U8020 (N_8020,N_7887,N_7843);
or U8021 (N_8021,N_7758,N_7580);
and U8022 (N_8022,N_7442,N_7026);
and U8023 (N_8023,N_7333,N_7611);
nor U8024 (N_8024,N_7547,N_7060);
nand U8025 (N_8025,N_7695,N_7865);
nor U8026 (N_8026,N_7098,N_7815);
nor U8027 (N_8027,N_7666,N_7349);
and U8028 (N_8028,N_7699,N_7392);
nand U8029 (N_8029,N_7270,N_7837);
and U8030 (N_8030,N_7733,N_7315);
and U8031 (N_8031,N_7445,N_7121);
or U8032 (N_8032,N_7901,N_7773);
and U8033 (N_8033,N_7717,N_7600);
and U8034 (N_8034,N_7670,N_7986);
nor U8035 (N_8035,N_7142,N_7932);
nand U8036 (N_8036,N_7852,N_7100);
nor U8037 (N_8037,N_7414,N_7799);
or U8038 (N_8038,N_7015,N_7701);
nor U8039 (N_8039,N_7503,N_7526);
and U8040 (N_8040,N_7757,N_7663);
or U8041 (N_8041,N_7453,N_7499);
xor U8042 (N_8042,N_7747,N_7898);
nor U8043 (N_8043,N_7783,N_7080);
nor U8044 (N_8044,N_7377,N_7356);
nand U8045 (N_8045,N_7275,N_7594);
and U8046 (N_8046,N_7381,N_7739);
or U8047 (N_8047,N_7016,N_7954);
nand U8048 (N_8048,N_7895,N_7544);
xnor U8049 (N_8049,N_7446,N_7926);
nor U8050 (N_8050,N_7147,N_7365);
nand U8051 (N_8051,N_7664,N_7124);
nand U8052 (N_8052,N_7199,N_7623);
and U8053 (N_8053,N_7688,N_7112);
nor U8054 (N_8054,N_7566,N_7330);
nor U8055 (N_8055,N_7960,N_7022);
and U8056 (N_8056,N_7448,N_7407);
nor U8057 (N_8057,N_7748,N_7849);
or U8058 (N_8058,N_7994,N_7172);
nand U8059 (N_8059,N_7494,N_7484);
nand U8060 (N_8060,N_7049,N_7181);
nand U8061 (N_8061,N_7386,N_7397);
and U8062 (N_8062,N_7078,N_7556);
nor U8063 (N_8063,N_7787,N_7317);
nand U8064 (N_8064,N_7668,N_7829);
nand U8065 (N_8065,N_7293,N_7366);
nor U8066 (N_8066,N_7576,N_7604);
nor U8067 (N_8067,N_7447,N_7608);
or U8068 (N_8068,N_7332,N_7568);
or U8069 (N_8069,N_7079,N_7292);
nor U8070 (N_8070,N_7949,N_7338);
and U8071 (N_8071,N_7310,N_7730);
and U8072 (N_8072,N_7055,N_7800);
nor U8073 (N_8073,N_7169,N_7584);
nor U8074 (N_8074,N_7665,N_7659);
and U8075 (N_8075,N_7327,N_7498);
or U8076 (N_8076,N_7200,N_7482);
nand U8077 (N_8077,N_7999,N_7583);
or U8078 (N_8078,N_7978,N_7367);
and U8079 (N_8079,N_7804,N_7158);
or U8080 (N_8080,N_7502,N_7213);
or U8081 (N_8081,N_7251,N_7712);
nor U8082 (N_8082,N_7391,N_7019);
and U8083 (N_8083,N_7593,N_7819);
nor U8084 (N_8084,N_7300,N_7864);
xor U8085 (N_8085,N_7486,N_7808);
or U8086 (N_8086,N_7045,N_7798);
nor U8087 (N_8087,N_7074,N_7025);
nand U8088 (N_8088,N_7959,N_7924);
nor U8089 (N_8089,N_7638,N_7579);
nor U8090 (N_8090,N_7878,N_7093);
or U8091 (N_8091,N_7255,N_7616);
or U8092 (N_8092,N_7925,N_7126);
or U8093 (N_8093,N_7020,N_7461);
and U8094 (N_8094,N_7229,N_7034);
nand U8095 (N_8095,N_7101,N_7032);
or U8096 (N_8096,N_7083,N_7910);
and U8097 (N_8097,N_7814,N_7490);
or U8098 (N_8098,N_7303,N_7643);
nand U8099 (N_8099,N_7048,N_7099);
nor U8100 (N_8100,N_7375,N_7627);
nand U8101 (N_8101,N_7420,N_7694);
and U8102 (N_8102,N_7288,N_7111);
or U8103 (N_8103,N_7676,N_7724);
or U8104 (N_8104,N_7191,N_7619);
or U8105 (N_8105,N_7094,N_7519);
nand U8106 (N_8106,N_7766,N_7769);
nand U8107 (N_8107,N_7212,N_7387);
xor U8108 (N_8108,N_7039,N_7529);
nand U8109 (N_8109,N_7687,N_7024);
nand U8110 (N_8110,N_7675,N_7294);
or U8111 (N_8111,N_7641,N_7388);
nand U8112 (N_8112,N_7072,N_7189);
nand U8113 (N_8113,N_7363,N_7248);
nand U8114 (N_8114,N_7533,N_7653);
or U8115 (N_8115,N_7150,N_7975);
or U8116 (N_8116,N_7462,N_7685);
or U8117 (N_8117,N_7329,N_7003);
and U8118 (N_8118,N_7995,N_7700);
nand U8119 (N_8119,N_7721,N_7869);
nand U8120 (N_8120,N_7308,N_7344);
nor U8121 (N_8121,N_7334,N_7803);
and U8122 (N_8122,N_7780,N_7192);
nor U8123 (N_8123,N_7913,N_7450);
nand U8124 (N_8124,N_7487,N_7430);
nand U8125 (N_8125,N_7259,N_7380);
nand U8126 (N_8126,N_7018,N_7817);
nand U8127 (N_8127,N_7120,N_7942);
and U8128 (N_8128,N_7122,N_7119);
nor U8129 (N_8129,N_7813,N_7969);
or U8130 (N_8130,N_7421,N_7137);
or U8131 (N_8131,N_7440,N_7920);
and U8132 (N_8132,N_7253,N_7007);
xor U8133 (N_8133,N_7419,N_7749);
or U8134 (N_8134,N_7649,N_7561);
and U8135 (N_8135,N_7847,N_7013);
or U8136 (N_8136,N_7469,N_7982);
nor U8137 (N_8137,N_7882,N_7046);
and U8138 (N_8138,N_7967,N_7173);
nor U8139 (N_8139,N_7834,N_7928);
nor U8140 (N_8140,N_7509,N_7422);
and U8141 (N_8141,N_7848,N_7417);
or U8142 (N_8142,N_7548,N_7915);
nand U8143 (N_8143,N_7639,N_7763);
nand U8144 (N_8144,N_7620,N_7642);
nand U8145 (N_8145,N_7632,N_7890);
or U8146 (N_8146,N_7698,N_7265);
nor U8147 (N_8147,N_7671,N_7984);
nor U8148 (N_8148,N_7467,N_7656);
or U8149 (N_8149,N_7514,N_7718);
and U8150 (N_8150,N_7939,N_7051);
nor U8151 (N_8151,N_7892,N_7170);
nand U8152 (N_8152,N_7297,N_7965);
and U8153 (N_8153,N_7410,N_7768);
nand U8154 (N_8154,N_7655,N_7236);
xor U8155 (N_8155,N_7821,N_7822);
nand U8156 (N_8156,N_7340,N_7056);
and U8157 (N_8157,N_7684,N_7746);
and U8158 (N_8158,N_7621,N_7412);
and U8159 (N_8159,N_7940,N_7631);
nor U8160 (N_8160,N_7776,N_7398);
or U8161 (N_8161,N_7057,N_7005);
or U8162 (N_8162,N_7515,N_7290);
nand U8163 (N_8163,N_7788,N_7283);
and U8164 (N_8164,N_7997,N_7006);
nor U8165 (N_8165,N_7538,N_7870);
and U8166 (N_8166,N_7581,N_7988);
or U8167 (N_8167,N_7737,N_7709);
nor U8168 (N_8168,N_7582,N_7035);
or U8169 (N_8169,N_7185,N_7601);
or U8170 (N_8170,N_7413,N_7596);
nand U8171 (N_8171,N_7411,N_7820);
nand U8172 (N_8172,N_7221,N_7672);
or U8173 (N_8173,N_7572,N_7985);
and U8174 (N_8174,N_7797,N_7465);
nand U8175 (N_8175,N_7577,N_7830);
and U8176 (N_8176,N_7304,N_7937);
xnor U8177 (N_8177,N_7341,N_7070);
or U8178 (N_8178,N_7402,N_7062);
xor U8179 (N_8179,N_7557,N_7337);
or U8180 (N_8180,N_7971,N_7203);
or U8181 (N_8181,N_7570,N_7745);
nor U8182 (N_8182,N_7862,N_7989);
and U8183 (N_8183,N_7610,N_7481);
nand U8184 (N_8184,N_7225,N_7851);
nor U8185 (N_8185,N_7753,N_7835);
nor U8186 (N_8186,N_7350,N_7722);
nor U8187 (N_8187,N_7563,N_7086);
nor U8188 (N_8188,N_7260,N_7107);
or U8189 (N_8189,N_7825,N_7618);
or U8190 (N_8190,N_7550,N_7194);
or U8191 (N_8191,N_7027,N_7727);
and U8192 (N_8192,N_7452,N_7991);
nor U8193 (N_8193,N_7795,N_7728);
and U8194 (N_8194,N_7723,N_7029);
nor U8195 (N_8195,N_7284,N_7634);
nor U8196 (N_8196,N_7472,N_7276);
nor U8197 (N_8197,N_7992,N_7370);
nor U8198 (N_8198,N_7853,N_7779);
nor U8199 (N_8199,N_7772,N_7599);
nand U8200 (N_8200,N_7661,N_7456);
and U8201 (N_8201,N_7873,N_7358);
and U8202 (N_8202,N_7307,N_7164);
and U8203 (N_8203,N_7084,N_7752);
nor U8204 (N_8204,N_7014,N_7416);
and U8205 (N_8205,N_7492,N_7648);
xnor U8206 (N_8206,N_7818,N_7681);
nand U8207 (N_8207,N_7824,N_7176);
or U8208 (N_8208,N_7560,N_7295);
nor U8209 (N_8209,N_7609,N_7188);
nor U8210 (N_8210,N_7360,N_7355);
nor U8211 (N_8211,N_7574,N_7109);
and U8212 (N_8212,N_7266,N_7385);
nand U8213 (N_8213,N_7952,N_7322);
nand U8214 (N_8214,N_7058,N_7697);
nor U8215 (N_8215,N_7426,N_7222);
xnor U8216 (N_8216,N_7517,N_7948);
nand U8217 (N_8217,N_7041,N_7838);
nand U8218 (N_8218,N_7277,N_7660);
or U8219 (N_8219,N_7961,N_7774);
or U8220 (N_8220,N_7371,N_7588);
nor U8221 (N_8221,N_7354,N_7807);
nand U8222 (N_8222,N_7883,N_7233);
or U8223 (N_8223,N_7943,N_7726);
nand U8224 (N_8224,N_7090,N_7161);
and U8225 (N_8225,N_7929,N_7996);
and U8226 (N_8226,N_7562,N_7934);
xnor U8227 (N_8227,N_7936,N_7974);
or U8228 (N_8228,N_7775,N_7393);
or U8229 (N_8229,N_7383,N_7647);
nand U8230 (N_8230,N_7302,N_7791);
or U8231 (N_8231,N_7918,N_7479);
nand U8232 (N_8232,N_7316,N_7127);
and U8233 (N_8233,N_7418,N_7081);
or U8234 (N_8234,N_7113,N_7801);
and U8235 (N_8235,N_7261,N_7425);
xnor U8236 (N_8236,N_7408,N_7597);
nor U8237 (N_8237,N_7108,N_7134);
and U8238 (N_8238,N_7624,N_7885);
or U8239 (N_8239,N_7289,N_7522);
or U8240 (N_8240,N_7673,N_7516);
or U8241 (N_8241,N_7979,N_7339);
or U8242 (N_8242,N_7714,N_7091);
nor U8243 (N_8243,N_7541,N_7021);
or U8244 (N_8244,N_7424,N_7657);
nand U8245 (N_8245,N_7778,N_7678);
and U8246 (N_8246,N_7497,N_7679);
nor U8247 (N_8247,N_7477,N_7252);
nor U8248 (N_8248,N_7458,N_7512);
nor U8249 (N_8249,N_7886,N_7811);
or U8250 (N_8250,N_7237,N_7470);
or U8251 (N_8251,N_7564,N_7513);
and U8252 (N_8252,N_7231,N_7175);
nor U8253 (N_8253,N_7951,N_7073);
nor U8254 (N_8254,N_7537,N_7287);
and U8255 (N_8255,N_7501,N_7927);
nor U8256 (N_8256,N_7163,N_7475);
nor U8257 (N_8257,N_7793,N_7612);
nand U8258 (N_8258,N_7941,N_7220);
nor U8259 (N_8259,N_7052,N_7794);
and U8260 (N_8260,N_7855,N_7434);
xnor U8261 (N_8261,N_7744,N_7917);
nand U8262 (N_8262,N_7038,N_7973);
and U8263 (N_8263,N_7211,N_7633);
xnor U8264 (N_8264,N_7323,N_7267);
xnor U8265 (N_8265,N_7162,N_7362);
or U8266 (N_8266,N_7364,N_7244);
or U8267 (N_8267,N_7919,N_7061);
nor U8268 (N_8268,N_7907,N_7806);
or U8269 (N_8269,N_7603,N_7536);
nand U8270 (N_8270,N_7796,N_7345);
nor U8271 (N_8271,N_7258,N_7493);
or U8272 (N_8272,N_7400,N_7646);
xor U8273 (N_8273,N_7899,N_7306);
nor U8274 (N_8274,N_7654,N_7399);
and U8275 (N_8275,N_7118,N_7353);
and U8276 (N_8276,N_7507,N_7947);
or U8277 (N_8277,N_7662,N_7357);
or U8278 (N_8278,N_7812,N_7789);
nand U8279 (N_8279,N_7549,N_7543);
nand U8280 (N_8280,N_7468,N_7770);
nor U8281 (N_8281,N_7809,N_7280);
or U8282 (N_8282,N_7184,N_7240);
nand U8283 (N_8283,N_7321,N_7802);
and U8284 (N_8284,N_7968,N_7858);
or U8285 (N_8285,N_7879,N_7630);
and U8286 (N_8286,N_7931,N_7204);
nand U8287 (N_8287,N_7382,N_7912);
and U8288 (N_8288,N_7586,N_7273);
and U8289 (N_8289,N_7651,N_7314);
and U8290 (N_8290,N_7152,N_7876);
nand U8291 (N_8291,N_7715,N_7553);
or U8292 (N_8292,N_7987,N_7914);
nand U8293 (N_8293,N_7245,N_7527);
nand U8294 (N_8294,N_7179,N_7554);
nand U8295 (N_8295,N_7077,N_7981);
or U8296 (N_8296,N_7218,N_7312);
and U8297 (N_8297,N_7488,N_7202);
and U8298 (N_8298,N_7299,N_7729);
and U8299 (N_8299,N_7652,N_7342);
nand U8300 (N_8300,N_7012,N_7208);
and U8301 (N_8301,N_7613,N_7075);
nand U8302 (N_8302,N_7841,N_7246);
and U8303 (N_8303,N_7428,N_7826);
and U8304 (N_8304,N_7742,N_7087);
nand U8305 (N_8305,N_7359,N_7324);
nand U8306 (N_8306,N_7884,N_7859);
and U8307 (N_8307,N_7781,N_7505);
nor U8308 (N_8308,N_7186,N_7219);
nor U8309 (N_8309,N_7703,N_7177);
nand U8310 (N_8310,N_7017,N_7990);
and U8311 (N_8311,N_7966,N_7944);
nor U8312 (N_8312,N_7767,N_7214);
and U8313 (N_8313,N_7318,N_7132);
or U8314 (N_8314,N_7506,N_7771);
or U8315 (N_8315,N_7963,N_7207);
nand U8316 (N_8316,N_7856,N_7071);
nand U8317 (N_8317,N_7154,N_7313);
or U8318 (N_8318,N_7319,N_7234);
nand U8319 (N_8319,N_7640,N_7592);
nand U8320 (N_8320,N_7110,N_7128);
nand U8321 (N_8321,N_7389,N_7922);
or U8322 (N_8322,N_7373,N_7023);
nand U8323 (N_8323,N_7827,N_7092);
and U8324 (N_8324,N_7508,N_7198);
and U8325 (N_8325,N_7249,N_7195);
and U8326 (N_8326,N_7531,N_7305);
nand U8327 (N_8327,N_7889,N_7066);
nand U8328 (N_8328,N_7478,N_7523);
and U8329 (N_8329,N_7254,N_7845);
and U8330 (N_8330,N_7704,N_7165);
nand U8331 (N_8331,N_7784,N_7614);
and U8332 (N_8332,N_7521,N_7875);
and U8333 (N_8333,N_7902,N_7063);
nor U8334 (N_8334,N_7130,N_7846);
and U8335 (N_8335,N_7140,N_7224);
nor U8336 (N_8336,N_7160,N_7136);
nand U8337 (N_8337,N_7950,N_7756);
xor U8338 (N_8338,N_7436,N_7635);
nor U8339 (N_8339,N_7285,N_7786);
nand U8340 (N_8340,N_7607,N_7532);
nor U8341 (N_8341,N_7369,N_7011);
nor U8342 (N_8342,N_7232,N_7953);
or U8343 (N_8343,N_7149,N_7291);
nor U8344 (N_8344,N_7565,N_7394);
and U8345 (N_8345,N_7031,N_7153);
or U8346 (N_8346,N_7053,N_7598);
nor U8347 (N_8347,N_7691,N_7650);
and U8348 (N_8348,N_7540,N_7534);
nand U8349 (N_8349,N_7956,N_7243);
or U8350 (N_8350,N_7861,N_7138);
nor U8351 (N_8351,N_7590,N_7278);
or U8352 (N_8352,N_7125,N_7692);
nor U8353 (N_8353,N_7009,N_7187);
nor U8354 (N_8354,N_7602,N_7880);
nor U8355 (N_8355,N_7464,N_7483);
and U8356 (N_8356,N_7201,N_7850);
nor U8357 (N_8357,N_7760,N_7764);
xor U8358 (N_8358,N_7658,N_7309);
nand U8359 (N_8359,N_7064,N_7765);
or U8360 (N_8360,N_7710,N_7591);
or U8361 (N_8361,N_7840,N_7347);
and U8362 (N_8362,N_7629,N_7713);
nand U8363 (N_8363,N_7168,N_7970);
nor U8364 (N_8364,N_7888,N_7043);
and U8365 (N_8365,N_7725,N_7104);
or U8366 (N_8366,N_7900,N_7945);
xnor U8367 (N_8367,N_7605,N_7792);
nand U8368 (N_8368,N_7972,N_7205);
nand U8369 (N_8369,N_7325,N_7677);
and U8370 (N_8370,N_7115,N_7433);
or U8371 (N_8371,N_7455,N_7615);
and U8372 (N_8372,N_7454,N_7114);
nand U8373 (N_8373,N_7872,N_7504);
nor U8374 (N_8374,N_7054,N_7690);
or U8375 (N_8375,N_7626,N_7832);
and U8376 (N_8376,N_7256,N_7050);
and U8377 (N_8377,N_7866,N_7155);
nor U8378 (N_8378,N_7683,N_7844);
and U8379 (N_8379,N_7933,N_7896);
nor U8380 (N_8380,N_7376,N_7520);
nand U8381 (N_8381,N_7938,N_7037);
nor U8382 (N_8382,N_7167,N_7669);
nor U8383 (N_8383,N_7867,N_7904);
and U8384 (N_8384,N_7816,N_7331);
and U8385 (N_8385,N_7511,N_7916);
nor U8386 (N_8386,N_7206,N_7500);
or U8387 (N_8387,N_7449,N_7068);
or U8388 (N_8388,N_7976,N_7065);
nand U8389 (N_8389,N_7595,N_7466);
or U8390 (N_8390,N_7443,N_7530);
nand U8391 (N_8391,N_7036,N_7559);
nand U8392 (N_8392,N_7178,N_7686);
or U8393 (N_8393,N_7575,N_7743);
nor U8394 (N_8394,N_7059,N_7437);
nand U8395 (N_8395,N_7301,N_7139);
nor U8396 (N_8396,N_7441,N_7298);
or U8397 (N_8397,N_7103,N_7871);
and U8398 (N_8398,N_7156,N_7209);
nand U8399 (N_8399,N_7854,N_7524);
and U8400 (N_8400,N_7196,N_7935);
and U8401 (N_8401,N_7286,N_7102);
nor U8402 (N_8402,N_7239,N_7719);
nand U8403 (N_8403,N_7116,N_7567);
or U8404 (N_8404,N_7088,N_7546);
and U8405 (N_8405,N_7343,N_7180);
or U8406 (N_8406,N_7558,N_7489);
nand U8407 (N_8407,N_7351,N_7711);
or U8408 (N_8408,N_7777,N_7495);
and U8409 (N_8409,N_7368,N_7636);
and U8410 (N_8410,N_7474,N_7183);
and U8411 (N_8411,N_7272,N_7190);
nand U8412 (N_8412,N_7197,N_7143);
or U8413 (N_8413,N_7089,N_7182);
nand U8414 (N_8414,N_7754,N_7117);
nand U8415 (N_8415,N_7734,N_7587);
nor U8416 (N_8416,N_7983,N_7958);
or U8417 (N_8417,N_7415,N_7491);
and U8418 (N_8418,N_7226,N_7042);
nor U8419 (N_8419,N_7047,N_7328);
nand U8420 (N_8420,N_7008,N_7439);
nor U8421 (N_8421,N_7268,N_7645);
or U8422 (N_8422,N_7998,N_7905);
nand U8423 (N_8423,N_7144,N_7762);
and U8424 (N_8424,N_7667,N_7379);
and U8425 (N_8425,N_7409,N_7457);
nand U8426 (N_8426,N_7217,N_7427);
or U8427 (N_8427,N_7569,N_7831);
or U8428 (N_8428,N_7460,N_7238);
nor U8429 (N_8429,N_7977,N_7263);
nand U8430 (N_8430,N_7761,N_7946);
and U8431 (N_8431,N_7573,N_7957);
nand U8432 (N_8432,N_7894,N_7839);
nand U8433 (N_8433,N_7326,N_7076);
nor U8434 (N_8434,N_7693,N_7897);
nor U8435 (N_8435,N_7028,N_7401);
and U8436 (N_8436,N_7708,N_7732);
nor U8437 (N_8437,N_7706,N_7644);
and U8438 (N_8438,N_7438,N_7740);
nor U8439 (N_8439,N_7625,N_7674);
and U8440 (N_8440,N_7874,N_7705);
and U8441 (N_8441,N_7159,N_7320);
nand U8442 (N_8442,N_7680,N_7403);
nand U8443 (N_8443,N_7868,N_7589);
and U8444 (N_8444,N_7955,N_7473);
xnor U8445 (N_8445,N_7622,N_7476);
or U8446 (N_8446,N_7282,N_7810);
or U8447 (N_8447,N_7860,N_7157);
nand U8448 (N_8448,N_7431,N_7145);
or U8449 (N_8449,N_7241,N_7750);
nor U8450 (N_8450,N_7738,N_7235);
or U8451 (N_8451,N_7395,N_7432);
xnor U8452 (N_8452,N_7881,N_7250);
nor U8453 (N_8453,N_7095,N_7707);
and U8454 (N_8454,N_7555,N_7404);
and U8455 (N_8455,N_7010,N_7230);
or U8456 (N_8456,N_7133,N_7131);
and U8457 (N_8457,N_7405,N_7210);
nand U8458 (N_8458,N_7891,N_7311);
nor U8459 (N_8459,N_7571,N_7545);
nor U8460 (N_8460,N_7141,N_7735);
nand U8461 (N_8461,N_7001,N_7044);
or U8462 (N_8462,N_7166,N_7525);
or U8463 (N_8463,N_7000,N_7471);
or U8464 (N_8464,N_7993,N_7463);
nor U8465 (N_8465,N_7148,N_7828);
and U8466 (N_8466,N_7720,N_7097);
or U8467 (N_8467,N_7346,N_7741);
and U8468 (N_8468,N_7485,N_7247);
nand U8469 (N_8469,N_7833,N_7129);
nand U8470 (N_8470,N_7911,N_7451);
or U8471 (N_8471,N_7105,N_7980);
nand U8472 (N_8472,N_7271,N_7528);
or U8473 (N_8473,N_7336,N_7930);
or U8474 (N_8474,N_7790,N_7637);
xor U8475 (N_8475,N_7429,N_7174);
or U8476 (N_8476,N_7842,N_7535);
or U8477 (N_8477,N_7348,N_7542);
xnor U8478 (N_8478,N_7281,N_7877);
nor U8479 (N_8479,N_7082,N_7551);
nand U8480 (N_8480,N_7228,N_7964);
and U8481 (N_8481,N_7836,N_7751);
and U8482 (N_8482,N_7903,N_7459);
and U8483 (N_8483,N_7384,N_7374);
nor U8484 (N_8484,N_7696,N_7030);
and U8485 (N_8485,N_7785,N_7923);
nand U8486 (N_8486,N_7617,N_7274);
nand U8487 (N_8487,N_7279,N_7378);
or U8488 (N_8488,N_7352,N_7480);
nor U8489 (N_8489,N_7223,N_7893);
or U8490 (N_8490,N_7731,N_7606);
nor U8491 (N_8491,N_7123,N_7406);
and U8492 (N_8492,N_7857,N_7921);
or U8493 (N_8493,N_7682,N_7257);
nor U8494 (N_8494,N_7782,N_7335);
and U8495 (N_8495,N_7689,N_7296);
and U8496 (N_8496,N_7423,N_7227);
and U8497 (N_8497,N_7759,N_7805);
nor U8498 (N_8498,N_7067,N_7002);
or U8499 (N_8499,N_7004,N_7578);
and U8500 (N_8500,N_7717,N_7088);
nand U8501 (N_8501,N_7353,N_7887);
nor U8502 (N_8502,N_7961,N_7835);
nor U8503 (N_8503,N_7487,N_7915);
nor U8504 (N_8504,N_7676,N_7226);
nand U8505 (N_8505,N_7812,N_7358);
and U8506 (N_8506,N_7401,N_7425);
nor U8507 (N_8507,N_7024,N_7206);
nand U8508 (N_8508,N_7729,N_7303);
or U8509 (N_8509,N_7346,N_7551);
nand U8510 (N_8510,N_7177,N_7820);
and U8511 (N_8511,N_7459,N_7359);
and U8512 (N_8512,N_7194,N_7097);
nor U8513 (N_8513,N_7581,N_7684);
nand U8514 (N_8514,N_7240,N_7884);
and U8515 (N_8515,N_7051,N_7443);
nor U8516 (N_8516,N_7745,N_7479);
or U8517 (N_8517,N_7059,N_7501);
or U8518 (N_8518,N_7540,N_7271);
nand U8519 (N_8519,N_7323,N_7174);
nand U8520 (N_8520,N_7332,N_7195);
nor U8521 (N_8521,N_7091,N_7359);
nand U8522 (N_8522,N_7510,N_7403);
nor U8523 (N_8523,N_7467,N_7791);
nand U8524 (N_8524,N_7551,N_7730);
or U8525 (N_8525,N_7471,N_7105);
nand U8526 (N_8526,N_7370,N_7075);
nor U8527 (N_8527,N_7794,N_7153);
or U8528 (N_8528,N_7256,N_7436);
or U8529 (N_8529,N_7904,N_7274);
or U8530 (N_8530,N_7847,N_7733);
nand U8531 (N_8531,N_7577,N_7620);
nor U8532 (N_8532,N_7314,N_7942);
nor U8533 (N_8533,N_7141,N_7252);
nand U8534 (N_8534,N_7739,N_7336);
and U8535 (N_8535,N_7447,N_7752);
or U8536 (N_8536,N_7251,N_7428);
and U8537 (N_8537,N_7786,N_7824);
and U8538 (N_8538,N_7725,N_7213);
or U8539 (N_8539,N_7457,N_7469);
nand U8540 (N_8540,N_7716,N_7332);
nor U8541 (N_8541,N_7840,N_7125);
or U8542 (N_8542,N_7747,N_7209);
xor U8543 (N_8543,N_7552,N_7789);
or U8544 (N_8544,N_7165,N_7632);
and U8545 (N_8545,N_7527,N_7608);
nor U8546 (N_8546,N_7146,N_7915);
and U8547 (N_8547,N_7549,N_7990);
nor U8548 (N_8548,N_7927,N_7065);
nand U8549 (N_8549,N_7661,N_7936);
or U8550 (N_8550,N_7074,N_7605);
and U8551 (N_8551,N_7623,N_7604);
or U8552 (N_8552,N_7952,N_7130);
and U8553 (N_8553,N_7265,N_7134);
and U8554 (N_8554,N_7508,N_7973);
nand U8555 (N_8555,N_7378,N_7948);
or U8556 (N_8556,N_7918,N_7175);
nor U8557 (N_8557,N_7928,N_7299);
or U8558 (N_8558,N_7251,N_7737);
nor U8559 (N_8559,N_7278,N_7838);
nand U8560 (N_8560,N_7012,N_7338);
and U8561 (N_8561,N_7016,N_7853);
and U8562 (N_8562,N_7009,N_7509);
and U8563 (N_8563,N_7844,N_7255);
nand U8564 (N_8564,N_7158,N_7014);
nor U8565 (N_8565,N_7407,N_7312);
and U8566 (N_8566,N_7577,N_7840);
and U8567 (N_8567,N_7885,N_7346);
nor U8568 (N_8568,N_7690,N_7899);
nor U8569 (N_8569,N_7749,N_7922);
and U8570 (N_8570,N_7426,N_7733);
or U8571 (N_8571,N_7870,N_7024);
and U8572 (N_8572,N_7530,N_7021);
and U8573 (N_8573,N_7230,N_7288);
nand U8574 (N_8574,N_7329,N_7000);
and U8575 (N_8575,N_7160,N_7774);
nor U8576 (N_8576,N_7819,N_7984);
nand U8577 (N_8577,N_7488,N_7000);
nand U8578 (N_8578,N_7765,N_7053);
and U8579 (N_8579,N_7480,N_7495);
and U8580 (N_8580,N_7071,N_7317);
nor U8581 (N_8581,N_7674,N_7467);
and U8582 (N_8582,N_7787,N_7505);
and U8583 (N_8583,N_7219,N_7075);
and U8584 (N_8584,N_7039,N_7943);
nand U8585 (N_8585,N_7128,N_7716);
nand U8586 (N_8586,N_7724,N_7123);
nor U8587 (N_8587,N_7042,N_7723);
nand U8588 (N_8588,N_7702,N_7804);
and U8589 (N_8589,N_7820,N_7585);
or U8590 (N_8590,N_7675,N_7284);
and U8591 (N_8591,N_7238,N_7901);
and U8592 (N_8592,N_7910,N_7847);
or U8593 (N_8593,N_7810,N_7528);
nand U8594 (N_8594,N_7542,N_7300);
and U8595 (N_8595,N_7344,N_7960);
xnor U8596 (N_8596,N_7247,N_7277);
nor U8597 (N_8597,N_7849,N_7655);
or U8598 (N_8598,N_7498,N_7356);
or U8599 (N_8599,N_7045,N_7816);
nand U8600 (N_8600,N_7689,N_7097);
or U8601 (N_8601,N_7663,N_7155);
nor U8602 (N_8602,N_7018,N_7567);
nor U8603 (N_8603,N_7386,N_7681);
or U8604 (N_8604,N_7720,N_7119);
nor U8605 (N_8605,N_7792,N_7987);
nor U8606 (N_8606,N_7414,N_7685);
nor U8607 (N_8607,N_7562,N_7697);
nor U8608 (N_8608,N_7917,N_7607);
or U8609 (N_8609,N_7243,N_7590);
and U8610 (N_8610,N_7230,N_7151);
nor U8611 (N_8611,N_7049,N_7394);
nand U8612 (N_8612,N_7410,N_7130);
and U8613 (N_8613,N_7342,N_7924);
or U8614 (N_8614,N_7079,N_7000);
or U8615 (N_8615,N_7049,N_7029);
or U8616 (N_8616,N_7554,N_7259);
nor U8617 (N_8617,N_7986,N_7983);
and U8618 (N_8618,N_7590,N_7995);
and U8619 (N_8619,N_7918,N_7599);
or U8620 (N_8620,N_7473,N_7687);
and U8621 (N_8621,N_7287,N_7352);
and U8622 (N_8622,N_7914,N_7631);
and U8623 (N_8623,N_7355,N_7335);
nor U8624 (N_8624,N_7349,N_7858);
nor U8625 (N_8625,N_7842,N_7296);
and U8626 (N_8626,N_7869,N_7283);
nand U8627 (N_8627,N_7201,N_7733);
nor U8628 (N_8628,N_7724,N_7288);
or U8629 (N_8629,N_7953,N_7425);
nand U8630 (N_8630,N_7823,N_7079);
nand U8631 (N_8631,N_7499,N_7469);
and U8632 (N_8632,N_7063,N_7985);
nor U8633 (N_8633,N_7544,N_7827);
and U8634 (N_8634,N_7738,N_7243);
nor U8635 (N_8635,N_7288,N_7599);
or U8636 (N_8636,N_7108,N_7964);
xnor U8637 (N_8637,N_7621,N_7597);
nor U8638 (N_8638,N_7162,N_7061);
and U8639 (N_8639,N_7929,N_7378);
nor U8640 (N_8640,N_7200,N_7341);
nor U8641 (N_8641,N_7043,N_7603);
nand U8642 (N_8642,N_7863,N_7672);
nand U8643 (N_8643,N_7742,N_7590);
nand U8644 (N_8644,N_7493,N_7398);
xor U8645 (N_8645,N_7053,N_7492);
or U8646 (N_8646,N_7661,N_7729);
or U8647 (N_8647,N_7914,N_7025);
xnor U8648 (N_8648,N_7384,N_7129);
nand U8649 (N_8649,N_7908,N_7544);
and U8650 (N_8650,N_7330,N_7745);
xor U8651 (N_8651,N_7263,N_7345);
and U8652 (N_8652,N_7591,N_7670);
and U8653 (N_8653,N_7223,N_7749);
and U8654 (N_8654,N_7585,N_7626);
and U8655 (N_8655,N_7566,N_7074);
nor U8656 (N_8656,N_7232,N_7778);
or U8657 (N_8657,N_7047,N_7501);
nand U8658 (N_8658,N_7869,N_7432);
nor U8659 (N_8659,N_7165,N_7642);
and U8660 (N_8660,N_7718,N_7781);
nor U8661 (N_8661,N_7115,N_7118);
nor U8662 (N_8662,N_7725,N_7861);
or U8663 (N_8663,N_7398,N_7189);
or U8664 (N_8664,N_7278,N_7584);
nand U8665 (N_8665,N_7825,N_7436);
or U8666 (N_8666,N_7874,N_7979);
or U8667 (N_8667,N_7804,N_7080);
or U8668 (N_8668,N_7038,N_7762);
and U8669 (N_8669,N_7418,N_7424);
and U8670 (N_8670,N_7727,N_7060);
or U8671 (N_8671,N_7429,N_7836);
nor U8672 (N_8672,N_7002,N_7795);
xor U8673 (N_8673,N_7977,N_7478);
or U8674 (N_8674,N_7880,N_7213);
nand U8675 (N_8675,N_7117,N_7995);
or U8676 (N_8676,N_7071,N_7319);
nand U8677 (N_8677,N_7024,N_7927);
nand U8678 (N_8678,N_7127,N_7813);
and U8679 (N_8679,N_7938,N_7642);
nor U8680 (N_8680,N_7745,N_7808);
nor U8681 (N_8681,N_7501,N_7614);
nor U8682 (N_8682,N_7979,N_7423);
nand U8683 (N_8683,N_7861,N_7489);
nor U8684 (N_8684,N_7647,N_7600);
and U8685 (N_8685,N_7686,N_7930);
and U8686 (N_8686,N_7621,N_7926);
nand U8687 (N_8687,N_7267,N_7637);
nand U8688 (N_8688,N_7387,N_7709);
and U8689 (N_8689,N_7653,N_7067);
or U8690 (N_8690,N_7066,N_7138);
nor U8691 (N_8691,N_7709,N_7137);
and U8692 (N_8692,N_7623,N_7694);
and U8693 (N_8693,N_7964,N_7846);
nand U8694 (N_8694,N_7516,N_7276);
or U8695 (N_8695,N_7191,N_7751);
nand U8696 (N_8696,N_7823,N_7710);
and U8697 (N_8697,N_7224,N_7677);
or U8698 (N_8698,N_7059,N_7663);
and U8699 (N_8699,N_7674,N_7838);
nand U8700 (N_8700,N_7277,N_7330);
or U8701 (N_8701,N_7916,N_7574);
nor U8702 (N_8702,N_7001,N_7543);
nor U8703 (N_8703,N_7140,N_7022);
nor U8704 (N_8704,N_7822,N_7763);
nor U8705 (N_8705,N_7480,N_7563);
nor U8706 (N_8706,N_7488,N_7760);
and U8707 (N_8707,N_7623,N_7855);
nor U8708 (N_8708,N_7555,N_7850);
nand U8709 (N_8709,N_7991,N_7858);
nand U8710 (N_8710,N_7944,N_7669);
nor U8711 (N_8711,N_7875,N_7621);
and U8712 (N_8712,N_7386,N_7321);
and U8713 (N_8713,N_7753,N_7467);
or U8714 (N_8714,N_7041,N_7620);
nor U8715 (N_8715,N_7238,N_7893);
and U8716 (N_8716,N_7199,N_7829);
nor U8717 (N_8717,N_7989,N_7864);
xor U8718 (N_8718,N_7129,N_7302);
and U8719 (N_8719,N_7637,N_7256);
nand U8720 (N_8720,N_7596,N_7389);
nand U8721 (N_8721,N_7822,N_7640);
or U8722 (N_8722,N_7823,N_7738);
and U8723 (N_8723,N_7751,N_7612);
and U8724 (N_8724,N_7144,N_7624);
nor U8725 (N_8725,N_7747,N_7893);
nand U8726 (N_8726,N_7065,N_7540);
or U8727 (N_8727,N_7595,N_7211);
or U8728 (N_8728,N_7093,N_7094);
nand U8729 (N_8729,N_7066,N_7393);
nand U8730 (N_8730,N_7603,N_7714);
nor U8731 (N_8731,N_7534,N_7614);
nor U8732 (N_8732,N_7074,N_7823);
nand U8733 (N_8733,N_7177,N_7375);
and U8734 (N_8734,N_7491,N_7447);
or U8735 (N_8735,N_7437,N_7266);
nor U8736 (N_8736,N_7622,N_7748);
nand U8737 (N_8737,N_7726,N_7724);
nor U8738 (N_8738,N_7338,N_7008);
nor U8739 (N_8739,N_7680,N_7473);
nor U8740 (N_8740,N_7487,N_7859);
nor U8741 (N_8741,N_7909,N_7672);
nand U8742 (N_8742,N_7387,N_7647);
or U8743 (N_8743,N_7933,N_7235);
or U8744 (N_8744,N_7232,N_7427);
nor U8745 (N_8745,N_7331,N_7687);
or U8746 (N_8746,N_7511,N_7456);
nor U8747 (N_8747,N_7185,N_7224);
nand U8748 (N_8748,N_7475,N_7915);
nand U8749 (N_8749,N_7271,N_7247);
nor U8750 (N_8750,N_7900,N_7130);
nor U8751 (N_8751,N_7244,N_7943);
or U8752 (N_8752,N_7132,N_7048);
nand U8753 (N_8753,N_7526,N_7980);
nor U8754 (N_8754,N_7066,N_7864);
and U8755 (N_8755,N_7531,N_7422);
nand U8756 (N_8756,N_7037,N_7608);
or U8757 (N_8757,N_7205,N_7107);
nor U8758 (N_8758,N_7058,N_7806);
nor U8759 (N_8759,N_7451,N_7799);
and U8760 (N_8760,N_7403,N_7354);
or U8761 (N_8761,N_7020,N_7710);
and U8762 (N_8762,N_7114,N_7491);
and U8763 (N_8763,N_7241,N_7464);
nor U8764 (N_8764,N_7397,N_7763);
nor U8765 (N_8765,N_7943,N_7095);
and U8766 (N_8766,N_7807,N_7216);
or U8767 (N_8767,N_7105,N_7810);
or U8768 (N_8768,N_7156,N_7862);
xnor U8769 (N_8769,N_7643,N_7336);
nor U8770 (N_8770,N_7035,N_7481);
and U8771 (N_8771,N_7618,N_7201);
nor U8772 (N_8772,N_7874,N_7158);
nand U8773 (N_8773,N_7275,N_7796);
nand U8774 (N_8774,N_7012,N_7040);
nand U8775 (N_8775,N_7585,N_7858);
and U8776 (N_8776,N_7402,N_7953);
or U8777 (N_8777,N_7728,N_7373);
or U8778 (N_8778,N_7386,N_7583);
or U8779 (N_8779,N_7489,N_7257);
or U8780 (N_8780,N_7290,N_7863);
nand U8781 (N_8781,N_7681,N_7464);
nor U8782 (N_8782,N_7102,N_7212);
and U8783 (N_8783,N_7707,N_7218);
nand U8784 (N_8784,N_7680,N_7685);
nand U8785 (N_8785,N_7788,N_7921);
or U8786 (N_8786,N_7939,N_7661);
or U8787 (N_8787,N_7872,N_7586);
nor U8788 (N_8788,N_7582,N_7027);
nor U8789 (N_8789,N_7674,N_7775);
nand U8790 (N_8790,N_7728,N_7995);
and U8791 (N_8791,N_7734,N_7883);
and U8792 (N_8792,N_7309,N_7770);
nor U8793 (N_8793,N_7429,N_7578);
nand U8794 (N_8794,N_7025,N_7193);
nand U8795 (N_8795,N_7528,N_7374);
nand U8796 (N_8796,N_7184,N_7196);
nor U8797 (N_8797,N_7133,N_7197);
nor U8798 (N_8798,N_7457,N_7410);
and U8799 (N_8799,N_7913,N_7486);
and U8800 (N_8800,N_7549,N_7725);
nor U8801 (N_8801,N_7913,N_7090);
or U8802 (N_8802,N_7315,N_7549);
or U8803 (N_8803,N_7348,N_7638);
and U8804 (N_8804,N_7882,N_7236);
nand U8805 (N_8805,N_7109,N_7378);
nor U8806 (N_8806,N_7264,N_7428);
nor U8807 (N_8807,N_7465,N_7520);
and U8808 (N_8808,N_7663,N_7689);
nor U8809 (N_8809,N_7983,N_7813);
nand U8810 (N_8810,N_7596,N_7179);
xnor U8811 (N_8811,N_7942,N_7808);
nand U8812 (N_8812,N_7543,N_7731);
nand U8813 (N_8813,N_7152,N_7022);
and U8814 (N_8814,N_7757,N_7686);
nor U8815 (N_8815,N_7349,N_7102);
or U8816 (N_8816,N_7429,N_7478);
nand U8817 (N_8817,N_7868,N_7618);
nand U8818 (N_8818,N_7758,N_7815);
nor U8819 (N_8819,N_7988,N_7601);
xor U8820 (N_8820,N_7489,N_7967);
nor U8821 (N_8821,N_7977,N_7416);
or U8822 (N_8822,N_7341,N_7315);
and U8823 (N_8823,N_7779,N_7153);
or U8824 (N_8824,N_7065,N_7813);
and U8825 (N_8825,N_7202,N_7389);
nor U8826 (N_8826,N_7259,N_7810);
or U8827 (N_8827,N_7951,N_7599);
and U8828 (N_8828,N_7289,N_7502);
and U8829 (N_8829,N_7586,N_7418);
and U8830 (N_8830,N_7663,N_7936);
nand U8831 (N_8831,N_7193,N_7149);
nor U8832 (N_8832,N_7488,N_7716);
nand U8833 (N_8833,N_7928,N_7306);
and U8834 (N_8834,N_7735,N_7628);
nor U8835 (N_8835,N_7296,N_7072);
nand U8836 (N_8836,N_7344,N_7525);
or U8837 (N_8837,N_7496,N_7031);
nor U8838 (N_8838,N_7558,N_7628);
and U8839 (N_8839,N_7655,N_7984);
and U8840 (N_8840,N_7019,N_7840);
nor U8841 (N_8841,N_7068,N_7347);
and U8842 (N_8842,N_7061,N_7261);
or U8843 (N_8843,N_7630,N_7858);
nor U8844 (N_8844,N_7584,N_7000);
or U8845 (N_8845,N_7788,N_7276);
nand U8846 (N_8846,N_7645,N_7103);
or U8847 (N_8847,N_7207,N_7450);
and U8848 (N_8848,N_7327,N_7734);
and U8849 (N_8849,N_7557,N_7622);
nor U8850 (N_8850,N_7697,N_7946);
nand U8851 (N_8851,N_7111,N_7430);
and U8852 (N_8852,N_7626,N_7541);
nand U8853 (N_8853,N_7355,N_7986);
and U8854 (N_8854,N_7128,N_7180);
and U8855 (N_8855,N_7451,N_7918);
and U8856 (N_8856,N_7038,N_7381);
and U8857 (N_8857,N_7423,N_7704);
and U8858 (N_8858,N_7318,N_7255);
and U8859 (N_8859,N_7413,N_7496);
nor U8860 (N_8860,N_7468,N_7987);
or U8861 (N_8861,N_7908,N_7791);
or U8862 (N_8862,N_7550,N_7264);
or U8863 (N_8863,N_7274,N_7163);
nor U8864 (N_8864,N_7837,N_7083);
and U8865 (N_8865,N_7749,N_7274);
nor U8866 (N_8866,N_7536,N_7458);
or U8867 (N_8867,N_7699,N_7742);
nand U8868 (N_8868,N_7543,N_7657);
and U8869 (N_8869,N_7310,N_7406);
nand U8870 (N_8870,N_7282,N_7468);
nor U8871 (N_8871,N_7308,N_7459);
and U8872 (N_8872,N_7748,N_7306);
nor U8873 (N_8873,N_7690,N_7287);
nor U8874 (N_8874,N_7798,N_7668);
nand U8875 (N_8875,N_7835,N_7490);
nor U8876 (N_8876,N_7029,N_7722);
nand U8877 (N_8877,N_7439,N_7625);
and U8878 (N_8878,N_7529,N_7061);
or U8879 (N_8879,N_7577,N_7449);
and U8880 (N_8880,N_7155,N_7115);
and U8881 (N_8881,N_7308,N_7560);
nand U8882 (N_8882,N_7863,N_7867);
nor U8883 (N_8883,N_7398,N_7582);
nand U8884 (N_8884,N_7664,N_7842);
nor U8885 (N_8885,N_7566,N_7462);
nand U8886 (N_8886,N_7337,N_7476);
nand U8887 (N_8887,N_7914,N_7515);
nand U8888 (N_8888,N_7050,N_7863);
nor U8889 (N_8889,N_7452,N_7064);
and U8890 (N_8890,N_7466,N_7338);
and U8891 (N_8891,N_7476,N_7599);
and U8892 (N_8892,N_7684,N_7760);
or U8893 (N_8893,N_7478,N_7752);
nand U8894 (N_8894,N_7540,N_7257);
nor U8895 (N_8895,N_7323,N_7456);
nor U8896 (N_8896,N_7438,N_7950);
or U8897 (N_8897,N_7371,N_7443);
or U8898 (N_8898,N_7648,N_7557);
nor U8899 (N_8899,N_7495,N_7072);
nor U8900 (N_8900,N_7584,N_7696);
and U8901 (N_8901,N_7036,N_7241);
nor U8902 (N_8902,N_7204,N_7883);
and U8903 (N_8903,N_7736,N_7423);
and U8904 (N_8904,N_7416,N_7856);
or U8905 (N_8905,N_7691,N_7639);
nand U8906 (N_8906,N_7841,N_7161);
nand U8907 (N_8907,N_7642,N_7032);
xor U8908 (N_8908,N_7234,N_7293);
and U8909 (N_8909,N_7462,N_7033);
or U8910 (N_8910,N_7905,N_7574);
nor U8911 (N_8911,N_7752,N_7913);
nand U8912 (N_8912,N_7537,N_7129);
nand U8913 (N_8913,N_7244,N_7225);
nor U8914 (N_8914,N_7032,N_7095);
nor U8915 (N_8915,N_7011,N_7321);
xor U8916 (N_8916,N_7406,N_7218);
or U8917 (N_8917,N_7637,N_7456);
or U8918 (N_8918,N_7300,N_7649);
xnor U8919 (N_8919,N_7857,N_7297);
nor U8920 (N_8920,N_7601,N_7886);
xnor U8921 (N_8921,N_7789,N_7779);
nand U8922 (N_8922,N_7385,N_7404);
and U8923 (N_8923,N_7232,N_7313);
nor U8924 (N_8924,N_7161,N_7108);
nor U8925 (N_8925,N_7791,N_7286);
nor U8926 (N_8926,N_7367,N_7444);
or U8927 (N_8927,N_7734,N_7650);
and U8928 (N_8928,N_7029,N_7350);
or U8929 (N_8929,N_7642,N_7822);
nor U8930 (N_8930,N_7216,N_7629);
or U8931 (N_8931,N_7427,N_7514);
nor U8932 (N_8932,N_7515,N_7193);
nor U8933 (N_8933,N_7703,N_7125);
nor U8934 (N_8934,N_7896,N_7963);
xor U8935 (N_8935,N_7665,N_7094);
nor U8936 (N_8936,N_7150,N_7197);
xnor U8937 (N_8937,N_7641,N_7881);
or U8938 (N_8938,N_7044,N_7333);
and U8939 (N_8939,N_7897,N_7448);
or U8940 (N_8940,N_7559,N_7055);
nand U8941 (N_8941,N_7041,N_7658);
or U8942 (N_8942,N_7731,N_7223);
and U8943 (N_8943,N_7966,N_7789);
nand U8944 (N_8944,N_7870,N_7626);
nand U8945 (N_8945,N_7843,N_7663);
or U8946 (N_8946,N_7230,N_7466);
nand U8947 (N_8947,N_7027,N_7274);
nor U8948 (N_8948,N_7769,N_7321);
or U8949 (N_8949,N_7480,N_7950);
nand U8950 (N_8950,N_7003,N_7404);
and U8951 (N_8951,N_7321,N_7185);
xor U8952 (N_8952,N_7536,N_7925);
and U8953 (N_8953,N_7926,N_7009);
nor U8954 (N_8954,N_7765,N_7436);
and U8955 (N_8955,N_7685,N_7517);
or U8956 (N_8956,N_7226,N_7023);
nand U8957 (N_8957,N_7902,N_7245);
nand U8958 (N_8958,N_7519,N_7243);
nand U8959 (N_8959,N_7723,N_7187);
nand U8960 (N_8960,N_7191,N_7437);
nor U8961 (N_8961,N_7343,N_7789);
and U8962 (N_8962,N_7717,N_7723);
xnor U8963 (N_8963,N_7124,N_7290);
and U8964 (N_8964,N_7027,N_7531);
and U8965 (N_8965,N_7193,N_7976);
nor U8966 (N_8966,N_7474,N_7186);
and U8967 (N_8967,N_7159,N_7161);
nor U8968 (N_8968,N_7950,N_7338);
and U8969 (N_8969,N_7102,N_7244);
nand U8970 (N_8970,N_7851,N_7303);
nor U8971 (N_8971,N_7728,N_7139);
nor U8972 (N_8972,N_7755,N_7721);
nand U8973 (N_8973,N_7822,N_7369);
or U8974 (N_8974,N_7402,N_7463);
nor U8975 (N_8975,N_7335,N_7252);
or U8976 (N_8976,N_7178,N_7507);
and U8977 (N_8977,N_7249,N_7393);
nand U8978 (N_8978,N_7530,N_7370);
or U8979 (N_8979,N_7773,N_7727);
or U8980 (N_8980,N_7153,N_7749);
nand U8981 (N_8981,N_7920,N_7881);
nand U8982 (N_8982,N_7988,N_7994);
nand U8983 (N_8983,N_7673,N_7115);
nand U8984 (N_8984,N_7410,N_7617);
or U8985 (N_8985,N_7318,N_7848);
and U8986 (N_8986,N_7617,N_7512);
nand U8987 (N_8987,N_7053,N_7318);
and U8988 (N_8988,N_7980,N_7791);
nand U8989 (N_8989,N_7072,N_7655);
xor U8990 (N_8990,N_7324,N_7297);
or U8991 (N_8991,N_7262,N_7472);
or U8992 (N_8992,N_7421,N_7694);
nor U8993 (N_8993,N_7246,N_7838);
or U8994 (N_8994,N_7892,N_7381);
and U8995 (N_8995,N_7345,N_7785);
nand U8996 (N_8996,N_7975,N_7244);
nor U8997 (N_8997,N_7908,N_7069);
nand U8998 (N_8998,N_7521,N_7308);
nand U8999 (N_8999,N_7930,N_7357);
and U9000 (N_9000,N_8161,N_8249);
nand U9001 (N_9001,N_8116,N_8135);
nor U9002 (N_9002,N_8827,N_8766);
nand U9003 (N_9003,N_8420,N_8687);
and U9004 (N_9004,N_8303,N_8950);
nor U9005 (N_9005,N_8921,N_8137);
and U9006 (N_9006,N_8009,N_8638);
or U9007 (N_9007,N_8835,N_8418);
and U9008 (N_9008,N_8098,N_8439);
or U9009 (N_9009,N_8389,N_8778);
nand U9010 (N_9010,N_8357,N_8901);
xor U9011 (N_9011,N_8524,N_8525);
and U9012 (N_9012,N_8772,N_8550);
nand U9013 (N_9013,N_8804,N_8539);
or U9014 (N_9014,N_8870,N_8682);
nor U9015 (N_9015,N_8604,N_8779);
or U9016 (N_9016,N_8654,N_8724);
or U9017 (N_9017,N_8500,N_8468);
or U9018 (N_9018,N_8898,N_8603);
or U9019 (N_9019,N_8690,N_8072);
and U9020 (N_9020,N_8636,N_8821);
nand U9021 (N_9021,N_8347,N_8973);
nor U9022 (N_9022,N_8353,N_8928);
nor U9023 (N_9023,N_8419,N_8570);
or U9024 (N_9024,N_8286,N_8554);
nand U9025 (N_9025,N_8120,N_8815);
and U9026 (N_9026,N_8018,N_8769);
nand U9027 (N_9027,N_8958,N_8021);
and U9028 (N_9028,N_8014,N_8482);
or U9029 (N_9029,N_8041,N_8894);
nor U9030 (N_9030,N_8872,N_8523);
nand U9031 (N_9031,N_8475,N_8071);
xnor U9032 (N_9032,N_8534,N_8093);
nand U9033 (N_9033,N_8794,N_8269);
nor U9034 (N_9034,N_8572,N_8226);
nand U9035 (N_9035,N_8885,N_8503);
and U9036 (N_9036,N_8774,N_8460);
nor U9037 (N_9037,N_8514,N_8734);
and U9038 (N_9038,N_8171,N_8229);
or U9039 (N_9039,N_8355,N_8810);
and U9040 (N_9040,N_8981,N_8732);
nor U9041 (N_9041,N_8531,N_8281);
nor U9042 (N_9042,N_8843,N_8753);
or U9043 (N_9043,N_8028,N_8092);
and U9044 (N_9044,N_8711,N_8264);
nand U9045 (N_9045,N_8624,N_8727);
nor U9046 (N_9046,N_8304,N_8702);
nor U9047 (N_9047,N_8469,N_8031);
or U9048 (N_9048,N_8719,N_8490);
and U9049 (N_9049,N_8549,N_8933);
nor U9050 (N_9050,N_8838,N_8956);
nand U9051 (N_9051,N_8090,N_8609);
nor U9052 (N_9052,N_8984,N_8723);
and U9053 (N_9053,N_8398,N_8217);
or U9054 (N_9054,N_8592,N_8785);
or U9055 (N_9055,N_8333,N_8083);
nand U9056 (N_9056,N_8813,N_8825);
and U9057 (N_9057,N_8218,N_8052);
nand U9058 (N_9058,N_8253,N_8105);
and U9059 (N_9059,N_8138,N_8075);
and U9060 (N_9060,N_8287,N_8438);
or U9061 (N_9061,N_8940,N_8081);
nor U9062 (N_9062,N_8240,N_8951);
nand U9063 (N_9063,N_8782,N_8430);
nor U9064 (N_9064,N_8507,N_8393);
and U9065 (N_9065,N_8803,N_8991);
nand U9066 (N_9066,N_8112,N_8095);
and U9067 (N_9067,N_8656,N_8833);
xnor U9068 (N_9068,N_8911,N_8074);
or U9069 (N_9069,N_8338,N_8808);
and U9070 (N_9070,N_8474,N_8372);
nand U9071 (N_9071,N_8150,N_8859);
and U9072 (N_9072,N_8521,N_8194);
or U9073 (N_9073,N_8513,N_8883);
nand U9074 (N_9074,N_8056,N_8849);
and U9075 (N_9075,N_8526,N_8713);
and U9076 (N_9076,N_8899,N_8718);
nand U9077 (N_9077,N_8458,N_8577);
and U9078 (N_9078,N_8557,N_8164);
or U9079 (N_9079,N_8392,N_8605);
nor U9080 (N_9080,N_8561,N_8729);
nor U9081 (N_9081,N_8446,N_8280);
nand U9082 (N_9082,N_8565,N_8325);
nand U9083 (N_9083,N_8851,N_8747);
nor U9084 (N_9084,N_8809,N_8427);
nand U9085 (N_9085,N_8027,N_8254);
or U9086 (N_9086,N_8348,N_8972);
and U9087 (N_9087,N_8457,N_8662);
and U9088 (N_9088,N_8387,N_8937);
or U9089 (N_9089,N_8587,N_8907);
nor U9090 (N_9090,N_8974,N_8674);
xor U9091 (N_9091,N_8154,N_8611);
nor U9092 (N_9092,N_8677,N_8967);
and U9093 (N_9093,N_8616,N_8332);
nor U9094 (N_9094,N_8001,N_8961);
nor U9095 (N_9095,N_8339,N_8118);
nor U9096 (N_9096,N_8932,N_8995);
and U9097 (N_9097,N_8544,N_8238);
nand U9098 (N_9098,N_8631,N_8764);
or U9099 (N_9099,N_8943,N_8672);
or U9100 (N_9100,N_8600,N_8011);
or U9101 (N_9101,N_8777,N_8910);
nor U9102 (N_9102,N_8228,N_8016);
nand U9103 (N_9103,N_8012,N_8757);
nand U9104 (N_9104,N_8990,N_8741);
nor U9105 (N_9105,N_8743,N_8294);
nand U9106 (N_9106,N_8936,N_8593);
or U9107 (N_9107,N_8265,N_8789);
nor U9108 (N_9108,N_8013,N_8395);
and U9109 (N_9109,N_8560,N_8767);
nor U9110 (N_9110,N_8874,N_8158);
nor U9111 (N_9111,N_8640,N_8415);
or U9112 (N_9112,N_8176,N_8046);
nor U9113 (N_9113,N_8296,N_8620);
nor U9114 (N_9114,N_8661,N_8520);
nor U9115 (N_9115,N_8407,N_8607);
nor U9116 (N_9116,N_8410,N_8752);
or U9117 (N_9117,N_8509,N_8220);
and U9118 (N_9118,N_8632,N_8136);
nand U9119 (N_9119,N_8517,N_8742);
or U9120 (N_9120,N_8246,N_8884);
xnor U9121 (N_9121,N_8165,N_8394);
and U9122 (N_9122,N_8391,N_8192);
or U9123 (N_9123,N_8431,N_8411);
nand U9124 (N_9124,N_8771,N_8856);
and U9125 (N_9125,N_8613,N_8447);
nor U9126 (N_9126,N_8660,N_8140);
nor U9127 (N_9127,N_8234,N_8614);
xnor U9128 (N_9128,N_8646,N_8643);
and U9129 (N_9129,N_8670,N_8222);
and U9130 (N_9130,N_8462,N_8519);
or U9131 (N_9131,N_8694,N_8379);
and U9132 (N_9132,N_8840,N_8080);
nand U9133 (N_9133,N_8553,N_8828);
xor U9134 (N_9134,N_8770,N_8184);
nor U9135 (N_9135,N_8814,N_8230);
nor U9136 (N_9136,N_8726,N_8902);
nand U9137 (N_9137,N_8309,N_8486);
and U9138 (N_9138,N_8979,N_8032);
nor U9139 (N_9139,N_8606,N_8584);
nand U9140 (N_9140,N_8848,N_8054);
and U9141 (N_9141,N_8139,N_8042);
and U9142 (N_9142,N_8867,N_8798);
and U9143 (N_9143,N_8893,N_8895);
or U9144 (N_9144,N_8963,N_8669);
nand U9145 (N_9145,N_8566,N_8793);
or U9146 (N_9146,N_8038,N_8417);
and U9147 (N_9147,N_8985,N_8231);
nand U9148 (N_9148,N_8683,N_8594);
nand U9149 (N_9149,N_8459,N_8705);
nand U9150 (N_9150,N_8652,N_8316);
or U9151 (N_9151,N_8084,N_8567);
nor U9152 (N_9152,N_8015,N_8877);
nand U9153 (N_9153,N_8295,N_8562);
and U9154 (N_9154,N_8059,N_8343);
or U9155 (N_9155,N_8225,N_8575);
nor U9156 (N_9156,N_8173,N_8598);
or U9157 (N_9157,N_8079,N_8436);
nor U9158 (N_9158,N_8920,N_8649);
nand U9159 (N_9159,N_8552,N_8679);
and U9160 (N_9160,N_8994,N_8927);
or U9161 (N_9161,N_8149,N_8002);
xnor U9162 (N_9162,N_8545,N_8706);
nor U9163 (N_9163,N_8388,N_8659);
and U9164 (N_9164,N_8077,N_8929);
or U9165 (N_9165,N_8712,N_8452);
or U9166 (N_9166,N_8630,N_8515);
nand U9167 (N_9167,N_8678,N_8744);
nand U9168 (N_9168,N_8700,N_8058);
xor U9169 (N_9169,N_8698,N_8276);
or U9170 (N_9170,N_8128,N_8908);
or U9171 (N_9171,N_8044,N_8471);
or U9172 (N_9172,N_8987,N_8917);
nand U9173 (N_9173,N_8982,N_8548);
and U9174 (N_9174,N_8998,N_8073);
nand U9175 (N_9175,N_8671,N_8257);
nor U9176 (N_9176,N_8461,N_8996);
or U9177 (N_9177,N_8914,N_8369);
and U9178 (N_9178,N_8209,N_8924);
or U9179 (N_9179,N_8761,N_8381);
or U9180 (N_9180,N_8107,N_8106);
or U9181 (N_9181,N_8615,N_8978);
and U9182 (N_9182,N_8125,N_8337);
nand U9183 (N_9183,N_8273,N_8201);
and U9184 (N_9184,N_8722,N_8335);
nand U9185 (N_9185,N_8426,N_8977);
xor U9186 (N_9186,N_8177,N_8290);
nor U9187 (N_9187,N_8836,N_8714);
nand U9188 (N_9188,N_8242,N_8181);
nor U9189 (N_9189,N_8454,N_8555);
and U9190 (N_9190,N_8875,N_8360);
and U9191 (N_9191,N_8024,N_8368);
or U9192 (N_9192,N_8935,N_8297);
nand U9193 (N_9193,N_8324,N_8196);
nand U9194 (N_9194,N_8506,N_8481);
nand U9195 (N_9195,N_8292,N_8829);
nand U9196 (N_9196,N_8658,N_8402);
nand U9197 (N_9197,N_8900,N_8288);
and U9198 (N_9198,N_8408,N_8183);
or U9199 (N_9199,N_8378,N_8628);
nand U9200 (N_9200,N_8302,N_8501);
or U9201 (N_9201,N_8617,N_8344);
and U9202 (N_9202,N_8146,N_8852);
nor U9203 (N_9203,N_8237,N_8170);
nor U9204 (N_9204,N_8760,N_8478);
or U9205 (N_9205,N_8413,N_8251);
or U9206 (N_9206,N_8445,N_8844);
and U9207 (N_9207,N_8113,N_8807);
nor U9208 (N_9208,N_8190,N_8608);
nor U9209 (N_9209,N_8350,N_8686);
or U9210 (N_9210,N_8377,N_8871);
or U9211 (N_9211,N_8094,N_8897);
and U9212 (N_9212,N_8868,N_8167);
nand U9213 (N_9213,N_8853,N_8941);
or U9214 (N_9214,N_8831,N_8494);
nand U9215 (N_9215,N_8863,N_8189);
and U9216 (N_9216,N_8876,N_8375);
nand U9217 (N_9217,N_8045,N_8980);
and U9218 (N_9218,N_8641,N_8285);
or U9219 (N_9219,N_8437,N_8925);
or U9220 (N_9220,N_8429,N_8055);
nor U9221 (N_9221,N_8299,N_8684);
nand U9222 (N_9222,N_8953,N_8114);
nand U9223 (N_9223,N_8571,N_8005);
nand U9224 (N_9224,N_8733,N_8959);
and U9225 (N_9225,N_8127,N_8076);
or U9226 (N_9226,N_8270,N_8213);
and U9227 (N_9227,N_8811,N_8108);
xor U9228 (N_9228,N_8409,N_8040);
nor U9229 (N_9229,N_8019,N_8905);
nor U9230 (N_9230,N_8971,N_8826);
nor U9231 (N_9231,N_8414,N_8653);
and U9232 (N_9232,N_8464,N_8330);
xnor U9233 (N_9233,N_8119,N_8799);
or U9234 (N_9234,N_8788,N_8354);
nand U9235 (N_9235,N_8992,N_8960);
nand U9236 (N_9236,N_8688,N_8952);
and U9237 (N_9237,N_8881,N_8730);
nor U9238 (N_9238,N_8147,N_8634);
and U9239 (N_9239,N_8745,N_8748);
nor U9240 (N_9240,N_8385,N_8358);
nor U9241 (N_9241,N_8896,N_8006);
nor U9242 (N_9242,N_8675,N_8647);
or U9243 (N_9243,N_8637,N_8882);
nor U9244 (N_9244,N_8585,N_8491);
nand U9245 (N_9245,N_8144,N_8948);
nand U9246 (N_9246,N_8252,N_8780);
or U9247 (N_9247,N_8017,N_8199);
and U9248 (N_9248,N_8195,N_8546);
nor U9249 (N_9249,N_8578,N_8866);
and U9250 (N_9250,N_8758,N_8432);
nand U9251 (N_9251,N_8180,N_8666);
or U9252 (N_9252,N_8708,N_8148);
nand U9253 (N_9253,N_8086,N_8440);
or U9254 (N_9254,N_8997,N_8168);
nor U9255 (N_9255,N_8612,N_8533);
nor U9256 (N_9256,N_8236,N_8340);
nand U9257 (N_9257,N_8131,N_8142);
nor U9258 (N_9258,N_8528,N_8942);
nor U9259 (N_9259,N_8421,N_8890);
or U9260 (N_9260,N_8004,N_8205);
or U9261 (N_9261,N_8716,N_8923);
nand U9262 (N_9262,N_8162,N_8122);
nor U9263 (N_9263,N_8435,N_8480);
nand U9264 (N_9264,N_8159,N_8823);
nand U9265 (N_9265,N_8663,N_8855);
and U9266 (N_9266,N_8858,N_8400);
or U9267 (N_9267,N_8256,N_8000);
and U9268 (N_9268,N_8166,N_8200);
and U9269 (N_9269,N_8068,N_8621);
nand U9270 (N_9270,N_8361,N_8709);
nor U9271 (N_9271,N_8370,N_8864);
xnor U9272 (N_9272,N_8371,N_8130);
xnor U9273 (N_9273,N_8484,N_8703);
nor U9274 (N_9274,N_8622,N_8488);
and U9275 (N_9275,N_8655,N_8223);
nand U9276 (N_9276,N_8219,N_8300);
nand U9277 (N_9277,N_8022,N_8078);
nand U9278 (N_9278,N_8913,N_8720);
or U9279 (N_9279,N_8644,N_8916);
nand U9280 (N_9280,N_8845,N_8541);
and U9281 (N_9281,N_8267,N_8047);
or U9282 (N_9282,N_8573,N_8126);
nor U9283 (N_9283,N_8097,N_8060);
nor U9284 (N_9284,N_8477,N_8062);
or U9285 (N_9285,N_8311,N_8336);
nor U9286 (N_9286,N_8352,N_8211);
nand U9287 (N_9287,N_8765,N_8441);
nand U9288 (N_9288,N_8839,N_8499);
and U9289 (N_9289,N_8988,N_8384);
nand U9290 (N_9290,N_8962,N_8160);
nand U9291 (N_9291,N_8989,N_8915);
and U9292 (N_9292,N_8854,N_8736);
or U9293 (N_9293,N_8100,N_8390);
nand U9294 (N_9294,N_8847,N_8543);
or U9295 (N_9295,N_8846,N_8918);
and U9296 (N_9296,N_8033,N_8401);
and U9297 (N_9297,N_8717,N_8132);
nand U9298 (N_9298,N_8197,N_8003);
nand U9299 (N_9299,N_8404,N_8102);
and U9300 (N_9300,N_8627,N_8824);
nor U9301 (N_9301,N_8029,N_8516);
nor U9302 (N_9302,N_8949,N_8087);
and U9303 (N_9303,N_8797,N_8185);
and U9304 (N_9304,N_8133,N_8695);
nor U9305 (N_9305,N_8103,N_8363);
nand U9306 (N_9306,N_8536,N_8317);
nor U9307 (N_9307,N_8096,N_8367);
nand U9308 (N_9308,N_8954,N_8955);
or U9309 (N_9309,N_8806,N_8559);
xnor U9310 (N_9310,N_8323,N_8629);
xnor U9311 (N_9311,N_8221,N_8049);
and U9312 (N_9312,N_8889,N_8243);
nor U9313 (N_9313,N_8245,N_8064);
and U9314 (N_9314,N_8244,N_8143);
or U9315 (N_9315,N_8817,N_8596);
or U9316 (N_9316,N_8676,N_8832);
nor U9317 (N_9317,N_8156,N_8939);
or U9318 (N_9318,N_8456,N_8403);
nand U9319 (N_9319,N_8558,N_8999);
nand U9320 (N_9320,N_8433,N_8293);
or U9321 (N_9321,N_8583,N_8063);
nor U9322 (N_9322,N_8473,N_8891);
nor U9323 (N_9323,N_8976,N_8291);
nand U9324 (N_9324,N_8235,N_8007);
nand U9325 (N_9325,N_8795,N_8424);
and U9326 (N_9326,N_8749,N_8787);
nor U9327 (N_9327,N_8830,N_8618);
nand U9328 (N_9328,N_8268,N_8822);
or U9329 (N_9329,N_8470,N_8057);
nand U9330 (N_9330,N_8210,N_8926);
nand U9331 (N_9331,N_8754,N_8775);
nor U9332 (N_9332,N_8065,N_8693);
nor U9333 (N_9333,N_8050,N_8837);
or U9334 (N_9334,N_8970,N_8667);
and U9335 (N_9335,N_8680,N_8715);
or U9336 (N_9336,N_8241,N_8023);
nor U9337 (N_9337,N_8443,N_8581);
or U9338 (N_9338,N_8673,N_8444);
or U9339 (N_9339,N_8463,N_8493);
and U9340 (N_9340,N_8314,N_8505);
and U9341 (N_9341,N_8564,N_8842);
and U9342 (N_9342,N_8530,N_8301);
xnor U9343 (N_9343,N_8104,N_8610);
or U9344 (N_9344,N_8476,N_8349);
or U9345 (N_9345,N_8639,N_8425);
xnor U9346 (N_9346,N_8356,N_8152);
nand U9347 (N_9347,N_8791,N_8756);
or U9348 (N_9348,N_8483,N_8318);
and U9349 (N_9349,N_8279,N_8965);
nand U9350 (N_9350,N_8738,N_8487);
nand U9351 (N_9351,N_8322,N_8495);
and U9352 (N_9352,N_8067,N_8039);
nor U9353 (N_9353,N_8373,N_8512);
or U9354 (N_9354,N_8651,N_8232);
or U9355 (N_9355,N_8048,N_8601);
nor U9356 (N_9356,N_8862,N_8380);
and U9357 (N_9357,N_8527,N_8153);
nand U9358 (N_9358,N_8448,N_8922);
or U9359 (N_9359,N_8880,N_8428);
nor U9360 (N_9360,N_8275,N_8969);
or U9361 (N_9361,N_8310,N_8986);
nand U9362 (N_9362,N_8597,N_8212);
and U9363 (N_9363,N_8163,N_8784);
and U9364 (N_9364,N_8819,N_8912);
or U9365 (N_9365,N_8586,N_8668);
or U9366 (N_9366,N_8664,N_8707);
or U9367 (N_9367,N_8043,N_8485);
xnor U9368 (N_9368,N_8271,N_8776);
nor U9369 (N_9369,N_8472,N_8283);
and U9370 (N_9370,N_8037,N_8931);
nor U9371 (N_9371,N_8633,N_8035);
nor U9372 (N_9372,N_8975,N_8315);
and U9373 (N_9373,N_8151,N_8869);
nor U9374 (N_9374,N_8945,N_8250);
nand U9375 (N_9375,N_8366,N_8258);
nand U9376 (N_9376,N_8650,N_8834);
nor U9377 (N_9377,N_8568,N_8328);
or U9378 (N_9378,N_8202,N_8091);
and U9379 (N_9379,N_8320,N_8903);
or U9380 (N_9380,N_8266,N_8701);
nand U9381 (N_9381,N_8069,N_8648);
or U9382 (N_9382,N_8203,N_8556);
and U9383 (N_9383,N_8510,N_8532);
nand U9384 (N_9384,N_8542,N_8642);
nor U9385 (N_9385,N_8964,N_8260);
or U9386 (N_9386,N_8860,N_8878);
nor U9387 (N_9387,N_8450,N_8547);
or U9388 (N_9388,N_8326,N_8115);
nor U9389 (N_9389,N_8026,N_8247);
or U9390 (N_9390,N_8865,N_8773);
or U9391 (N_9391,N_8790,N_8262);
nor U9392 (N_9392,N_8053,N_8175);
and U9393 (N_9393,N_8820,N_8537);
nor U9394 (N_9394,N_8759,N_8331);
and U9395 (N_9395,N_8579,N_8227);
nor U9396 (N_9396,N_8697,N_8492);
or U9397 (N_9397,N_8365,N_8551);
nor U9398 (N_9398,N_8312,N_8191);
nor U9399 (N_9399,N_8689,N_8983);
or U9400 (N_9400,N_8182,N_8207);
nor U9401 (N_9401,N_8802,N_8938);
and U9402 (N_9402,N_8498,N_8416);
or U9403 (N_9403,N_8319,N_8298);
or U9404 (N_9404,N_8216,N_8904);
and U9405 (N_9405,N_8599,N_8351);
nand U9406 (N_9406,N_8313,N_8342);
nor U9407 (N_9407,N_8511,N_8763);
and U9408 (N_9408,N_8781,N_8645);
nor U9409 (N_9409,N_8259,N_8088);
nor U9410 (N_9410,N_8085,N_8272);
or U9411 (N_9411,N_8934,N_8239);
and U9412 (N_9412,N_8178,N_8755);
nand U9413 (N_9413,N_8187,N_8214);
and U9414 (N_9414,N_8740,N_8591);
and U9415 (N_9415,N_8451,N_8957);
and U9416 (N_9416,N_8930,N_8215);
nor U9417 (N_9417,N_8329,N_8224);
nand U9418 (N_9418,N_8502,N_8540);
nand U9419 (N_9419,N_8696,N_8919);
nor U9420 (N_9420,N_8796,N_8282);
and U9421 (N_9421,N_8169,N_8233);
and U9422 (N_9422,N_8725,N_8812);
nand U9423 (N_9423,N_8850,N_8665);
nand U9424 (N_9424,N_8345,N_8625);
nor U9425 (N_9425,N_8816,N_8861);
nand U9426 (N_9426,N_8946,N_8307);
nor U9427 (N_9427,N_8206,N_8685);
nand U9428 (N_9428,N_8841,N_8465);
nor U9429 (N_9429,N_8479,N_8442);
nand U9430 (N_9430,N_8186,N_8423);
nor U9431 (N_9431,N_8449,N_8422);
and U9432 (N_9432,N_8563,N_8750);
and U9433 (N_9433,N_8188,N_8386);
and U9434 (N_9434,N_8082,N_8801);
and U9435 (N_9435,N_8359,N_8731);
nand U9436 (N_9436,N_8051,N_8582);
nor U9437 (N_9437,N_8751,N_8101);
nand U9438 (N_9438,N_8590,N_8362);
nand U9439 (N_9439,N_8574,N_8595);
nor U9440 (N_9440,N_8274,N_8248);
or U9441 (N_9441,N_8879,N_8602);
nor U9442 (N_9442,N_8327,N_8121);
or U9443 (N_9443,N_8522,N_8099);
or U9444 (N_9444,N_8145,N_8396);
or U9445 (N_9445,N_8061,N_8735);
nor U9446 (N_9446,N_8489,N_8466);
and U9447 (N_9447,N_8623,N_8434);
nor U9448 (N_9448,N_8508,N_8589);
nor U9449 (N_9449,N_8947,N_8036);
nor U9450 (N_9450,N_8886,N_8635);
or U9451 (N_9451,N_8497,N_8383);
or U9452 (N_9452,N_8364,N_8405);
and U9453 (N_9453,N_8786,N_8681);
and U9454 (N_9454,N_8496,N_8030);
nand U9455 (N_9455,N_8341,N_8157);
nor U9456 (N_9456,N_8020,N_8768);
and U9457 (N_9457,N_8070,N_8619);
or U9458 (N_9458,N_8376,N_8968);
nor U9459 (N_9459,N_8109,N_8800);
nand U9460 (N_9460,N_8818,N_8576);
nor U9461 (N_9461,N_8569,N_8737);
nand U9462 (N_9462,N_8699,N_8657);
or U9463 (N_9463,N_8382,N_8008);
nor U9464 (N_9464,N_8399,N_8704);
nor U9465 (N_9465,N_8277,N_8334);
or U9466 (N_9466,N_8746,N_8467);
or U9467 (N_9467,N_8944,N_8529);
and U9468 (N_9468,N_8034,N_8805);
and U9469 (N_9469,N_8117,N_8289);
nand U9470 (N_9470,N_8111,N_8346);
nor U9471 (N_9471,N_8193,N_8993);
nor U9472 (N_9472,N_8179,N_8089);
or U9473 (N_9473,N_8906,N_8025);
or U9474 (N_9474,N_8010,N_8888);
nand U9475 (N_9475,N_8305,N_8308);
nor U9476 (N_9476,N_8284,N_8504);
nand U9477 (N_9477,N_8124,N_8535);
nor U9478 (N_9478,N_8321,N_8174);
nor U9479 (N_9479,N_8397,N_8538);
or U9480 (N_9480,N_8762,N_8255);
or U9481 (N_9481,N_8406,N_8066);
or U9482 (N_9482,N_8208,N_8739);
and U9483 (N_9483,N_8892,N_8374);
or U9484 (N_9484,N_8412,N_8204);
nor U9485 (N_9485,N_8728,N_8966);
nor U9486 (N_9486,N_8909,N_8134);
or U9487 (N_9487,N_8141,N_8691);
nor U9488 (N_9488,N_8692,N_8887);
and U9489 (N_9489,N_8110,N_8261);
nor U9490 (N_9490,N_8129,N_8626);
nand U9491 (N_9491,N_8123,N_8721);
nand U9492 (N_9492,N_8518,N_8710);
nor U9493 (N_9493,N_8873,N_8278);
nor U9494 (N_9494,N_8263,N_8792);
or U9495 (N_9495,N_8580,N_8306);
nand U9496 (N_9496,N_8172,N_8453);
or U9497 (N_9497,N_8155,N_8857);
and U9498 (N_9498,N_8455,N_8198);
nor U9499 (N_9499,N_8783,N_8588);
nand U9500 (N_9500,N_8933,N_8551);
nor U9501 (N_9501,N_8198,N_8319);
and U9502 (N_9502,N_8536,N_8152);
nor U9503 (N_9503,N_8071,N_8600);
or U9504 (N_9504,N_8330,N_8958);
and U9505 (N_9505,N_8578,N_8008);
or U9506 (N_9506,N_8784,N_8407);
and U9507 (N_9507,N_8504,N_8196);
or U9508 (N_9508,N_8267,N_8075);
and U9509 (N_9509,N_8984,N_8289);
nor U9510 (N_9510,N_8328,N_8282);
or U9511 (N_9511,N_8190,N_8212);
and U9512 (N_9512,N_8915,N_8214);
nand U9513 (N_9513,N_8056,N_8344);
nand U9514 (N_9514,N_8186,N_8314);
nor U9515 (N_9515,N_8079,N_8710);
nor U9516 (N_9516,N_8124,N_8880);
or U9517 (N_9517,N_8817,N_8275);
nand U9518 (N_9518,N_8569,N_8662);
nand U9519 (N_9519,N_8564,N_8793);
or U9520 (N_9520,N_8978,N_8965);
nor U9521 (N_9521,N_8154,N_8539);
and U9522 (N_9522,N_8728,N_8574);
nor U9523 (N_9523,N_8208,N_8813);
nor U9524 (N_9524,N_8510,N_8328);
and U9525 (N_9525,N_8719,N_8532);
nand U9526 (N_9526,N_8495,N_8334);
or U9527 (N_9527,N_8747,N_8334);
nor U9528 (N_9528,N_8270,N_8171);
or U9529 (N_9529,N_8452,N_8236);
nor U9530 (N_9530,N_8168,N_8257);
nand U9531 (N_9531,N_8241,N_8868);
nand U9532 (N_9532,N_8487,N_8819);
and U9533 (N_9533,N_8776,N_8028);
and U9534 (N_9534,N_8856,N_8080);
nor U9535 (N_9535,N_8325,N_8349);
or U9536 (N_9536,N_8065,N_8860);
and U9537 (N_9537,N_8946,N_8374);
and U9538 (N_9538,N_8523,N_8423);
or U9539 (N_9539,N_8058,N_8474);
and U9540 (N_9540,N_8072,N_8221);
nor U9541 (N_9541,N_8991,N_8240);
or U9542 (N_9542,N_8457,N_8750);
and U9543 (N_9543,N_8637,N_8783);
or U9544 (N_9544,N_8361,N_8470);
nand U9545 (N_9545,N_8862,N_8238);
xor U9546 (N_9546,N_8384,N_8679);
or U9547 (N_9547,N_8763,N_8383);
and U9548 (N_9548,N_8870,N_8667);
xor U9549 (N_9549,N_8711,N_8988);
nand U9550 (N_9550,N_8722,N_8717);
nand U9551 (N_9551,N_8949,N_8246);
nor U9552 (N_9552,N_8062,N_8883);
or U9553 (N_9553,N_8232,N_8681);
and U9554 (N_9554,N_8031,N_8593);
nand U9555 (N_9555,N_8086,N_8563);
and U9556 (N_9556,N_8304,N_8285);
nand U9557 (N_9557,N_8562,N_8289);
nor U9558 (N_9558,N_8885,N_8951);
nor U9559 (N_9559,N_8488,N_8846);
nor U9560 (N_9560,N_8859,N_8717);
or U9561 (N_9561,N_8878,N_8540);
nor U9562 (N_9562,N_8299,N_8575);
and U9563 (N_9563,N_8047,N_8632);
nand U9564 (N_9564,N_8852,N_8411);
or U9565 (N_9565,N_8091,N_8522);
nor U9566 (N_9566,N_8284,N_8696);
or U9567 (N_9567,N_8253,N_8568);
or U9568 (N_9568,N_8409,N_8283);
and U9569 (N_9569,N_8675,N_8005);
and U9570 (N_9570,N_8867,N_8250);
or U9571 (N_9571,N_8354,N_8100);
nor U9572 (N_9572,N_8619,N_8967);
nor U9573 (N_9573,N_8380,N_8242);
and U9574 (N_9574,N_8099,N_8989);
nand U9575 (N_9575,N_8029,N_8937);
and U9576 (N_9576,N_8719,N_8233);
or U9577 (N_9577,N_8518,N_8897);
or U9578 (N_9578,N_8070,N_8010);
nor U9579 (N_9579,N_8775,N_8702);
nand U9580 (N_9580,N_8542,N_8315);
and U9581 (N_9581,N_8527,N_8539);
and U9582 (N_9582,N_8821,N_8890);
nand U9583 (N_9583,N_8744,N_8309);
nor U9584 (N_9584,N_8181,N_8924);
or U9585 (N_9585,N_8836,N_8971);
and U9586 (N_9586,N_8791,N_8432);
xnor U9587 (N_9587,N_8231,N_8737);
nand U9588 (N_9588,N_8580,N_8596);
or U9589 (N_9589,N_8670,N_8209);
and U9590 (N_9590,N_8678,N_8880);
and U9591 (N_9591,N_8807,N_8608);
nor U9592 (N_9592,N_8969,N_8511);
nand U9593 (N_9593,N_8010,N_8531);
nor U9594 (N_9594,N_8088,N_8362);
nand U9595 (N_9595,N_8639,N_8194);
and U9596 (N_9596,N_8843,N_8832);
and U9597 (N_9597,N_8981,N_8301);
or U9598 (N_9598,N_8678,N_8407);
nand U9599 (N_9599,N_8747,N_8013);
nor U9600 (N_9600,N_8544,N_8726);
xnor U9601 (N_9601,N_8121,N_8375);
nor U9602 (N_9602,N_8016,N_8786);
nor U9603 (N_9603,N_8541,N_8948);
and U9604 (N_9604,N_8851,N_8118);
xnor U9605 (N_9605,N_8845,N_8963);
nor U9606 (N_9606,N_8422,N_8655);
nor U9607 (N_9607,N_8954,N_8503);
or U9608 (N_9608,N_8135,N_8755);
or U9609 (N_9609,N_8924,N_8737);
or U9610 (N_9610,N_8622,N_8464);
nor U9611 (N_9611,N_8421,N_8979);
and U9612 (N_9612,N_8721,N_8941);
nand U9613 (N_9613,N_8749,N_8750);
and U9614 (N_9614,N_8452,N_8648);
and U9615 (N_9615,N_8609,N_8324);
or U9616 (N_9616,N_8691,N_8916);
and U9617 (N_9617,N_8509,N_8525);
nand U9618 (N_9618,N_8311,N_8316);
or U9619 (N_9619,N_8879,N_8169);
nand U9620 (N_9620,N_8850,N_8361);
and U9621 (N_9621,N_8700,N_8989);
and U9622 (N_9622,N_8781,N_8610);
and U9623 (N_9623,N_8106,N_8497);
nor U9624 (N_9624,N_8042,N_8637);
nor U9625 (N_9625,N_8433,N_8641);
nor U9626 (N_9626,N_8039,N_8912);
and U9627 (N_9627,N_8518,N_8736);
nor U9628 (N_9628,N_8274,N_8185);
nand U9629 (N_9629,N_8636,N_8162);
or U9630 (N_9630,N_8787,N_8807);
or U9631 (N_9631,N_8923,N_8479);
nand U9632 (N_9632,N_8334,N_8715);
and U9633 (N_9633,N_8121,N_8775);
or U9634 (N_9634,N_8663,N_8111);
xor U9635 (N_9635,N_8502,N_8968);
or U9636 (N_9636,N_8246,N_8175);
and U9637 (N_9637,N_8285,N_8227);
nor U9638 (N_9638,N_8822,N_8026);
nor U9639 (N_9639,N_8293,N_8889);
nor U9640 (N_9640,N_8722,N_8652);
nand U9641 (N_9641,N_8477,N_8322);
and U9642 (N_9642,N_8287,N_8968);
and U9643 (N_9643,N_8683,N_8173);
and U9644 (N_9644,N_8907,N_8196);
nor U9645 (N_9645,N_8314,N_8954);
nand U9646 (N_9646,N_8944,N_8427);
nor U9647 (N_9647,N_8320,N_8562);
and U9648 (N_9648,N_8256,N_8026);
nand U9649 (N_9649,N_8468,N_8233);
or U9650 (N_9650,N_8299,N_8402);
nand U9651 (N_9651,N_8099,N_8032);
or U9652 (N_9652,N_8071,N_8761);
nor U9653 (N_9653,N_8425,N_8932);
and U9654 (N_9654,N_8644,N_8193);
or U9655 (N_9655,N_8914,N_8533);
nand U9656 (N_9656,N_8152,N_8209);
nor U9657 (N_9657,N_8136,N_8039);
nand U9658 (N_9658,N_8711,N_8320);
and U9659 (N_9659,N_8804,N_8835);
and U9660 (N_9660,N_8988,N_8697);
nor U9661 (N_9661,N_8199,N_8479);
or U9662 (N_9662,N_8042,N_8402);
nor U9663 (N_9663,N_8433,N_8222);
nor U9664 (N_9664,N_8951,N_8146);
or U9665 (N_9665,N_8041,N_8416);
nand U9666 (N_9666,N_8494,N_8576);
nor U9667 (N_9667,N_8413,N_8964);
or U9668 (N_9668,N_8418,N_8180);
nand U9669 (N_9669,N_8888,N_8942);
and U9670 (N_9670,N_8242,N_8109);
and U9671 (N_9671,N_8713,N_8710);
xnor U9672 (N_9672,N_8289,N_8395);
nand U9673 (N_9673,N_8872,N_8652);
nand U9674 (N_9674,N_8595,N_8082);
nand U9675 (N_9675,N_8091,N_8682);
or U9676 (N_9676,N_8482,N_8036);
nand U9677 (N_9677,N_8154,N_8741);
or U9678 (N_9678,N_8357,N_8830);
and U9679 (N_9679,N_8945,N_8001);
nand U9680 (N_9680,N_8186,N_8252);
nor U9681 (N_9681,N_8670,N_8851);
and U9682 (N_9682,N_8659,N_8200);
nor U9683 (N_9683,N_8244,N_8387);
nand U9684 (N_9684,N_8272,N_8980);
nor U9685 (N_9685,N_8830,N_8223);
nand U9686 (N_9686,N_8959,N_8820);
and U9687 (N_9687,N_8765,N_8841);
and U9688 (N_9688,N_8937,N_8227);
nand U9689 (N_9689,N_8361,N_8806);
nor U9690 (N_9690,N_8051,N_8388);
nor U9691 (N_9691,N_8011,N_8647);
and U9692 (N_9692,N_8314,N_8634);
or U9693 (N_9693,N_8609,N_8355);
nand U9694 (N_9694,N_8049,N_8394);
and U9695 (N_9695,N_8198,N_8958);
nand U9696 (N_9696,N_8809,N_8933);
nand U9697 (N_9697,N_8233,N_8627);
nand U9698 (N_9698,N_8736,N_8935);
nor U9699 (N_9699,N_8846,N_8022);
and U9700 (N_9700,N_8122,N_8945);
and U9701 (N_9701,N_8918,N_8077);
and U9702 (N_9702,N_8864,N_8751);
or U9703 (N_9703,N_8087,N_8876);
and U9704 (N_9704,N_8006,N_8361);
xor U9705 (N_9705,N_8925,N_8609);
or U9706 (N_9706,N_8166,N_8704);
nand U9707 (N_9707,N_8425,N_8068);
or U9708 (N_9708,N_8188,N_8661);
or U9709 (N_9709,N_8130,N_8264);
nand U9710 (N_9710,N_8101,N_8477);
nor U9711 (N_9711,N_8245,N_8749);
and U9712 (N_9712,N_8340,N_8660);
nor U9713 (N_9713,N_8444,N_8685);
or U9714 (N_9714,N_8196,N_8800);
or U9715 (N_9715,N_8115,N_8123);
nand U9716 (N_9716,N_8459,N_8788);
or U9717 (N_9717,N_8972,N_8299);
and U9718 (N_9718,N_8812,N_8804);
and U9719 (N_9719,N_8600,N_8040);
nand U9720 (N_9720,N_8864,N_8521);
or U9721 (N_9721,N_8884,N_8742);
and U9722 (N_9722,N_8536,N_8098);
nor U9723 (N_9723,N_8060,N_8480);
or U9724 (N_9724,N_8778,N_8602);
nand U9725 (N_9725,N_8717,N_8204);
nor U9726 (N_9726,N_8250,N_8346);
nand U9727 (N_9727,N_8056,N_8732);
nand U9728 (N_9728,N_8892,N_8752);
nor U9729 (N_9729,N_8916,N_8060);
or U9730 (N_9730,N_8878,N_8621);
or U9731 (N_9731,N_8722,N_8419);
nor U9732 (N_9732,N_8466,N_8873);
nand U9733 (N_9733,N_8416,N_8917);
and U9734 (N_9734,N_8347,N_8115);
or U9735 (N_9735,N_8122,N_8786);
nand U9736 (N_9736,N_8247,N_8187);
nor U9737 (N_9737,N_8560,N_8181);
nand U9738 (N_9738,N_8231,N_8787);
nor U9739 (N_9739,N_8601,N_8188);
nor U9740 (N_9740,N_8488,N_8136);
nand U9741 (N_9741,N_8006,N_8282);
and U9742 (N_9742,N_8574,N_8497);
or U9743 (N_9743,N_8694,N_8136);
nor U9744 (N_9744,N_8719,N_8083);
nor U9745 (N_9745,N_8389,N_8666);
nor U9746 (N_9746,N_8900,N_8836);
nor U9747 (N_9747,N_8699,N_8294);
and U9748 (N_9748,N_8159,N_8665);
nor U9749 (N_9749,N_8523,N_8243);
nor U9750 (N_9750,N_8789,N_8297);
xnor U9751 (N_9751,N_8408,N_8781);
or U9752 (N_9752,N_8983,N_8169);
and U9753 (N_9753,N_8743,N_8826);
nand U9754 (N_9754,N_8276,N_8219);
or U9755 (N_9755,N_8647,N_8922);
or U9756 (N_9756,N_8469,N_8570);
and U9757 (N_9757,N_8319,N_8813);
nor U9758 (N_9758,N_8493,N_8193);
nand U9759 (N_9759,N_8422,N_8613);
nand U9760 (N_9760,N_8095,N_8040);
and U9761 (N_9761,N_8232,N_8198);
xor U9762 (N_9762,N_8578,N_8155);
and U9763 (N_9763,N_8086,N_8320);
or U9764 (N_9764,N_8251,N_8006);
or U9765 (N_9765,N_8018,N_8052);
or U9766 (N_9766,N_8772,N_8747);
or U9767 (N_9767,N_8346,N_8743);
nor U9768 (N_9768,N_8911,N_8587);
or U9769 (N_9769,N_8300,N_8189);
nor U9770 (N_9770,N_8964,N_8518);
nor U9771 (N_9771,N_8215,N_8157);
nor U9772 (N_9772,N_8126,N_8352);
nand U9773 (N_9773,N_8454,N_8797);
and U9774 (N_9774,N_8037,N_8026);
and U9775 (N_9775,N_8270,N_8414);
nand U9776 (N_9776,N_8928,N_8376);
or U9777 (N_9777,N_8279,N_8799);
nor U9778 (N_9778,N_8374,N_8538);
or U9779 (N_9779,N_8678,N_8546);
nand U9780 (N_9780,N_8272,N_8453);
and U9781 (N_9781,N_8561,N_8631);
or U9782 (N_9782,N_8120,N_8707);
nor U9783 (N_9783,N_8522,N_8348);
xor U9784 (N_9784,N_8376,N_8176);
nand U9785 (N_9785,N_8177,N_8192);
or U9786 (N_9786,N_8445,N_8829);
nor U9787 (N_9787,N_8062,N_8738);
or U9788 (N_9788,N_8820,N_8400);
xnor U9789 (N_9789,N_8207,N_8138);
or U9790 (N_9790,N_8816,N_8928);
nor U9791 (N_9791,N_8900,N_8652);
and U9792 (N_9792,N_8117,N_8966);
nand U9793 (N_9793,N_8296,N_8061);
nand U9794 (N_9794,N_8172,N_8919);
or U9795 (N_9795,N_8832,N_8384);
or U9796 (N_9796,N_8666,N_8964);
or U9797 (N_9797,N_8588,N_8006);
or U9798 (N_9798,N_8344,N_8276);
and U9799 (N_9799,N_8359,N_8651);
nor U9800 (N_9800,N_8404,N_8467);
or U9801 (N_9801,N_8054,N_8768);
nand U9802 (N_9802,N_8916,N_8080);
nand U9803 (N_9803,N_8657,N_8039);
nor U9804 (N_9804,N_8729,N_8512);
nor U9805 (N_9805,N_8518,N_8873);
nand U9806 (N_9806,N_8152,N_8861);
nand U9807 (N_9807,N_8526,N_8777);
nand U9808 (N_9808,N_8125,N_8576);
nand U9809 (N_9809,N_8363,N_8305);
and U9810 (N_9810,N_8148,N_8133);
nor U9811 (N_9811,N_8413,N_8547);
xnor U9812 (N_9812,N_8872,N_8269);
xnor U9813 (N_9813,N_8182,N_8084);
nand U9814 (N_9814,N_8516,N_8411);
nor U9815 (N_9815,N_8470,N_8221);
and U9816 (N_9816,N_8684,N_8180);
and U9817 (N_9817,N_8275,N_8584);
nor U9818 (N_9818,N_8609,N_8136);
nand U9819 (N_9819,N_8898,N_8138);
and U9820 (N_9820,N_8632,N_8111);
or U9821 (N_9821,N_8382,N_8598);
nand U9822 (N_9822,N_8789,N_8202);
nor U9823 (N_9823,N_8805,N_8684);
or U9824 (N_9824,N_8569,N_8830);
nand U9825 (N_9825,N_8146,N_8945);
nor U9826 (N_9826,N_8739,N_8243);
or U9827 (N_9827,N_8766,N_8315);
nand U9828 (N_9828,N_8895,N_8225);
xnor U9829 (N_9829,N_8094,N_8193);
nand U9830 (N_9830,N_8361,N_8669);
nand U9831 (N_9831,N_8721,N_8616);
and U9832 (N_9832,N_8755,N_8901);
or U9833 (N_9833,N_8691,N_8289);
nand U9834 (N_9834,N_8060,N_8041);
nand U9835 (N_9835,N_8232,N_8015);
nand U9836 (N_9836,N_8139,N_8227);
nand U9837 (N_9837,N_8202,N_8920);
xnor U9838 (N_9838,N_8127,N_8367);
xnor U9839 (N_9839,N_8526,N_8999);
nor U9840 (N_9840,N_8976,N_8483);
or U9841 (N_9841,N_8072,N_8650);
or U9842 (N_9842,N_8429,N_8653);
nand U9843 (N_9843,N_8864,N_8617);
and U9844 (N_9844,N_8612,N_8172);
nand U9845 (N_9845,N_8863,N_8205);
nand U9846 (N_9846,N_8394,N_8345);
nand U9847 (N_9847,N_8116,N_8888);
and U9848 (N_9848,N_8545,N_8764);
or U9849 (N_9849,N_8282,N_8038);
nand U9850 (N_9850,N_8243,N_8809);
nor U9851 (N_9851,N_8508,N_8686);
and U9852 (N_9852,N_8073,N_8282);
or U9853 (N_9853,N_8793,N_8091);
or U9854 (N_9854,N_8386,N_8226);
nor U9855 (N_9855,N_8771,N_8607);
nor U9856 (N_9856,N_8570,N_8485);
or U9857 (N_9857,N_8850,N_8736);
nand U9858 (N_9858,N_8681,N_8865);
or U9859 (N_9859,N_8507,N_8024);
and U9860 (N_9860,N_8736,N_8220);
nand U9861 (N_9861,N_8416,N_8317);
nand U9862 (N_9862,N_8802,N_8840);
and U9863 (N_9863,N_8989,N_8957);
nor U9864 (N_9864,N_8055,N_8953);
nand U9865 (N_9865,N_8275,N_8727);
and U9866 (N_9866,N_8665,N_8786);
xor U9867 (N_9867,N_8992,N_8076);
nor U9868 (N_9868,N_8346,N_8809);
and U9869 (N_9869,N_8619,N_8245);
and U9870 (N_9870,N_8160,N_8445);
nand U9871 (N_9871,N_8298,N_8530);
and U9872 (N_9872,N_8138,N_8444);
nor U9873 (N_9873,N_8299,N_8630);
or U9874 (N_9874,N_8404,N_8844);
xnor U9875 (N_9875,N_8197,N_8609);
nor U9876 (N_9876,N_8303,N_8472);
nor U9877 (N_9877,N_8586,N_8992);
nor U9878 (N_9878,N_8816,N_8079);
or U9879 (N_9879,N_8160,N_8143);
nand U9880 (N_9880,N_8687,N_8972);
nand U9881 (N_9881,N_8518,N_8248);
and U9882 (N_9882,N_8513,N_8988);
nand U9883 (N_9883,N_8222,N_8259);
or U9884 (N_9884,N_8759,N_8106);
nand U9885 (N_9885,N_8006,N_8530);
xnor U9886 (N_9886,N_8667,N_8702);
or U9887 (N_9887,N_8165,N_8025);
nand U9888 (N_9888,N_8665,N_8542);
and U9889 (N_9889,N_8949,N_8579);
nor U9890 (N_9890,N_8051,N_8412);
nor U9891 (N_9891,N_8810,N_8123);
nor U9892 (N_9892,N_8583,N_8483);
nand U9893 (N_9893,N_8087,N_8402);
and U9894 (N_9894,N_8734,N_8204);
nand U9895 (N_9895,N_8390,N_8043);
nand U9896 (N_9896,N_8522,N_8841);
or U9897 (N_9897,N_8500,N_8825);
nor U9898 (N_9898,N_8152,N_8031);
nor U9899 (N_9899,N_8648,N_8200);
or U9900 (N_9900,N_8623,N_8348);
or U9901 (N_9901,N_8957,N_8194);
or U9902 (N_9902,N_8935,N_8802);
or U9903 (N_9903,N_8500,N_8987);
and U9904 (N_9904,N_8310,N_8720);
nand U9905 (N_9905,N_8158,N_8891);
xnor U9906 (N_9906,N_8552,N_8338);
nor U9907 (N_9907,N_8184,N_8775);
nor U9908 (N_9908,N_8950,N_8135);
or U9909 (N_9909,N_8472,N_8083);
nor U9910 (N_9910,N_8414,N_8894);
nor U9911 (N_9911,N_8301,N_8843);
or U9912 (N_9912,N_8315,N_8661);
nor U9913 (N_9913,N_8834,N_8361);
nand U9914 (N_9914,N_8240,N_8539);
or U9915 (N_9915,N_8352,N_8476);
xor U9916 (N_9916,N_8517,N_8383);
and U9917 (N_9917,N_8846,N_8019);
nor U9918 (N_9918,N_8291,N_8785);
or U9919 (N_9919,N_8553,N_8207);
nand U9920 (N_9920,N_8960,N_8507);
nand U9921 (N_9921,N_8585,N_8329);
and U9922 (N_9922,N_8051,N_8208);
or U9923 (N_9923,N_8647,N_8498);
nor U9924 (N_9924,N_8508,N_8737);
nor U9925 (N_9925,N_8456,N_8331);
nor U9926 (N_9926,N_8167,N_8371);
and U9927 (N_9927,N_8027,N_8762);
nor U9928 (N_9928,N_8674,N_8695);
nand U9929 (N_9929,N_8695,N_8960);
nor U9930 (N_9930,N_8110,N_8806);
nand U9931 (N_9931,N_8180,N_8257);
or U9932 (N_9932,N_8878,N_8765);
nor U9933 (N_9933,N_8552,N_8627);
and U9934 (N_9934,N_8329,N_8301);
nor U9935 (N_9935,N_8229,N_8519);
nor U9936 (N_9936,N_8896,N_8826);
nand U9937 (N_9937,N_8117,N_8735);
and U9938 (N_9938,N_8994,N_8646);
and U9939 (N_9939,N_8660,N_8079);
nand U9940 (N_9940,N_8974,N_8456);
or U9941 (N_9941,N_8034,N_8161);
and U9942 (N_9942,N_8309,N_8985);
nand U9943 (N_9943,N_8684,N_8984);
nand U9944 (N_9944,N_8097,N_8704);
nand U9945 (N_9945,N_8364,N_8655);
and U9946 (N_9946,N_8379,N_8197);
nor U9947 (N_9947,N_8811,N_8073);
or U9948 (N_9948,N_8834,N_8647);
nand U9949 (N_9949,N_8373,N_8993);
nand U9950 (N_9950,N_8839,N_8391);
nand U9951 (N_9951,N_8183,N_8413);
nor U9952 (N_9952,N_8505,N_8574);
and U9953 (N_9953,N_8392,N_8207);
nor U9954 (N_9954,N_8607,N_8589);
nand U9955 (N_9955,N_8057,N_8967);
or U9956 (N_9956,N_8911,N_8094);
xnor U9957 (N_9957,N_8140,N_8898);
or U9958 (N_9958,N_8217,N_8166);
nand U9959 (N_9959,N_8317,N_8648);
nor U9960 (N_9960,N_8463,N_8698);
or U9961 (N_9961,N_8128,N_8536);
nor U9962 (N_9962,N_8477,N_8324);
and U9963 (N_9963,N_8284,N_8173);
and U9964 (N_9964,N_8496,N_8111);
and U9965 (N_9965,N_8729,N_8395);
or U9966 (N_9966,N_8982,N_8150);
nand U9967 (N_9967,N_8544,N_8248);
nand U9968 (N_9968,N_8244,N_8380);
or U9969 (N_9969,N_8782,N_8502);
or U9970 (N_9970,N_8059,N_8408);
or U9971 (N_9971,N_8854,N_8627);
and U9972 (N_9972,N_8769,N_8346);
nand U9973 (N_9973,N_8252,N_8027);
or U9974 (N_9974,N_8471,N_8355);
nor U9975 (N_9975,N_8851,N_8214);
nor U9976 (N_9976,N_8242,N_8579);
nor U9977 (N_9977,N_8736,N_8758);
and U9978 (N_9978,N_8334,N_8772);
or U9979 (N_9979,N_8729,N_8609);
or U9980 (N_9980,N_8101,N_8901);
or U9981 (N_9981,N_8503,N_8008);
nand U9982 (N_9982,N_8640,N_8295);
and U9983 (N_9983,N_8855,N_8686);
or U9984 (N_9984,N_8326,N_8925);
nand U9985 (N_9985,N_8267,N_8477);
nand U9986 (N_9986,N_8867,N_8778);
and U9987 (N_9987,N_8894,N_8196);
nor U9988 (N_9988,N_8484,N_8409);
or U9989 (N_9989,N_8448,N_8165);
nand U9990 (N_9990,N_8312,N_8434);
nor U9991 (N_9991,N_8184,N_8790);
nor U9992 (N_9992,N_8864,N_8092);
or U9993 (N_9993,N_8124,N_8741);
nor U9994 (N_9994,N_8755,N_8987);
and U9995 (N_9995,N_8389,N_8342);
and U9996 (N_9996,N_8126,N_8564);
or U9997 (N_9997,N_8594,N_8672);
nand U9998 (N_9998,N_8508,N_8371);
and U9999 (N_9999,N_8684,N_8567);
or UO_0 (O_0,N_9117,N_9786);
xnor UO_1 (O_1,N_9413,N_9725);
and UO_2 (O_2,N_9817,N_9184);
and UO_3 (O_3,N_9854,N_9255);
xor UO_4 (O_4,N_9186,N_9459);
or UO_5 (O_5,N_9703,N_9095);
and UO_6 (O_6,N_9365,N_9839);
xnor UO_7 (O_7,N_9000,N_9237);
or UO_8 (O_8,N_9168,N_9400);
nand UO_9 (O_9,N_9264,N_9081);
or UO_10 (O_10,N_9316,N_9105);
nor UO_11 (O_11,N_9661,N_9579);
nand UO_12 (O_12,N_9017,N_9630);
and UO_13 (O_13,N_9140,N_9007);
nor UO_14 (O_14,N_9450,N_9405);
and UO_15 (O_15,N_9730,N_9647);
or UO_16 (O_16,N_9559,N_9215);
and UO_17 (O_17,N_9021,N_9241);
xor UO_18 (O_18,N_9808,N_9918);
nand UO_19 (O_19,N_9260,N_9844);
nor UO_20 (O_20,N_9120,N_9843);
nand UO_21 (O_21,N_9401,N_9609);
nor UO_22 (O_22,N_9093,N_9691);
or UO_23 (O_23,N_9479,N_9284);
and UO_24 (O_24,N_9207,N_9537);
nor UO_25 (O_25,N_9980,N_9009);
nand UO_26 (O_26,N_9269,N_9865);
nand UO_27 (O_27,N_9272,N_9209);
or UO_28 (O_28,N_9288,N_9673);
nor UO_29 (O_29,N_9353,N_9952);
or UO_30 (O_30,N_9753,N_9884);
xnor UO_31 (O_31,N_9030,N_9664);
nor UO_32 (O_32,N_9623,N_9951);
or UO_33 (O_33,N_9467,N_9885);
nor UO_34 (O_34,N_9682,N_9738);
nand UO_35 (O_35,N_9086,N_9495);
nand UO_36 (O_36,N_9228,N_9666);
or UO_37 (O_37,N_9261,N_9350);
and UO_38 (O_38,N_9718,N_9438);
nor UO_39 (O_39,N_9769,N_9655);
nor UO_40 (O_40,N_9115,N_9205);
nand UO_41 (O_41,N_9285,N_9897);
nor UO_42 (O_42,N_9462,N_9799);
and UO_43 (O_43,N_9028,N_9315);
nand UO_44 (O_44,N_9301,N_9942);
xor UO_45 (O_45,N_9988,N_9204);
nor UO_46 (O_46,N_9530,N_9571);
nand UO_47 (O_47,N_9158,N_9022);
or UO_48 (O_48,N_9581,N_9181);
nor UO_49 (O_49,N_9742,N_9464);
or UO_50 (O_50,N_9779,N_9757);
or UO_51 (O_51,N_9573,N_9814);
nand UO_52 (O_52,N_9858,N_9832);
or UO_53 (O_53,N_9616,N_9524);
nor UO_54 (O_54,N_9922,N_9517);
or UO_55 (O_55,N_9054,N_9624);
nand UO_56 (O_56,N_9826,N_9877);
or UO_57 (O_57,N_9445,N_9034);
or UO_58 (O_58,N_9793,N_9398);
or UO_59 (O_59,N_9454,N_9046);
nor UO_60 (O_60,N_9455,N_9834);
or UO_61 (O_61,N_9411,N_9185);
and UO_62 (O_62,N_9110,N_9441);
or UO_63 (O_63,N_9855,N_9368);
xor UO_64 (O_64,N_9613,N_9809);
nor UO_65 (O_65,N_9866,N_9302);
or UO_66 (O_66,N_9972,N_9849);
nor UO_67 (O_67,N_9035,N_9641);
nor UO_68 (O_68,N_9695,N_9882);
and UO_69 (O_69,N_9615,N_9389);
and UO_70 (O_70,N_9138,N_9783);
nand UO_71 (O_71,N_9578,N_9699);
xor UO_72 (O_72,N_9088,N_9919);
nand UO_73 (O_73,N_9935,N_9429);
nand UO_74 (O_74,N_9121,N_9056);
nand UO_75 (O_75,N_9582,N_9370);
nor UO_76 (O_76,N_9653,N_9824);
nor UO_77 (O_77,N_9483,N_9561);
and UO_78 (O_78,N_9506,N_9903);
and UO_79 (O_79,N_9577,N_9887);
nor UO_80 (O_80,N_9881,N_9500);
and UO_81 (O_81,N_9690,N_9688);
xor UO_82 (O_82,N_9823,N_9060);
nand UO_83 (O_83,N_9475,N_9554);
nor UO_84 (O_84,N_9279,N_9852);
and UO_85 (O_85,N_9700,N_9078);
nor UO_86 (O_86,N_9902,N_9446);
nand UO_87 (O_87,N_9491,N_9827);
and UO_88 (O_88,N_9011,N_9702);
or UO_89 (O_89,N_9126,N_9617);
and UO_90 (O_90,N_9199,N_9280);
and UO_91 (O_91,N_9558,N_9289);
nor UO_92 (O_92,N_9962,N_9262);
or UO_93 (O_93,N_9175,N_9190);
or UO_94 (O_94,N_9473,N_9864);
and UO_95 (O_95,N_9715,N_9515);
and UO_96 (O_96,N_9274,N_9178);
or UO_97 (O_97,N_9087,N_9201);
nand UO_98 (O_98,N_9342,N_9380);
nand UO_99 (O_99,N_9632,N_9258);
nand UO_100 (O_100,N_9239,N_9541);
or UO_101 (O_101,N_9679,N_9328);
or UO_102 (O_102,N_9929,N_9476);
nor UO_103 (O_103,N_9780,N_9969);
nand UO_104 (O_104,N_9434,N_9543);
or UO_105 (O_105,N_9132,N_9904);
and UO_106 (O_106,N_9176,N_9869);
and UO_107 (O_107,N_9638,N_9644);
nor UO_108 (O_108,N_9755,N_9364);
nor UO_109 (O_109,N_9901,N_9414);
and UO_110 (O_110,N_9440,N_9777);
nor UO_111 (O_111,N_9708,N_9512);
nand UO_112 (O_112,N_9296,N_9133);
or UO_113 (O_113,N_9820,N_9229);
and UO_114 (O_114,N_9155,N_9409);
nand UO_115 (O_115,N_9842,N_9016);
and UO_116 (O_116,N_9967,N_9125);
and UO_117 (O_117,N_9090,N_9719);
nor UO_118 (O_118,N_9310,N_9698);
and UO_119 (O_119,N_9905,N_9195);
and UO_120 (O_120,N_9442,N_9164);
nand UO_121 (O_121,N_9539,N_9568);
or UO_122 (O_122,N_9714,N_9565);
xor UO_123 (O_123,N_9489,N_9658);
nand UO_124 (O_124,N_9815,N_9361);
nand UO_125 (O_125,N_9367,N_9527);
nand UO_126 (O_126,N_9580,N_9430);
or UO_127 (O_127,N_9047,N_9914);
or UO_128 (O_128,N_9183,N_9841);
and UO_129 (O_129,N_9569,N_9928);
nand UO_130 (O_130,N_9044,N_9576);
and UO_131 (O_131,N_9068,N_9064);
or UO_132 (O_132,N_9925,N_9751);
nand UO_133 (O_133,N_9618,N_9676);
nand UO_134 (O_134,N_9012,N_9896);
nor UO_135 (O_135,N_9135,N_9743);
and UO_136 (O_136,N_9509,N_9329);
nor UO_137 (O_137,N_9979,N_9340);
and UO_138 (O_138,N_9998,N_9266);
or UO_139 (O_139,N_9785,N_9354);
nor UO_140 (O_140,N_9193,N_9231);
and UO_141 (O_141,N_9927,N_9831);
nand UO_142 (O_142,N_9739,N_9163);
or UO_143 (O_143,N_9895,N_9701);
nor UO_144 (O_144,N_9888,N_9298);
nor UO_145 (O_145,N_9546,N_9249);
nand UO_146 (O_146,N_9294,N_9493);
or UO_147 (O_147,N_9382,N_9829);
nor UO_148 (O_148,N_9776,N_9657);
nand UO_149 (O_149,N_9394,N_9331);
nand UO_150 (O_150,N_9234,N_9482);
nand UO_151 (O_151,N_9308,N_9520);
or UO_152 (O_152,N_9307,N_9795);
nor UO_153 (O_153,N_9734,N_9911);
or UO_154 (O_154,N_9511,N_9069);
nand UO_155 (O_155,N_9122,N_9744);
nand UO_156 (O_156,N_9908,N_9924);
or UO_157 (O_157,N_9497,N_9319);
nor UO_158 (O_158,N_9694,N_9416);
and UO_159 (O_159,N_9423,N_9639);
nand UO_160 (O_160,N_9667,N_9073);
nand UO_161 (O_161,N_9989,N_9723);
nand UO_162 (O_162,N_9847,N_9388);
nand UO_163 (O_163,N_9084,N_9800);
and UO_164 (O_164,N_9244,N_9299);
nor UO_165 (O_165,N_9259,N_9202);
or UO_166 (O_166,N_9290,N_9246);
and UO_167 (O_167,N_9782,N_9505);
or UO_168 (O_168,N_9396,N_9216);
and UO_169 (O_169,N_9642,N_9548);
nand UO_170 (O_170,N_9381,N_9993);
or UO_171 (O_171,N_9355,N_9304);
and UO_172 (O_172,N_9226,N_9188);
and UO_173 (O_173,N_9981,N_9620);
and UO_174 (O_174,N_9456,N_9650);
or UO_175 (O_175,N_9070,N_9949);
or UO_176 (O_176,N_9363,N_9148);
nand UO_177 (O_177,N_9521,N_9312);
nand UO_178 (O_178,N_9798,N_9336);
or UO_179 (O_179,N_9161,N_9663);
nor UO_180 (O_180,N_9614,N_9648);
nor UO_181 (O_181,N_9092,N_9151);
nor UO_182 (O_182,N_9759,N_9094);
nand UO_183 (O_183,N_9139,N_9391);
nor UO_184 (O_184,N_9420,N_9461);
or UO_185 (O_185,N_9604,N_9592);
nor UO_186 (O_186,N_9850,N_9544);
and UO_187 (O_187,N_9242,N_9930);
nor UO_188 (O_188,N_9061,N_9263);
and UO_189 (O_189,N_9732,N_9619);
nor UO_190 (O_190,N_9225,N_9439);
or UO_191 (O_191,N_9662,N_9886);
or UO_192 (O_192,N_9480,N_9529);
nor UO_193 (O_193,N_9102,N_9560);
and UO_194 (O_194,N_9504,N_9983);
nor UO_195 (O_195,N_9322,N_9737);
nand UO_196 (O_196,N_9421,N_9099);
and UO_197 (O_197,N_9254,N_9080);
nand UO_198 (O_198,N_9253,N_9538);
xor UO_199 (O_199,N_9145,N_9545);
nor UO_200 (O_200,N_9174,N_9124);
or UO_201 (O_201,N_9404,N_9451);
nand UO_202 (O_202,N_9670,N_9567);
nor UO_203 (O_203,N_9196,N_9003);
and UO_204 (O_204,N_9874,N_9142);
and UO_205 (O_205,N_9360,N_9096);
nor UO_206 (O_206,N_9055,N_9303);
nand UO_207 (O_207,N_9646,N_9032);
xnor UO_208 (O_208,N_9941,N_9863);
and UO_209 (O_209,N_9977,N_9306);
nor UO_210 (O_210,N_9819,N_9171);
xnor UO_211 (O_211,N_9051,N_9830);
nor UO_212 (O_212,N_9945,N_9157);
nand UO_213 (O_213,N_9966,N_9503);
and UO_214 (O_214,N_9318,N_9077);
nand UO_215 (O_215,N_9432,N_9348);
and UO_216 (O_216,N_9950,N_9214);
nand UO_217 (O_217,N_9933,N_9343);
nor UO_218 (O_218,N_9267,N_9805);
nor UO_219 (O_219,N_9760,N_9603);
or UO_220 (O_220,N_9013,N_9526);
or UO_221 (O_221,N_9344,N_9337);
or UO_222 (O_222,N_9106,N_9997);
nor UO_223 (O_223,N_9518,N_9057);
and UO_224 (O_224,N_9627,N_9477);
or UO_225 (O_225,N_9075,N_9453);
and UO_226 (O_226,N_9019,N_9740);
xnor UO_227 (O_227,N_9856,N_9079);
and UO_228 (O_228,N_9407,N_9369);
and UO_229 (O_229,N_9297,N_9510);
or UO_230 (O_230,N_9704,N_9167);
nand UO_231 (O_231,N_9633,N_9023);
and UO_232 (O_232,N_9923,N_9802);
nand UO_233 (O_233,N_9478,N_9066);
and UO_234 (O_234,N_9346,N_9341);
nand UO_235 (O_235,N_9458,N_9426);
and UO_236 (O_236,N_9268,N_9716);
nor UO_237 (O_237,N_9300,N_9484);
or UO_238 (O_238,N_9083,N_9376);
and UO_239 (O_239,N_9940,N_9562);
nand UO_240 (O_240,N_9098,N_9909);
or UO_241 (O_241,N_9778,N_9602);
nor UO_242 (O_242,N_9996,N_9020);
and UO_243 (O_243,N_9496,N_9774);
and UO_244 (O_244,N_9883,N_9722);
and UO_245 (O_245,N_9425,N_9251);
and UO_246 (O_246,N_9871,N_9042);
nor UO_247 (O_247,N_9248,N_9665);
or UO_248 (O_248,N_9194,N_9292);
and UO_249 (O_249,N_9472,N_9835);
nand UO_250 (O_250,N_9837,N_9878);
nand UO_251 (O_251,N_9756,N_9457);
or UO_252 (O_252,N_9970,N_9867);
xor UO_253 (O_253,N_9833,N_9052);
nand UO_254 (O_254,N_9920,N_9797);
or UO_255 (O_255,N_9975,N_9851);
or UO_256 (O_256,N_9766,N_9921);
and UO_257 (O_257,N_9089,N_9408);
or UO_258 (O_258,N_9123,N_9072);
or UO_259 (O_259,N_9103,N_9213);
nor UO_260 (O_260,N_9956,N_9492);
and UO_261 (O_261,N_9198,N_9550);
and UO_262 (O_262,N_9696,N_9433);
nand UO_263 (O_263,N_9727,N_9724);
nand UO_264 (O_264,N_9533,N_9470);
and UO_265 (O_265,N_9377,N_9427);
nand UO_266 (O_266,N_9861,N_9490);
and UO_267 (O_267,N_9452,N_9948);
nor UO_268 (O_268,N_9485,N_9705);
nor UO_269 (O_269,N_9392,N_9351);
nor UO_270 (O_270,N_9137,N_9801);
nor UO_271 (O_271,N_9265,N_9900);
nor UO_272 (O_272,N_9384,N_9711);
and UO_273 (O_273,N_9685,N_9965);
and UO_274 (O_274,N_9374,N_9008);
nor UO_275 (O_275,N_9605,N_9435);
or UO_276 (O_276,N_9177,N_9208);
or UO_277 (O_277,N_9397,N_9610);
nor UO_278 (O_278,N_9502,N_9059);
or UO_279 (O_279,N_9811,N_9053);
nand UO_280 (O_280,N_9223,N_9984);
nor UO_281 (O_281,N_9295,N_9323);
or UO_282 (O_282,N_9612,N_9807);
nor UO_283 (O_283,N_9041,N_9065);
nand UO_284 (O_284,N_9160,N_9649);
nor UO_285 (O_285,N_9812,N_9747);
and UO_286 (O_286,N_9912,N_9062);
nor UO_287 (O_287,N_9460,N_9848);
nor UO_288 (O_288,N_9222,N_9781);
and UO_289 (O_289,N_9386,N_9516);
and UO_290 (O_290,N_9036,N_9031);
nor UO_291 (O_291,N_9587,N_9631);
nor UO_292 (O_292,N_9906,N_9217);
nor UO_293 (O_293,N_9806,N_9211);
nor UO_294 (O_294,N_9588,N_9447);
nand UO_295 (O_295,N_9957,N_9845);
nand UO_296 (O_296,N_9735,N_9002);
nor UO_297 (O_297,N_9995,N_9557);
nor UO_298 (O_298,N_9210,N_9890);
nand UO_299 (O_299,N_9936,N_9219);
or UO_300 (O_300,N_9551,N_9687);
and UO_301 (O_301,N_9278,N_9330);
or UO_302 (O_302,N_9628,N_9282);
or UO_303 (O_303,N_9963,N_9974);
nand UO_304 (O_304,N_9487,N_9444);
nand UO_305 (O_305,N_9127,N_9748);
nand UO_306 (O_306,N_9383,N_9689);
nor UO_307 (O_307,N_9270,N_9333);
nand UO_308 (O_308,N_9788,N_9027);
xor UO_309 (O_309,N_9403,N_9893);
and UO_310 (O_310,N_9118,N_9422);
and UO_311 (O_311,N_9314,N_9170);
and UO_312 (O_312,N_9335,N_9230);
or UO_313 (O_313,N_9736,N_9136);
nand UO_314 (O_314,N_9507,N_9758);
or UO_315 (O_315,N_9166,N_9471);
nor UO_316 (O_316,N_9597,N_9169);
and UO_317 (O_317,N_9555,N_9156);
nor UO_318 (O_318,N_9325,N_9607);
nor UO_319 (O_319,N_9660,N_9321);
or UO_320 (O_320,N_9352,N_9987);
or UO_321 (O_321,N_9221,N_9712);
nand UO_322 (O_322,N_9324,N_9729);
or UO_323 (O_323,N_9393,N_9358);
or UO_324 (O_324,N_9356,N_9953);
nor UO_325 (O_325,N_9172,N_9668);
nand UO_326 (O_326,N_9192,N_9317);
nor UO_327 (O_327,N_9693,N_9860);
and UO_328 (O_328,N_9119,N_9540);
and UO_329 (O_329,N_9591,N_9173);
and UO_330 (O_330,N_9764,N_9236);
and UO_331 (O_331,N_9143,N_9144);
nand UO_332 (O_332,N_9710,N_9273);
nand UO_333 (O_333,N_9100,N_9672);
nor UO_334 (O_334,N_9074,N_9049);
nor UO_335 (O_335,N_9773,N_9978);
nand UO_336 (O_336,N_9153,N_9752);
nor UO_337 (O_337,N_9415,N_9982);
nor UO_338 (O_338,N_9349,N_9224);
nor UO_339 (O_339,N_9992,N_9566);
or UO_340 (O_340,N_9043,N_9286);
and UO_341 (O_341,N_9271,N_9481);
and UO_342 (O_342,N_9050,N_9625);
nand UO_343 (O_343,N_9754,N_9402);
nor UO_344 (O_344,N_9959,N_9366);
or UO_345 (O_345,N_9645,N_9534);
or UO_346 (O_346,N_9549,N_9746);
nand UO_347 (O_347,N_9899,N_9575);
nor UO_348 (O_348,N_9240,N_9134);
nor UO_349 (O_349,N_9147,N_9519);
nor UO_350 (O_350,N_9709,N_9939);
xnor UO_351 (O_351,N_9165,N_9390);
or UO_352 (O_352,N_9678,N_9488);
nand UO_353 (O_353,N_9180,N_9513);
and UO_354 (O_354,N_9250,N_9654);
and UO_355 (O_355,N_9233,N_9626);
or UO_356 (O_356,N_9916,N_9220);
and UO_357 (O_357,N_9958,N_9825);
or UO_358 (O_358,N_9775,N_9332);
or UO_359 (O_359,N_9634,N_9436);
nand UO_360 (O_360,N_9671,N_9113);
nand UO_361 (O_361,N_9001,N_9821);
nand UO_362 (O_362,N_9463,N_9733);
xnor UO_363 (O_363,N_9787,N_9621);
nor UO_364 (O_364,N_9311,N_9071);
and UO_365 (O_365,N_9907,N_9018);
or UO_366 (O_366,N_9154,N_9412);
or UO_367 (O_367,N_9067,N_9629);
nand UO_368 (O_368,N_9063,N_9584);
and UO_369 (O_369,N_9846,N_9686);
nand UO_370 (O_370,N_9589,N_9287);
nor UO_371 (O_371,N_9608,N_9971);
nand UO_372 (O_372,N_9385,N_9994);
nor UO_373 (O_373,N_9596,N_9857);
and UO_374 (O_374,N_9431,N_9033);
nand UO_375 (O_375,N_9585,N_9347);
and UO_376 (O_376,N_9960,N_9943);
xor UO_377 (O_377,N_9891,N_9437);
nor UO_378 (O_378,N_9728,N_9564);
and UO_379 (O_379,N_9656,N_9150);
or UO_380 (O_380,N_9037,N_9599);
nor UO_381 (O_381,N_9683,N_9359);
or UO_382 (O_382,N_9570,N_9468);
nor UO_383 (O_383,N_9859,N_9130);
or UO_384 (O_384,N_9010,N_9418);
and UO_385 (O_385,N_9556,N_9761);
or UO_386 (O_386,N_9961,N_9309);
nor UO_387 (O_387,N_9111,N_9889);
nand UO_388 (O_388,N_9991,N_9892);
and UO_389 (O_389,N_9720,N_9600);
nand UO_390 (O_390,N_9362,N_9378);
or UO_391 (O_391,N_9771,N_9006);
nor UO_392 (O_392,N_9552,N_9999);
nor UO_393 (O_393,N_9191,N_9112);
and UO_394 (O_394,N_9636,N_9828);
and UO_395 (O_395,N_9305,N_9104);
or UO_396 (O_396,N_9637,N_9796);
xor UO_397 (O_397,N_9024,N_9880);
nand UO_398 (O_398,N_9652,N_9097);
or UO_399 (O_399,N_9474,N_9697);
or UO_400 (O_400,N_9466,N_9531);
and UO_401 (O_401,N_9680,N_9320);
nor UO_402 (O_402,N_9706,N_9276);
nand UO_403 (O_403,N_9762,N_9651);
nand UO_404 (O_404,N_9536,N_9146);
and UO_405 (O_405,N_9792,N_9238);
and UO_406 (O_406,N_9327,N_9873);
and UO_407 (O_407,N_9179,N_9257);
nand UO_408 (O_408,N_9108,N_9937);
nor UO_409 (O_409,N_9938,N_9227);
or UO_410 (O_410,N_9091,N_9313);
nor UO_411 (O_411,N_9014,N_9640);
nand UO_412 (O_412,N_9944,N_9622);
nand UO_413 (O_413,N_9976,N_9107);
nor UO_414 (O_414,N_9593,N_9528);
nand UO_415 (O_415,N_9731,N_9932);
and UO_416 (O_416,N_9116,N_9525);
nand UO_417 (O_417,N_9508,N_9553);
nor UO_418 (O_418,N_9954,N_9045);
or UO_419 (O_419,N_9810,N_9868);
nand UO_420 (O_420,N_9721,N_9252);
nand UO_421 (O_421,N_9522,N_9514);
xnor UO_422 (O_422,N_9419,N_9399);
or UO_423 (O_423,N_9040,N_9443);
nor UO_424 (O_424,N_9523,N_9082);
or UO_425 (O_425,N_9898,N_9813);
and UO_426 (O_426,N_9058,N_9535);
and UO_427 (O_427,N_9726,N_9542);
and UO_428 (O_428,N_9375,N_9334);
or UO_429 (O_429,N_9256,N_9931);
or UO_430 (O_430,N_9373,N_9595);
nand UO_431 (O_431,N_9345,N_9659);
xnor UO_432 (O_432,N_9428,N_9692);
or UO_433 (O_433,N_9338,N_9547);
or UO_434 (O_434,N_9293,N_9494);
and UO_435 (O_435,N_9790,N_9501);
nand UO_436 (O_436,N_9749,N_9159);
nor UO_437 (O_437,N_9406,N_9674);
or UO_438 (O_438,N_9448,N_9277);
nor UO_439 (O_439,N_9677,N_9946);
nor UO_440 (O_440,N_9598,N_9934);
and UO_441 (O_441,N_9128,N_9926);
or UO_442 (O_442,N_9870,N_9187);
and UO_443 (O_443,N_9767,N_9149);
or UO_444 (O_444,N_9131,N_9590);
nor UO_445 (O_445,N_9741,N_9853);
or UO_446 (O_446,N_9372,N_9770);
nand UO_447 (O_447,N_9275,N_9029);
or UO_448 (O_448,N_9339,N_9410);
nor UO_449 (O_449,N_9004,N_9486);
nand UO_450 (O_450,N_9985,N_9283);
or UO_451 (O_451,N_9469,N_9745);
or UO_452 (O_452,N_9152,N_9371);
and UO_453 (O_453,N_9794,N_9765);
nor UO_454 (O_454,N_9707,N_9182);
or UO_455 (O_455,N_9838,N_9910);
or UO_456 (O_456,N_9594,N_9281);
or UO_457 (O_457,N_9606,N_9964);
nand UO_458 (O_458,N_9218,N_9326);
nand UO_459 (O_459,N_9684,N_9818);
and UO_460 (O_460,N_9235,N_9669);
nor UO_461 (O_461,N_9681,N_9915);
or UO_462 (O_462,N_9200,N_9498);
and UO_463 (O_463,N_9822,N_9245);
and UO_464 (O_464,N_9109,N_9417);
or UO_465 (O_465,N_9039,N_9076);
or UO_466 (O_466,N_9387,N_9424);
or UO_467 (O_467,N_9872,N_9203);
nand UO_468 (O_468,N_9015,N_9968);
nand UO_469 (O_469,N_9876,N_9291);
nand UO_470 (O_470,N_9197,N_9038);
and UO_471 (O_471,N_9601,N_9465);
and UO_472 (O_472,N_9955,N_9840);
nor UO_473 (O_473,N_9247,N_9913);
or UO_474 (O_474,N_9816,N_9532);
and UO_475 (O_475,N_9973,N_9085);
or UO_476 (O_476,N_9499,N_9048);
nand UO_477 (O_477,N_9206,N_9611);
nor UO_478 (O_478,N_9232,N_9141);
xor UO_479 (O_479,N_9803,N_9572);
and UO_480 (O_480,N_9635,N_9025);
and UO_481 (O_481,N_9586,N_9917);
or UO_482 (O_482,N_9212,N_9643);
or UO_483 (O_483,N_9379,N_9713);
nand UO_484 (O_484,N_9947,N_9101);
nand UO_485 (O_485,N_9763,N_9875);
and UO_486 (O_486,N_9879,N_9114);
nor UO_487 (O_487,N_9768,N_9784);
nand UO_488 (O_488,N_9005,N_9395);
or UO_489 (O_489,N_9189,N_9836);
nand UO_490 (O_490,N_9862,N_9772);
or UO_491 (O_491,N_9026,N_9804);
or UO_492 (O_492,N_9791,N_9357);
nor UO_493 (O_493,N_9675,N_9243);
nand UO_494 (O_494,N_9986,N_9574);
nor UO_495 (O_495,N_9717,N_9583);
or UO_496 (O_496,N_9563,N_9750);
nand UO_497 (O_497,N_9990,N_9894);
or UO_498 (O_498,N_9449,N_9129);
and UO_499 (O_499,N_9789,N_9162);
nor UO_500 (O_500,N_9619,N_9502);
nor UO_501 (O_501,N_9406,N_9832);
nand UO_502 (O_502,N_9833,N_9116);
and UO_503 (O_503,N_9797,N_9841);
nand UO_504 (O_504,N_9862,N_9457);
nand UO_505 (O_505,N_9563,N_9530);
or UO_506 (O_506,N_9871,N_9315);
nand UO_507 (O_507,N_9715,N_9011);
nor UO_508 (O_508,N_9604,N_9164);
and UO_509 (O_509,N_9459,N_9198);
nand UO_510 (O_510,N_9525,N_9685);
or UO_511 (O_511,N_9900,N_9683);
and UO_512 (O_512,N_9645,N_9169);
nand UO_513 (O_513,N_9792,N_9733);
nand UO_514 (O_514,N_9780,N_9912);
and UO_515 (O_515,N_9142,N_9584);
nand UO_516 (O_516,N_9456,N_9541);
and UO_517 (O_517,N_9770,N_9239);
or UO_518 (O_518,N_9282,N_9439);
nor UO_519 (O_519,N_9117,N_9710);
nor UO_520 (O_520,N_9821,N_9221);
nand UO_521 (O_521,N_9168,N_9423);
and UO_522 (O_522,N_9543,N_9073);
xor UO_523 (O_523,N_9016,N_9676);
nor UO_524 (O_524,N_9696,N_9230);
nor UO_525 (O_525,N_9296,N_9713);
and UO_526 (O_526,N_9152,N_9051);
or UO_527 (O_527,N_9737,N_9541);
or UO_528 (O_528,N_9231,N_9510);
or UO_529 (O_529,N_9143,N_9829);
nor UO_530 (O_530,N_9093,N_9086);
or UO_531 (O_531,N_9437,N_9750);
nand UO_532 (O_532,N_9382,N_9918);
and UO_533 (O_533,N_9841,N_9617);
nand UO_534 (O_534,N_9237,N_9439);
or UO_535 (O_535,N_9809,N_9042);
nand UO_536 (O_536,N_9347,N_9669);
nor UO_537 (O_537,N_9655,N_9970);
and UO_538 (O_538,N_9856,N_9523);
and UO_539 (O_539,N_9645,N_9059);
nor UO_540 (O_540,N_9692,N_9120);
or UO_541 (O_541,N_9607,N_9119);
or UO_542 (O_542,N_9472,N_9681);
and UO_543 (O_543,N_9783,N_9582);
or UO_544 (O_544,N_9114,N_9630);
or UO_545 (O_545,N_9566,N_9312);
and UO_546 (O_546,N_9415,N_9210);
or UO_547 (O_547,N_9691,N_9573);
or UO_548 (O_548,N_9485,N_9493);
and UO_549 (O_549,N_9011,N_9339);
nand UO_550 (O_550,N_9345,N_9596);
nor UO_551 (O_551,N_9733,N_9473);
xnor UO_552 (O_552,N_9289,N_9343);
and UO_553 (O_553,N_9537,N_9067);
and UO_554 (O_554,N_9307,N_9463);
or UO_555 (O_555,N_9148,N_9662);
and UO_556 (O_556,N_9152,N_9916);
and UO_557 (O_557,N_9547,N_9118);
nor UO_558 (O_558,N_9366,N_9295);
or UO_559 (O_559,N_9821,N_9815);
nor UO_560 (O_560,N_9615,N_9311);
nor UO_561 (O_561,N_9817,N_9177);
or UO_562 (O_562,N_9847,N_9269);
nor UO_563 (O_563,N_9269,N_9491);
nand UO_564 (O_564,N_9611,N_9096);
xnor UO_565 (O_565,N_9728,N_9332);
nor UO_566 (O_566,N_9408,N_9067);
and UO_567 (O_567,N_9496,N_9005);
and UO_568 (O_568,N_9131,N_9947);
nand UO_569 (O_569,N_9865,N_9072);
nor UO_570 (O_570,N_9932,N_9096);
or UO_571 (O_571,N_9478,N_9051);
nor UO_572 (O_572,N_9686,N_9298);
nand UO_573 (O_573,N_9324,N_9240);
nor UO_574 (O_574,N_9317,N_9124);
nor UO_575 (O_575,N_9600,N_9532);
nand UO_576 (O_576,N_9872,N_9437);
nand UO_577 (O_577,N_9043,N_9357);
and UO_578 (O_578,N_9982,N_9288);
nand UO_579 (O_579,N_9881,N_9610);
nand UO_580 (O_580,N_9231,N_9310);
nor UO_581 (O_581,N_9247,N_9108);
or UO_582 (O_582,N_9349,N_9786);
and UO_583 (O_583,N_9060,N_9117);
or UO_584 (O_584,N_9299,N_9693);
and UO_585 (O_585,N_9580,N_9527);
or UO_586 (O_586,N_9632,N_9461);
or UO_587 (O_587,N_9754,N_9853);
and UO_588 (O_588,N_9782,N_9467);
and UO_589 (O_589,N_9994,N_9166);
nand UO_590 (O_590,N_9535,N_9808);
nand UO_591 (O_591,N_9028,N_9761);
and UO_592 (O_592,N_9120,N_9551);
and UO_593 (O_593,N_9528,N_9312);
or UO_594 (O_594,N_9974,N_9720);
nand UO_595 (O_595,N_9519,N_9107);
or UO_596 (O_596,N_9124,N_9623);
nand UO_597 (O_597,N_9346,N_9172);
and UO_598 (O_598,N_9653,N_9893);
or UO_599 (O_599,N_9651,N_9616);
nor UO_600 (O_600,N_9500,N_9570);
and UO_601 (O_601,N_9055,N_9514);
nand UO_602 (O_602,N_9778,N_9030);
nor UO_603 (O_603,N_9027,N_9903);
nor UO_604 (O_604,N_9730,N_9429);
nor UO_605 (O_605,N_9078,N_9673);
and UO_606 (O_606,N_9964,N_9724);
nand UO_607 (O_607,N_9414,N_9716);
nand UO_608 (O_608,N_9069,N_9453);
and UO_609 (O_609,N_9568,N_9151);
and UO_610 (O_610,N_9121,N_9506);
nand UO_611 (O_611,N_9875,N_9444);
nand UO_612 (O_612,N_9969,N_9342);
nand UO_613 (O_613,N_9914,N_9495);
or UO_614 (O_614,N_9205,N_9462);
and UO_615 (O_615,N_9913,N_9945);
or UO_616 (O_616,N_9972,N_9923);
nor UO_617 (O_617,N_9706,N_9052);
nor UO_618 (O_618,N_9531,N_9578);
and UO_619 (O_619,N_9178,N_9352);
and UO_620 (O_620,N_9114,N_9368);
nor UO_621 (O_621,N_9983,N_9474);
nor UO_622 (O_622,N_9664,N_9280);
nand UO_623 (O_623,N_9958,N_9434);
and UO_624 (O_624,N_9075,N_9403);
nand UO_625 (O_625,N_9857,N_9026);
nand UO_626 (O_626,N_9879,N_9682);
or UO_627 (O_627,N_9577,N_9151);
nor UO_628 (O_628,N_9181,N_9481);
xor UO_629 (O_629,N_9158,N_9672);
and UO_630 (O_630,N_9947,N_9941);
nand UO_631 (O_631,N_9529,N_9252);
nor UO_632 (O_632,N_9753,N_9541);
and UO_633 (O_633,N_9943,N_9005);
or UO_634 (O_634,N_9503,N_9262);
nand UO_635 (O_635,N_9173,N_9901);
nand UO_636 (O_636,N_9382,N_9956);
and UO_637 (O_637,N_9395,N_9597);
nand UO_638 (O_638,N_9541,N_9525);
and UO_639 (O_639,N_9481,N_9851);
and UO_640 (O_640,N_9037,N_9848);
and UO_641 (O_641,N_9906,N_9035);
nand UO_642 (O_642,N_9828,N_9540);
nor UO_643 (O_643,N_9467,N_9154);
and UO_644 (O_644,N_9357,N_9620);
nor UO_645 (O_645,N_9373,N_9255);
and UO_646 (O_646,N_9074,N_9298);
xor UO_647 (O_647,N_9557,N_9120);
and UO_648 (O_648,N_9767,N_9151);
nor UO_649 (O_649,N_9764,N_9453);
nor UO_650 (O_650,N_9934,N_9931);
nor UO_651 (O_651,N_9227,N_9612);
nand UO_652 (O_652,N_9069,N_9825);
or UO_653 (O_653,N_9791,N_9477);
nor UO_654 (O_654,N_9707,N_9402);
and UO_655 (O_655,N_9022,N_9634);
or UO_656 (O_656,N_9615,N_9394);
or UO_657 (O_657,N_9520,N_9113);
or UO_658 (O_658,N_9952,N_9838);
nand UO_659 (O_659,N_9902,N_9974);
nand UO_660 (O_660,N_9340,N_9480);
nand UO_661 (O_661,N_9334,N_9738);
or UO_662 (O_662,N_9744,N_9399);
nor UO_663 (O_663,N_9498,N_9089);
and UO_664 (O_664,N_9828,N_9561);
and UO_665 (O_665,N_9178,N_9239);
or UO_666 (O_666,N_9415,N_9929);
or UO_667 (O_667,N_9901,N_9882);
and UO_668 (O_668,N_9118,N_9484);
nand UO_669 (O_669,N_9438,N_9551);
or UO_670 (O_670,N_9423,N_9121);
nor UO_671 (O_671,N_9476,N_9673);
and UO_672 (O_672,N_9751,N_9442);
xor UO_673 (O_673,N_9008,N_9797);
and UO_674 (O_674,N_9747,N_9566);
and UO_675 (O_675,N_9379,N_9191);
nor UO_676 (O_676,N_9870,N_9933);
or UO_677 (O_677,N_9767,N_9286);
nor UO_678 (O_678,N_9308,N_9692);
and UO_679 (O_679,N_9795,N_9181);
or UO_680 (O_680,N_9345,N_9884);
nand UO_681 (O_681,N_9236,N_9362);
and UO_682 (O_682,N_9069,N_9986);
or UO_683 (O_683,N_9491,N_9484);
and UO_684 (O_684,N_9177,N_9089);
nor UO_685 (O_685,N_9579,N_9361);
nand UO_686 (O_686,N_9939,N_9294);
or UO_687 (O_687,N_9636,N_9768);
and UO_688 (O_688,N_9029,N_9721);
and UO_689 (O_689,N_9639,N_9305);
nor UO_690 (O_690,N_9137,N_9451);
nand UO_691 (O_691,N_9480,N_9777);
and UO_692 (O_692,N_9020,N_9448);
nor UO_693 (O_693,N_9962,N_9149);
and UO_694 (O_694,N_9356,N_9892);
and UO_695 (O_695,N_9495,N_9618);
and UO_696 (O_696,N_9542,N_9353);
nor UO_697 (O_697,N_9280,N_9293);
and UO_698 (O_698,N_9673,N_9392);
and UO_699 (O_699,N_9864,N_9895);
nor UO_700 (O_700,N_9519,N_9195);
or UO_701 (O_701,N_9964,N_9190);
or UO_702 (O_702,N_9504,N_9372);
nor UO_703 (O_703,N_9979,N_9683);
or UO_704 (O_704,N_9505,N_9026);
and UO_705 (O_705,N_9193,N_9513);
or UO_706 (O_706,N_9635,N_9118);
and UO_707 (O_707,N_9609,N_9255);
and UO_708 (O_708,N_9558,N_9919);
and UO_709 (O_709,N_9361,N_9022);
or UO_710 (O_710,N_9355,N_9916);
or UO_711 (O_711,N_9712,N_9194);
nor UO_712 (O_712,N_9924,N_9708);
and UO_713 (O_713,N_9259,N_9052);
nor UO_714 (O_714,N_9612,N_9628);
and UO_715 (O_715,N_9912,N_9546);
and UO_716 (O_716,N_9804,N_9550);
or UO_717 (O_717,N_9092,N_9676);
and UO_718 (O_718,N_9703,N_9340);
nand UO_719 (O_719,N_9775,N_9557);
nor UO_720 (O_720,N_9774,N_9988);
and UO_721 (O_721,N_9619,N_9981);
nor UO_722 (O_722,N_9786,N_9528);
or UO_723 (O_723,N_9716,N_9838);
and UO_724 (O_724,N_9374,N_9153);
nor UO_725 (O_725,N_9102,N_9917);
and UO_726 (O_726,N_9535,N_9673);
nor UO_727 (O_727,N_9132,N_9907);
or UO_728 (O_728,N_9746,N_9805);
nand UO_729 (O_729,N_9045,N_9558);
nor UO_730 (O_730,N_9821,N_9969);
or UO_731 (O_731,N_9010,N_9013);
nand UO_732 (O_732,N_9165,N_9216);
nor UO_733 (O_733,N_9281,N_9643);
nand UO_734 (O_734,N_9707,N_9978);
or UO_735 (O_735,N_9226,N_9568);
and UO_736 (O_736,N_9139,N_9308);
or UO_737 (O_737,N_9232,N_9532);
and UO_738 (O_738,N_9715,N_9085);
and UO_739 (O_739,N_9317,N_9744);
or UO_740 (O_740,N_9988,N_9497);
nand UO_741 (O_741,N_9108,N_9097);
and UO_742 (O_742,N_9259,N_9951);
nand UO_743 (O_743,N_9530,N_9704);
xnor UO_744 (O_744,N_9319,N_9624);
nor UO_745 (O_745,N_9779,N_9702);
and UO_746 (O_746,N_9664,N_9425);
or UO_747 (O_747,N_9440,N_9788);
nand UO_748 (O_748,N_9873,N_9989);
nand UO_749 (O_749,N_9193,N_9370);
xnor UO_750 (O_750,N_9073,N_9163);
or UO_751 (O_751,N_9495,N_9746);
or UO_752 (O_752,N_9202,N_9018);
nor UO_753 (O_753,N_9612,N_9955);
nand UO_754 (O_754,N_9968,N_9583);
and UO_755 (O_755,N_9196,N_9591);
nand UO_756 (O_756,N_9442,N_9714);
xor UO_757 (O_757,N_9968,N_9600);
or UO_758 (O_758,N_9999,N_9821);
nor UO_759 (O_759,N_9599,N_9558);
and UO_760 (O_760,N_9788,N_9113);
and UO_761 (O_761,N_9516,N_9963);
or UO_762 (O_762,N_9160,N_9364);
nand UO_763 (O_763,N_9785,N_9402);
nor UO_764 (O_764,N_9485,N_9411);
xnor UO_765 (O_765,N_9079,N_9118);
and UO_766 (O_766,N_9962,N_9438);
nand UO_767 (O_767,N_9190,N_9594);
nor UO_768 (O_768,N_9075,N_9320);
nand UO_769 (O_769,N_9676,N_9481);
nand UO_770 (O_770,N_9802,N_9089);
nor UO_771 (O_771,N_9565,N_9025);
or UO_772 (O_772,N_9636,N_9800);
nand UO_773 (O_773,N_9441,N_9120);
nand UO_774 (O_774,N_9004,N_9976);
nor UO_775 (O_775,N_9820,N_9198);
nor UO_776 (O_776,N_9019,N_9253);
nand UO_777 (O_777,N_9700,N_9902);
or UO_778 (O_778,N_9597,N_9454);
or UO_779 (O_779,N_9336,N_9730);
nand UO_780 (O_780,N_9366,N_9473);
nor UO_781 (O_781,N_9414,N_9995);
nand UO_782 (O_782,N_9174,N_9349);
and UO_783 (O_783,N_9343,N_9326);
and UO_784 (O_784,N_9804,N_9644);
xnor UO_785 (O_785,N_9827,N_9452);
and UO_786 (O_786,N_9761,N_9537);
or UO_787 (O_787,N_9369,N_9455);
or UO_788 (O_788,N_9879,N_9206);
and UO_789 (O_789,N_9762,N_9910);
nand UO_790 (O_790,N_9244,N_9415);
or UO_791 (O_791,N_9056,N_9579);
or UO_792 (O_792,N_9980,N_9144);
nand UO_793 (O_793,N_9070,N_9846);
nor UO_794 (O_794,N_9046,N_9608);
and UO_795 (O_795,N_9764,N_9667);
or UO_796 (O_796,N_9607,N_9694);
or UO_797 (O_797,N_9861,N_9368);
or UO_798 (O_798,N_9338,N_9941);
nor UO_799 (O_799,N_9664,N_9034);
or UO_800 (O_800,N_9420,N_9842);
and UO_801 (O_801,N_9406,N_9906);
nor UO_802 (O_802,N_9495,N_9463);
nand UO_803 (O_803,N_9647,N_9492);
and UO_804 (O_804,N_9054,N_9253);
nand UO_805 (O_805,N_9726,N_9167);
nor UO_806 (O_806,N_9453,N_9566);
nand UO_807 (O_807,N_9169,N_9638);
nand UO_808 (O_808,N_9507,N_9604);
nand UO_809 (O_809,N_9217,N_9396);
nor UO_810 (O_810,N_9723,N_9717);
or UO_811 (O_811,N_9723,N_9015);
and UO_812 (O_812,N_9883,N_9150);
or UO_813 (O_813,N_9795,N_9560);
and UO_814 (O_814,N_9759,N_9111);
and UO_815 (O_815,N_9148,N_9022);
nand UO_816 (O_816,N_9182,N_9682);
nand UO_817 (O_817,N_9233,N_9362);
nor UO_818 (O_818,N_9626,N_9458);
and UO_819 (O_819,N_9899,N_9797);
nor UO_820 (O_820,N_9500,N_9518);
nand UO_821 (O_821,N_9620,N_9750);
or UO_822 (O_822,N_9699,N_9729);
or UO_823 (O_823,N_9591,N_9185);
nor UO_824 (O_824,N_9952,N_9139);
and UO_825 (O_825,N_9410,N_9582);
nand UO_826 (O_826,N_9280,N_9925);
nor UO_827 (O_827,N_9023,N_9378);
and UO_828 (O_828,N_9954,N_9850);
nor UO_829 (O_829,N_9203,N_9873);
nand UO_830 (O_830,N_9374,N_9506);
nand UO_831 (O_831,N_9915,N_9255);
nand UO_832 (O_832,N_9644,N_9539);
nand UO_833 (O_833,N_9183,N_9804);
nor UO_834 (O_834,N_9489,N_9764);
nor UO_835 (O_835,N_9525,N_9253);
nor UO_836 (O_836,N_9561,N_9490);
nand UO_837 (O_837,N_9693,N_9354);
and UO_838 (O_838,N_9939,N_9091);
or UO_839 (O_839,N_9503,N_9265);
nor UO_840 (O_840,N_9661,N_9779);
nor UO_841 (O_841,N_9527,N_9254);
and UO_842 (O_842,N_9220,N_9252);
or UO_843 (O_843,N_9309,N_9742);
xor UO_844 (O_844,N_9908,N_9557);
xor UO_845 (O_845,N_9568,N_9671);
and UO_846 (O_846,N_9412,N_9434);
nand UO_847 (O_847,N_9162,N_9986);
and UO_848 (O_848,N_9342,N_9886);
or UO_849 (O_849,N_9259,N_9534);
nand UO_850 (O_850,N_9146,N_9557);
xnor UO_851 (O_851,N_9010,N_9909);
and UO_852 (O_852,N_9051,N_9792);
or UO_853 (O_853,N_9801,N_9824);
nor UO_854 (O_854,N_9987,N_9344);
nor UO_855 (O_855,N_9060,N_9587);
and UO_856 (O_856,N_9982,N_9135);
nor UO_857 (O_857,N_9476,N_9231);
or UO_858 (O_858,N_9805,N_9024);
or UO_859 (O_859,N_9995,N_9994);
nor UO_860 (O_860,N_9403,N_9267);
nand UO_861 (O_861,N_9932,N_9704);
and UO_862 (O_862,N_9601,N_9246);
nor UO_863 (O_863,N_9757,N_9900);
or UO_864 (O_864,N_9768,N_9225);
or UO_865 (O_865,N_9576,N_9447);
nand UO_866 (O_866,N_9508,N_9214);
nand UO_867 (O_867,N_9175,N_9114);
and UO_868 (O_868,N_9959,N_9147);
nor UO_869 (O_869,N_9553,N_9489);
and UO_870 (O_870,N_9666,N_9707);
or UO_871 (O_871,N_9199,N_9652);
nand UO_872 (O_872,N_9141,N_9361);
nand UO_873 (O_873,N_9970,N_9669);
or UO_874 (O_874,N_9663,N_9211);
xnor UO_875 (O_875,N_9730,N_9113);
and UO_876 (O_876,N_9650,N_9930);
or UO_877 (O_877,N_9370,N_9783);
nor UO_878 (O_878,N_9476,N_9219);
and UO_879 (O_879,N_9455,N_9712);
xnor UO_880 (O_880,N_9043,N_9508);
nor UO_881 (O_881,N_9764,N_9364);
and UO_882 (O_882,N_9165,N_9953);
nand UO_883 (O_883,N_9648,N_9159);
nand UO_884 (O_884,N_9570,N_9853);
and UO_885 (O_885,N_9092,N_9499);
xor UO_886 (O_886,N_9888,N_9713);
xor UO_887 (O_887,N_9503,N_9715);
and UO_888 (O_888,N_9764,N_9207);
nand UO_889 (O_889,N_9585,N_9139);
nand UO_890 (O_890,N_9757,N_9926);
and UO_891 (O_891,N_9460,N_9502);
or UO_892 (O_892,N_9701,N_9750);
nand UO_893 (O_893,N_9079,N_9639);
nor UO_894 (O_894,N_9055,N_9670);
and UO_895 (O_895,N_9776,N_9727);
or UO_896 (O_896,N_9591,N_9468);
nand UO_897 (O_897,N_9090,N_9400);
and UO_898 (O_898,N_9052,N_9103);
nor UO_899 (O_899,N_9984,N_9437);
or UO_900 (O_900,N_9868,N_9560);
nand UO_901 (O_901,N_9759,N_9261);
nand UO_902 (O_902,N_9824,N_9040);
nor UO_903 (O_903,N_9866,N_9343);
nor UO_904 (O_904,N_9395,N_9901);
nor UO_905 (O_905,N_9755,N_9568);
nor UO_906 (O_906,N_9125,N_9226);
nand UO_907 (O_907,N_9035,N_9165);
xnor UO_908 (O_908,N_9602,N_9412);
and UO_909 (O_909,N_9913,N_9960);
nand UO_910 (O_910,N_9443,N_9015);
or UO_911 (O_911,N_9431,N_9859);
nor UO_912 (O_912,N_9589,N_9540);
xnor UO_913 (O_913,N_9508,N_9826);
and UO_914 (O_914,N_9896,N_9909);
nor UO_915 (O_915,N_9690,N_9786);
or UO_916 (O_916,N_9628,N_9024);
nand UO_917 (O_917,N_9555,N_9686);
nand UO_918 (O_918,N_9739,N_9539);
nand UO_919 (O_919,N_9229,N_9417);
and UO_920 (O_920,N_9125,N_9475);
nor UO_921 (O_921,N_9905,N_9996);
nand UO_922 (O_922,N_9079,N_9358);
nor UO_923 (O_923,N_9410,N_9066);
nor UO_924 (O_924,N_9752,N_9989);
and UO_925 (O_925,N_9014,N_9368);
and UO_926 (O_926,N_9627,N_9617);
and UO_927 (O_927,N_9783,N_9346);
xor UO_928 (O_928,N_9610,N_9560);
and UO_929 (O_929,N_9281,N_9207);
and UO_930 (O_930,N_9737,N_9941);
nor UO_931 (O_931,N_9329,N_9887);
nand UO_932 (O_932,N_9936,N_9010);
nor UO_933 (O_933,N_9877,N_9129);
or UO_934 (O_934,N_9589,N_9783);
or UO_935 (O_935,N_9934,N_9551);
and UO_936 (O_936,N_9654,N_9632);
nand UO_937 (O_937,N_9104,N_9965);
nand UO_938 (O_938,N_9884,N_9859);
or UO_939 (O_939,N_9595,N_9764);
or UO_940 (O_940,N_9707,N_9174);
or UO_941 (O_941,N_9483,N_9324);
nand UO_942 (O_942,N_9347,N_9670);
or UO_943 (O_943,N_9115,N_9034);
or UO_944 (O_944,N_9461,N_9782);
nand UO_945 (O_945,N_9652,N_9701);
or UO_946 (O_946,N_9338,N_9998);
nand UO_947 (O_947,N_9488,N_9513);
and UO_948 (O_948,N_9362,N_9218);
nor UO_949 (O_949,N_9154,N_9563);
and UO_950 (O_950,N_9434,N_9202);
and UO_951 (O_951,N_9973,N_9257);
or UO_952 (O_952,N_9443,N_9125);
nor UO_953 (O_953,N_9940,N_9100);
or UO_954 (O_954,N_9685,N_9131);
nand UO_955 (O_955,N_9924,N_9780);
xor UO_956 (O_956,N_9803,N_9817);
or UO_957 (O_957,N_9603,N_9216);
or UO_958 (O_958,N_9688,N_9889);
nand UO_959 (O_959,N_9520,N_9238);
nor UO_960 (O_960,N_9340,N_9638);
or UO_961 (O_961,N_9400,N_9251);
nor UO_962 (O_962,N_9000,N_9401);
nand UO_963 (O_963,N_9407,N_9503);
or UO_964 (O_964,N_9785,N_9057);
nand UO_965 (O_965,N_9213,N_9878);
and UO_966 (O_966,N_9814,N_9357);
or UO_967 (O_967,N_9159,N_9835);
nor UO_968 (O_968,N_9683,N_9058);
or UO_969 (O_969,N_9744,N_9871);
or UO_970 (O_970,N_9507,N_9181);
and UO_971 (O_971,N_9594,N_9616);
and UO_972 (O_972,N_9792,N_9694);
and UO_973 (O_973,N_9435,N_9478);
or UO_974 (O_974,N_9961,N_9739);
nor UO_975 (O_975,N_9809,N_9017);
and UO_976 (O_976,N_9243,N_9226);
or UO_977 (O_977,N_9827,N_9772);
and UO_978 (O_978,N_9578,N_9295);
or UO_979 (O_979,N_9503,N_9158);
and UO_980 (O_980,N_9695,N_9884);
nand UO_981 (O_981,N_9595,N_9433);
or UO_982 (O_982,N_9782,N_9099);
or UO_983 (O_983,N_9633,N_9997);
nor UO_984 (O_984,N_9488,N_9401);
or UO_985 (O_985,N_9142,N_9309);
and UO_986 (O_986,N_9330,N_9410);
and UO_987 (O_987,N_9710,N_9451);
and UO_988 (O_988,N_9813,N_9910);
and UO_989 (O_989,N_9614,N_9847);
or UO_990 (O_990,N_9474,N_9591);
nor UO_991 (O_991,N_9296,N_9981);
and UO_992 (O_992,N_9200,N_9495);
nand UO_993 (O_993,N_9525,N_9870);
or UO_994 (O_994,N_9957,N_9017);
nand UO_995 (O_995,N_9552,N_9825);
nand UO_996 (O_996,N_9087,N_9634);
or UO_997 (O_997,N_9659,N_9149);
nand UO_998 (O_998,N_9250,N_9002);
or UO_999 (O_999,N_9555,N_9197);
or UO_1000 (O_1000,N_9219,N_9677);
or UO_1001 (O_1001,N_9308,N_9819);
nor UO_1002 (O_1002,N_9114,N_9701);
nand UO_1003 (O_1003,N_9654,N_9886);
and UO_1004 (O_1004,N_9677,N_9795);
and UO_1005 (O_1005,N_9954,N_9867);
or UO_1006 (O_1006,N_9422,N_9419);
nand UO_1007 (O_1007,N_9721,N_9177);
and UO_1008 (O_1008,N_9353,N_9302);
or UO_1009 (O_1009,N_9096,N_9551);
or UO_1010 (O_1010,N_9140,N_9341);
or UO_1011 (O_1011,N_9689,N_9137);
nor UO_1012 (O_1012,N_9409,N_9410);
and UO_1013 (O_1013,N_9828,N_9213);
nor UO_1014 (O_1014,N_9073,N_9189);
and UO_1015 (O_1015,N_9723,N_9625);
and UO_1016 (O_1016,N_9271,N_9926);
and UO_1017 (O_1017,N_9410,N_9571);
nand UO_1018 (O_1018,N_9663,N_9223);
nor UO_1019 (O_1019,N_9471,N_9058);
or UO_1020 (O_1020,N_9131,N_9689);
and UO_1021 (O_1021,N_9841,N_9621);
nand UO_1022 (O_1022,N_9711,N_9114);
nor UO_1023 (O_1023,N_9138,N_9409);
nand UO_1024 (O_1024,N_9435,N_9615);
xor UO_1025 (O_1025,N_9702,N_9972);
nand UO_1026 (O_1026,N_9841,N_9492);
nand UO_1027 (O_1027,N_9841,N_9952);
nor UO_1028 (O_1028,N_9376,N_9392);
nand UO_1029 (O_1029,N_9331,N_9684);
and UO_1030 (O_1030,N_9241,N_9250);
and UO_1031 (O_1031,N_9193,N_9996);
nor UO_1032 (O_1032,N_9029,N_9933);
or UO_1033 (O_1033,N_9857,N_9818);
nor UO_1034 (O_1034,N_9241,N_9130);
nand UO_1035 (O_1035,N_9202,N_9971);
nand UO_1036 (O_1036,N_9640,N_9176);
nand UO_1037 (O_1037,N_9006,N_9661);
and UO_1038 (O_1038,N_9890,N_9181);
and UO_1039 (O_1039,N_9874,N_9700);
nor UO_1040 (O_1040,N_9786,N_9189);
nand UO_1041 (O_1041,N_9439,N_9978);
and UO_1042 (O_1042,N_9981,N_9544);
nand UO_1043 (O_1043,N_9572,N_9762);
and UO_1044 (O_1044,N_9515,N_9426);
nor UO_1045 (O_1045,N_9033,N_9285);
or UO_1046 (O_1046,N_9392,N_9861);
nand UO_1047 (O_1047,N_9975,N_9018);
nor UO_1048 (O_1048,N_9365,N_9241);
and UO_1049 (O_1049,N_9937,N_9228);
or UO_1050 (O_1050,N_9848,N_9865);
or UO_1051 (O_1051,N_9839,N_9991);
xor UO_1052 (O_1052,N_9151,N_9274);
nor UO_1053 (O_1053,N_9836,N_9024);
or UO_1054 (O_1054,N_9103,N_9002);
or UO_1055 (O_1055,N_9466,N_9330);
or UO_1056 (O_1056,N_9667,N_9525);
nor UO_1057 (O_1057,N_9131,N_9565);
nand UO_1058 (O_1058,N_9235,N_9540);
nor UO_1059 (O_1059,N_9912,N_9130);
and UO_1060 (O_1060,N_9727,N_9634);
nand UO_1061 (O_1061,N_9145,N_9596);
and UO_1062 (O_1062,N_9708,N_9738);
and UO_1063 (O_1063,N_9559,N_9916);
nand UO_1064 (O_1064,N_9620,N_9922);
nand UO_1065 (O_1065,N_9426,N_9846);
nand UO_1066 (O_1066,N_9988,N_9510);
nand UO_1067 (O_1067,N_9828,N_9961);
nand UO_1068 (O_1068,N_9838,N_9548);
nand UO_1069 (O_1069,N_9628,N_9004);
xnor UO_1070 (O_1070,N_9130,N_9488);
nor UO_1071 (O_1071,N_9307,N_9078);
xnor UO_1072 (O_1072,N_9815,N_9599);
nor UO_1073 (O_1073,N_9992,N_9460);
or UO_1074 (O_1074,N_9312,N_9620);
nor UO_1075 (O_1075,N_9584,N_9978);
and UO_1076 (O_1076,N_9165,N_9254);
and UO_1077 (O_1077,N_9295,N_9521);
nor UO_1078 (O_1078,N_9535,N_9029);
and UO_1079 (O_1079,N_9813,N_9386);
and UO_1080 (O_1080,N_9918,N_9478);
nor UO_1081 (O_1081,N_9883,N_9652);
nand UO_1082 (O_1082,N_9041,N_9608);
nand UO_1083 (O_1083,N_9111,N_9009);
or UO_1084 (O_1084,N_9213,N_9449);
nand UO_1085 (O_1085,N_9117,N_9362);
nor UO_1086 (O_1086,N_9010,N_9147);
or UO_1087 (O_1087,N_9980,N_9161);
and UO_1088 (O_1088,N_9042,N_9659);
nor UO_1089 (O_1089,N_9693,N_9924);
and UO_1090 (O_1090,N_9782,N_9188);
nand UO_1091 (O_1091,N_9924,N_9827);
nand UO_1092 (O_1092,N_9194,N_9740);
and UO_1093 (O_1093,N_9415,N_9471);
nand UO_1094 (O_1094,N_9367,N_9297);
and UO_1095 (O_1095,N_9157,N_9928);
nand UO_1096 (O_1096,N_9519,N_9906);
nor UO_1097 (O_1097,N_9062,N_9757);
or UO_1098 (O_1098,N_9777,N_9633);
and UO_1099 (O_1099,N_9259,N_9840);
nand UO_1100 (O_1100,N_9897,N_9122);
nand UO_1101 (O_1101,N_9538,N_9592);
or UO_1102 (O_1102,N_9421,N_9498);
nor UO_1103 (O_1103,N_9824,N_9147);
nor UO_1104 (O_1104,N_9418,N_9703);
nor UO_1105 (O_1105,N_9706,N_9330);
nand UO_1106 (O_1106,N_9125,N_9825);
and UO_1107 (O_1107,N_9968,N_9730);
and UO_1108 (O_1108,N_9404,N_9478);
nand UO_1109 (O_1109,N_9361,N_9498);
or UO_1110 (O_1110,N_9607,N_9853);
nand UO_1111 (O_1111,N_9092,N_9627);
nor UO_1112 (O_1112,N_9326,N_9190);
nand UO_1113 (O_1113,N_9641,N_9455);
nand UO_1114 (O_1114,N_9085,N_9819);
nor UO_1115 (O_1115,N_9131,N_9543);
nor UO_1116 (O_1116,N_9617,N_9686);
nor UO_1117 (O_1117,N_9906,N_9742);
and UO_1118 (O_1118,N_9542,N_9332);
nor UO_1119 (O_1119,N_9040,N_9251);
and UO_1120 (O_1120,N_9819,N_9488);
nor UO_1121 (O_1121,N_9002,N_9538);
nand UO_1122 (O_1122,N_9268,N_9651);
nand UO_1123 (O_1123,N_9181,N_9098);
or UO_1124 (O_1124,N_9304,N_9462);
and UO_1125 (O_1125,N_9910,N_9722);
and UO_1126 (O_1126,N_9160,N_9853);
nand UO_1127 (O_1127,N_9403,N_9967);
nor UO_1128 (O_1128,N_9681,N_9752);
nor UO_1129 (O_1129,N_9313,N_9657);
nand UO_1130 (O_1130,N_9139,N_9920);
and UO_1131 (O_1131,N_9448,N_9812);
nand UO_1132 (O_1132,N_9507,N_9355);
and UO_1133 (O_1133,N_9969,N_9667);
and UO_1134 (O_1134,N_9599,N_9309);
nand UO_1135 (O_1135,N_9524,N_9683);
and UO_1136 (O_1136,N_9395,N_9171);
nand UO_1137 (O_1137,N_9609,N_9739);
and UO_1138 (O_1138,N_9522,N_9311);
nor UO_1139 (O_1139,N_9406,N_9910);
nand UO_1140 (O_1140,N_9337,N_9981);
nand UO_1141 (O_1141,N_9502,N_9424);
or UO_1142 (O_1142,N_9110,N_9873);
and UO_1143 (O_1143,N_9316,N_9992);
nor UO_1144 (O_1144,N_9980,N_9583);
nor UO_1145 (O_1145,N_9325,N_9646);
nand UO_1146 (O_1146,N_9509,N_9464);
or UO_1147 (O_1147,N_9949,N_9079);
nand UO_1148 (O_1148,N_9828,N_9836);
nor UO_1149 (O_1149,N_9593,N_9006);
or UO_1150 (O_1150,N_9060,N_9430);
nor UO_1151 (O_1151,N_9617,N_9260);
nor UO_1152 (O_1152,N_9543,N_9786);
or UO_1153 (O_1153,N_9160,N_9248);
nor UO_1154 (O_1154,N_9279,N_9481);
nor UO_1155 (O_1155,N_9435,N_9243);
nand UO_1156 (O_1156,N_9963,N_9535);
and UO_1157 (O_1157,N_9568,N_9088);
nor UO_1158 (O_1158,N_9242,N_9974);
and UO_1159 (O_1159,N_9621,N_9431);
and UO_1160 (O_1160,N_9224,N_9853);
nor UO_1161 (O_1161,N_9010,N_9741);
nor UO_1162 (O_1162,N_9083,N_9886);
and UO_1163 (O_1163,N_9726,N_9506);
and UO_1164 (O_1164,N_9860,N_9559);
nand UO_1165 (O_1165,N_9670,N_9695);
or UO_1166 (O_1166,N_9485,N_9062);
and UO_1167 (O_1167,N_9197,N_9226);
and UO_1168 (O_1168,N_9203,N_9404);
or UO_1169 (O_1169,N_9735,N_9153);
nand UO_1170 (O_1170,N_9676,N_9268);
nand UO_1171 (O_1171,N_9352,N_9713);
nor UO_1172 (O_1172,N_9509,N_9568);
nand UO_1173 (O_1173,N_9146,N_9662);
or UO_1174 (O_1174,N_9220,N_9705);
and UO_1175 (O_1175,N_9225,N_9992);
or UO_1176 (O_1176,N_9506,N_9204);
nor UO_1177 (O_1177,N_9816,N_9089);
and UO_1178 (O_1178,N_9461,N_9039);
nand UO_1179 (O_1179,N_9094,N_9693);
or UO_1180 (O_1180,N_9898,N_9521);
nand UO_1181 (O_1181,N_9532,N_9706);
nor UO_1182 (O_1182,N_9271,N_9998);
or UO_1183 (O_1183,N_9525,N_9147);
nor UO_1184 (O_1184,N_9055,N_9693);
and UO_1185 (O_1185,N_9743,N_9411);
or UO_1186 (O_1186,N_9550,N_9596);
nor UO_1187 (O_1187,N_9726,N_9306);
or UO_1188 (O_1188,N_9762,N_9242);
or UO_1189 (O_1189,N_9284,N_9680);
nand UO_1190 (O_1190,N_9241,N_9268);
nor UO_1191 (O_1191,N_9803,N_9806);
and UO_1192 (O_1192,N_9884,N_9267);
or UO_1193 (O_1193,N_9843,N_9633);
nand UO_1194 (O_1194,N_9940,N_9905);
or UO_1195 (O_1195,N_9901,N_9144);
and UO_1196 (O_1196,N_9645,N_9095);
nor UO_1197 (O_1197,N_9596,N_9894);
nand UO_1198 (O_1198,N_9011,N_9996);
nor UO_1199 (O_1199,N_9089,N_9646);
nand UO_1200 (O_1200,N_9833,N_9128);
or UO_1201 (O_1201,N_9885,N_9306);
nor UO_1202 (O_1202,N_9875,N_9807);
nand UO_1203 (O_1203,N_9689,N_9328);
nor UO_1204 (O_1204,N_9672,N_9388);
and UO_1205 (O_1205,N_9506,N_9821);
nand UO_1206 (O_1206,N_9429,N_9899);
nand UO_1207 (O_1207,N_9845,N_9041);
nand UO_1208 (O_1208,N_9027,N_9288);
nand UO_1209 (O_1209,N_9713,N_9465);
xnor UO_1210 (O_1210,N_9845,N_9894);
nor UO_1211 (O_1211,N_9333,N_9673);
nand UO_1212 (O_1212,N_9119,N_9139);
nand UO_1213 (O_1213,N_9210,N_9277);
nor UO_1214 (O_1214,N_9956,N_9349);
and UO_1215 (O_1215,N_9337,N_9017);
or UO_1216 (O_1216,N_9606,N_9789);
nand UO_1217 (O_1217,N_9300,N_9063);
nor UO_1218 (O_1218,N_9669,N_9960);
and UO_1219 (O_1219,N_9782,N_9307);
xor UO_1220 (O_1220,N_9025,N_9804);
nor UO_1221 (O_1221,N_9558,N_9793);
nor UO_1222 (O_1222,N_9096,N_9413);
or UO_1223 (O_1223,N_9002,N_9403);
nand UO_1224 (O_1224,N_9152,N_9783);
or UO_1225 (O_1225,N_9902,N_9041);
nor UO_1226 (O_1226,N_9411,N_9578);
nand UO_1227 (O_1227,N_9241,N_9535);
nor UO_1228 (O_1228,N_9775,N_9349);
or UO_1229 (O_1229,N_9405,N_9318);
nor UO_1230 (O_1230,N_9152,N_9466);
and UO_1231 (O_1231,N_9495,N_9466);
or UO_1232 (O_1232,N_9564,N_9271);
and UO_1233 (O_1233,N_9490,N_9039);
nand UO_1234 (O_1234,N_9433,N_9873);
nor UO_1235 (O_1235,N_9939,N_9208);
nor UO_1236 (O_1236,N_9997,N_9789);
nor UO_1237 (O_1237,N_9615,N_9031);
nor UO_1238 (O_1238,N_9213,N_9290);
and UO_1239 (O_1239,N_9444,N_9359);
and UO_1240 (O_1240,N_9230,N_9493);
and UO_1241 (O_1241,N_9133,N_9299);
and UO_1242 (O_1242,N_9716,N_9975);
nor UO_1243 (O_1243,N_9608,N_9581);
nand UO_1244 (O_1244,N_9276,N_9423);
nor UO_1245 (O_1245,N_9710,N_9132);
or UO_1246 (O_1246,N_9508,N_9181);
or UO_1247 (O_1247,N_9971,N_9304);
nand UO_1248 (O_1248,N_9529,N_9465);
nand UO_1249 (O_1249,N_9849,N_9433);
nand UO_1250 (O_1250,N_9317,N_9115);
or UO_1251 (O_1251,N_9364,N_9925);
and UO_1252 (O_1252,N_9398,N_9301);
xnor UO_1253 (O_1253,N_9866,N_9516);
and UO_1254 (O_1254,N_9764,N_9325);
nand UO_1255 (O_1255,N_9571,N_9459);
or UO_1256 (O_1256,N_9234,N_9026);
or UO_1257 (O_1257,N_9060,N_9213);
nand UO_1258 (O_1258,N_9976,N_9302);
nor UO_1259 (O_1259,N_9124,N_9741);
nor UO_1260 (O_1260,N_9869,N_9113);
and UO_1261 (O_1261,N_9585,N_9882);
nor UO_1262 (O_1262,N_9594,N_9648);
nand UO_1263 (O_1263,N_9352,N_9070);
nand UO_1264 (O_1264,N_9074,N_9697);
or UO_1265 (O_1265,N_9607,N_9730);
nand UO_1266 (O_1266,N_9190,N_9493);
nor UO_1267 (O_1267,N_9593,N_9799);
or UO_1268 (O_1268,N_9036,N_9373);
or UO_1269 (O_1269,N_9470,N_9327);
nor UO_1270 (O_1270,N_9645,N_9702);
nor UO_1271 (O_1271,N_9532,N_9150);
nor UO_1272 (O_1272,N_9876,N_9774);
nand UO_1273 (O_1273,N_9457,N_9204);
nor UO_1274 (O_1274,N_9035,N_9744);
and UO_1275 (O_1275,N_9478,N_9111);
nand UO_1276 (O_1276,N_9949,N_9376);
and UO_1277 (O_1277,N_9411,N_9784);
and UO_1278 (O_1278,N_9386,N_9884);
or UO_1279 (O_1279,N_9238,N_9170);
nand UO_1280 (O_1280,N_9910,N_9384);
and UO_1281 (O_1281,N_9399,N_9645);
nand UO_1282 (O_1282,N_9925,N_9451);
or UO_1283 (O_1283,N_9125,N_9949);
nor UO_1284 (O_1284,N_9233,N_9786);
nor UO_1285 (O_1285,N_9276,N_9523);
nand UO_1286 (O_1286,N_9447,N_9254);
and UO_1287 (O_1287,N_9330,N_9144);
nand UO_1288 (O_1288,N_9658,N_9211);
or UO_1289 (O_1289,N_9633,N_9836);
nor UO_1290 (O_1290,N_9427,N_9157);
and UO_1291 (O_1291,N_9055,N_9396);
nand UO_1292 (O_1292,N_9950,N_9732);
nor UO_1293 (O_1293,N_9719,N_9257);
xnor UO_1294 (O_1294,N_9096,N_9865);
and UO_1295 (O_1295,N_9909,N_9926);
nand UO_1296 (O_1296,N_9380,N_9092);
nor UO_1297 (O_1297,N_9965,N_9370);
nor UO_1298 (O_1298,N_9047,N_9310);
and UO_1299 (O_1299,N_9776,N_9480);
or UO_1300 (O_1300,N_9320,N_9846);
and UO_1301 (O_1301,N_9226,N_9012);
nor UO_1302 (O_1302,N_9450,N_9142);
or UO_1303 (O_1303,N_9282,N_9898);
nor UO_1304 (O_1304,N_9764,N_9260);
and UO_1305 (O_1305,N_9665,N_9986);
nand UO_1306 (O_1306,N_9380,N_9585);
nor UO_1307 (O_1307,N_9949,N_9916);
and UO_1308 (O_1308,N_9939,N_9781);
or UO_1309 (O_1309,N_9278,N_9308);
nand UO_1310 (O_1310,N_9402,N_9683);
and UO_1311 (O_1311,N_9935,N_9436);
nand UO_1312 (O_1312,N_9769,N_9312);
xnor UO_1313 (O_1313,N_9203,N_9657);
nand UO_1314 (O_1314,N_9202,N_9801);
nor UO_1315 (O_1315,N_9890,N_9081);
xor UO_1316 (O_1316,N_9472,N_9029);
and UO_1317 (O_1317,N_9184,N_9002);
nor UO_1318 (O_1318,N_9523,N_9517);
nand UO_1319 (O_1319,N_9303,N_9221);
xor UO_1320 (O_1320,N_9671,N_9090);
nand UO_1321 (O_1321,N_9175,N_9013);
or UO_1322 (O_1322,N_9816,N_9888);
nor UO_1323 (O_1323,N_9099,N_9643);
and UO_1324 (O_1324,N_9243,N_9699);
xnor UO_1325 (O_1325,N_9814,N_9704);
nand UO_1326 (O_1326,N_9776,N_9636);
nor UO_1327 (O_1327,N_9967,N_9676);
nand UO_1328 (O_1328,N_9959,N_9440);
nor UO_1329 (O_1329,N_9840,N_9031);
nor UO_1330 (O_1330,N_9996,N_9889);
or UO_1331 (O_1331,N_9284,N_9090);
or UO_1332 (O_1332,N_9571,N_9319);
nand UO_1333 (O_1333,N_9454,N_9798);
and UO_1334 (O_1334,N_9026,N_9272);
nor UO_1335 (O_1335,N_9261,N_9086);
and UO_1336 (O_1336,N_9671,N_9894);
and UO_1337 (O_1337,N_9075,N_9744);
and UO_1338 (O_1338,N_9751,N_9136);
and UO_1339 (O_1339,N_9632,N_9764);
nand UO_1340 (O_1340,N_9694,N_9815);
or UO_1341 (O_1341,N_9225,N_9755);
and UO_1342 (O_1342,N_9323,N_9690);
and UO_1343 (O_1343,N_9396,N_9786);
nand UO_1344 (O_1344,N_9974,N_9276);
nor UO_1345 (O_1345,N_9594,N_9986);
and UO_1346 (O_1346,N_9950,N_9059);
nor UO_1347 (O_1347,N_9035,N_9073);
or UO_1348 (O_1348,N_9828,N_9482);
nand UO_1349 (O_1349,N_9220,N_9131);
nand UO_1350 (O_1350,N_9912,N_9085);
or UO_1351 (O_1351,N_9137,N_9674);
nand UO_1352 (O_1352,N_9698,N_9768);
nand UO_1353 (O_1353,N_9930,N_9178);
nor UO_1354 (O_1354,N_9456,N_9131);
nand UO_1355 (O_1355,N_9121,N_9228);
nand UO_1356 (O_1356,N_9141,N_9318);
nor UO_1357 (O_1357,N_9828,N_9480);
nand UO_1358 (O_1358,N_9539,N_9572);
nand UO_1359 (O_1359,N_9964,N_9894);
nor UO_1360 (O_1360,N_9144,N_9599);
nor UO_1361 (O_1361,N_9665,N_9725);
nor UO_1362 (O_1362,N_9923,N_9049);
or UO_1363 (O_1363,N_9500,N_9649);
nand UO_1364 (O_1364,N_9833,N_9121);
and UO_1365 (O_1365,N_9677,N_9509);
and UO_1366 (O_1366,N_9697,N_9420);
nand UO_1367 (O_1367,N_9404,N_9320);
nor UO_1368 (O_1368,N_9398,N_9842);
or UO_1369 (O_1369,N_9884,N_9005);
nor UO_1370 (O_1370,N_9565,N_9550);
and UO_1371 (O_1371,N_9742,N_9388);
nand UO_1372 (O_1372,N_9119,N_9600);
and UO_1373 (O_1373,N_9032,N_9129);
xor UO_1374 (O_1374,N_9555,N_9991);
or UO_1375 (O_1375,N_9524,N_9544);
or UO_1376 (O_1376,N_9051,N_9643);
nor UO_1377 (O_1377,N_9961,N_9008);
nand UO_1378 (O_1378,N_9768,N_9604);
nand UO_1379 (O_1379,N_9094,N_9229);
nor UO_1380 (O_1380,N_9436,N_9865);
nor UO_1381 (O_1381,N_9235,N_9188);
nand UO_1382 (O_1382,N_9268,N_9961);
and UO_1383 (O_1383,N_9112,N_9593);
nand UO_1384 (O_1384,N_9378,N_9235);
nor UO_1385 (O_1385,N_9732,N_9273);
nor UO_1386 (O_1386,N_9903,N_9712);
or UO_1387 (O_1387,N_9065,N_9708);
nand UO_1388 (O_1388,N_9267,N_9363);
nand UO_1389 (O_1389,N_9959,N_9900);
and UO_1390 (O_1390,N_9322,N_9327);
nor UO_1391 (O_1391,N_9753,N_9479);
nor UO_1392 (O_1392,N_9813,N_9185);
nand UO_1393 (O_1393,N_9139,N_9885);
and UO_1394 (O_1394,N_9789,N_9102);
nor UO_1395 (O_1395,N_9547,N_9711);
and UO_1396 (O_1396,N_9340,N_9716);
or UO_1397 (O_1397,N_9379,N_9079);
nand UO_1398 (O_1398,N_9058,N_9895);
nor UO_1399 (O_1399,N_9134,N_9126);
nor UO_1400 (O_1400,N_9491,N_9436);
nor UO_1401 (O_1401,N_9029,N_9685);
or UO_1402 (O_1402,N_9400,N_9890);
or UO_1403 (O_1403,N_9964,N_9382);
or UO_1404 (O_1404,N_9897,N_9610);
or UO_1405 (O_1405,N_9055,N_9355);
or UO_1406 (O_1406,N_9885,N_9431);
xnor UO_1407 (O_1407,N_9554,N_9387);
and UO_1408 (O_1408,N_9556,N_9170);
nand UO_1409 (O_1409,N_9175,N_9804);
and UO_1410 (O_1410,N_9805,N_9866);
and UO_1411 (O_1411,N_9236,N_9204);
xor UO_1412 (O_1412,N_9254,N_9354);
or UO_1413 (O_1413,N_9950,N_9461);
nand UO_1414 (O_1414,N_9975,N_9664);
xnor UO_1415 (O_1415,N_9292,N_9334);
or UO_1416 (O_1416,N_9970,N_9042);
nand UO_1417 (O_1417,N_9202,N_9784);
nand UO_1418 (O_1418,N_9167,N_9140);
and UO_1419 (O_1419,N_9348,N_9923);
and UO_1420 (O_1420,N_9608,N_9849);
nor UO_1421 (O_1421,N_9392,N_9996);
nor UO_1422 (O_1422,N_9282,N_9662);
and UO_1423 (O_1423,N_9727,N_9893);
nor UO_1424 (O_1424,N_9929,N_9475);
nand UO_1425 (O_1425,N_9346,N_9179);
and UO_1426 (O_1426,N_9076,N_9066);
nor UO_1427 (O_1427,N_9630,N_9719);
nor UO_1428 (O_1428,N_9904,N_9112);
or UO_1429 (O_1429,N_9604,N_9136);
or UO_1430 (O_1430,N_9547,N_9912);
and UO_1431 (O_1431,N_9545,N_9647);
nor UO_1432 (O_1432,N_9107,N_9654);
nand UO_1433 (O_1433,N_9846,N_9012);
nand UO_1434 (O_1434,N_9188,N_9630);
nor UO_1435 (O_1435,N_9333,N_9416);
nand UO_1436 (O_1436,N_9267,N_9482);
nor UO_1437 (O_1437,N_9142,N_9719);
or UO_1438 (O_1438,N_9313,N_9456);
and UO_1439 (O_1439,N_9442,N_9626);
nor UO_1440 (O_1440,N_9400,N_9758);
nor UO_1441 (O_1441,N_9485,N_9179);
nor UO_1442 (O_1442,N_9495,N_9505);
nand UO_1443 (O_1443,N_9935,N_9368);
nand UO_1444 (O_1444,N_9458,N_9613);
nand UO_1445 (O_1445,N_9232,N_9795);
nand UO_1446 (O_1446,N_9100,N_9586);
or UO_1447 (O_1447,N_9072,N_9884);
nand UO_1448 (O_1448,N_9911,N_9434);
nor UO_1449 (O_1449,N_9333,N_9019);
or UO_1450 (O_1450,N_9030,N_9231);
nor UO_1451 (O_1451,N_9191,N_9984);
nor UO_1452 (O_1452,N_9761,N_9533);
and UO_1453 (O_1453,N_9481,N_9620);
nor UO_1454 (O_1454,N_9851,N_9179);
or UO_1455 (O_1455,N_9328,N_9422);
and UO_1456 (O_1456,N_9277,N_9800);
nand UO_1457 (O_1457,N_9998,N_9255);
nand UO_1458 (O_1458,N_9155,N_9160);
or UO_1459 (O_1459,N_9922,N_9191);
and UO_1460 (O_1460,N_9555,N_9599);
and UO_1461 (O_1461,N_9435,N_9427);
or UO_1462 (O_1462,N_9469,N_9079);
nand UO_1463 (O_1463,N_9147,N_9888);
or UO_1464 (O_1464,N_9945,N_9515);
or UO_1465 (O_1465,N_9738,N_9151);
or UO_1466 (O_1466,N_9903,N_9149);
or UO_1467 (O_1467,N_9470,N_9073);
or UO_1468 (O_1468,N_9130,N_9411);
nor UO_1469 (O_1469,N_9493,N_9198);
or UO_1470 (O_1470,N_9651,N_9556);
nor UO_1471 (O_1471,N_9964,N_9607);
nor UO_1472 (O_1472,N_9434,N_9715);
nand UO_1473 (O_1473,N_9897,N_9676);
and UO_1474 (O_1474,N_9180,N_9797);
or UO_1475 (O_1475,N_9174,N_9430);
and UO_1476 (O_1476,N_9192,N_9613);
nand UO_1477 (O_1477,N_9547,N_9874);
and UO_1478 (O_1478,N_9151,N_9097);
and UO_1479 (O_1479,N_9501,N_9608);
and UO_1480 (O_1480,N_9372,N_9911);
or UO_1481 (O_1481,N_9128,N_9623);
xnor UO_1482 (O_1482,N_9463,N_9103);
nand UO_1483 (O_1483,N_9014,N_9623);
nor UO_1484 (O_1484,N_9038,N_9420);
or UO_1485 (O_1485,N_9294,N_9104);
and UO_1486 (O_1486,N_9930,N_9088);
and UO_1487 (O_1487,N_9735,N_9659);
nand UO_1488 (O_1488,N_9554,N_9463);
and UO_1489 (O_1489,N_9193,N_9650);
nor UO_1490 (O_1490,N_9146,N_9816);
nor UO_1491 (O_1491,N_9375,N_9491);
nor UO_1492 (O_1492,N_9872,N_9100);
and UO_1493 (O_1493,N_9098,N_9373);
nor UO_1494 (O_1494,N_9628,N_9805);
nor UO_1495 (O_1495,N_9285,N_9052);
and UO_1496 (O_1496,N_9284,N_9865);
nor UO_1497 (O_1497,N_9972,N_9212);
nand UO_1498 (O_1498,N_9296,N_9817);
and UO_1499 (O_1499,N_9933,N_9214);
endmodule