module basic_500_3000_500_3_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_248,In_168);
or U1 (N_1,In_266,In_27);
and U2 (N_2,In_123,In_471);
nand U3 (N_3,In_86,In_399);
nor U4 (N_4,In_146,In_137);
nor U5 (N_5,In_259,In_379);
nand U6 (N_6,In_384,In_331);
nand U7 (N_7,In_439,In_374);
or U8 (N_8,In_285,In_268);
nand U9 (N_9,In_148,In_232);
nor U10 (N_10,In_30,In_192);
and U11 (N_11,In_116,In_205);
or U12 (N_12,In_250,In_244);
or U13 (N_13,In_185,In_241);
or U14 (N_14,In_286,In_154);
nor U15 (N_15,In_180,In_108);
nand U16 (N_16,In_56,In_187);
nor U17 (N_17,In_103,In_219);
and U18 (N_18,In_173,In_448);
nor U19 (N_19,In_59,In_310);
nor U20 (N_20,In_412,In_63);
nand U21 (N_21,In_386,In_243);
nand U22 (N_22,In_179,In_363);
nand U23 (N_23,In_453,In_409);
nor U24 (N_24,In_304,In_438);
and U25 (N_25,In_70,In_92);
and U26 (N_26,In_306,In_383);
and U27 (N_27,In_80,In_258);
nor U28 (N_28,In_196,In_329);
nor U29 (N_29,In_493,In_323);
nor U30 (N_30,In_177,In_368);
and U31 (N_31,In_396,In_12);
and U32 (N_32,In_54,In_475);
or U33 (N_33,In_72,In_201);
or U34 (N_34,In_25,In_382);
or U35 (N_35,In_182,In_288);
and U36 (N_36,In_98,In_89);
or U37 (N_37,In_58,In_37);
and U38 (N_38,In_94,In_195);
or U39 (N_39,In_193,In_169);
nor U40 (N_40,In_407,In_324);
and U41 (N_41,In_320,In_121);
or U42 (N_42,In_176,In_361);
and U43 (N_43,In_473,In_351);
nand U44 (N_44,In_356,In_111);
nand U45 (N_45,In_47,In_492);
or U46 (N_46,In_208,In_230);
and U47 (N_47,In_334,In_155);
nand U48 (N_48,In_341,In_387);
nor U49 (N_49,In_408,In_314);
or U50 (N_50,In_450,In_283);
and U51 (N_51,In_255,In_378);
or U52 (N_52,In_494,In_353);
or U53 (N_53,In_367,In_274);
and U54 (N_54,In_434,In_484);
or U55 (N_55,In_117,In_23);
or U56 (N_56,In_488,In_242);
and U57 (N_57,In_444,In_313);
or U58 (N_58,In_60,In_11);
and U59 (N_59,In_470,In_252);
nand U60 (N_60,In_78,In_385);
nand U61 (N_61,In_156,In_391);
or U62 (N_62,In_370,In_401);
nand U63 (N_63,In_17,In_495);
and U64 (N_64,In_433,In_332);
nand U65 (N_65,In_104,In_490);
nand U66 (N_66,In_45,In_393);
nor U67 (N_67,In_263,In_298);
and U68 (N_68,In_411,In_191);
nand U69 (N_69,In_429,In_218);
or U70 (N_70,In_337,In_499);
nand U71 (N_71,In_50,In_315);
nand U72 (N_72,In_120,In_199);
and U73 (N_73,In_394,In_97);
xnor U74 (N_74,In_464,In_7);
nor U75 (N_75,In_321,In_481);
nor U76 (N_76,In_2,In_280);
xor U77 (N_77,In_90,In_152);
or U78 (N_78,In_64,In_57);
xnor U79 (N_79,In_40,In_22);
nor U80 (N_80,In_373,In_46);
or U81 (N_81,In_364,In_486);
nor U82 (N_82,In_144,In_333);
nand U83 (N_83,In_188,In_247);
and U84 (N_84,In_294,In_153);
and U85 (N_85,In_85,In_431);
nor U86 (N_86,In_222,In_100);
and U87 (N_87,In_372,In_139);
or U88 (N_88,In_61,In_442);
nand U89 (N_89,In_102,In_451);
and U90 (N_90,In_99,In_212);
nor U91 (N_91,In_319,In_261);
nor U92 (N_92,In_480,In_307);
nor U93 (N_93,In_260,In_145);
and U94 (N_94,In_34,In_295);
nor U95 (N_95,In_308,In_41);
or U96 (N_96,In_140,In_389);
or U97 (N_97,In_381,In_462);
and U98 (N_98,In_81,In_149);
and U99 (N_99,In_126,In_71);
or U100 (N_100,In_106,In_210);
or U101 (N_101,In_238,In_457);
and U102 (N_102,In_265,In_269);
nor U103 (N_103,In_427,In_198);
nand U104 (N_104,In_234,In_466);
nor U105 (N_105,In_416,In_69);
nand U106 (N_106,In_456,In_335);
and U107 (N_107,In_380,In_282);
and U108 (N_108,In_419,In_18);
or U109 (N_109,In_175,In_327);
nand U110 (N_110,In_115,In_33);
or U111 (N_111,In_352,In_209);
or U112 (N_112,In_421,In_297);
nor U113 (N_113,In_91,In_236);
or U114 (N_114,In_340,In_114);
or U115 (N_115,In_62,In_132);
and U116 (N_116,In_240,In_231);
or U117 (N_117,In_4,In_472);
or U118 (N_118,In_21,In_432);
and U119 (N_119,In_204,In_299);
or U120 (N_120,In_257,In_5);
and U121 (N_121,In_423,In_425);
nand U122 (N_122,In_157,In_77);
and U123 (N_123,In_485,In_38);
or U124 (N_124,In_73,In_461);
nor U125 (N_125,In_312,In_66);
and U126 (N_126,In_403,In_253);
or U127 (N_127,In_42,In_53);
nor U128 (N_128,In_211,In_107);
or U129 (N_129,In_362,In_184);
nor U130 (N_130,In_36,In_402);
xor U131 (N_131,In_122,In_227);
nand U132 (N_132,In_213,In_96);
nor U133 (N_133,In_405,In_328);
nor U134 (N_134,In_326,In_13);
nand U135 (N_135,In_482,In_136);
or U136 (N_136,In_440,In_371);
or U137 (N_137,In_161,In_68);
or U138 (N_138,In_221,In_330);
nand U139 (N_139,In_437,In_489);
and U140 (N_140,In_455,In_93);
or U141 (N_141,In_134,In_51);
xor U142 (N_142,In_460,In_118);
and U143 (N_143,In_147,In_127);
nand U144 (N_144,In_343,In_14);
or U145 (N_145,In_84,In_430);
nand U146 (N_146,In_477,In_366);
and U147 (N_147,In_181,In_246);
nor U148 (N_148,In_200,In_296);
or U149 (N_149,In_26,In_67);
nand U150 (N_150,In_422,In_135);
nand U151 (N_151,In_491,In_281);
and U152 (N_152,In_101,In_113);
and U153 (N_153,In_158,In_262);
nand U154 (N_154,In_251,In_487);
and U155 (N_155,In_224,In_16);
or U156 (N_156,In_48,In_357);
and U157 (N_157,In_325,In_170);
or U158 (N_158,In_76,In_128);
or U159 (N_159,In_390,In_150);
nand U160 (N_160,In_428,In_95);
nand U161 (N_161,In_354,In_28);
nand U162 (N_162,In_317,In_498);
or U163 (N_163,In_239,In_349);
and U164 (N_164,In_8,In_254);
or U165 (N_165,In_459,In_83);
nor U166 (N_166,In_74,In_141);
nor U167 (N_167,In_31,In_418);
or U168 (N_168,In_88,In_468);
and U169 (N_169,In_377,In_164);
nor U170 (N_170,In_9,In_483);
nor U171 (N_171,In_465,In_369);
or U172 (N_172,In_226,In_476);
nor U173 (N_173,In_216,In_497);
and U174 (N_174,In_479,In_225);
and U175 (N_175,In_206,In_395);
or U176 (N_176,In_131,In_342);
nand U177 (N_177,In_124,In_138);
or U178 (N_178,In_130,In_375);
nand U179 (N_179,In_183,In_49);
nand U180 (N_180,In_223,In_249);
or U181 (N_181,In_435,In_10);
and U182 (N_182,In_309,In_229);
or U183 (N_183,In_233,In_458);
nand U184 (N_184,In_336,In_478);
nor U185 (N_185,In_119,In_398);
nand U186 (N_186,In_267,In_197);
nor U187 (N_187,In_365,In_322);
or U188 (N_188,In_125,In_275);
nor U189 (N_189,In_186,In_469);
and U190 (N_190,In_443,In_463);
and U191 (N_191,In_346,In_348);
or U192 (N_192,In_43,In_347);
nand U193 (N_193,In_190,In_358);
and U194 (N_194,In_279,In_467);
and U195 (N_195,In_142,In_24);
nand U196 (N_196,In_291,In_165);
nand U197 (N_197,In_109,In_178);
and U198 (N_198,In_276,In_32);
nor U199 (N_199,In_441,In_163);
nand U200 (N_200,In_110,In_446);
nand U201 (N_201,In_65,In_151);
and U202 (N_202,In_167,In_454);
or U203 (N_203,In_290,In_406);
nand U204 (N_204,In_75,In_447);
nand U205 (N_205,In_355,In_194);
or U206 (N_206,In_245,In_162);
or U207 (N_207,In_0,In_289);
and U208 (N_208,In_174,In_452);
and U209 (N_209,In_293,In_278);
or U210 (N_210,In_413,In_360);
nor U211 (N_211,In_424,In_20);
nor U212 (N_212,In_284,In_376);
or U213 (N_213,In_305,In_207);
and U214 (N_214,In_270,In_6);
and U215 (N_215,In_129,In_303);
and U216 (N_216,In_39,In_79);
nand U217 (N_217,In_417,In_35);
nor U218 (N_218,In_414,In_44);
or U219 (N_219,In_228,In_400);
nor U220 (N_220,In_474,In_301);
or U221 (N_221,In_133,In_449);
or U222 (N_222,In_311,In_189);
or U223 (N_223,In_237,In_235);
or U224 (N_224,In_445,In_1);
nor U225 (N_225,In_292,In_277);
or U226 (N_226,In_171,In_159);
nor U227 (N_227,In_82,In_496);
nand U228 (N_228,In_436,In_215);
or U229 (N_229,In_359,In_338);
or U230 (N_230,In_426,In_410);
nor U231 (N_231,In_316,In_160);
nor U232 (N_232,In_392,In_29);
nor U233 (N_233,In_339,In_143);
or U234 (N_234,In_272,In_273);
and U235 (N_235,In_3,In_397);
nand U236 (N_236,In_344,In_388);
and U237 (N_237,In_264,In_15);
nor U238 (N_238,In_420,In_172);
nand U239 (N_239,In_300,In_214);
nand U240 (N_240,In_203,In_166);
and U241 (N_241,In_55,In_52);
nand U242 (N_242,In_105,In_19);
and U243 (N_243,In_256,In_302);
and U244 (N_244,In_415,In_217);
nor U245 (N_245,In_220,In_404);
or U246 (N_246,In_87,In_350);
and U247 (N_247,In_202,In_112);
nand U248 (N_248,In_318,In_271);
nor U249 (N_249,In_287,In_345);
or U250 (N_250,In_277,In_377);
and U251 (N_251,In_63,In_369);
or U252 (N_252,In_220,In_19);
or U253 (N_253,In_21,In_339);
and U254 (N_254,In_236,In_51);
nor U255 (N_255,In_303,In_176);
nor U256 (N_256,In_3,In_465);
nor U257 (N_257,In_166,In_391);
or U258 (N_258,In_287,In_84);
nor U259 (N_259,In_298,In_82);
or U260 (N_260,In_291,In_339);
nor U261 (N_261,In_211,In_167);
and U262 (N_262,In_347,In_453);
nand U263 (N_263,In_256,In_31);
or U264 (N_264,In_334,In_498);
nand U265 (N_265,In_267,In_70);
nor U266 (N_266,In_246,In_144);
nor U267 (N_267,In_465,In_481);
nand U268 (N_268,In_226,In_327);
nor U269 (N_269,In_266,In_179);
nor U270 (N_270,In_4,In_53);
nor U271 (N_271,In_177,In_495);
and U272 (N_272,In_72,In_155);
and U273 (N_273,In_338,In_200);
and U274 (N_274,In_73,In_25);
nand U275 (N_275,In_235,In_184);
and U276 (N_276,In_145,In_34);
and U277 (N_277,In_137,In_11);
nand U278 (N_278,In_244,In_271);
nand U279 (N_279,In_437,In_163);
and U280 (N_280,In_349,In_486);
nand U281 (N_281,In_267,In_440);
nand U282 (N_282,In_288,In_321);
and U283 (N_283,In_195,In_248);
nand U284 (N_284,In_156,In_196);
nand U285 (N_285,In_137,In_66);
nand U286 (N_286,In_242,In_470);
and U287 (N_287,In_474,In_235);
and U288 (N_288,In_353,In_198);
or U289 (N_289,In_61,In_290);
and U290 (N_290,In_380,In_430);
nor U291 (N_291,In_482,In_432);
nand U292 (N_292,In_496,In_438);
nand U293 (N_293,In_73,In_112);
or U294 (N_294,In_372,In_484);
nor U295 (N_295,In_24,In_418);
and U296 (N_296,In_48,In_136);
nand U297 (N_297,In_462,In_32);
nand U298 (N_298,In_318,In_230);
nor U299 (N_299,In_171,In_365);
nand U300 (N_300,In_380,In_162);
nand U301 (N_301,In_17,In_289);
nor U302 (N_302,In_498,In_314);
nor U303 (N_303,In_405,In_91);
and U304 (N_304,In_136,In_3);
nand U305 (N_305,In_263,In_59);
nand U306 (N_306,In_427,In_325);
or U307 (N_307,In_494,In_294);
nor U308 (N_308,In_165,In_109);
nand U309 (N_309,In_463,In_417);
and U310 (N_310,In_43,In_298);
and U311 (N_311,In_464,In_203);
or U312 (N_312,In_202,In_243);
and U313 (N_313,In_217,In_177);
nor U314 (N_314,In_434,In_52);
or U315 (N_315,In_459,In_60);
or U316 (N_316,In_213,In_442);
or U317 (N_317,In_244,In_448);
and U318 (N_318,In_274,In_181);
and U319 (N_319,In_432,In_202);
nand U320 (N_320,In_209,In_325);
nand U321 (N_321,In_162,In_392);
or U322 (N_322,In_270,In_79);
nand U323 (N_323,In_177,In_122);
nor U324 (N_324,In_223,In_202);
nor U325 (N_325,In_288,In_89);
or U326 (N_326,In_477,In_480);
and U327 (N_327,In_41,In_61);
nand U328 (N_328,In_91,In_473);
or U329 (N_329,In_187,In_2);
nor U330 (N_330,In_86,In_413);
nand U331 (N_331,In_16,In_42);
or U332 (N_332,In_247,In_57);
and U333 (N_333,In_28,In_25);
nor U334 (N_334,In_189,In_2);
nand U335 (N_335,In_315,In_256);
nand U336 (N_336,In_27,In_107);
nor U337 (N_337,In_194,In_7);
nand U338 (N_338,In_224,In_407);
or U339 (N_339,In_295,In_30);
nor U340 (N_340,In_240,In_213);
nand U341 (N_341,In_244,In_451);
and U342 (N_342,In_23,In_375);
nand U343 (N_343,In_475,In_327);
and U344 (N_344,In_147,In_159);
nand U345 (N_345,In_440,In_467);
nand U346 (N_346,In_409,In_139);
and U347 (N_347,In_455,In_177);
or U348 (N_348,In_363,In_215);
nor U349 (N_349,In_306,In_489);
and U350 (N_350,In_388,In_19);
or U351 (N_351,In_233,In_285);
nand U352 (N_352,In_336,In_484);
or U353 (N_353,In_224,In_173);
and U354 (N_354,In_117,In_445);
and U355 (N_355,In_98,In_305);
nor U356 (N_356,In_299,In_366);
nor U357 (N_357,In_464,In_465);
nand U358 (N_358,In_350,In_366);
nand U359 (N_359,In_192,In_359);
nor U360 (N_360,In_91,In_29);
and U361 (N_361,In_468,In_127);
and U362 (N_362,In_115,In_383);
nor U363 (N_363,In_175,In_18);
and U364 (N_364,In_43,In_110);
nor U365 (N_365,In_65,In_230);
nor U366 (N_366,In_160,In_91);
nand U367 (N_367,In_430,In_485);
nand U368 (N_368,In_130,In_66);
and U369 (N_369,In_364,In_35);
and U370 (N_370,In_28,In_214);
nand U371 (N_371,In_220,In_371);
nor U372 (N_372,In_140,In_136);
or U373 (N_373,In_486,In_78);
nor U374 (N_374,In_85,In_139);
and U375 (N_375,In_458,In_170);
or U376 (N_376,In_434,In_364);
nand U377 (N_377,In_312,In_34);
and U378 (N_378,In_334,In_302);
nand U379 (N_379,In_489,In_107);
and U380 (N_380,In_1,In_43);
or U381 (N_381,In_161,In_409);
nand U382 (N_382,In_329,In_90);
nor U383 (N_383,In_348,In_402);
and U384 (N_384,In_305,In_9);
nand U385 (N_385,In_51,In_250);
and U386 (N_386,In_340,In_315);
nor U387 (N_387,In_244,In_337);
and U388 (N_388,In_328,In_240);
or U389 (N_389,In_456,In_460);
nor U390 (N_390,In_259,In_171);
nand U391 (N_391,In_82,In_99);
nor U392 (N_392,In_241,In_14);
nand U393 (N_393,In_66,In_176);
nor U394 (N_394,In_355,In_141);
and U395 (N_395,In_189,In_52);
or U396 (N_396,In_146,In_474);
nor U397 (N_397,In_457,In_432);
nor U398 (N_398,In_484,In_62);
nand U399 (N_399,In_401,In_95);
nor U400 (N_400,In_289,In_164);
or U401 (N_401,In_281,In_419);
nor U402 (N_402,In_285,In_274);
or U403 (N_403,In_461,In_243);
or U404 (N_404,In_256,In_260);
nand U405 (N_405,In_76,In_155);
or U406 (N_406,In_337,In_59);
and U407 (N_407,In_107,In_323);
and U408 (N_408,In_460,In_161);
nand U409 (N_409,In_211,In_135);
nor U410 (N_410,In_132,In_50);
or U411 (N_411,In_128,In_445);
nor U412 (N_412,In_481,In_446);
nand U413 (N_413,In_312,In_230);
nor U414 (N_414,In_297,In_88);
or U415 (N_415,In_429,In_411);
nand U416 (N_416,In_325,In_430);
nand U417 (N_417,In_14,In_335);
or U418 (N_418,In_448,In_344);
nor U419 (N_419,In_443,In_363);
nor U420 (N_420,In_359,In_90);
and U421 (N_421,In_361,In_465);
nand U422 (N_422,In_397,In_317);
nand U423 (N_423,In_283,In_294);
or U424 (N_424,In_444,In_364);
nor U425 (N_425,In_275,In_269);
and U426 (N_426,In_300,In_95);
and U427 (N_427,In_297,In_407);
and U428 (N_428,In_400,In_405);
and U429 (N_429,In_336,In_446);
or U430 (N_430,In_250,In_46);
and U431 (N_431,In_379,In_123);
nand U432 (N_432,In_149,In_113);
nand U433 (N_433,In_342,In_192);
or U434 (N_434,In_156,In_261);
and U435 (N_435,In_260,In_25);
nor U436 (N_436,In_429,In_224);
nand U437 (N_437,In_281,In_250);
and U438 (N_438,In_349,In_278);
or U439 (N_439,In_142,In_446);
and U440 (N_440,In_342,In_132);
nand U441 (N_441,In_328,In_222);
or U442 (N_442,In_70,In_193);
nor U443 (N_443,In_257,In_434);
and U444 (N_444,In_214,In_347);
nor U445 (N_445,In_134,In_155);
nand U446 (N_446,In_249,In_99);
and U447 (N_447,In_57,In_185);
or U448 (N_448,In_400,In_248);
nor U449 (N_449,In_200,In_463);
nand U450 (N_450,In_487,In_285);
and U451 (N_451,In_305,In_343);
or U452 (N_452,In_43,In_3);
and U453 (N_453,In_28,In_179);
and U454 (N_454,In_486,In_384);
and U455 (N_455,In_364,In_220);
or U456 (N_456,In_104,In_133);
nand U457 (N_457,In_332,In_440);
nand U458 (N_458,In_82,In_272);
or U459 (N_459,In_15,In_294);
or U460 (N_460,In_292,In_30);
nand U461 (N_461,In_69,In_54);
nor U462 (N_462,In_497,In_137);
nand U463 (N_463,In_21,In_269);
or U464 (N_464,In_259,In_34);
nand U465 (N_465,In_236,In_24);
or U466 (N_466,In_187,In_336);
or U467 (N_467,In_333,In_49);
and U468 (N_468,In_387,In_216);
or U469 (N_469,In_271,In_442);
nand U470 (N_470,In_14,In_320);
and U471 (N_471,In_309,In_126);
nand U472 (N_472,In_117,In_492);
nor U473 (N_473,In_419,In_247);
or U474 (N_474,In_407,In_290);
or U475 (N_475,In_385,In_305);
or U476 (N_476,In_94,In_72);
nand U477 (N_477,In_142,In_6);
nor U478 (N_478,In_97,In_35);
nor U479 (N_479,In_488,In_134);
and U480 (N_480,In_450,In_40);
nor U481 (N_481,In_378,In_381);
or U482 (N_482,In_300,In_5);
xor U483 (N_483,In_135,In_188);
nor U484 (N_484,In_366,In_68);
or U485 (N_485,In_401,In_478);
nor U486 (N_486,In_461,In_29);
and U487 (N_487,In_153,In_394);
nor U488 (N_488,In_8,In_54);
nor U489 (N_489,In_226,In_1);
nand U490 (N_490,In_251,In_268);
nor U491 (N_491,In_287,In_237);
nand U492 (N_492,In_399,In_295);
nor U493 (N_493,In_77,In_74);
nor U494 (N_494,In_174,In_127);
nand U495 (N_495,In_424,In_82);
and U496 (N_496,In_469,In_136);
nor U497 (N_497,In_16,In_32);
nand U498 (N_498,In_482,In_224);
or U499 (N_499,In_24,In_323);
or U500 (N_500,In_207,In_280);
nor U501 (N_501,In_419,In_439);
and U502 (N_502,In_352,In_388);
or U503 (N_503,In_125,In_94);
and U504 (N_504,In_266,In_74);
or U505 (N_505,In_438,In_156);
or U506 (N_506,In_18,In_136);
or U507 (N_507,In_149,In_32);
nand U508 (N_508,In_292,In_354);
nor U509 (N_509,In_190,In_472);
nor U510 (N_510,In_198,In_212);
or U511 (N_511,In_85,In_167);
nor U512 (N_512,In_20,In_217);
or U513 (N_513,In_423,In_492);
nor U514 (N_514,In_157,In_261);
nor U515 (N_515,In_347,In_54);
and U516 (N_516,In_97,In_371);
or U517 (N_517,In_405,In_441);
or U518 (N_518,In_414,In_161);
and U519 (N_519,In_23,In_255);
nand U520 (N_520,In_220,In_190);
and U521 (N_521,In_143,In_293);
nand U522 (N_522,In_17,In_211);
or U523 (N_523,In_65,In_456);
or U524 (N_524,In_191,In_97);
nor U525 (N_525,In_360,In_39);
or U526 (N_526,In_35,In_285);
or U527 (N_527,In_355,In_39);
xor U528 (N_528,In_50,In_332);
or U529 (N_529,In_356,In_350);
and U530 (N_530,In_172,In_82);
nor U531 (N_531,In_327,In_290);
nor U532 (N_532,In_339,In_222);
nand U533 (N_533,In_321,In_198);
and U534 (N_534,In_55,In_216);
nor U535 (N_535,In_28,In_111);
or U536 (N_536,In_78,In_276);
nand U537 (N_537,In_329,In_239);
nand U538 (N_538,In_48,In_460);
nand U539 (N_539,In_107,In_366);
nand U540 (N_540,In_264,In_458);
nor U541 (N_541,In_430,In_159);
xor U542 (N_542,In_413,In_316);
and U543 (N_543,In_361,In_486);
and U544 (N_544,In_391,In_14);
and U545 (N_545,In_474,In_350);
and U546 (N_546,In_11,In_400);
and U547 (N_547,In_283,In_50);
nand U548 (N_548,In_462,In_391);
nor U549 (N_549,In_62,In_194);
or U550 (N_550,In_135,In_95);
nor U551 (N_551,In_186,In_55);
and U552 (N_552,In_344,In_439);
or U553 (N_553,In_296,In_26);
nand U554 (N_554,In_376,In_325);
nand U555 (N_555,In_223,In_423);
xor U556 (N_556,In_31,In_144);
nor U557 (N_557,In_409,In_47);
or U558 (N_558,In_89,In_353);
nand U559 (N_559,In_262,In_133);
nand U560 (N_560,In_69,In_315);
nor U561 (N_561,In_173,In_260);
or U562 (N_562,In_187,In_307);
nand U563 (N_563,In_211,In_312);
nor U564 (N_564,In_206,In_122);
or U565 (N_565,In_13,In_454);
nand U566 (N_566,In_75,In_421);
nand U567 (N_567,In_267,In_277);
or U568 (N_568,In_10,In_451);
and U569 (N_569,In_191,In_93);
nor U570 (N_570,In_36,In_417);
nor U571 (N_571,In_394,In_495);
nor U572 (N_572,In_436,In_155);
nand U573 (N_573,In_152,In_417);
or U574 (N_574,In_427,In_4);
and U575 (N_575,In_249,In_422);
or U576 (N_576,In_44,In_28);
nand U577 (N_577,In_64,In_12);
nor U578 (N_578,In_332,In_10);
nor U579 (N_579,In_75,In_80);
nand U580 (N_580,In_153,In_327);
and U581 (N_581,In_414,In_78);
or U582 (N_582,In_448,In_289);
and U583 (N_583,In_144,In_251);
nor U584 (N_584,In_450,In_211);
nor U585 (N_585,In_338,In_37);
nand U586 (N_586,In_28,In_99);
nor U587 (N_587,In_52,In_19);
nand U588 (N_588,In_169,In_441);
nand U589 (N_589,In_409,In_231);
or U590 (N_590,In_418,In_303);
and U591 (N_591,In_291,In_231);
nor U592 (N_592,In_284,In_382);
and U593 (N_593,In_263,In_287);
nor U594 (N_594,In_332,In_496);
or U595 (N_595,In_351,In_42);
or U596 (N_596,In_153,In_112);
or U597 (N_597,In_9,In_311);
and U598 (N_598,In_383,In_177);
or U599 (N_599,In_127,In_239);
or U600 (N_600,In_399,In_284);
nor U601 (N_601,In_107,In_122);
or U602 (N_602,In_288,In_311);
nand U603 (N_603,In_30,In_103);
or U604 (N_604,In_122,In_244);
nand U605 (N_605,In_209,In_147);
nor U606 (N_606,In_250,In_165);
nor U607 (N_607,In_36,In_388);
or U608 (N_608,In_122,In_33);
and U609 (N_609,In_193,In_141);
or U610 (N_610,In_401,In_448);
or U611 (N_611,In_96,In_145);
xor U612 (N_612,In_173,In_455);
or U613 (N_613,In_3,In_429);
and U614 (N_614,In_127,In_335);
nor U615 (N_615,In_201,In_427);
or U616 (N_616,In_346,In_304);
nor U617 (N_617,In_418,In_389);
nand U618 (N_618,In_72,In_37);
or U619 (N_619,In_54,In_185);
or U620 (N_620,In_436,In_492);
nand U621 (N_621,In_397,In_207);
nand U622 (N_622,In_413,In_479);
nand U623 (N_623,In_177,In_373);
or U624 (N_624,In_467,In_282);
nor U625 (N_625,In_408,In_147);
nor U626 (N_626,In_223,In_209);
nand U627 (N_627,In_107,In_236);
nor U628 (N_628,In_310,In_277);
or U629 (N_629,In_179,In_191);
or U630 (N_630,In_38,In_454);
nor U631 (N_631,In_297,In_35);
nand U632 (N_632,In_21,In_97);
or U633 (N_633,In_108,In_203);
nand U634 (N_634,In_316,In_474);
nor U635 (N_635,In_22,In_170);
nor U636 (N_636,In_210,In_250);
xnor U637 (N_637,In_392,In_121);
nand U638 (N_638,In_367,In_187);
nand U639 (N_639,In_61,In_230);
or U640 (N_640,In_21,In_160);
nand U641 (N_641,In_443,In_465);
or U642 (N_642,In_346,In_340);
and U643 (N_643,In_416,In_165);
and U644 (N_644,In_337,In_287);
and U645 (N_645,In_328,In_298);
nand U646 (N_646,In_118,In_400);
nand U647 (N_647,In_314,In_167);
nor U648 (N_648,In_144,In_319);
or U649 (N_649,In_10,In_313);
and U650 (N_650,In_151,In_387);
nand U651 (N_651,In_283,In_218);
nor U652 (N_652,In_19,In_403);
nor U653 (N_653,In_462,In_147);
and U654 (N_654,In_369,In_306);
nand U655 (N_655,In_76,In_15);
or U656 (N_656,In_173,In_387);
and U657 (N_657,In_346,In_222);
nand U658 (N_658,In_255,In_367);
or U659 (N_659,In_52,In_253);
nor U660 (N_660,In_306,In_441);
nand U661 (N_661,In_405,In_316);
or U662 (N_662,In_381,In_238);
or U663 (N_663,In_119,In_331);
and U664 (N_664,In_171,In_160);
and U665 (N_665,In_450,In_75);
and U666 (N_666,In_434,In_466);
and U667 (N_667,In_322,In_128);
nor U668 (N_668,In_366,In_99);
nor U669 (N_669,In_383,In_358);
nor U670 (N_670,In_432,In_12);
nand U671 (N_671,In_125,In_232);
nor U672 (N_672,In_2,In_9);
xor U673 (N_673,In_131,In_130);
nand U674 (N_674,In_270,In_68);
or U675 (N_675,In_352,In_476);
and U676 (N_676,In_205,In_16);
nand U677 (N_677,In_386,In_61);
or U678 (N_678,In_138,In_50);
nand U679 (N_679,In_419,In_223);
or U680 (N_680,In_392,In_12);
and U681 (N_681,In_53,In_466);
and U682 (N_682,In_345,In_397);
and U683 (N_683,In_189,In_177);
and U684 (N_684,In_394,In_404);
nand U685 (N_685,In_384,In_402);
nand U686 (N_686,In_489,In_436);
and U687 (N_687,In_483,In_211);
and U688 (N_688,In_23,In_185);
or U689 (N_689,In_398,In_409);
and U690 (N_690,In_239,In_457);
nand U691 (N_691,In_87,In_489);
xor U692 (N_692,In_183,In_331);
nor U693 (N_693,In_47,In_267);
and U694 (N_694,In_499,In_200);
nor U695 (N_695,In_333,In_160);
and U696 (N_696,In_26,In_131);
or U697 (N_697,In_326,In_146);
nand U698 (N_698,In_32,In_441);
nand U699 (N_699,In_200,In_495);
nor U700 (N_700,In_438,In_272);
nor U701 (N_701,In_483,In_316);
nor U702 (N_702,In_12,In_354);
or U703 (N_703,In_179,In_364);
or U704 (N_704,In_123,In_425);
nand U705 (N_705,In_485,In_138);
or U706 (N_706,In_165,In_185);
and U707 (N_707,In_398,In_469);
and U708 (N_708,In_31,In_331);
nand U709 (N_709,In_335,In_298);
nand U710 (N_710,In_165,In_401);
nor U711 (N_711,In_440,In_233);
nor U712 (N_712,In_487,In_413);
nor U713 (N_713,In_457,In_289);
nor U714 (N_714,In_173,In_336);
and U715 (N_715,In_486,In_248);
or U716 (N_716,In_423,In_433);
nor U717 (N_717,In_331,In_453);
nand U718 (N_718,In_412,In_242);
or U719 (N_719,In_285,In_21);
or U720 (N_720,In_325,In_190);
nor U721 (N_721,In_453,In_44);
nand U722 (N_722,In_459,In_40);
nor U723 (N_723,In_436,In_62);
or U724 (N_724,In_166,In_482);
or U725 (N_725,In_380,In_406);
and U726 (N_726,In_78,In_165);
nand U727 (N_727,In_484,In_496);
and U728 (N_728,In_139,In_72);
or U729 (N_729,In_90,In_164);
nor U730 (N_730,In_465,In_69);
or U731 (N_731,In_391,In_275);
nand U732 (N_732,In_427,In_484);
and U733 (N_733,In_144,In_284);
nor U734 (N_734,In_180,In_26);
nor U735 (N_735,In_374,In_141);
or U736 (N_736,In_110,In_95);
or U737 (N_737,In_468,In_443);
and U738 (N_738,In_242,In_385);
nor U739 (N_739,In_30,In_16);
or U740 (N_740,In_476,In_105);
nand U741 (N_741,In_201,In_460);
nor U742 (N_742,In_150,In_39);
nand U743 (N_743,In_394,In_238);
nand U744 (N_744,In_182,In_29);
and U745 (N_745,In_92,In_102);
nor U746 (N_746,In_227,In_471);
nor U747 (N_747,In_21,In_221);
nor U748 (N_748,In_65,In_192);
nand U749 (N_749,In_134,In_97);
or U750 (N_750,In_327,In_53);
or U751 (N_751,In_123,In_336);
nand U752 (N_752,In_92,In_300);
nor U753 (N_753,In_283,In_421);
and U754 (N_754,In_224,In_324);
and U755 (N_755,In_404,In_388);
or U756 (N_756,In_46,In_427);
nor U757 (N_757,In_89,In_425);
nor U758 (N_758,In_270,In_209);
nand U759 (N_759,In_170,In_107);
nor U760 (N_760,In_470,In_342);
or U761 (N_761,In_436,In_238);
nand U762 (N_762,In_353,In_150);
nand U763 (N_763,In_86,In_411);
nor U764 (N_764,In_0,In_195);
nor U765 (N_765,In_89,In_464);
nor U766 (N_766,In_49,In_186);
or U767 (N_767,In_11,In_74);
or U768 (N_768,In_7,In_16);
or U769 (N_769,In_446,In_343);
nor U770 (N_770,In_127,In_111);
or U771 (N_771,In_256,In_190);
nor U772 (N_772,In_390,In_295);
and U773 (N_773,In_237,In_391);
or U774 (N_774,In_23,In_429);
and U775 (N_775,In_300,In_369);
nor U776 (N_776,In_165,In_280);
nor U777 (N_777,In_384,In_153);
nand U778 (N_778,In_129,In_261);
nand U779 (N_779,In_275,In_19);
or U780 (N_780,In_449,In_299);
nor U781 (N_781,In_123,In_136);
nand U782 (N_782,In_408,In_489);
or U783 (N_783,In_403,In_343);
xor U784 (N_784,In_209,In_220);
nand U785 (N_785,In_323,In_378);
nor U786 (N_786,In_249,In_381);
nor U787 (N_787,In_294,In_393);
and U788 (N_788,In_245,In_413);
nand U789 (N_789,In_289,In_187);
or U790 (N_790,In_227,In_242);
nand U791 (N_791,In_268,In_300);
nor U792 (N_792,In_141,In_197);
and U793 (N_793,In_210,In_490);
or U794 (N_794,In_282,In_216);
and U795 (N_795,In_208,In_296);
or U796 (N_796,In_354,In_339);
nand U797 (N_797,In_267,In_332);
and U798 (N_798,In_158,In_122);
nand U799 (N_799,In_480,In_184);
or U800 (N_800,In_445,In_451);
and U801 (N_801,In_214,In_186);
nand U802 (N_802,In_352,In_248);
nand U803 (N_803,In_303,In_37);
or U804 (N_804,In_425,In_166);
or U805 (N_805,In_453,In_374);
nand U806 (N_806,In_435,In_319);
nor U807 (N_807,In_337,In_336);
or U808 (N_808,In_302,In_339);
nor U809 (N_809,In_127,In_71);
nand U810 (N_810,In_44,In_322);
xnor U811 (N_811,In_149,In_219);
nor U812 (N_812,In_121,In_423);
and U813 (N_813,In_449,In_218);
nand U814 (N_814,In_173,In_14);
and U815 (N_815,In_334,In_45);
nor U816 (N_816,In_319,In_458);
and U817 (N_817,In_343,In_436);
nor U818 (N_818,In_266,In_147);
and U819 (N_819,In_267,In_45);
and U820 (N_820,In_172,In_16);
and U821 (N_821,In_102,In_473);
and U822 (N_822,In_11,In_230);
or U823 (N_823,In_129,In_60);
or U824 (N_824,In_342,In_113);
nor U825 (N_825,In_62,In_305);
or U826 (N_826,In_414,In_425);
and U827 (N_827,In_432,In_356);
and U828 (N_828,In_455,In_256);
nand U829 (N_829,In_440,In_89);
nand U830 (N_830,In_412,In_145);
nand U831 (N_831,In_113,In_51);
nor U832 (N_832,In_460,In_225);
nand U833 (N_833,In_204,In_402);
nor U834 (N_834,In_391,In_494);
and U835 (N_835,In_225,In_118);
or U836 (N_836,In_422,In_85);
and U837 (N_837,In_136,In_457);
nor U838 (N_838,In_424,In_59);
or U839 (N_839,In_202,In_35);
and U840 (N_840,In_33,In_415);
nor U841 (N_841,In_220,In_321);
or U842 (N_842,In_92,In_329);
and U843 (N_843,In_318,In_9);
and U844 (N_844,In_264,In_268);
nor U845 (N_845,In_329,In_76);
nand U846 (N_846,In_499,In_475);
or U847 (N_847,In_385,In_468);
and U848 (N_848,In_136,In_370);
nand U849 (N_849,In_484,In_253);
or U850 (N_850,In_203,In_291);
xor U851 (N_851,In_188,In_197);
and U852 (N_852,In_228,In_35);
nand U853 (N_853,In_469,In_146);
nand U854 (N_854,In_92,In_78);
or U855 (N_855,In_432,In_33);
and U856 (N_856,In_116,In_276);
and U857 (N_857,In_274,In_1);
and U858 (N_858,In_495,In_96);
or U859 (N_859,In_247,In_267);
or U860 (N_860,In_68,In_336);
nor U861 (N_861,In_219,In_164);
and U862 (N_862,In_248,In_71);
or U863 (N_863,In_97,In_458);
and U864 (N_864,In_465,In_478);
or U865 (N_865,In_226,In_335);
nand U866 (N_866,In_204,In_18);
nor U867 (N_867,In_21,In_348);
and U868 (N_868,In_193,In_55);
nand U869 (N_869,In_185,In_424);
nor U870 (N_870,In_181,In_485);
and U871 (N_871,In_253,In_143);
nor U872 (N_872,In_297,In_166);
or U873 (N_873,In_143,In_483);
and U874 (N_874,In_280,In_332);
or U875 (N_875,In_216,In_156);
or U876 (N_876,In_385,In_434);
nand U877 (N_877,In_308,In_474);
or U878 (N_878,In_110,In_365);
or U879 (N_879,In_188,In_433);
or U880 (N_880,In_129,In_46);
or U881 (N_881,In_474,In_78);
nor U882 (N_882,In_127,In_369);
or U883 (N_883,In_61,In_253);
nor U884 (N_884,In_235,In_441);
or U885 (N_885,In_455,In_258);
nand U886 (N_886,In_473,In_128);
nand U887 (N_887,In_490,In_456);
nand U888 (N_888,In_49,In_352);
and U889 (N_889,In_295,In_486);
or U890 (N_890,In_398,In_379);
nand U891 (N_891,In_350,In_314);
nor U892 (N_892,In_242,In_254);
nor U893 (N_893,In_130,In_317);
or U894 (N_894,In_361,In_420);
and U895 (N_895,In_61,In_150);
or U896 (N_896,In_355,In_431);
or U897 (N_897,In_235,In_231);
nor U898 (N_898,In_72,In_366);
xnor U899 (N_899,In_351,In_215);
or U900 (N_900,In_471,In_327);
and U901 (N_901,In_387,In_464);
or U902 (N_902,In_402,In_85);
xor U903 (N_903,In_109,In_382);
and U904 (N_904,In_424,In_25);
nor U905 (N_905,In_118,In_38);
xnor U906 (N_906,In_482,In_323);
xor U907 (N_907,In_329,In_37);
nor U908 (N_908,In_81,In_114);
and U909 (N_909,In_336,In_220);
or U910 (N_910,In_192,In_219);
or U911 (N_911,In_424,In_62);
nor U912 (N_912,In_80,In_459);
nor U913 (N_913,In_202,In_386);
nor U914 (N_914,In_378,In_117);
and U915 (N_915,In_73,In_400);
and U916 (N_916,In_96,In_397);
and U917 (N_917,In_324,In_68);
or U918 (N_918,In_240,In_94);
and U919 (N_919,In_344,In_235);
or U920 (N_920,In_373,In_376);
or U921 (N_921,In_18,In_15);
and U922 (N_922,In_380,In_232);
nor U923 (N_923,In_218,In_244);
nand U924 (N_924,In_381,In_137);
and U925 (N_925,In_177,In_152);
nand U926 (N_926,In_113,In_92);
nor U927 (N_927,In_382,In_309);
and U928 (N_928,In_6,In_413);
nor U929 (N_929,In_134,In_246);
and U930 (N_930,In_296,In_94);
nand U931 (N_931,In_278,In_314);
nand U932 (N_932,In_307,In_186);
and U933 (N_933,In_304,In_340);
nand U934 (N_934,In_359,In_40);
and U935 (N_935,In_110,In_482);
nor U936 (N_936,In_353,In_481);
nand U937 (N_937,In_211,In_128);
nand U938 (N_938,In_291,In_66);
and U939 (N_939,In_272,In_295);
nand U940 (N_940,In_286,In_135);
nand U941 (N_941,In_481,In_14);
xnor U942 (N_942,In_469,In_497);
or U943 (N_943,In_266,In_300);
or U944 (N_944,In_465,In_295);
nand U945 (N_945,In_315,In_68);
nor U946 (N_946,In_404,In_427);
nand U947 (N_947,In_387,In_469);
nor U948 (N_948,In_84,In_118);
or U949 (N_949,In_354,In_213);
or U950 (N_950,In_82,In_384);
and U951 (N_951,In_121,In_442);
nand U952 (N_952,In_492,In_284);
nor U953 (N_953,In_35,In_351);
or U954 (N_954,In_384,In_316);
nor U955 (N_955,In_445,In_184);
nand U956 (N_956,In_66,In_261);
nor U957 (N_957,In_482,In_411);
and U958 (N_958,In_157,In_177);
or U959 (N_959,In_143,In_338);
nand U960 (N_960,In_166,In_29);
and U961 (N_961,In_265,In_471);
nor U962 (N_962,In_411,In_127);
and U963 (N_963,In_20,In_219);
nor U964 (N_964,In_170,In_124);
nor U965 (N_965,In_207,In_475);
or U966 (N_966,In_443,In_95);
xnor U967 (N_967,In_318,In_413);
and U968 (N_968,In_395,In_320);
nand U969 (N_969,In_419,In_132);
and U970 (N_970,In_162,In_385);
nand U971 (N_971,In_327,In_497);
and U972 (N_972,In_75,In_424);
nor U973 (N_973,In_166,In_169);
nand U974 (N_974,In_115,In_130);
nor U975 (N_975,In_295,In_82);
and U976 (N_976,In_121,In_120);
nand U977 (N_977,In_192,In_32);
nand U978 (N_978,In_384,In_199);
or U979 (N_979,In_429,In_98);
or U980 (N_980,In_375,In_236);
nand U981 (N_981,In_442,In_462);
or U982 (N_982,In_121,In_492);
nand U983 (N_983,In_145,In_266);
nand U984 (N_984,In_424,In_350);
or U985 (N_985,In_275,In_389);
nor U986 (N_986,In_73,In_119);
nand U987 (N_987,In_90,In_432);
nand U988 (N_988,In_84,In_162);
or U989 (N_989,In_485,In_361);
or U990 (N_990,In_59,In_278);
nor U991 (N_991,In_42,In_91);
nor U992 (N_992,In_400,In_4);
nand U993 (N_993,In_263,In_302);
nor U994 (N_994,In_242,In_276);
or U995 (N_995,In_454,In_174);
nor U996 (N_996,In_240,In_191);
or U997 (N_997,In_274,In_254);
and U998 (N_998,In_488,In_384);
nand U999 (N_999,In_397,In_1);
nand U1000 (N_1000,N_530,N_539);
and U1001 (N_1001,N_481,N_763);
and U1002 (N_1002,N_918,N_653);
and U1003 (N_1003,N_292,N_181);
nand U1004 (N_1004,N_11,N_981);
and U1005 (N_1005,N_355,N_625);
and U1006 (N_1006,N_694,N_671);
nor U1007 (N_1007,N_430,N_632);
or U1008 (N_1008,N_478,N_318);
or U1009 (N_1009,N_865,N_161);
nand U1010 (N_1010,N_412,N_484);
or U1011 (N_1011,N_913,N_647);
nand U1012 (N_1012,N_39,N_84);
or U1013 (N_1013,N_483,N_980);
or U1014 (N_1014,N_63,N_819);
or U1015 (N_1015,N_184,N_725);
and U1016 (N_1016,N_234,N_958);
and U1017 (N_1017,N_868,N_49);
nand U1018 (N_1018,N_482,N_891);
nor U1019 (N_1019,N_660,N_629);
nor U1020 (N_1020,N_263,N_453);
nor U1021 (N_1021,N_662,N_202);
and U1022 (N_1022,N_427,N_343);
and U1023 (N_1023,N_390,N_152);
nand U1024 (N_1024,N_515,N_875);
or U1025 (N_1025,N_902,N_406);
nor U1026 (N_1026,N_414,N_247);
nand U1027 (N_1027,N_450,N_762);
or U1028 (N_1028,N_719,N_567);
or U1029 (N_1029,N_947,N_726);
or U1030 (N_1030,N_603,N_806);
nor U1031 (N_1031,N_907,N_335);
nor U1032 (N_1032,N_702,N_999);
nand U1033 (N_1033,N_559,N_943);
nand U1034 (N_1034,N_644,N_945);
and U1035 (N_1035,N_168,N_407);
or U1036 (N_1036,N_944,N_51);
nand U1037 (N_1037,N_342,N_87);
nor U1038 (N_1038,N_142,N_27);
nand U1039 (N_1039,N_790,N_900);
nand U1040 (N_1040,N_445,N_315);
and U1041 (N_1041,N_86,N_976);
nor U1042 (N_1042,N_133,N_587);
or U1043 (N_1043,N_48,N_788);
nand U1044 (N_1044,N_909,N_737);
and U1045 (N_1045,N_322,N_731);
nor U1046 (N_1046,N_700,N_30);
or U1047 (N_1047,N_800,N_718);
or U1048 (N_1048,N_523,N_639);
nor U1049 (N_1049,N_245,N_13);
nor U1050 (N_1050,N_62,N_616);
nand U1051 (N_1051,N_753,N_498);
and U1052 (N_1052,N_104,N_882);
nand U1053 (N_1053,N_962,N_151);
nand U1054 (N_1054,N_334,N_906);
and U1055 (N_1055,N_733,N_823);
nor U1056 (N_1056,N_6,N_768);
and U1057 (N_1057,N_735,N_77);
or U1058 (N_1058,N_465,N_985);
nor U1059 (N_1059,N_249,N_821);
nor U1060 (N_1060,N_712,N_393);
or U1061 (N_1061,N_120,N_618);
nor U1062 (N_1062,N_827,N_112);
and U1063 (N_1063,N_929,N_29);
nor U1064 (N_1064,N_40,N_818);
or U1065 (N_1065,N_71,N_396);
or U1066 (N_1066,N_187,N_248);
or U1067 (N_1067,N_764,N_670);
and U1068 (N_1068,N_989,N_912);
nand U1069 (N_1069,N_423,N_828);
or U1070 (N_1070,N_717,N_138);
and U1071 (N_1071,N_885,N_488);
nor U1072 (N_1072,N_887,N_535);
or U1073 (N_1073,N_287,N_750);
and U1074 (N_1074,N_941,N_919);
nand U1075 (N_1075,N_449,N_429);
nor U1076 (N_1076,N_198,N_507);
and U1077 (N_1077,N_46,N_123);
nor U1078 (N_1078,N_233,N_746);
or U1079 (N_1079,N_744,N_643);
nand U1080 (N_1080,N_37,N_172);
nand U1081 (N_1081,N_417,N_610);
or U1082 (N_1082,N_389,N_816);
nor U1083 (N_1083,N_959,N_373);
and U1084 (N_1084,N_16,N_103);
and U1085 (N_1085,N_739,N_770);
nor U1086 (N_1086,N_192,N_131);
nor U1087 (N_1087,N_923,N_676);
and U1088 (N_1088,N_808,N_226);
nand U1089 (N_1089,N_748,N_973);
or U1090 (N_1090,N_419,N_574);
and U1091 (N_1091,N_297,N_877);
and U1092 (N_1092,N_107,N_765);
and U1093 (N_1093,N_967,N_119);
or U1094 (N_1094,N_99,N_128);
nor U1095 (N_1095,N_214,N_338);
nand U1096 (N_1096,N_640,N_117);
nor U1097 (N_1097,N_599,N_398);
nor U1098 (N_1098,N_328,N_269);
nor U1099 (N_1099,N_946,N_873);
and U1100 (N_1100,N_475,N_490);
nor U1101 (N_1101,N_4,N_74);
or U1102 (N_1102,N_9,N_223);
nand U1103 (N_1103,N_794,N_311);
nor U1104 (N_1104,N_513,N_312);
and U1105 (N_1105,N_924,N_309);
nor U1106 (N_1106,N_303,N_88);
nand U1107 (N_1107,N_296,N_47);
nor U1108 (N_1108,N_841,N_997);
xor U1109 (N_1109,N_569,N_651);
nor U1110 (N_1110,N_705,N_837);
and U1111 (N_1111,N_583,N_26);
nor U1112 (N_1112,N_562,N_815);
nor U1113 (N_1113,N_635,N_914);
nor U1114 (N_1114,N_791,N_145);
or U1115 (N_1115,N_504,N_479);
and U1116 (N_1116,N_463,N_969);
or U1117 (N_1117,N_261,N_938);
or U1118 (N_1118,N_502,N_810);
nand U1119 (N_1119,N_55,N_345);
nand U1120 (N_1120,N_560,N_302);
and U1121 (N_1121,N_211,N_863);
and U1122 (N_1122,N_391,N_301);
and U1123 (N_1123,N_934,N_421);
nor U1124 (N_1124,N_687,N_352);
and U1125 (N_1125,N_260,N_447);
nand U1126 (N_1126,N_267,N_520);
or U1127 (N_1127,N_136,N_455);
and U1128 (N_1128,N_114,N_850);
and U1129 (N_1129,N_171,N_774);
nand U1130 (N_1130,N_540,N_991);
nor U1131 (N_1131,N_22,N_313);
and U1132 (N_1132,N_456,N_408);
xor U1133 (N_1133,N_758,N_283);
nor U1134 (N_1134,N_109,N_21);
or U1135 (N_1135,N_771,N_156);
nand U1136 (N_1136,N_521,N_575);
nand U1137 (N_1137,N_403,N_232);
and U1138 (N_1138,N_295,N_505);
or U1139 (N_1139,N_272,N_489);
and U1140 (N_1140,N_711,N_205);
nor U1141 (N_1141,N_221,N_265);
or U1142 (N_1142,N_217,N_709);
nand U1143 (N_1143,N_52,N_494);
and U1144 (N_1144,N_372,N_582);
nand U1145 (N_1145,N_874,N_693);
nand U1146 (N_1146,N_704,N_473);
nor U1147 (N_1147,N_243,N_208);
and U1148 (N_1148,N_655,N_164);
xor U1149 (N_1149,N_444,N_369);
nor U1150 (N_1150,N_72,N_820);
and U1151 (N_1151,N_91,N_111);
nand U1152 (N_1152,N_387,N_85);
nor U1153 (N_1153,N_833,N_952);
nand U1154 (N_1154,N_305,N_978);
nand U1155 (N_1155,N_351,N_314);
or U1156 (N_1156,N_802,N_749);
nor U1157 (N_1157,N_201,N_224);
or U1158 (N_1158,N_732,N_341);
nand U1159 (N_1159,N_206,N_317);
nor U1160 (N_1160,N_708,N_80);
or U1161 (N_1161,N_817,N_856);
or U1162 (N_1162,N_386,N_320);
or U1163 (N_1163,N_404,N_491);
nand U1164 (N_1164,N_781,N_94);
and U1165 (N_1165,N_755,N_593);
nand U1166 (N_1166,N_975,N_385);
nand U1167 (N_1167,N_257,N_664);
nand U1168 (N_1168,N_858,N_751);
or U1169 (N_1169,N_195,N_552);
nor U1170 (N_1170,N_282,N_888);
and U1171 (N_1171,N_319,N_852);
and U1172 (N_1172,N_778,N_415);
nor U1173 (N_1173,N_571,N_411);
nor U1174 (N_1174,N_754,N_641);
or U1175 (N_1175,N_799,N_880);
and U1176 (N_1176,N_101,N_499);
or U1177 (N_1177,N_225,N_554);
and U1178 (N_1178,N_663,N_501);
and U1179 (N_1179,N_12,N_59);
or U1180 (N_1180,N_689,N_547);
nor U1181 (N_1181,N_595,N_920);
and U1182 (N_1182,N_596,N_200);
and U1183 (N_1183,N_327,N_125);
or U1184 (N_1184,N_273,N_592);
and U1185 (N_1185,N_961,N_35);
and U1186 (N_1186,N_966,N_96);
xor U1187 (N_1187,N_124,N_154);
and U1188 (N_1188,N_987,N_558);
nor U1189 (N_1189,N_957,N_988);
nand U1190 (N_1190,N_843,N_76);
and U1191 (N_1191,N_127,N_264);
nand U1192 (N_1192,N_310,N_650);
and U1193 (N_1193,N_878,N_165);
or U1194 (N_1194,N_374,N_426);
and U1195 (N_1195,N_609,N_684);
xor U1196 (N_1196,N_139,N_908);
nand U1197 (N_1197,N_715,N_840);
nor U1198 (N_1198,N_678,N_5);
nand U1199 (N_1199,N_446,N_691);
nand U1200 (N_1200,N_178,N_543);
and U1201 (N_1201,N_759,N_734);
xnor U1202 (N_1202,N_646,N_326);
and U1203 (N_1203,N_935,N_23);
nor U1204 (N_1204,N_576,N_626);
or U1205 (N_1205,N_228,N_948);
or U1206 (N_1206,N_75,N_25);
and U1207 (N_1207,N_548,N_578);
and U1208 (N_1208,N_155,N_382);
nor U1209 (N_1209,N_306,N_531);
nand U1210 (N_1210,N_8,N_986);
or U1211 (N_1211,N_497,N_469);
nor U1212 (N_1212,N_285,N_402);
or U1213 (N_1213,N_207,N_238);
and U1214 (N_1214,N_370,N_50);
or U1215 (N_1215,N_937,N_604);
and U1216 (N_1216,N_814,N_537);
nand U1217 (N_1217,N_955,N_714);
nor U1218 (N_1218,N_1,N_174);
nand U1219 (N_1219,N_400,N_784);
nor U1220 (N_1220,N_364,N_363);
nand U1221 (N_1221,N_798,N_602);
or U1222 (N_1222,N_897,N_97);
or U1223 (N_1223,N_33,N_607);
or U1224 (N_1224,N_92,N_996);
or U1225 (N_1225,N_332,N_274);
nand U1226 (N_1226,N_579,N_425);
nand U1227 (N_1227,N_896,N_358);
or U1228 (N_1228,N_106,N_679);
and U1229 (N_1229,N_801,N_876);
and U1230 (N_1230,N_786,N_826);
or U1231 (N_1231,N_685,N_573);
or U1232 (N_1232,N_190,N_659);
or U1233 (N_1233,N_621,N_254);
nor U1234 (N_1234,N_19,N_835);
xnor U1235 (N_1235,N_901,N_340);
nand U1236 (N_1236,N_433,N_300);
and U1237 (N_1237,N_89,N_471);
nor U1238 (N_1238,N_448,N_276);
nor U1239 (N_1239,N_204,N_728);
nand U1240 (N_1240,N_510,N_898);
nor U1241 (N_1241,N_69,N_894);
and U1242 (N_1242,N_251,N_658);
or U1243 (N_1243,N_468,N_3);
nor U1244 (N_1244,N_682,N_636);
nand U1245 (N_1245,N_506,N_782);
and U1246 (N_1246,N_825,N_144);
nand U1247 (N_1247,N_931,N_974);
nor U1248 (N_1248,N_927,N_461);
or U1249 (N_1249,N_730,N_839);
or U1250 (N_1250,N_525,N_278);
nor U1251 (N_1251,N_42,N_527);
or U1252 (N_1252,N_118,N_44);
and U1253 (N_1253,N_886,N_157);
nor U1254 (N_1254,N_173,N_665);
xnor U1255 (N_1255,N_255,N_93);
and U1256 (N_1256,N_60,N_162);
and U1257 (N_1257,N_699,N_928);
and U1258 (N_1258,N_968,N_995);
nor U1259 (N_1259,N_443,N_964);
and U1260 (N_1260,N_323,N_108);
nand U1261 (N_1261,N_805,N_581);
and U1262 (N_1262,N_724,N_881);
nand U1263 (N_1263,N_526,N_321);
or U1264 (N_1264,N_851,N_707);
nand U1265 (N_1265,N_235,N_434);
or U1266 (N_1266,N_533,N_182);
nor U1267 (N_1267,N_477,N_410);
or U1268 (N_1268,N_409,N_31);
nor U1269 (N_1269,N_600,N_102);
nor U1270 (N_1270,N_67,N_992);
and U1271 (N_1271,N_793,N_727);
nand U1272 (N_1272,N_516,N_167);
nand U1273 (N_1273,N_683,N_209);
nor U1274 (N_1274,N_696,N_736);
or U1275 (N_1275,N_557,N_803);
or U1276 (N_1276,N_842,N_422);
and U1277 (N_1277,N_698,N_54);
or U1278 (N_1278,N_633,N_509);
or U1279 (N_1279,N_706,N_695);
nand U1280 (N_1280,N_492,N_472);
and U1281 (N_1281,N_681,N_18);
xnor U1282 (N_1282,N_541,N_889);
nand U1283 (N_1283,N_413,N_418);
or U1284 (N_1284,N_384,N_28);
or U1285 (N_1285,N_776,N_7);
and U1286 (N_1286,N_553,N_242);
or U1287 (N_1287,N_916,N_892);
and U1288 (N_1288,N_847,N_0);
nor U1289 (N_1289,N_652,N_220);
or U1290 (N_1290,N_110,N_230);
and U1291 (N_1291,N_487,N_637);
nor U1292 (N_1292,N_316,N_809);
and U1293 (N_1293,N_137,N_667);
and U1294 (N_1294,N_258,N_738);
or U1295 (N_1295,N_859,N_550);
nor U1296 (N_1296,N_388,N_831);
and U1297 (N_1297,N_237,N_349);
nand U1298 (N_1298,N_135,N_792);
and U1299 (N_1299,N_360,N_910);
nand U1300 (N_1300,N_457,N_241);
nor U1301 (N_1301,N_722,N_20);
nand U1302 (N_1302,N_532,N_972);
nand U1303 (N_1303,N_890,N_512);
or U1304 (N_1304,N_741,N_756);
or U1305 (N_1305,N_307,N_377);
and U1306 (N_1306,N_555,N_942);
xor U1307 (N_1307,N_862,N_518);
and U1308 (N_1308,N_729,N_486);
and U1309 (N_1309,N_115,N_769);
nand U1310 (N_1310,N_713,N_848);
nor U1311 (N_1311,N_572,N_866);
and U1312 (N_1312,N_304,N_534);
and U1313 (N_1313,N_361,N_170);
and U1314 (N_1314,N_522,N_379);
nand U1315 (N_1315,N_657,N_116);
and U1316 (N_1316,N_546,N_933);
nand U1317 (N_1317,N_993,N_517);
or U1318 (N_1318,N_65,N_288);
nor U1319 (N_1319,N_614,N_939);
nor U1320 (N_1320,N_467,N_246);
nand U1321 (N_1321,N_857,N_45);
nand U1322 (N_1322,N_846,N_395);
nand U1323 (N_1323,N_284,N_917);
nand U1324 (N_1324,N_982,N_812);
and U1325 (N_1325,N_542,N_844);
nand U1326 (N_1326,N_435,N_963);
nor U1327 (N_1327,N_971,N_150);
or U1328 (N_1328,N_464,N_675);
and U1329 (N_1329,N_197,N_199);
and U1330 (N_1330,N_775,N_867);
nor U1331 (N_1331,N_325,N_869);
and U1332 (N_1332,N_371,N_141);
and U1333 (N_1333,N_796,N_879);
nand U1334 (N_1334,N_466,N_397);
nor U1335 (N_1335,N_564,N_983);
nand U1336 (N_1336,N_291,N_495);
nor U1337 (N_1337,N_745,N_742);
nor U1338 (N_1338,N_280,N_367);
and U1339 (N_1339,N_766,N_606);
or U1340 (N_1340,N_854,N_346);
or U1341 (N_1341,N_915,N_905);
or U1342 (N_1342,N_281,N_723);
nor U1343 (N_1343,N_813,N_143);
nor U1344 (N_1344,N_638,N_797);
nand U1345 (N_1345,N_872,N_777);
or U1346 (N_1346,N_210,N_68);
or U1347 (N_1347,N_271,N_493);
or U1348 (N_1348,N_613,N_252);
nand U1349 (N_1349,N_589,N_420);
nand U1350 (N_1350,N_203,N_615);
or U1351 (N_1351,N_259,N_591);
nor U1352 (N_1352,N_376,N_380);
or U1353 (N_1353,N_381,N_836);
and U1354 (N_1354,N_462,N_105);
nor U1355 (N_1355,N_950,N_268);
nand U1356 (N_1356,N_392,N_36);
nand U1357 (N_1357,N_611,N_761);
or U1358 (N_1358,N_563,N_936);
or U1359 (N_1359,N_34,N_838);
or U1360 (N_1360,N_286,N_474);
nand U1361 (N_1361,N_686,N_921);
nand U1362 (N_1362,N_953,N_503);
nor U1363 (N_1363,N_132,N_357);
nand U1364 (N_1364,N_146,N_324);
nand U1365 (N_1365,N_645,N_15);
or U1366 (N_1366,N_747,N_216);
nand U1367 (N_1367,N_965,N_185);
and U1368 (N_1368,N_470,N_331);
nor U1369 (N_1369,N_416,N_218);
nand U1370 (N_1370,N_439,N_64);
or U1371 (N_1371,N_903,N_951);
and U1372 (N_1372,N_148,N_870);
and U1373 (N_1373,N_624,N_979);
nand U1374 (N_1374,N_43,N_960);
or U1375 (N_1375,N_549,N_824);
nand U1376 (N_1376,N_811,N_368);
or U1377 (N_1377,N_612,N_126);
xor U1378 (N_1378,N_634,N_122);
nand U1379 (N_1379,N_294,N_436);
or U1380 (N_1380,N_459,N_690);
xnor U1381 (N_1381,N_787,N_191);
or U1382 (N_1382,N_590,N_853);
and U1383 (N_1383,N_956,N_990);
nand U1384 (N_1384,N_716,N_849);
or U1385 (N_1385,N_783,N_56);
nor U1386 (N_1386,N_95,N_38);
and U1387 (N_1387,N_551,N_720);
nor U1388 (N_1388,N_186,N_177);
nor U1389 (N_1389,N_767,N_884);
and U1390 (N_1390,N_163,N_688);
or U1391 (N_1391,N_855,N_622);
and U1392 (N_1392,N_236,N_757);
and U1393 (N_1393,N_519,N_864);
and U1394 (N_1394,N_290,N_785);
and U1395 (N_1395,N_925,N_262);
or U1396 (N_1396,N_597,N_773);
nor U1397 (N_1397,N_932,N_61);
nor U1398 (N_1398,N_860,N_772);
and U1399 (N_1399,N_375,N_437);
and U1400 (N_1400,N_356,N_586);
and U1401 (N_1401,N_147,N_710);
nand U1402 (N_1402,N_438,N_188);
or U1403 (N_1403,N_212,N_353);
or U1404 (N_1404,N_79,N_451);
nor U1405 (N_1405,N_588,N_529);
and U1406 (N_1406,N_480,N_442);
or U1407 (N_1407,N_175,N_366);
nand U1408 (N_1408,N_954,N_289);
nor U1409 (N_1409,N_90,N_53);
or U1410 (N_1410,N_70,N_183);
nand U1411 (N_1411,N_500,N_807);
nor U1412 (N_1412,N_893,N_703);
xor U1413 (N_1413,N_779,N_630);
nor U1414 (N_1414,N_672,N_78);
nor U1415 (N_1415,N_619,N_424);
or U1416 (N_1416,N_160,N_601);
or U1417 (N_1417,N_904,N_405);
nor U1418 (N_1418,N_219,N_428);
nor U1419 (N_1419,N_832,N_176);
nor U1420 (N_1420,N_524,N_354);
or U1421 (N_1421,N_795,N_496);
nand U1422 (N_1422,N_460,N_570);
nand U1423 (N_1423,N_344,N_485);
and U1424 (N_1424,N_677,N_441);
and U1425 (N_1425,N_83,N_140);
and U1426 (N_1426,N_674,N_10);
and U1427 (N_1427,N_394,N_347);
nand U1428 (N_1428,N_511,N_584);
or U1429 (N_1429,N_538,N_594);
nand U1430 (N_1430,N_58,N_158);
or U1431 (N_1431,N_365,N_608);
or U1432 (N_1432,N_627,N_949);
and U1433 (N_1433,N_279,N_256);
or U1434 (N_1434,N_277,N_82);
nand U1435 (N_1435,N_545,N_829);
nand U1436 (N_1436,N_654,N_565);
or U1437 (N_1437,N_930,N_830);
xnor U1438 (N_1438,N_922,N_508);
or U1439 (N_1439,N_244,N_180);
or U1440 (N_1440,N_668,N_130);
nor U1441 (N_1441,N_431,N_166);
nand U1442 (N_1442,N_159,N_348);
or U1443 (N_1443,N_454,N_193);
nand U1444 (N_1444,N_977,N_760);
nor U1445 (N_1445,N_580,N_926);
or U1446 (N_1446,N_66,N_266);
nor U1447 (N_1447,N_899,N_432);
nand U1448 (N_1448,N_81,N_14);
or U1449 (N_1449,N_743,N_440);
or U1450 (N_1450,N_649,N_528);
nand U1451 (N_1451,N_32,N_189);
or U1452 (N_1452,N_631,N_362);
nand U1453 (N_1453,N_359,N_669);
and U1454 (N_1454,N_229,N_100);
nand U1455 (N_1455,N_661,N_605);
nor U1456 (N_1456,N_458,N_336);
and U1457 (N_1457,N_231,N_293);
nand U1458 (N_1458,N_642,N_617);
and U1459 (N_1459,N_701,N_994);
nand U1460 (N_1460,N_250,N_215);
or U1461 (N_1461,N_861,N_383);
nand U1462 (N_1462,N_620,N_845);
nor U1463 (N_1463,N_623,N_721);
and U1464 (N_1464,N_213,N_298);
nand U1465 (N_1465,N_561,N_598);
and U1466 (N_1466,N_149,N_113);
nor U1467 (N_1467,N_692,N_308);
and U1468 (N_1468,N_57,N_275);
nor U1469 (N_1469,N_780,N_998);
and U1470 (N_1470,N_911,N_804);
and U1471 (N_1471,N_536,N_98);
and U1472 (N_1472,N_227,N_239);
nor U1473 (N_1473,N_194,N_2);
and U1474 (N_1474,N_452,N_401);
nand U1475 (N_1475,N_568,N_544);
nor U1476 (N_1476,N_834,N_656);
nor U1477 (N_1477,N_270,N_330);
nor U1478 (N_1478,N_253,N_169);
nor U1479 (N_1479,N_333,N_73);
or U1480 (N_1480,N_740,N_24);
and U1481 (N_1481,N_329,N_940);
and U1482 (N_1482,N_153,N_895);
or U1483 (N_1483,N_350,N_697);
nor U1484 (N_1484,N_299,N_121);
or U1485 (N_1485,N_17,N_222);
nor U1486 (N_1486,N_129,N_673);
nand U1487 (N_1487,N_476,N_970);
or U1488 (N_1488,N_378,N_789);
nor U1489 (N_1489,N_984,N_752);
nand U1490 (N_1490,N_337,N_41);
nand U1491 (N_1491,N_628,N_179);
and U1492 (N_1492,N_577,N_399);
nand U1493 (N_1493,N_556,N_196);
or U1494 (N_1494,N_680,N_566);
and U1495 (N_1495,N_648,N_339);
nand U1496 (N_1496,N_514,N_871);
xnor U1497 (N_1497,N_666,N_822);
or U1498 (N_1498,N_585,N_883);
nand U1499 (N_1499,N_134,N_240);
and U1500 (N_1500,N_788,N_982);
nor U1501 (N_1501,N_664,N_877);
or U1502 (N_1502,N_695,N_259);
nor U1503 (N_1503,N_711,N_68);
or U1504 (N_1504,N_509,N_974);
nand U1505 (N_1505,N_599,N_42);
nand U1506 (N_1506,N_388,N_39);
xnor U1507 (N_1507,N_176,N_32);
nor U1508 (N_1508,N_872,N_945);
nand U1509 (N_1509,N_939,N_787);
or U1510 (N_1510,N_268,N_893);
xor U1511 (N_1511,N_71,N_98);
nor U1512 (N_1512,N_689,N_327);
nand U1513 (N_1513,N_907,N_141);
nand U1514 (N_1514,N_338,N_495);
nor U1515 (N_1515,N_417,N_191);
nand U1516 (N_1516,N_269,N_335);
nor U1517 (N_1517,N_81,N_502);
nand U1518 (N_1518,N_457,N_440);
or U1519 (N_1519,N_434,N_779);
nor U1520 (N_1520,N_95,N_917);
nand U1521 (N_1521,N_561,N_922);
xor U1522 (N_1522,N_59,N_393);
or U1523 (N_1523,N_154,N_549);
nor U1524 (N_1524,N_581,N_535);
nand U1525 (N_1525,N_771,N_467);
nand U1526 (N_1526,N_937,N_945);
and U1527 (N_1527,N_311,N_485);
nand U1528 (N_1528,N_282,N_904);
nor U1529 (N_1529,N_942,N_35);
or U1530 (N_1530,N_331,N_899);
nand U1531 (N_1531,N_239,N_301);
and U1532 (N_1532,N_823,N_570);
or U1533 (N_1533,N_593,N_682);
and U1534 (N_1534,N_927,N_136);
and U1535 (N_1535,N_906,N_327);
and U1536 (N_1536,N_719,N_341);
nor U1537 (N_1537,N_32,N_794);
and U1538 (N_1538,N_152,N_275);
or U1539 (N_1539,N_515,N_702);
nand U1540 (N_1540,N_419,N_554);
xnor U1541 (N_1541,N_69,N_587);
nor U1542 (N_1542,N_255,N_50);
or U1543 (N_1543,N_747,N_421);
nor U1544 (N_1544,N_369,N_160);
or U1545 (N_1545,N_367,N_182);
or U1546 (N_1546,N_813,N_740);
or U1547 (N_1547,N_828,N_580);
xor U1548 (N_1548,N_549,N_673);
or U1549 (N_1549,N_777,N_764);
and U1550 (N_1550,N_932,N_331);
or U1551 (N_1551,N_353,N_193);
nand U1552 (N_1552,N_874,N_532);
or U1553 (N_1553,N_599,N_701);
or U1554 (N_1554,N_825,N_918);
nor U1555 (N_1555,N_151,N_78);
or U1556 (N_1556,N_416,N_636);
nor U1557 (N_1557,N_807,N_348);
and U1558 (N_1558,N_130,N_405);
nor U1559 (N_1559,N_18,N_102);
nor U1560 (N_1560,N_168,N_420);
nor U1561 (N_1561,N_374,N_94);
or U1562 (N_1562,N_569,N_719);
or U1563 (N_1563,N_55,N_344);
nand U1564 (N_1564,N_13,N_687);
nor U1565 (N_1565,N_359,N_411);
nand U1566 (N_1566,N_6,N_822);
nand U1567 (N_1567,N_763,N_998);
nor U1568 (N_1568,N_498,N_166);
and U1569 (N_1569,N_68,N_754);
nand U1570 (N_1570,N_34,N_926);
and U1571 (N_1571,N_438,N_14);
nand U1572 (N_1572,N_304,N_704);
or U1573 (N_1573,N_966,N_334);
or U1574 (N_1574,N_671,N_7);
nand U1575 (N_1575,N_401,N_86);
nand U1576 (N_1576,N_992,N_876);
nor U1577 (N_1577,N_295,N_381);
and U1578 (N_1578,N_647,N_180);
nor U1579 (N_1579,N_922,N_461);
and U1580 (N_1580,N_170,N_793);
nand U1581 (N_1581,N_386,N_332);
nand U1582 (N_1582,N_343,N_744);
nor U1583 (N_1583,N_535,N_699);
or U1584 (N_1584,N_586,N_474);
nand U1585 (N_1585,N_49,N_284);
nor U1586 (N_1586,N_48,N_209);
nor U1587 (N_1587,N_788,N_490);
and U1588 (N_1588,N_45,N_823);
nor U1589 (N_1589,N_408,N_903);
and U1590 (N_1590,N_121,N_893);
nand U1591 (N_1591,N_992,N_440);
and U1592 (N_1592,N_936,N_276);
nor U1593 (N_1593,N_438,N_714);
nand U1594 (N_1594,N_659,N_655);
nor U1595 (N_1595,N_438,N_829);
or U1596 (N_1596,N_27,N_875);
or U1597 (N_1597,N_128,N_977);
nand U1598 (N_1598,N_763,N_810);
nor U1599 (N_1599,N_783,N_979);
and U1600 (N_1600,N_626,N_640);
and U1601 (N_1601,N_288,N_235);
nor U1602 (N_1602,N_493,N_935);
nand U1603 (N_1603,N_253,N_531);
nor U1604 (N_1604,N_944,N_275);
nand U1605 (N_1605,N_671,N_609);
or U1606 (N_1606,N_446,N_851);
nor U1607 (N_1607,N_644,N_418);
nor U1608 (N_1608,N_39,N_143);
or U1609 (N_1609,N_380,N_411);
and U1610 (N_1610,N_706,N_626);
or U1611 (N_1611,N_743,N_314);
nand U1612 (N_1612,N_443,N_118);
nor U1613 (N_1613,N_175,N_590);
nand U1614 (N_1614,N_770,N_921);
or U1615 (N_1615,N_832,N_893);
or U1616 (N_1616,N_376,N_862);
and U1617 (N_1617,N_293,N_108);
nor U1618 (N_1618,N_701,N_486);
nand U1619 (N_1619,N_408,N_12);
and U1620 (N_1620,N_555,N_377);
and U1621 (N_1621,N_517,N_670);
and U1622 (N_1622,N_847,N_941);
nand U1623 (N_1623,N_445,N_695);
nor U1624 (N_1624,N_776,N_270);
nor U1625 (N_1625,N_447,N_131);
nand U1626 (N_1626,N_67,N_772);
and U1627 (N_1627,N_159,N_730);
or U1628 (N_1628,N_162,N_569);
and U1629 (N_1629,N_724,N_78);
nand U1630 (N_1630,N_334,N_183);
or U1631 (N_1631,N_330,N_933);
nand U1632 (N_1632,N_16,N_159);
nand U1633 (N_1633,N_216,N_70);
nor U1634 (N_1634,N_101,N_698);
or U1635 (N_1635,N_260,N_668);
and U1636 (N_1636,N_940,N_330);
nand U1637 (N_1637,N_521,N_776);
nor U1638 (N_1638,N_340,N_409);
nor U1639 (N_1639,N_979,N_218);
and U1640 (N_1640,N_991,N_485);
or U1641 (N_1641,N_629,N_998);
and U1642 (N_1642,N_183,N_151);
nor U1643 (N_1643,N_324,N_748);
nor U1644 (N_1644,N_854,N_13);
or U1645 (N_1645,N_307,N_87);
nor U1646 (N_1646,N_431,N_619);
nor U1647 (N_1647,N_36,N_823);
nand U1648 (N_1648,N_507,N_85);
nand U1649 (N_1649,N_382,N_92);
nor U1650 (N_1650,N_885,N_435);
or U1651 (N_1651,N_11,N_164);
or U1652 (N_1652,N_96,N_804);
and U1653 (N_1653,N_418,N_684);
and U1654 (N_1654,N_775,N_728);
or U1655 (N_1655,N_945,N_622);
and U1656 (N_1656,N_725,N_158);
nand U1657 (N_1657,N_690,N_994);
nand U1658 (N_1658,N_347,N_423);
nor U1659 (N_1659,N_680,N_68);
nand U1660 (N_1660,N_653,N_838);
nor U1661 (N_1661,N_993,N_641);
nor U1662 (N_1662,N_96,N_571);
nor U1663 (N_1663,N_346,N_503);
and U1664 (N_1664,N_48,N_259);
nand U1665 (N_1665,N_713,N_372);
nor U1666 (N_1666,N_279,N_662);
or U1667 (N_1667,N_174,N_524);
or U1668 (N_1668,N_106,N_949);
nor U1669 (N_1669,N_427,N_874);
nand U1670 (N_1670,N_492,N_593);
or U1671 (N_1671,N_806,N_544);
nor U1672 (N_1672,N_268,N_971);
nand U1673 (N_1673,N_755,N_15);
or U1674 (N_1674,N_167,N_864);
nand U1675 (N_1675,N_974,N_86);
and U1676 (N_1676,N_834,N_473);
nor U1677 (N_1677,N_80,N_454);
nor U1678 (N_1678,N_87,N_435);
and U1679 (N_1679,N_816,N_226);
or U1680 (N_1680,N_806,N_891);
nor U1681 (N_1681,N_994,N_227);
and U1682 (N_1682,N_78,N_324);
and U1683 (N_1683,N_462,N_634);
and U1684 (N_1684,N_477,N_170);
nor U1685 (N_1685,N_688,N_188);
nand U1686 (N_1686,N_124,N_3);
nor U1687 (N_1687,N_834,N_801);
nand U1688 (N_1688,N_787,N_259);
or U1689 (N_1689,N_911,N_811);
nor U1690 (N_1690,N_206,N_976);
and U1691 (N_1691,N_889,N_134);
or U1692 (N_1692,N_488,N_178);
or U1693 (N_1693,N_415,N_722);
and U1694 (N_1694,N_587,N_610);
nand U1695 (N_1695,N_453,N_212);
and U1696 (N_1696,N_886,N_821);
nand U1697 (N_1697,N_879,N_565);
or U1698 (N_1698,N_525,N_117);
xor U1699 (N_1699,N_901,N_483);
nor U1700 (N_1700,N_781,N_827);
and U1701 (N_1701,N_737,N_608);
xnor U1702 (N_1702,N_877,N_311);
nand U1703 (N_1703,N_96,N_711);
and U1704 (N_1704,N_64,N_356);
or U1705 (N_1705,N_831,N_673);
nand U1706 (N_1706,N_188,N_133);
or U1707 (N_1707,N_599,N_971);
nor U1708 (N_1708,N_231,N_247);
nor U1709 (N_1709,N_546,N_433);
and U1710 (N_1710,N_950,N_103);
and U1711 (N_1711,N_880,N_120);
or U1712 (N_1712,N_306,N_191);
and U1713 (N_1713,N_778,N_770);
nor U1714 (N_1714,N_91,N_854);
and U1715 (N_1715,N_954,N_208);
nor U1716 (N_1716,N_472,N_724);
and U1717 (N_1717,N_150,N_139);
nor U1718 (N_1718,N_925,N_336);
and U1719 (N_1719,N_263,N_233);
nand U1720 (N_1720,N_165,N_757);
nand U1721 (N_1721,N_246,N_411);
nor U1722 (N_1722,N_759,N_56);
nor U1723 (N_1723,N_675,N_70);
nor U1724 (N_1724,N_560,N_759);
or U1725 (N_1725,N_838,N_85);
and U1726 (N_1726,N_93,N_652);
nand U1727 (N_1727,N_12,N_823);
nor U1728 (N_1728,N_287,N_713);
nand U1729 (N_1729,N_625,N_515);
and U1730 (N_1730,N_451,N_340);
or U1731 (N_1731,N_638,N_430);
nand U1732 (N_1732,N_150,N_800);
nor U1733 (N_1733,N_474,N_86);
nor U1734 (N_1734,N_741,N_901);
nor U1735 (N_1735,N_475,N_878);
and U1736 (N_1736,N_974,N_803);
nand U1737 (N_1737,N_892,N_842);
nand U1738 (N_1738,N_583,N_394);
and U1739 (N_1739,N_205,N_437);
nor U1740 (N_1740,N_159,N_752);
nand U1741 (N_1741,N_854,N_380);
nor U1742 (N_1742,N_695,N_178);
nor U1743 (N_1743,N_482,N_804);
or U1744 (N_1744,N_459,N_470);
and U1745 (N_1745,N_35,N_107);
nor U1746 (N_1746,N_925,N_763);
and U1747 (N_1747,N_599,N_558);
nand U1748 (N_1748,N_518,N_956);
and U1749 (N_1749,N_982,N_201);
or U1750 (N_1750,N_324,N_661);
nor U1751 (N_1751,N_75,N_57);
or U1752 (N_1752,N_751,N_955);
nor U1753 (N_1753,N_120,N_806);
and U1754 (N_1754,N_714,N_861);
and U1755 (N_1755,N_121,N_949);
nand U1756 (N_1756,N_120,N_56);
or U1757 (N_1757,N_146,N_925);
or U1758 (N_1758,N_561,N_34);
nand U1759 (N_1759,N_466,N_359);
or U1760 (N_1760,N_715,N_507);
nand U1761 (N_1761,N_24,N_884);
nand U1762 (N_1762,N_207,N_611);
or U1763 (N_1763,N_352,N_418);
and U1764 (N_1764,N_857,N_174);
nor U1765 (N_1765,N_570,N_28);
nor U1766 (N_1766,N_885,N_66);
nor U1767 (N_1767,N_806,N_408);
and U1768 (N_1768,N_977,N_608);
and U1769 (N_1769,N_741,N_412);
and U1770 (N_1770,N_62,N_263);
nor U1771 (N_1771,N_97,N_267);
nor U1772 (N_1772,N_316,N_874);
xnor U1773 (N_1773,N_22,N_653);
or U1774 (N_1774,N_696,N_288);
nand U1775 (N_1775,N_478,N_466);
and U1776 (N_1776,N_149,N_400);
nand U1777 (N_1777,N_516,N_169);
or U1778 (N_1778,N_174,N_42);
or U1779 (N_1779,N_635,N_889);
nand U1780 (N_1780,N_968,N_795);
or U1781 (N_1781,N_413,N_26);
or U1782 (N_1782,N_273,N_162);
or U1783 (N_1783,N_460,N_351);
nand U1784 (N_1784,N_881,N_365);
xnor U1785 (N_1785,N_332,N_333);
nand U1786 (N_1786,N_535,N_571);
and U1787 (N_1787,N_413,N_661);
nor U1788 (N_1788,N_510,N_824);
and U1789 (N_1789,N_15,N_428);
and U1790 (N_1790,N_711,N_270);
nand U1791 (N_1791,N_277,N_975);
nand U1792 (N_1792,N_378,N_914);
or U1793 (N_1793,N_519,N_678);
or U1794 (N_1794,N_256,N_46);
or U1795 (N_1795,N_967,N_336);
nand U1796 (N_1796,N_634,N_165);
nor U1797 (N_1797,N_680,N_261);
or U1798 (N_1798,N_91,N_496);
nor U1799 (N_1799,N_548,N_111);
and U1800 (N_1800,N_504,N_487);
or U1801 (N_1801,N_490,N_909);
nand U1802 (N_1802,N_973,N_573);
and U1803 (N_1803,N_88,N_182);
nand U1804 (N_1804,N_993,N_501);
nor U1805 (N_1805,N_141,N_920);
nor U1806 (N_1806,N_447,N_224);
or U1807 (N_1807,N_560,N_658);
nand U1808 (N_1808,N_27,N_743);
nor U1809 (N_1809,N_572,N_46);
and U1810 (N_1810,N_769,N_305);
nor U1811 (N_1811,N_483,N_72);
or U1812 (N_1812,N_147,N_655);
or U1813 (N_1813,N_782,N_184);
nand U1814 (N_1814,N_691,N_180);
and U1815 (N_1815,N_54,N_794);
or U1816 (N_1816,N_965,N_9);
and U1817 (N_1817,N_513,N_65);
nor U1818 (N_1818,N_298,N_817);
or U1819 (N_1819,N_239,N_648);
nor U1820 (N_1820,N_77,N_466);
nor U1821 (N_1821,N_45,N_818);
and U1822 (N_1822,N_470,N_648);
or U1823 (N_1823,N_680,N_621);
or U1824 (N_1824,N_836,N_935);
or U1825 (N_1825,N_312,N_417);
nor U1826 (N_1826,N_222,N_514);
nand U1827 (N_1827,N_145,N_832);
and U1828 (N_1828,N_104,N_368);
nor U1829 (N_1829,N_300,N_73);
and U1830 (N_1830,N_39,N_374);
nand U1831 (N_1831,N_718,N_246);
nand U1832 (N_1832,N_335,N_725);
and U1833 (N_1833,N_829,N_878);
nor U1834 (N_1834,N_756,N_378);
nand U1835 (N_1835,N_999,N_375);
and U1836 (N_1836,N_58,N_348);
and U1837 (N_1837,N_257,N_319);
and U1838 (N_1838,N_717,N_562);
and U1839 (N_1839,N_305,N_128);
nor U1840 (N_1840,N_87,N_531);
nor U1841 (N_1841,N_43,N_64);
and U1842 (N_1842,N_51,N_741);
nand U1843 (N_1843,N_274,N_168);
nand U1844 (N_1844,N_851,N_593);
nand U1845 (N_1845,N_574,N_771);
and U1846 (N_1846,N_343,N_922);
and U1847 (N_1847,N_222,N_310);
and U1848 (N_1848,N_287,N_488);
nand U1849 (N_1849,N_20,N_452);
or U1850 (N_1850,N_890,N_602);
nor U1851 (N_1851,N_105,N_212);
nand U1852 (N_1852,N_82,N_603);
or U1853 (N_1853,N_119,N_166);
nor U1854 (N_1854,N_697,N_874);
nor U1855 (N_1855,N_147,N_406);
or U1856 (N_1856,N_499,N_758);
nand U1857 (N_1857,N_455,N_705);
nand U1858 (N_1858,N_638,N_818);
nor U1859 (N_1859,N_766,N_756);
nor U1860 (N_1860,N_102,N_270);
or U1861 (N_1861,N_540,N_362);
or U1862 (N_1862,N_353,N_852);
and U1863 (N_1863,N_615,N_477);
nand U1864 (N_1864,N_17,N_710);
nor U1865 (N_1865,N_845,N_143);
and U1866 (N_1866,N_782,N_715);
nand U1867 (N_1867,N_503,N_256);
nand U1868 (N_1868,N_654,N_102);
or U1869 (N_1869,N_900,N_61);
and U1870 (N_1870,N_157,N_856);
or U1871 (N_1871,N_264,N_14);
nand U1872 (N_1872,N_9,N_851);
and U1873 (N_1873,N_593,N_999);
xor U1874 (N_1874,N_674,N_616);
and U1875 (N_1875,N_157,N_181);
and U1876 (N_1876,N_45,N_47);
nor U1877 (N_1877,N_536,N_370);
nand U1878 (N_1878,N_780,N_912);
nand U1879 (N_1879,N_270,N_290);
or U1880 (N_1880,N_995,N_965);
nand U1881 (N_1881,N_547,N_995);
nor U1882 (N_1882,N_547,N_107);
nand U1883 (N_1883,N_20,N_945);
nand U1884 (N_1884,N_819,N_238);
or U1885 (N_1885,N_900,N_605);
or U1886 (N_1886,N_988,N_828);
nor U1887 (N_1887,N_406,N_915);
and U1888 (N_1888,N_419,N_142);
and U1889 (N_1889,N_430,N_399);
nand U1890 (N_1890,N_143,N_107);
and U1891 (N_1891,N_626,N_583);
nor U1892 (N_1892,N_30,N_756);
nor U1893 (N_1893,N_948,N_210);
or U1894 (N_1894,N_538,N_869);
or U1895 (N_1895,N_739,N_472);
nor U1896 (N_1896,N_759,N_474);
nor U1897 (N_1897,N_649,N_234);
nand U1898 (N_1898,N_194,N_616);
nor U1899 (N_1899,N_410,N_28);
and U1900 (N_1900,N_949,N_370);
and U1901 (N_1901,N_797,N_454);
xnor U1902 (N_1902,N_625,N_670);
nor U1903 (N_1903,N_233,N_384);
or U1904 (N_1904,N_421,N_523);
or U1905 (N_1905,N_991,N_344);
or U1906 (N_1906,N_783,N_246);
and U1907 (N_1907,N_44,N_521);
nand U1908 (N_1908,N_255,N_88);
nor U1909 (N_1909,N_390,N_1);
nor U1910 (N_1910,N_574,N_488);
nand U1911 (N_1911,N_483,N_547);
or U1912 (N_1912,N_686,N_653);
nand U1913 (N_1913,N_909,N_617);
and U1914 (N_1914,N_257,N_913);
or U1915 (N_1915,N_816,N_531);
or U1916 (N_1916,N_270,N_874);
nor U1917 (N_1917,N_377,N_927);
nand U1918 (N_1918,N_39,N_22);
and U1919 (N_1919,N_583,N_686);
and U1920 (N_1920,N_237,N_208);
or U1921 (N_1921,N_368,N_970);
nor U1922 (N_1922,N_533,N_313);
and U1923 (N_1923,N_634,N_914);
nand U1924 (N_1924,N_166,N_869);
nor U1925 (N_1925,N_177,N_539);
nor U1926 (N_1926,N_415,N_513);
nand U1927 (N_1927,N_32,N_172);
or U1928 (N_1928,N_20,N_959);
nand U1929 (N_1929,N_617,N_206);
nand U1930 (N_1930,N_621,N_960);
or U1931 (N_1931,N_240,N_63);
or U1932 (N_1932,N_849,N_468);
nor U1933 (N_1933,N_673,N_807);
and U1934 (N_1934,N_53,N_598);
nor U1935 (N_1935,N_422,N_224);
or U1936 (N_1936,N_661,N_684);
or U1937 (N_1937,N_771,N_572);
or U1938 (N_1938,N_775,N_290);
nor U1939 (N_1939,N_904,N_549);
and U1940 (N_1940,N_670,N_28);
and U1941 (N_1941,N_811,N_232);
or U1942 (N_1942,N_850,N_252);
or U1943 (N_1943,N_967,N_25);
and U1944 (N_1944,N_602,N_46);
and U1945 (N_1945,N_343,N_675);
nor U1946 (N_1946,N_651,N_432);
nand U1947 (N_1947,N_536,N_694);
and U1948 (N_1948,N_994,N_956);
and U1949 (N_1949,N_944,N_654);
nand U1950 (N_1950,N_33,N_546);
and U1951 (N_1951,N_634,N_710);
nor U1952 (N_1952,N_346,N_990);
nand U1953 (N_1953,N_151,N_880);
or U1954 (N_1954,N_229,N_290);
or U1955 (N_1955,N_680,N_122);
and U1956 (N_1956,N_440,N_450);
nor U1957 (N_1957,N_116,N_836);
nand U1958 (N_1958,N_906,N_837);
and U1959 (N_1959,N_739,N_721);
and U1960 (N_1960,N_470,N_263);
nor U1961 (N_1961,N_85,N_617);
and U1962 (N_1962,N_884,N_471);
or U1963 (N_1963,N_99,N_712);
and U1964 (N_1964,N_809,N_674);
or U1965 (N_1965,N_47,N_348);
nand U1966 (N_1966,N_552,N_622);
or U1967 (N_1967,N_785,N_689);
nor U1968 (N_1968,N_23,N_116);
nor U1969 (N_1969,N_578,N_744);
and U1970 (N_1970,N_777,N_879);
xnor U1971 (N_1971,N_693,N_733);
nor U1972 (N_1972,N_585,N_391);
nand U1973 (N_1973,N_537,N_871);
or U1974 (N_1974,N_175,N_113);
or U1975 (N_1975,N_928,N_74);
nor U1976 (N_1976,N_977,N_27);
nor U1977 (N_1977,N_993,N_362);
nor U1978 (N_1978,N_229,N_949);
nor U1979 (N_1979,N_384,N_815);
or U1980 (N_1980,N_521,N_511);
nand U1981 (N_1981,N_171,N_284);
nand U1982 (N_1982,N_732,N_846);
nand U1983 (N_1983,N_287,N_250);
and U1984 (N_1984,N_689,N_167);
and U1985 (N_1985,N_731,N_471);
nand U1986 (N_1986,N_154,N_93);
nand U1987 (N_1987,N_805,N_374);
or U1988 (N_1988,N_806,N_358);
or U1989 (N_1989,N_752,N_72);
nor U1990 (N_1990,N_864,N_697);
nor U1991 (N_1991,N_617,N_604);
nor U1992 (N_1992,N_772,N_129);
nand U1993 (N_1993,N_345,N_190);
nor U1994 (N_1994,N_135,N_172);
or U1995 (N_1995,N_368,N_644);
or U1996 (N_1996,N_933,N_890);
nand U1997 (N_1997,N_471,N_779);
and U1998 (N_1998,N_374,N_286);
or U1999 (N_1999,N_365,N_358);
or U2000 (N_2000,N_1835,N_1887);
nor U2001 (N_2001,N_1191,N_1581);
and U2002 (N_2002,N_1998,N_1413);
or U2003 (N_2003,N_1931,N_1484);
or U2004 (N_2004,N_1288,N_1159);
and U2005 (N_2005,N_1181,N_1759);
or U2006 (N_2006,N_1678,N_1302);
nor U2007 (N_2007,N_1874,N_1505);
nor U2008 (N_2008,N_1824,N_1025);
nand U2009 (N_2009,N_1662,N_1008);
and U2010 (N_2010,N_1730,N_1882);
nand U2011 (N_2011,N_1431,N_1233);
or U2012 (N_2012,N_1347,N_1753);
or U2013 (N_2013,N_1775,N_1208);
nor U2014 (N_2014,N_1490,N_1984);
nor U2015 (N_2015,N_1833,N_1111);
or U2016 (N_2016,N_1647,N_1176);
or U2017 (N_2017,N_1544,N_1488);
and U2018 (N_2018,N_1661,N_1022);
nand U2019 (N_2019,N_1818,N_1764);
nor U2020 (N_2020,N_1690,N_1986);
and U2021 (N_2021,N_1628,N_1183);
nand U2022 (N_2022,N_1865,N_1018);
nor U2023 (N_2023,N_1124,N_1923);
nor U2024 (N_2024,N_1382,N_1058);
and U2025 (N_2025,N_1259,N_1851);
nor U2026 (N_2026,N_1061,N_1040);
nand U2027 (N_2027,N_1175,N_1449);
or U2028 (N_2028,N_1687,N_1305);
nand U2029 (N_2029,N_1593,N_1618);
nand U2030 (N_2030,N_1954,N_1798);
or U2031 (N_2031,N_1322,N_1781);
or U2032 (N_2032,N_1079,N_1357);
nand U2033 (N_2033,N_1763,N_1486);
or U2034 (N_2034,N_1467,N_1161);
and U2035 (N_2035,N_1979,N_1260);
nand U2036 (N_2036,N_1434,N_1335);
and U2037 (N_2037,N_1318,N_1095);
or U2038 (N_2038,N_1767,N_1749);
nor U2039 (N_2039,N_1920,N_1658);
or U2040 (N_2040,N_1837,N_1757);
nor U2041 (N_2041,N_1190,N_1027);
or U2042 (N_2042,N_1090,N_1418);
nand U2043 (N_2043,N_1209,N_1586);
and U2044 (N_2044,N_1797,N_1733);
or U2045 (N_2045,N_1212,N_1555);
nor U2046 (N_2046,N_1199,N_1068);
nor U2047 (N_2047,N_1044,N_1439);
or U2048 (N_2048,N_1359,N_1745);
or U2049 (N_2049,N_1063,N_1724);
nand U2050 (N_2050,N_1007,N_1522);
and U2051 (N_2051,N_1165,N_1067);
nand U2052 (N_2052,N_1453,N_1813);
and U2053 (N_2053,N_1584,N_1126);
or U2054 (N_2054,N_1545,N_1185);
and U2055 (N_2055,N_1683,N_1392);
and U2056 (N_2056,N_1978,N_1541);
nand U2057 (N_2057,N_1535,N_1939);
and U2058 (N_2058,N_1747,N_1228);
nand U2059 (N_2059,N_1150,N_1908);
or U2060 (N_2060,N_1346,N_1692);
nand U2061 (N_2061,N_1620,N_1670);
nand U2062 (N_2062,N_1600,N_1719);
nand U2063 (N_2063,N_1447,N_1668);
nand U2064 (N_2064,N_1677,N_1356);
nand U2065 (N_2065,N_1354,N_1187);
xor U2066 (N_2066,N_1560,N_1353);
nor U2067 (N_2067,N_1222,N_1086);
or U2068 (N_2068,N_1765,N_1870);
and U2069 (N_2069,N_1868,N_1147);
or U2070 (N_2070,N_1533,N_1846);
and U2071 (N_2071,N_1529,N_1458);
nor U2072 (N_2072,N_1223,N_1229);
nand U2073 (N_2073,N_1959,N_1031);
nor U2074 (N_2074,N_1009,N_1646);
or U2075 (N_2075,N_1799,N_1910);
or U2076 (N_2076,N_1982,N_1091);
or U2077 (N_2077,N_1784,N_1700);
nor U2078 (N_2078,N_1601,N_1475);
or U2079 (N_2079,N_1705,N_1078);
nand U2080 (N_2080,N_1549,N_1613);
and U2081 (N_2081,N_1045,N_1000);
nor U2082 (N_2082,N_1215,N_1917);
and U2083 (N_2083,N_1497,N_1950);
or U2084 (N_2084,N_1178,N_1246);
nor U2085 (N_2085,N_1239,N_1129);
nor U2086 (N_2086,N_1139,N_1242);
nor U2087 (N_2087,N_1526,N_1153);
and U2088 (N_2088,N_1904,N_1788);
nor U2089 (N_2089,N_1992,N_1831);
and U2090 (N_2090,N_1438,N_1023);
and U2091 (N_2091,N_1587,N_1213);
or U2092 (N_2092,N_1214,N_1550);
nor U2093 (N_2093,N_1862,N_1196);
and U2094 (N_2094,N_1750,N_1463);
and U2095 (N_2095,N_1743,N_1036);
or U2096 (N_2096,N_1368,N_1103);
or U2097 (N_2097,N_1961,N_1399);
and U2098 (N_2098,N_1925,N_1274);
nor U2099 (N_2099,N_1240,N_1729);
nor U2100 (N_2100,N_1388,N_1532);
or U2101 (N_2101,N_1660,N_1047);
and U2102 (N_2102,N_1930,N_1245);
and U2103 (N_2103,N_1531,N_1226);
nand U2104 (N_2104,N_1446,N_1174);
or U2105 (N_2105,N_1599,N_1442);
nand U2106 (N_2106,N_1944,N_1070);
and U2107 (N_2107,N_1460,N_1182);
and U2108 (N_2108,N_1012,N_1946);
nor U2109 (N_2109,N_1732,N_1348);
nand U2110 (N_2110,N_1366,N_1790);
nor U2111 (N_2111,N_1911,N_1097);
nand U2112 (N_2112,N_1616,N_1372);
or U2113 (N_2113,N_1207,N_1928);
xor U2114 (N_2114,N_1756,N_1666);
nand U2115 (N_2115,N_1574,N_1970);
nand U2116 (N_2116,N_1723,N_1989);
nor U2117 (N_2117,N_1496,N_1462);
and U2118 (N_2118,N_1332,N_1945);
nand U2119 (N_2119,N_1247,N_1117);
and U2120 (N_2120,N_1663,N_1643);
or U2121 (N_2121,N_1156,N_1316);
nor U2122 (N_2122,N_1268,N_1146);
or U2123 (N_2123,N_1426,N_1411);
or U2124 (N_2124,N_1594,N_1440);
and U2125 (N_2125,N_1107,N_1128);
or U2126 (N_2126,N_1282,N_1738);
nand U2127 (N_2127,N_1468,N_1610);
nand U2128 (N_2128,N_1958,N_1717);
and U2129 (N_2129,N_1679,N_1546);
nor U2130 (N_2130,N_1755,N_1115);
nand U2131 (N_2131,N_1841,N_1867);
nor U2132 (N_2132,N_1971,N_1901);
nor U2133 (N_2133,N_1471,N_1256);
nor U2134 (N_2134,N_1397,N_1514);
nand U2135 (N_2135,N_1807,N_1200);
nor U2136 (N_2136,N_1886,N_1402);
nand U2137 (N_2137,N_1029,N_1375);
nor U2138 (N_2138,N_1381,N_1404);
nand U2139 (N_2139,N_1337,N_1977);
nand U2140 (N_2140,N_1880,N_1748);
nor U2141 (N_2141,N_1433,N_1121);
nand U2142 (N_2142,N_1585,N_1850);
nor U2143 (N_2143,N_1675,N_1441);
nand U2144 (N_2144,N_1016,N_1273);
or U2145 (N_2145,N_1626,N_1391);
and U2146 (N_2146,N_1151,N_1452);
nand U2147 (N_2147,N_1605,N_1374);
nand U2148 (N_2148,N_1983,N_1590);
or U2149 (N_2149,N_1030,N_1508);
and U2150 (N_2150,N_1563,N_1639);
and U2151 (N_2151,N_1667,N_1100);
or U2152 (N_2152,N_1548,N_1427);
or U2153 (N_2153,N_1137,N_1326);
nand U2154 (N_2154,N_1843,N_1297);
and U2155 (N_2155,N_1792,N_1263);
and U2156 (N_2156,N_1480,N_1783);
nor U2157 (N_2157,N_1021,N_1448);
nor U2158 (N_2158,N_1518,N_1125);
nand U2159 (N_2159,N_1855,N_1527);
nor U2160 (N_2160,N_1949,N_1361);
and U2161 (N_2161,N_1470,N_1596);
and U2162 (N_2162,N_1665,N_1506);
nand U2163 (N_2163,N_1445,N_1564);
or U2164 (N_2164,N_1774,N_1823);
nand U2165 (N_2165,N_1644,N_1808);
nand U2166 (N_2166,N_1217,N_1154);
or U2167 (N_2167,N_1968,N_1325);
nor U2168 (N_2168,N_1580,N_1055);
nor U2169 (N_2169,N_1973,N_1157);
and U2170 (N_2170,N_1652,N_1511);
nand U2171 (N_2171,N_1845,N_1811);
nand U2172 (N_2172,N_1004,N_1052);
or U2173 (N_2173,N_1312,N_1393);
nor U2174 (N_2174,N_1281,N_1192);
nor U2175 (N_2175,N_1279,N_1951);
nor U2176 (N_2176,N_1669,N_1876);
and U2177 (N_2177,N_1019,N_1990);
nor U2178 (N_2178,N_1803,N_1524);
nand U2179 (N_2179,N_1791,N_1894);
and U2180 (N_2180,N_1889,N_1994);
nand U2181 (N_2181,N_1487,N_1349);
or U2182 (N_2182,N_1884,N_1474);
and U2183 (N_2183,N_1311,N_1503);
nor U2184 (N_2184,N_1410,N_1809);
nand U2185 (N_2185,N_1037,N_1048);
or U2186 (N_2186,N_1231,N_1712);
and U2187 (N_2187,N_1572,N_1559);
nor U2188 (N_2188,N_1686,N_1341);
and U2189 (N_2189,N_1557,N_1164);
nand U2190 (N_2190,N_1947,N_1542);
or U2191 (N_2191,N_1454,N_1144);
nand U2192 (N_2192,N_1543,N_1081);
nor U2193 (N_2193,N_1583,N_1276);
nand U2194 (N_2194,N_1500,N_1477);
and U2195 (N_2195,N_1856,N_1872);
nand U2196 (N_2196,N_1362,N_1697);
xnor U2197 (N_2197,N_1530,N_1725);
and U2198 (N_2198,N_1857,N_1822);
and U2199 (N_2199,N_1424,N_1254);
or U2200 (N_2200,N_1033,N_1266);
nand U2201 (N_2201,N_1493,N_1109);
nand U2202 (N_2202,N_1782,N_1331);
xor U2203 (N_2203,N_1751,N_1933);
nor U2204 (N_2204,N_1547,N_1345);
nand U2205 (N_2205,N_1769,N_1094);
or U2206 (N_2206,N_1011,N_1069);
or U2207 (N_2207,N_1829,N_1744);
and U2208 (N_2208,N_1976,N_1777);
and U2209 (N_2209,N_1119,N_1575);
nand U2210 (N_2210,N_1849,N_1333);
nand U2211 (N_2211,N_1272,N_1659);
or U2212 (N_2212,N_1786,N_1737);
nand U2213 (N_2213,N_1953,N_1836);
nor U2214 (N_2214,N_1172,N_1597);
and U2215 (N_2215,N_1386,N_1428);
nor U2216 (N_2216,N_1307,N_1510);
nand U2217 (N_2217,N_1234,N_1934);
nand U2218 (N_2218,N_1026,N_1980);
or U2219 (N_2219,N_1974,N_1170);
nor U2220 (N_2220,N_1376,N_1948);
nand U2221 (N_2221,N_1378,N_1017);
nor U2222 (N_2222,N_1623,N_1132);
nor U2223 (N_2223,N_1364,N_1918);
nor U2224 (N_2224,N_1568,N_1895);
xor U2225 (N_2225,N_1827,N_1414);
nand U2226 (N_2226,N_1006,N_1770);
or U2227 (N_2227,N_1221,N_1906);
nor U2228 (N_2228,N_1385,N_1878);
nand U2229 (N_2229,N_1089,N_1936);
or U2230 (N_2230,N_1203,N_1721);
or U2231 (N_2231,N_1450,N_1932);
and U2232 (N_2232,N_1010,N_1360);
nor U2233 (N_2233,N_1735,N_1625);
nand U2234 (N_2234,N_1415,N_1863);
nand U2235 (N_2235,N_1380,N_1525);
and U2236 (N_2236,N_1269,N_1056);
nand U2237 (N_2237,N_1778,N_1299);
nand U2238 (N_2238,N_1598,N_1720);
nand U2239 (N_2239,N_1145,N_1975);
nor U2240 (N_2240,N_1820,N_1236);
nand U2241 (N_2241,N_1672,N_1105);
and U2242 (N_2242,N_1840,N_1842);
nand U2243 (N_2243,N_1704,N_1334);
nor U2244 (N_2244,N_1162,N_1432);
or U2245 (N_2245,N_1141,N_1059);
or U2246 (N_2246,N_1962,N_1320);
or U2247 (N_2247,N_1379,N_1194);
and U2248 (N_2248,N_1285,N_1230);
or U2249 (N_2249,N_1520,N_1395);
and U2250 (N_2250,N_1892,N_1065);
nor U2251 (N_2251,N_1714,N_1873);
and U2252 (N_2252,N_1921,N_1869);
nor U2253 (N_2253,N_1166,N_1314);
and U2254 (N_2254,N_1812,N_1631);
or U2255 (N_2255,N_1891,N_1645);
or U2256 (N_2256,N_1796,N_1654);
nor U2257 (N_2257,N_1638,N_1177);
nand U2258 (N_2258,N_1768,N_1607);
nand U2259 (N_2259,N_1815,N_1186);
nor U2260 (N_2260,N_1996,N_1671);
nor U2261 (N_2261,N_1534,N_1567);
nor U2262 (N_2262,N_1993,N_1942);
nor U2263 (N_2263,N_1495,N_1821);
nand U2264 (N_2264,N_1123,N_1403);
and U2265 (N_2265,N_1336,N_1425);
nand U2266 (N_2266,N_1830,N_1826);
nor U2267 (N_2267,N_1800,N_1972);
or U2268 (N_2268,N_1509,N_1758);
nand U2269 (N_2269,N_1512,N_1502);
or U2270 (N_2270,N_1636,N_1429);
or U2271 (N_2271,N_1020,N_1922);
or U2272 (N_2272,N_1773,N_1401);
or U2273 (N_2273,N_1680,N_1637);
and U2274 (N_2274,N_1028,N_1198);
nand U2275 (N_2275,N_1966,N_1664);
nor U2276 (N_2276,N_1875,N_1396);
and U2277 (N_2277,N_1595,N_1848);
and U2278 (N_2278,N_1491,N_1267);
and U2279 (N_2279,N_1789,N_1417);
nand U2280 (N_2280,N_1131,N_1612);
or U2281 (N_2281,N_1472,N_1140);
or U2282 (N_2282,N_1795,N_1540);
nand U2283 (N_2283,N_1085,N_1787);
nor U2284 (N_2284,N_1801,N_1991);
and U2285 (N_2285,N_1168,N_1854);
or U2286 (N_2286,N_1113,N_1746);
nor U2287 (N_2287,N_1816,N_1709);
nor U2288 (N_2288,N_1343,N_1776);
nand U2289 (N_2289,N_1148,N_1519);
and U2290 (N_2290,N_1005,N_1630);
and U2291 (N_2291,N_1363,N_1455);
nand U2292 (N_2292,N_1571,N_1114);
and U2293 (N_2293,N_1780,N_1499);
or U2294 (N_2294,N_1814,N_1466);
nor U2295 (N_2295,N_1825,N_1451);
nand U2296 (N_2296,N_1250,N_1398);
nor U2297 (N_2297,N_1369,N_1435);
or U2298 (N_2298,N_1860,N_1469);
nand U2299 (N_2299,N_1066,N_1038);
and U2300 (N_2300,N_1309,N_1561);
or U2301 (N_2301,N_1573,N_1566);
nand U2302 (N_2302,N_1915,N_1110);
nor U2303 (N_2303,N_1400,N_1604);
nand U2304 (N_2304,N_1193,N_1112);
nor U2305 (N_2305,N_1766,N_1999);
or U2306 (N_2306,N_1219,N_1265);
nor U2307 (N_2307,N_1308,N_1804);
or U2308 (N_2308,N_1002,N_1298);
and U2309 (N_2309,N_1558,N_1576);
or U2310 (N_2310,N_1539,N_1409);
or U2311 (N_2311,N_1551,N_1722);
nand U2312 (N_2312,N_1073,N_1960);
nand U2313 (N_2313,N_1858,N_1290);
and U2314 (N_2314,N_1676,N_1352);
nor U2315 (N_2315,N_1706,N_1489);
xnor U2316 (N_2316,N_1914,N_1050);
and U2317 (N_2317,N_1853,N_1554);
nor U2318 (N_2318,N_1899,N_1762);
nor U2319 (N_2319,N_1252,N_1003);
nor U2320 (N_2320,N_1365,N_1304);
or U2321 (N_2321,N_1080,N_1286);
or U2322 (N_2322,N_1035,N_1701);
nor U2323 (N_2323,N_1955,N_1698);
and U2324 (N_2324,N_1464,N_1351);
and U2325 (N_2325,N_1528,N_1997);
nor U2326 (N_2326,N_1941,N_1935);
and U2327 (N_2327,N_1014,N_1929);
nor U2328 (N_2328,N_1189,N_1591);
or U2329 (N_2329,N_1708,N_1926);
and U2330 (N_2330,N_1118,N_1088);
nor U2331 (N_2331,N_1553,N_1339);
and U2332 (N_2332,N_1046,N_1981);
nand U2333 (N_2333,N_1909,N_1210);
nor U2334 (N_2334,N_1377,N_1578);
nor U2335 (N_2335,N_1498,N_1127);
nand U2336 (N_2336,N_1275,N_1713);
nand U2337 (N_2337,N_1405,N_1695);
and U2338 (N_2338,N_1350,N_1437);
nand U2339 (N_2339,N_1674,N_1513);
nand U2340 (N_2340,N_1741,N_1093);
nand U2341 (N_2341,N_1943,N_1479);
nand U2342 (N_2342,N_1995,N_1793);
or U2343 (N_2343,N_1054,N_1130);
xor U2344 (N_2344,N_1373,N_1293);
nor U2345 (N_2345,N_1802,N_1328);
nor U2346 (N_2346,N_1280,N_1171);
nand U2347 (N_2347,N_1456,N_1120);
nor U2348 (N_2348,N_1270,N_1552);
or U2349 (N_2349,N_1327,N_1641);
nor U2350 (N_2350,N_1443,N_1062);
nor U2351 (N_2351,N_1284,N_1060);
nand U2352 (N_2352,N_1754,N_1102);
and U2353 (N_2353,N_1682,N_1220);
or U2354 (N_2354,N_1071,N_1481);
and U2355 (N_2355,N_1742,N_1390);
nor U2356 (N_2356,N_1696,N_1883);
nand U2357 (N_2357,N_1383,N_1938);
and U2358 (N_2358,N_1394,N_1232);
or U2359 (N_2359,N_1370,N_1303);
nor U2360 (N_2360,N_1430,N_1734);
nor U2361 (N_2361,N_1206,N_1642);
nand U2362 (N_2362,N_1485,N_1785);
nand U2363 (N_2363,N_1300,N_1261);
and U2364 (N_2364,N_1913,N_1416);
or U2365 (N_2365,N_1579,N_1098);
nor U2366 (N_2366,N_1819,N_1627);
or U2367 (N_2367,N_1740,N_1963);
or U2368 (N_2368,N_1890,N_1838);
xnor U2369 (N_2369,N_1885,N_1483);
and U2370 (N_2370,N_1839,N_1294);
nand U2371 (N_2371,N_1478,N_1716);
and U2372 (N_2372,N_1122,N_1444);
nand U2373 (N_2373,N_1371,N_1204);
or U2374 (N_2374,N_1255,N_1688);
and U2375 (N_2375,N_1916,N_1707);
and U2376 (N_2376,N_1202,N_1956);
nand U2377 (N_2377,N_1847,N_1406);
nor U2378 (N_2378,N_1049,N_1728);
nor U2379 (N_2379,N_1957,N_1108);
or U2380 (N_2380,N_1051,N_1138);
and U2381 (N_2381,N_1278,N_1106);
nand U2382 (N_2382,N_1076,N_1099);
or U2383 (N_2383,N_1726,N_1650);
nor U2384 (N_2384,N_1699,N_1492);
nor U2385 (N_2385,N_1459,N_1969);
nor U2386 (N_2386,N_1609,N_1606);
and U2387 (N_2387,N_1633,N_1731);
nand U2388 (N_2388,N_1258,N_1087);
and U2389 (N_2389,N_1237,N_1898);
xnor U2390 (N_2390,N_1169,N_1521);
or U2391 (N_2391,N_1565,N_1702);
or U2392 (N_2392,N_1893,N_1201);
nor U2393 (N_2393,N_1422,N_1965);
and U2394 (N_2394,N_1834,N_1752);
and U2395 (N_2395,N_1163,N_1494);
nor U2396 (N_2396,N_1879,N_1900);
xor U2397 (N_2397,N_1864,N_1866);
nand U2398 (N_2398,N_1691,N_1589);
and U2399 (N_2399,N_1817,N_1224);
nand U2400 (N_2400,N_1152,N_1024);
and U2401 (N_2401,N_1315,N_1238);
or U2402 (N_2402,N_1727,N_1718);
nor U2403 (N_2403,N_1629,N_1216);
and U2404 (N_2404,N_1075,N_1640);
nor U2405 (N_2405,N_1501,N_1064);
nand U2406 (N_2406,N_1324,N_1101);
or U2407 (N_2407,N_1582,N_1407);
nor U2408 (N_2408,N_1227,N_1912);
nor U2409 (N_2409,N_1828,N_1461);
and U2410 (N_2410,N_1473,N_1538);
nand U2411 (N_2411,N_1158,N_1603);
or U2412 (N_2412,N_1436,N_1881);
nand U2413 (N_2413,N_1602,N_1805);
or U2414 (N_2414,N_1635,N_1985);
and U2415 (N_2415,N_1877,N_1861);
nor U2416 (N_2416,N_1632,N_1257);
and U2417 (N_2417,N_1077,N_1736);
nand U2418 (N_2418,N_1423,N_1096);
or U2419 (N_2419,N_1624,N_1218);
nor U2420 (N_2420,N_1771,N_1319);
nor U2421 (N_2421,N_1317,N_1615);
or U2422 (N_2422,N_1408,N_1907);
nand U2423 (N_2423,N_1412,N_1136);
nor U2424 (N_2424,N_1251,N_1330);
nand U2425 (N_2425,N_1384,N_1358);
or U2426 (N_2426,N_1072,N_1355);
and U2427 (N_2427,N_1180,N_1241);
and U2428 (N_2428,N_1634,N_1173);
nand U2429 (N_2429,N_1211,N_1032);
xnor U2430 (N_2430,N_1287,N_1244);
nand U2431 (N_2431,N_1516,N_1367);
nand U2432 (N_2432,N_1689,N_1457);
nor U2433 (N_2433,N_1041,N_1556);
and U2434 (N_2434,N_1937,N_1619);
nor U2435 (N_2435,N_1262,N_1592);
nor U2436 (N_2436,N_1897,N_1482);
or U2437 (N_2437,N_1015,N_1684);
and U2438 (N_2438,N_1536,N_1082);
nor U2439 (N_2439,N_1042,N_1651);
nand U2440 (N_2440,N_1249,N_1243);
nand U2441 (N_2441,N_1179,N_1656);
or U2442 (N_2442,N_1517,N_1084);
nor U2443 (N_2443,N_1739,N_1905);
and U2444 (N_2444,N_1611,N_1338);
nor U2445 (N_2445,N_1760,N_1142);
and U2446 (N_2446,N_1655,N_1340);
nand U2447 (N_2447,N_1859,N_1092);
nand U2448 (N_2448,N_1420,N_1653);
or U2449 (N_2449,N_1155,N_1621);
or U2450 (N_2450,N_1283,N_1924);
or U2451 (N_2451,N_1083,N_1039);
and U2452 (N_2452,N_1988,N_1761);
and U2453 (N_2453,N_1323,N_1135);
nand U2454 (N_2454,N_1964,N_1710);
or U2455 (N_2455,N_1577,N_1034);
or U2456 (N_2456,N_1149,N_1648);
or U2457 (N_2457,N_1306,N_1888);
and U2458 (N_2458,N_1188,N_1225);
and U2459 (N_2459,N_1507,N_1344);
and U2460 (N_2460,N_1329,N_1523);
and U2461 (N_2461,N_1342,N_1184);
nand U2462 (N_2462,N_1504,N_1074);
or U2463 (N_2463,N_1711,N_1053);
and U2464 (N_2464,N_1608,N_1001);
nor U2465 (N_2465,N_1515,N_1235);
or U2466 (N_2466,N_1617,N_1321);
and U2467 (N_2467,N_1537,N_1419);
and U2468 (N_2468,N_1927,N_1703);
or U2469 (N_2469,N_1562,N_1143);
nand U2470 (N_2470,N_1779,N_1794);
nor U2471 (N_2471,N_1871,N_1104);
and U2472 (N_2472,N_1902,N_1271);
nor U2473 (N_2473,N_1310,N_1614);
nand U2474 (N_2474,N_1952,N_1253);
or U2475 (N_2475,N_1476,N_1622);
and U2476 (N_2476,N_1301,N_1810);
and U2477 (N_2477,N_1296,N_1570);
nor U2478 (N_2478,N_1292,N_1133);
and U2479 (N_2479,N_1919,N_1013);
nand U2480 (N_2480,N_1673,N_1772);
nand U2481 (N_2481,N_1057,N_1195);
or U2482 (N_2482,N_1313,N_1387);
and U2483 (N_2483,N_1569,N_1806);
and U2484 (N_2484,N_1197,N_1160);
and U2485 (N_2485,N_1649,N_1852);
and U2486 (N_2486,N_1940,N_1291);
and U2487 (N_2487,N_1896,N_1465);
nand U2488 (N_2488,N_1264,N_1277);
nor U2489 (N_2489,N_1588,N_1693);
nand U2490 (N_2490,N_1832,N_1167);
nand U2491 (N_2491,N_1205,N_1694);
nor U2492 (N_2492,N_1715,N_1657);
or U2493 (N_2493,N_1116,N_1421);
and U2494 (N_2494,N_1134,N_1987);
and U2495 (N_2495,N_1043,N_1903);
and U2496 (N_2496,N_1685,N_1295);
nand U2497 (N_2497,N_1967,N_1389);
nand U2498 (N_2498,N_1681,N_1844);
and U2499 (N_2499,N_1248,N_1289);
or U2500 (N_2500,N_1592,N_1587);
and U2501 (N_2501,N_1029,N_1899);
nor U2502 (N_2502,N_1399,N_1576);
or U2503 (N_2503,N_1803,N_1692);
nand U2504 (N_2504,N_1029,N_1437);
nor U2505 (N_2505,N_1078,N_1884);
nand U2506 (N_2506,N_1983,N_1667);
and U2507 (N_2507,N_1355,N_1673);
nand U2508 (N_2508,N_1935,N_1598);
nor U2509 (N_2509,N_1690,N_1858);
nor U2510 (N_2510,N_1105,N_1249);
and U2511 (N_2511,N_1638,N_1680);
nor U2512 (N_2512,N_1860,N_1003);
or U2513 (N_2513,N_1329,N_1592);
or U2514 (N_2514,N_1046,N_1470);
nand U2515 (N_2515,N_1354,N_1063);
and U2516 (N_2516,N_1959,N_1162);
nor U2517 (N_2517,N_1002,N_1828);
nor U2518 (N_2518,N_1256,N_1517);
nand U2519 (N_2519,N_1609,N_1571);
nand U2520 (N_2520,N_1758,N_1594);
or U2521 (N_2521,N_1310,N_1247);
and U2522 (N_2522,N_1563,N_1108);
nor U2523 (N_2523,N_1536,N_1491);
or U2524 (N_2524,N_1309,N_1808);
and U2525 (N_2525,N_1565,N_1835);
nand U2526 (N_2526,N_1626,N_1646);
nor U2527 (N_2527,N_1793,N_1923);
nand U2528 (N_2528,N_1429,N_1391);
and U2529 (N_2529,N_1896,N_1060);
nor U2530 (N_2530,N_1748,N_1791);
nor U2531 (N_2531,N_1137,N_1303);
and U2532 (N_2532,N_1664,N_1804);
and U2533 (N_2533,N_1533,N_1535);
nand U2534 (N_2534,N_1571,N_1963);
or U2535 (N_2535,N_1523,N_1382);
or U2536 (N_2536,N_1136,N_1331);
and U2537 (N_2537,N_1280,N_1089);
or U2538 (N_2538,N_1366,N_1844);
nor U2539 (N_2539,N_1810,N_1299);
nor U2540 (N_2540,N_1867,N_1336);
and U2541 (N_2541,N_1941,N_1700);
nor U2542 (N_2542,N_1567,N_1853);
or U2543 (N_2543,N_1953,N_1070);
nor U2544 (N_2544,N_1191,N_1185);
nor U2545 (N_2545,N_1604,N_1794);
or U2546 (N_2546,N_1540,N_1597);
and U2547 (N_2547,N_1136,N_1524);
nand U2548 (N_2548,N_1807,N_1253);
xor U2549 (N_2549,N_1481,N_1487);
nand U2550 (N_2550,N_1109,N_1914);
and U2551 (N_2551,N_1741,N_1232);
and U2552 (N_2552,N_1068,N_1259);
nand U2553 (N_2553,N_1973,N_1034);
or U2554 (N_2554,N_1160,N_1638);
nand U2555 (N_2555,N_1764,N_1156);
and U2556 (N_2556,N_1051,N_1681);
nand U2557 (N_2557,N_1334,N_1919);
or U2558 (N_2558,N_1821,N_1871);
nand U2559 (N_2559,N_1124,N_1856);
nand U2560 (N_2560,N_1295,N_1931);
nor U2561 (N_2561,N_1826,N_1781);
nand U2562 (N_2562,N_1001,N_1120);
nand U2563 (N_2563,N_1551,N_1700);
or U2564 (N_2564,N_1880,N_1503);
and U2565 (N_2565,N_1870,N_1836);
nand U2566 (N_2566,N_1671,N_1222);
or U2567 (N_2567,N_1314,N_1553);
and U2568 (N_2568,N_1721,N_1599);
nor U2569 (N_2569,N_1016,N_1343);
and U2570 (N_2570,N_1799,N_1101);
or U2571 (N_2571,N_1456,N_1989);
nor U2572 (N_2572,N_1186,N_1576);
or U2573 (N_2573,N_1044,N_1010);
or U2574 (N_2574,N_1464,N_1020);
and U2575 (N_2575,N_1252,N_1002);
or U2576 (N_2576,N_1258,N_1826);
nand U2577 (N_2577,N_1248,N_1290);
xor U2578 (N_2578,N_1944,N_1991);
and U2579 (N_2579,N_1192,N_1218);
and U2580 (N_2580,N_1982,N_1574);
or U2581 (N_2581,N_1501,N_1215);
nand U2582 (N_2582,N_1271,N_1980);
nor U2583 (N_2583,N_1623,N_1082);
nand U2584 (N_2584,N_1339,N_1921);
and U2585 (N_2585,N_1726,N_1927);
nand U2586 (N_2586,N_1030,N_1013);
nand U2587 (N_2587,N_1860,N_1487);
and U2588 (N_2588,N_1208,N_1689);
or U2589 (N_2589,N_1518,N_1891);
or U2590 (N_2590,N_1670,N_1257);
and U2591 (N_2591,N_1520,N_1569);
nand U2592 (N_2592,N_1743,N_1639);
or U2593 (N_2593,N_1584,N_1173);
and U2594 (N_2594,N_1365,N_1729);
nor U2595 (N_2595,N_1698,N_1199);
and U2596 (N_2596,N_1238,N_1787);
and U2597 (N_2597,N_1944,N_1242);
nand U2598 (N_2598,N_1663,N_1276);
nand U2599 (N_2599,N_1840,N_1120);
or U2600 (N_2600,N_1931,N_1721);
or U2601 (N_2601,N_1770,N_1011);
nand U2602 (N_2602,N_1081,N_1396);
nor U2603 (N_2603,N_1053,N_1578);
nor U2604 (N_2604,N_1354,N_1373);
nand U2605 (N_2605,N_1564,N_1952);
nand U2606 (N_2606,N_1276,N_1033);
nor U2607 (N_2607,N_1686,N_1543);
or U2608 (N_2608,N_1637,N_1728);
nand U2609 (N_2609,N_1461,N_1378);
or U2610 (N_2610,N_1798,N_1373);
nand U2611 (N_2611,N_1086,N_1140);
nor U2612 (N_2612,N_1848,N_1656);
nand U2613 (N_2613,N_1294,N_1354);
and U2614 (N_2614,N_1893,N_1568);
and U2615 (N_2615,N_1319,N_1959);
nor U2616 (N_2616,N_1047,N_1522);
nor U2617 (N_2617,N_1127,N_1424);
nor U2618 (N_2618,N_1876,N_1213);
and U2619 (N_2619,N_1948,N_1169);
nand U2620 (N_2620,N_1284,N_1217);
and U2621 (N_2621,N_1273,N_1772);
nor U2622 (N_2622,N_1317,N_1571);
and U2623 (N_2623,N_1997,N_1121);
nor U2624 (N_2624,N_1631,N_1442);
nor U2625 (N_2625,N_1183,N_1509);
and U2626 (N_2626,N_1558,N_1781);
and U2627 (N_2627,N_1720,N_1055);
or U2628 (N_2628,N_1701,N_1824);
or U2629 (N_2629,N_1278,N_1074);
nor U2630 (N_2630,N_1046,N_1132);
nor U2631 (N_2631,N_1015,N_1404);
nor U2632 (N_2632,N_1351,N_1752);
nor U2633 (N_2633,N_1885,N_1949);
and U2634 (N_2634,N_1348,N_1542);
nor U2635 (N_2635,N_1102,N_1424);
nand U2636 (N_2636,N_1382,N_1057);
or U2637 (N_2637,N_1405,N_1756);
nand U2638 (N_2638,N_1015,N_1232);
nor U2639 (N_2639,N_1213,N_1538);
or U2640 (N_2640,N_1506,N_1801);
nor U2641 (N_2641,N_1939,N_1654);
nand U2642 (N_2642,N_1881,N_1192);
and U2643 (N_2643,N_1835,N_1436);
nor U2644 (N_2644,N_1116,N_1980);
and U2645 (N_2645,N_1887,N_1947);
and U2646 (N_2646,N_1475,N_1624);
nor U2647 (N_2647,N_1801,N_1464);
or U2648 (N_2648,N_1931,N_1537);
nor U2649 (N_2649,N_1460,N_1681);
nor U2650 (N_2650,N_1361,N_1832);
or U2651 (N_2651,N_1759,N_1519);
or U2652 (N_2652,N_1014,N_1191);
nand U2653 (N_2653,N_1345,N_1228);
and U2654 (N_2654,N_1190,N_1820);
nor U2655 (N_2655,N_1371,N_1852);
or U2656 (N_2656,N_1890,N_1834);
and U2657 (N_2657,N_1638,N_1305);
or U2658 (N_2658,N_1501,N_1760);
and U2659 (N_2659,N_1571,N_1942);
or U2660 (N_2660,N_1965,N_1391);
and U2661 (N_2661,N_1795,N_1920);
and U2662 (N_2662,N_1401,N_1447);
nor U2663 (N_2663,N_1709,N_1773);
nor U2664 (N_2664,N_1110,N_1370);
or U2665 (N_2665,N_1505,N_1290);
and U2666 (N_2666,N_1051,N_1271);
or U2667 (N_2667,N_1560,N_1125);
or U2668 (N_2668,N_1551,N_1979);
nand U2669 (N_2669,N_1188,N_1950);
nor U2670 (N_2670,N_1916,N_1570);
nand U2671 (N_2671,N_1758,N_1739);
and U2672 (N_2672,N_1500,N_1417);
or U2673 (N_2673,N_1303,N_1707);
or U2674 (N_2674,N_1699,N_1260);
nor U2675 (N_2675,N_1447,N_1032);
nand U2676 (N_2676,N_1396,N_1287);
nor U2677 (N_2677,N_1608,N_1288);
or U2678 (N_2678,N_1584,N_1668);
or U2679 (N_2679,N_1566,N_1329);
and U2680 (N_2680,N_1359,N_1023);
nor U2681 (N_2681,N_1336,N_1267);
and U2682 (N_2682,N_1001,N_1614);
or U2683 (N_2683,N_1485,N_1274);
and U2684 (N_2684,N_1862,N_1000);
nand U2685 (N_2685,N_1376,N_1697);
nand U2686 (N_2686,N_1702,N_1687);
or U2687 (N_2687,N_1656,N_1426);
nand U2688 (N_2688,N_1801,N_1144);
or U2689 (N_2689,N_1900,N_1209);
nor U2690 (N_2690,N_1591,N_1557);
and U2691 (N_2691,N_1352,N_1762);
nand U2692 (N_2692,N_1781,N_1317);
or U2693 (N_2693,N_1699,N_1165);
or U2694 (N_2694,N_1882,N_1955);
or U2695 (N_2695,N_1449,N_1151);
nor U2696 (N_2696,N_1226,N_1047);
or U2697 (N_2697,N_1792,N_1088);
nand U2698 (N_2698,N_1454,N_1705);
and U2699 (N_2699,N_1950,N_1765);
or U2700 (N_2700,N_1409,N_1367);
or U2701 (N_2701,N_1664,N_1024);
nor U2702 (N_2702,N_1032,N_1714);
or U2703 (N_2703,N_1609,N_1517);
nor U2704 (N_2704,N_1598,N_1374);
nor U2705 (N_2705,N_1373,N_1352);
nand U2706 (N_2706,N_1961,N_1587);
nor U2707 (N_2707,N_1915,N_1232);
or U2708 (N_2708,N_1184,N_1299);
and U2709 (N_2709,N_1018,N_1171);
nand U2710 (N_2710,N_1375,N_1018);
nor U2711 (N_2711,N_1421,N_1708);
and U2712 (N_2712,N_1000,N_1979);
nor U2713 (N_2713,N_1101,N_1873);
nor U2714 (N_2714,N_1828,N_1080);
and U2715 (N_2715,N_1970,N_1221);
nand U2716 (N_2716,N_1754,N_1045);
and U2717 (N_2717,N_1410,N_1870);
nand U2718 (N_2718,N_1948,N_1297);
nand U2719 (N_2719,N_1594,N_1324);
nor U2720 (N_2720,N_1808,N_1105);
nand U2721 (N_2721,N_1955,N_1984);
or U2722 (N_2722,N_1251,N_1679);
nand U2723 (N_2723,N_1405,N_1937);
nand U2724 (N_2724,N_1343,N_1404);
or U2725 (N_2725,N_1869,N_1537);
nand U2726 (N_2726,N_1271,N_1921);
or U2727 (N_2727,N_1537,N_1920);
or U2728 (N_2728,N_1692,N_1784);
or U2729 (N_2729,N_1374,N_1467);
or U2730 (N_2730,N_1112,N_1668);
nand U2731 (N_2731,N_1460,N_1523);
and U2732 (N_2732,N_1287,N_1670);
nand U2733 (N_2733,N_1764,N_1126);
nand U2734 (N_2734,N_1595,N_1217);
or U2735 (N_2735,N_1562,N_1239);
or U2736 (N_2736,N_1528,N_1118);
nor U2737 (N_2737,N_1042,N_1276);
nor U2738 (N_2738,N_1560,N_1386);
and U2739 (N_2739,N_1681,N_1040);
or U2740 (N_2740,N_1762,N_1024);
nand U2741 (N_2741,N_1531,N_1110);
nor U2742 (N_2742,N_1676,N_1380);
nand U2743 (N_2743,N_1037,N_1030);
nor U2744 (N_2744,N_1164,N_1521);
or U2745 (N_2745,N_1807,N_1652);
and U2746 (N_2746,N_1467,N_1574);
nand U2747 (N_2747,N_1802,N_1539);
or U2748 (N_2748,N_1596,N_1387);
nand U2749 (N_2749,N_1872,N_1877);
and U2750 (N_2750,N_1199,N_1885);
or U2751 (N_2751,N_1498,N_1968);
nor U2752 (N_2752,N_1981,N_1958);
or U2753 (N_2753,N_1776,N_1971);
nor U2754 (N_2754,N_1310,N_1819);
nand U2755 (N_2755,N_1553,N_1811);
nor U2756 (N_2756,N_1022,N_1714);
nand U2757 (N_2757,N_1702,N_1852);
nand U2758 (N_2758,N_1368,N_1128);
and U2759 (N_2759,N_1433,N_1826);
and U2760 (N_2760,N_1214,N_1039);
nand U2761 (N_2761,N_1744,N_1458);
nor U2762 (N_2762,N_1999,N_1913);
nor U2763 (N_2763,N_1276,N_1077);
or U2764 (N_2764,N_1943,N_1384);
nand U2765 (N_2765,N_1598,N_1366);
nand U2766 (N_2766,N_1814,N_1933);
nand U2767 (N_2767,N_1867,N_1095);
or U2768 (N_2768,N_1055,N_1417);
nor U2769 (N_2769,N_1973,N_1636);
or U2770 (N_2770,N_1350,N_1213);
nor U2771 (N_2771,N_1294,N_1399);
and U2772 (N_2772,N_1777,N_1766);
and U2773 (N_2773,N_1484,N_1775);
or U2774 (N_2774,N_1074,N_1230);
nand U2775 (N_2775,N_1744,N_1451);
or U2776 (N_2776,N_1851,N_1686);
nor U2777 (N_2777,N_1991,N_1827);
nor U2778 (N_2778,N_1930,N_1933);
or U2779 (N_2779,N_1736,N_1141);
or U2780 (N_2780,N_1729,N_1170);
nand U2781 (N_2781,N_1665,N_1853);
and U2782 (N_2782,N_1004,N_1967);
and U2783 (N_2783,N_1283,N_1383);
and U2784 (N_2784,N_1102,N_1483);
nor U2785 (N_2785,N_1195,N_1634);
and U2786 (N_2786,N_1633,N_1655);
or U2787 (N_2787,N_1377,N_1986);
nand U2788 (N_2788,N_1643,N_1820);
and U2789 (N_2789,N_1539,N_1725);
and U2790 (N_2790,N_1579,N_1489);
nor U2791 (N_2791,N_1027,N_1808);
or U2792 (N_2792,N_1226,N_1729);
nand U2793 (N_2793,N_1709,N_1554);
and U2794 (N_2794,N_1375,N_1333);
or U2795 (N_2795,N_1448,N_1191);
or U2796 (N_2796,N_1836,N_1361);
and U2797 (N_2797,N_1654,N_1118);
or U2798 (N_2798,N_1638,N_1321);
nand U2799 (N_2799,N_1901,N_1551);
nor U2800 (N_2800,N_1791,N_1312);
nand U2801 (N_2801,N_1282,N_1400);
nor U2802 (N_2802,N_1595,N_1266);
nand U2803 (N_2803,N_1114,N_1230);
or U2804 (N_2804,N_1695,N_1368);
nor U2805 (N_2805,N_1219,N_1891);
and U2806 (N_2806,N_1270,N_1723);
and U2807 (N_2807,N_1789,N_1446);
or U2808 (N_2808,N_1503,N_1439);
nor U2809 (N_2809,N_1137,N_1855);
or U2810 (N_2810,N_1985,N_1243);
and U2811 (N_2811,N_1830,N_1459);
nor U2812 (N_2812,N_1315,N_1117);
nor U2813 (N_2813,N_1914,N_1673);
xor U2814 (N_2814,N_1779,N_1177);
and U2815 (N_2815,N_1815,N_1023);
and U2816 (N_2816,N_1667,N_1536);
or U2817 (N_2817,N_1757,N_1561);
or U2818 (N_2818,N_1674,N_1791);
or U2819 (N_2819,N_1633,N_1148);
and U2820 (N_2820,N_1784,N_1550);
nand U2821 (N_2821,N_1864,N_1465);
xor U2822 (N_2822,N_1102,N_1169);
nor U2823 (N_2823,N_1319,N_1806);
nor U2824 (N_2824,N_1373,N_1740);
nand U2825 (N_2825,N_1805,N_1674);
or U2826 (N_2826,N_1529,N_1319);
and U2827 (N_2827,N_1687,N_1286);
nand U2828 (N_2828,N_1155,N_1424);
and U2829 (N_2829,N_1589,N_1487);
and U2830 (N_2830,N_1256,N_1482);
and U2831 (N_2831,N_1445,N_1523);
nor U2832 (N_2832,N_1641,N_1324);
or U2833 (N_2833,N_1058,N_1911);
nand U2834 (N_2834,N_1505,N_1336);
and U2835 (N_2835,N_1776,N_1166);
and U2836 (N_2836,N_1888,N_1982);
nor U2837 (N_2837,N_1166,N_1478);
nand U2838 (N_2838,N_1289,N_1818);
nand U2839 (N_2839,N_1955,N_1028);
nand U2840 (N_2840,N_1955,N_1041);
and U2841 (N_2841,N_1504,N_1934);
nor U2842 (N_2842,N_1804,N_1827);
or U2843 (N_2843,N_1587,N_1210);
nor U2844 (N_2844,N_1285,N_1986);
and U2845 (N_2845,N_1793,N_1818);
and U2846 (N_2846,N_1021,N_1833);
or U2847 (N_2847,N_1307,N_1088);
nand U2848 (N_2848,N_1387,N_1602);
and U2849 (N_2849,N_1074,N_1835);
nand U2850 (N_2850,N_1517,N_1727);
and U2851 (N_2851,N_1780,N_1220);
nor U2852 (N_2852,N_1003,N_1930);
nor U2853 (N_2853,N_1355,N_1944);
nor U2854 (N_2854,N_1588,N_1447);
and U2855 (N_2855,N_1562,N_1826);
nor U2856 (N_2856,N_1911,N_1478);
nand U2857 (N_2857,N_1656,N_1921);
nor U2858 (N_2858,N_1892,N_1411);
and U2859 (N_2859,N_1812,N_1378);
or U2860 (N_2860,N_1350,N_1884);
and U2861 (N_2861,N_1293,N_1351);
or U2862 (N_2862,N_1123,N_1178);
or U2863 (N_2863,N_1793,N_1967);
and U2864 (N_2864,N_1926,N_1694);
or U2865 (N_2865,N_1314,N_1603);
or U2866 (N_2866,N_1521,N_1380);
nor U2867 (N_2867,N_1695,N_1269);
nand U2868 (N_2868,N_1175,N_1884);
and U2869 (N_2869,N_1211,N_1727);
or U2870 (N_2870,N_1073,N_1825);
nor U2871 (N_2871,N_1256,N_1358);
or U2872 (N_2872,N_1281,N_1116);
nand U2873 (N_2873,N_1177,N_1688);
and U2874 (N_2874,N_1174,N_1957);
nor U2875 (N_2875,N_1776,N_1099);
nor U2876 (N_2876,N_1632,N_1179);
or U2877 (N_2877,N_1166,N_1756);
nand U2878 (N_2878,N_1835,N_1971);
nand U2879 (N_2879,N_1492,N_1250);
nand U2880 (N_2880,N_1892,N_1741);
nor U2881 (N_2881,N_1178,N_1670);
and U2882 (N_2882,N_1170,N_1243);
nand U2883 (N_2883,N_1140,N_1499);
nand U2884 (N_2884,N_1351,N_1068);
nor U2885 (N_2885,N_1545,N_1231);
nor U2886 (N_2886,N_1203,N_1720);
or U2887 (N_2887,N_1798,N_1693);
and U2888 (N_2888,N_1438,N_1809);
and U2889 (N_2889,N_1053,N_1650);
nand U2890 (N_2890,N_1565,N_1242);
nand U2891 (N_2891,N_1798,N_1222);
nand U2892 (N_2892,N_1580,N_1863);
nand U2893 (N_2893,N_1933,N_1085);
nand U2894 (N_2894,N_1367,N_1227);
nor U2895 (N_2895,N_1194,N_1279);
nor U2896 (N_2896,N_1242,N_1044);
and U2897 (N_2897,N_1825,N_1324);
and U2898 (N_2898,N_1832,N_1713);
nand U2899 (N_2899,N_1769,N_1878);
and U2900 (N_2900,N_1379,N_1819);
nor U2901 (N_2901,N_1385,N_1730);
or U2902 (N_2902,N_1193,N_1859);
nor U2903 (N_2903,N_1778,N_1249);
nor U2904 (N_2904,N_1499,N_1116);
xor U2905 (N_2905,N_1559,N_1523);
nor U2906 (N_2906,N_1324,N_1075);
nand U2907 (N_2907,N_1076,N_1554);
and U2908 (N_2908,N_1167,N_1472);
and U2909 (N_2909,N_1294,N_1536);
and U2910 (N_2910,N_1961,N_1172);
or U2911 (N_2911,N_1049,N_1667);
nand U2912 (N_2912,N_1447,N_1618);
or U2913 (N_2913,N_1084,N_1976);
nand U2914 (N_2914,N_1344,N_1970);
or U2915 (N_2915,N_1706,N_1378);
nor U2916 (N_2916,N_1160,N_1114);
or U2917 (N_2917,N_1233,N_1661);
nor U2918 (N_2918,N_1964,N_1016);
nor U2919 (N_2919,N_1311,N_1985);
nand U2920 (N_2920,N_1037,N_1025);
nor U2921 (N_2921,N_1571,N_1187);
or U2922 (N_2922,N_1234,N_1631);
nand U2923 (N_2923,N_1071,N_1300);
nand U2924 (N_2924,N_1731,N_1850);
nor U2925 (N_2925,N_1759,N_1359);
nand U2926 (N_2926,N_1299,N_1490);
or U2927 (N_2927,N_1173,N_1919);
xor U2928 (N_2928,N_1211,N_1642);
nand U2929 (N_2929,N_1552,N_1774);
nor U2930 (N_2930,N_1771,N_1021);
nor U2931 (N_2931,N_1485,N_1710);
nand U2932 (N_2932,N_1897,N_1371);
nor U2933 (N_2933,N_1686,N_1196);
nor U2934 (N_2934,N_1734,N_1992);
or U2935 (N_2935,N_1209,N_1950);
or U2936 (N_2936,N_1083,N_1205);
and U2937 (N_2937,N_1723,N_1179);
nor U2938 (N_2938,N_1162,N_1334);
and U2939 (N_2939,N_1903,N_1699);
nand U2940 (N_2940,N_1749,N_1137);
nor U2941 (N_2941,N_1701,N_1334);
nand U2942 (N_2942,N_1534,N_1891);
nor U2943 (N_2943,N_1675,N_1803);
and U2944 (N_2944,N_1484,N_1887);
and U2945 (N_2945,N_1007,N_1235);
xnor U2946 (N_2946,N_1911,N_1578);
nor U2947 (N_2947,N_1845,N_1163);
and U2948 (N_2948,N_1534,N_1754);
or U2949 (N_2949,N_1784,N_1785);
nand U2950 (N_2950,N_1835,N_1341);
or U2951 (N_2951,N_1725,N_1106);
and U2952 (N_2952,N_1528,N_1596);
or U2953 (N_2953,N_1369,N_1703);
nor U2954 (N_2954,N_1685,N_1678);
nand U2955 (N_2955,N_1626,N_1287);
nor U2956 (N_2956,N_1225,N_1612);
and U2957 (N_2957,N_1063,N_1477);
nand U2958 (N_2958,N_1719,N_1830);
or U2959 (N_2959,N_1746,N_1258);
and U2960 (N_2960,N_1321,N_1888);
nor U2961 (N_2961,N_1001,N_1204);
or U2962 (N_2962,N_1163,N_1770);
nor U2963 (N_2963,N_1116,N_1088);
or U2964 (N_2964,N_1998,N_1287);
or U2965 (N_2965,N_1502,N_1530);
nor U2966 (N_2966,N_1041,N_1127);
nor U2967 (N_2967,N_1460,N_1462);
or U2968 (N_2968,N_1685,N_1356);
and U2969 (N_2969,N_1280,N_1589);
and U2970 (N_2970,N_1579,N_1701);
nor U2971 (N_2971,N_1800,N_1898);
or U2972 (N_2972,N_1394,N_1703);
or U2973 (N_2973,N_1121,N_1048);
or U2974 (N_2974,N_1370,N_1524);
nand U2975 (N_2975,N_1609,N_1670);
nand U2976 (N_2976,N_1769,N_1180);
nor U2977 (N_2977,N_1911,N_1356);
nor U2978 (N_2978,N_1756,N_1964);
nor U2979 (N_2979,N_1761,N_1983);
or U2980 (N_2980,N_1092,N_1538);
or U2981 (N_2981,N_1862,N_1325);
nor U2982 (N_2982,N_1265,N_1586);
and U2983 (N_2983,N_1613,N_1764);
nand U2984 (N_2984,N_1138,N_1892);
xnor U2985 (N_2985,N_1531,N_1489);
nor U2986 (N_2986,N_1810,N_1215);
or U2987 (N_2987,N_1080,N_1091);
nor U2988 (N_2988,N_1882,N_1454);
nand U2989 (N_2989,N_1238,N_1890);
and U2990 (N_2990,N_1302,N_1150);
nand U2991 (N_2991,N_1300,N_1481);
and U2992 (N_2992,N_1489,N_1799);
or U2993 (N_2993,N_1166,N_1926);
and U2994 (N_2994,N_1570,N_1272);
or U2995 (N_2995,N_1464,N_1294);
nor U2996 (N_2996,N_1944,N_1034);
nor U2997 (N_2997,N_1468,N_1510);
and U2998 (N_2998,N_1965,N_1217);
nor U2999 (N_2999,N_1977,N_1408);
or UO_0 (O_0,N_2513,N_2032);
and UO_1 (O_1,N_2658,N_2896);
nand UO_2 (O_2,N_2935,N_2069);
nor UO_3 (O_3,N_2694,N_2537);
or UO_4 (O_4,N_2979,N_2618);
or UO_5 (O_5,N_2597,N_2973);
nand UO_6 (O_6,N_2278,N_2053);
or UO_7 (O_7,N_2595,N_2055);
and UO_8 (O_8,N_2811,N_2028);
nand UO_9 (O_9,N_2961,N_2668);
or UO_10 (O_10,N_2713,N_2615);
or UO_11 (O_11,N_2066,N_2575);
nor UO_12 (O_12,N_2981,N_2490);
nand UO_13 (O_13,N_2628,N_2566);
nand UO_14 (O_14,N_2106,N_2315);
or UO_15 (O_15,N_2698,N_2621);
and UO_16 (O_16,N_2437,N_2962);
or UO_17 (O_17,N_2888,N_2988);
nand UO_18 (O_18,N_2378,N_2840);
or UO_19 (O_19,N_2910,N_2275);
nand UO_20 (O_20,N_2655,N_2890);
and UO_21 (O_21,N_2031,N_2281);
or UO_22 (O_22,N_2284,N_2306);
and UO_23 (O_23,N_2605,N_2602);
or UO_24 (O_24,N_2159,N_2276);
xnor UO_25 (O_25,N_2571,N_2419);
nor UO_26 (O_26,N_2849,N_2380);
or UO_27 (O_27,N_2594,N_2555);
nand UO_28 (O_28,N_2895,N_2051);
nand UO_29 (O_29,N_2416,N_2057);
or UO_30 (O_30,N_2309,N_2360);
nor UO_31 (O_31,N_2936,N_2868);
nand UO_32 (O_32,N_2090,N_2004);
or UO_33 (O_33,N_2877,N_2227);
or UO_34 (O_34,N_2706,N_2984);
nand UO_35 (O_35,N_2608,N_2785);
and UO_36 (O_36,N_2815,N_2643);
nor UO_37 (O_37,N_2287,N_2906);
nand UO_38 (O_38,N_2348,N_2806);
nor UO_39 (O_39,N_2182,N_2238);
nor UO_40 (O_40,N_2716,N_2253);
nand UO_41 (O_41,N_2146,N_2909);
and UO_42 (O_42,N_2230,N_2314);
or UO_43 (O_43,N_2781,N_2249);
nor UO_44 (O_44,N_2952,N_2383);
and UO_45 (O_45,N_2688,N_2510);
and UO_46 (O_46,N_2542,N_2019);
nand UO_47 (O_47,N_2679,N_2955);
nand UO_48 (O_48,N_2258,N_2385);
or UO_49 (O_49,N_2374,N_2234);
nor UO_50 (O_50,N_2963,N_2285);
and UO_51 (O_51,N_2394,N_2947);
nor UO_52 (O_52,N_2300,N_2659);
and UO_53 (O_53,N_2558,N_2612);
and UO_54 (O_54,N_2082,N_2439);
nor UO_55 (O_55,N_2722,N_2010);
nor UO_56 (O_56,N_2587,N_2465);
or UO_57 (O_57,N_2538,N_2012);
or UO_58 (O_58,N_2755,N_2908);
nand UO_59 (O_59,N_2593,N_2732);
or UO_60 (O_60,N_2903,N_2519);
nand UO_61 (O_61,N_2544,N_2451);
or UO_62 (O_62,N_2173,N_2350);
nand UO_63 (O_63,N_2714,N_2407);
nor UO_64 (O_64,N_2990,N_2746);
and UO_65 (O_65,N_2479,N_2289);
nand UO_66 (O_66,N_2844,N_2855);
or UO_67 (O_67,N_2393,N_2637);
xnor UO_68 (O_68,N_2837,N_2398);
and UO_69 (O_69,N_2632,N_2072);
nand UO_70 (O_70,N_2842,N_2665);
and UO_71 (O_71,N_2681,N_2183);
nand UO_72 (O_72,N_2968,N_2929);
nand UO_73 (O_73,N_2081,N_2100);
nand UO_74 (O_74,N_2241,N_2015);
and UO_75 (O_75,N_2812,N_2911);
nand UO_76 (O_76,N_2466,N_2279);
nor UO_77 (O_77,N_2550,N_2181);
nor UO_78 (O_78,N_2307,N_2945);
or UO_79 (O_79,N_2109,N_2860);
nand UO_80 (O_80,N_2491,N_2431);
nand UO_81 (O_81,N_2187,N_2196);
nor UO_82 (O_82,N_2726,N_2404);
or UO_83 (O_83,N_2740,N_2782);
or UO_84 (O_84,N_2718,N_2695);
nand UO_85 (O_85,N_2344,N_2447);
and UO_86 (O_86,N_2677,N_2273);
and UO_87 (O_87,N_2559,N_2129);
nand UO_88 (O_88,N_2789,N_2453);
and UO_89 (O_89,N_2166,N_2515);
or UO_90 (O_90,N_2891,N_2356);
nor UO_91 (O_91,N_2124,N_2867);
nor UO_92 (O_92,N_2195,N_2500);
and UO_93 (O_93,N_2369,N_2108);
nand UO_94 (O_94,N_2770,N_2017);
or UO_95 (O_95,N_2112,N_2145);
nor UO_96 (O_96,N_2531,N_2304);
and UO_97 (O_97,N_2921,N_2020);
or UO_98 (O_98,N_2156,N_2399);
or UO_99 (O_99,N_2687,N_2172);
and UO_100 (O_100,N_2636,N_2841);
and UO_101 (O_101,N_2682,N_2366);
nand UO_102 (O_102,N_2633,N_2452);
nor UO_103 (O_103,N_2678,N_2128);
or UO_104 (O_104,N_2331,N_2950);
and UO_105 (O_105,N_2590,N_2016);
nand UO_106 (O_106,N_2879,N_2684);
and UO_107 (O_107,N_2126,N_2581);
nand UO_108 (O_108,N_2846,N_2324);
nand UO_109 (O_109,N_2949,N_2268);
or UO_110 (O_110,N_2352,N_2926);
or UO_111 (O_111,N_2420,N_2556);
or UO_112 (O_112,N_2730,N_2756);
and UO_113 (O_113,N_2335,N_2354);
and UO_114 (O_114,N_2778,N_2332);
nor UO_115 (O_115,N_2574,N_2983);
nand UO_116 (O_116,N_2960,N_2074);
nor UO_117 (O_117,N_2235,N_2036);
or UO_118 (O_118,N_2430,N_2325);
or UO_119 (O_119,N_2414,N_2522);
nor UO_120 (O_120,N_2232,N_2553);
nand UO_121 (O_121,N_2613,N_2824);
or UO_122 (O_122,N_2080,N_2345);
or UO_123 (O_123,N_2303,N_2462);
or UO_124 (O_124,N_2093,N_2830);
nor UO_125 (O_125,N_2110,N_2767);
or UO_126 (O_126,N_2614,N_2362);
and UO_127 (O_127,N_2673,N_2623);
nand UO_128 (O_128,N_2599,N_2833);
nand UO_129 (O_129,N_2991,N_2798);
or UO_130 (O_130,N_2889,N_2858);
or UO_131 (O_131,N_2436,N_2246);
and UO_132 (O_132,N_2905,N_2390);
or UO_133 (O_133,N_2944,N_2337);
nand UO_134 (O_134,N_2167,N_2266);
nor UO_135 (O_135,N_2517,N_2863);
nand UO_136 (O_136,N_2835,N_2242);
nor UO_137 (O_137,N_2475,N_2153);
and UO_138 (O_138,N_2804,N_2155);
nor UO_139 (O_139,N_2922,N_2058);
xnor UO_140 (O_140,N_2790,N_2121);
or UO_141 (O_141,N_2675,N_2381);
nand UO_142 (O_142,N_2663,N_2045);
and UO_143 (O_143,N_2996,N_2271);
and UO_144 (O_144,N_2334,N_2330);
and UO_145 (O_145,N_2758,N_2191);
nand UO_146 (O_146,N_2305,N_2193);
nor UO_147 (O_147,N_2577,N_2715);
and UO_148 (O_148,N_2799,N_2788);
nor UO_149 (O_149,N_2464,N_2083);
and UO_150 (O_150,N_2854,N_2367);
nand UO_151 (O_151,N_2711,N_2839);
nand UO_152 (O_152,N_2070,N_2986);
or UO_153 (O_153,N_2697,N_2073);
nor UO_154 (O_154,N_2586,N_2987);
nand UO_155 (O_155,N_2161,N_2493);
nand UO_156 (O_156,N_2967,N_2138);
and UO_157 (O_157,N_2099,N_2619);
and UO_158 (O_158,N_2104,N_2794);
or UO_159 (O_159,N_2122,N_2934);
nor UO_160 (O_160,N_2939,N_2180);
and UO_161 (O_161,N_2818,N_2027);
nor UO_162 (O_162,N_2805,N_2223);
or UO_163 (O_163,N_2518,N_2079);
or UO_164 (O_164,N_2511,N_2194);
or UO_165 (O_165,N_2030,N_2410);
or UO_166 (O_166,N_2208,N_2293);
nand UO_167 (O_167,N_2876,N_2213);
or UO_168 (O_168,N_2872,N_2894);
or UO_169 (O_169,N_2139,N_2443);
and UO_170 (O_170,N_2470,N_2568);
and UO_171 (O_171,N_2954,N_2002);
xor UO_172 (O_172,N_2919,N_2064);
or UO_173 (O_173,N_2869,N_2469);
nor UO_174 (O_174,N_2282,N_2429);
or UO_175 (O_175,N_2918,N_2257);
and UO_176 (O_176,N_2759,N_2168);
nand UO_177 (O_177,N_2251,N_2904);
nand UO_178 (O_178,N_2657,N_2664);
or UO_179 (O_179,N_2426,N_2338);
or UO_180 (O_180,N_2527,N_2137);
or UO_181 (O_181,N_2739,N_2297);
or UO_182 (O_182,N_2907,N_2813);
nor UO_183 (O_183,N_2576,N_2084);
nand UO_184 (O_184,N_2496,N_2188);
and UO_185 (O_185,N_2319,N_2499);
nor UO_186 (O_186,N_2993,N_2358);
nand UO_187 (O_187,N_2578,N_2528);
nor UO_188 (O_188,N_2737,N_2545);
nand UO_189 (O_189,N_2006,N_2492);
and UO_190 (O_190,N_2205,N_2065);
and UO_191 (O_191,N_2603,N_2512);
nand UO_192 (O_192,N_2088,N_2202);
nor UO_193 (O_193,N_2260,N_2320);
or UO_194 (O_194,N_2539,N_2647);
and UO_195 (O_195,N_2717,N_2976);
or UO_196 (O_196,N_2047,N_2371);
nand UO_197 (O_197,N_2389,N_2119);
nor UO_198 (O_198,N_2765,N_2728);
nand UO_199 (O_199,N_2724,N_2795);
and UO_200 (O_200,N_2397,N_2572);
nand UO_201 (O_201,N_2580,N_2977);
nor UO_202 (O_202,N_2411,N_2913);
nand UO_203 (O_203,N_2827,N_2440);
or UO_204 (O_204,N_2783,N_2834);
nand UO_205 (O_205,N_2843,N_2434);
and UO_206 (O_206,N_2741,N_2086);
and UO_207 (O_207,N_2828,N_2206);
or UO_208 (O_208,N_2766,N_2541);
and UO_209 (O_209,N_2482,N_2822);
and UO_210 (O_210,N_2725,N_2772);
nand UO_211 (O_211,N_2263,N_2920);
nor UO_212 (O_212,N_2685,N_2807);
and UO_213 (O_213,N_2269,N_2900);
or UO_214 (O_214,N_2120,N_2485);
nand UO_215 (O_215,N_2561,N_2630);
nand UO_216 (O_216,N_2532,N_2209);
and UO_217 (O_217,N_2240,N_2745);
or UO_218 (O_218,N_2588,N_2933);
or UO_219 (O_219,N_2005,N_2095);
or UO_220 (O_220,N_2417,N_2925);
xnor UO_221 (O_221,N_2771,N_2326);
and UO_222 (O_222,N_2308,N_2113);
nor UO_223 (O_223,N_2038,N_2940);
and UO_224 (O_224,N_2671,N_2132);
nor UO_225 (O_225,N_2874,N_2884);
nand UO_226 (O_226,N_2856,N_2007);
or UO_227 (O_227,N_2264,N_2642);
nor UO_228 (O_228,N_2583,N_2731);
and UO_229 (O_229,N_2892,N_2916);
and UO_230 (O_230,N_2964,N_2547);
and UO_231 (O_231,N_2025,N_2768);
and UO_232 (O_232,N_2254,N_2185);
and UO_233 (O_233,N_2301,N_2762);
nand UO_234 (O_234,N_2942,N_2078);
or UO_235 (O_235,N_2042,N_2102);
nor UO_236 (O_236,N_2503,N_2226);
nand UO_237 (O_237,N_2565,N_2956);
and UO_238 (O_238,N_2525,N_2409);
nand UO_239 (O_239,N_2401,N_2640);
and UO_240 (O_240,N_2885,N_2814);
and UO_241 (O_241,N_2870,N_2039);
or UO_242 (O_242,N_2857,N_2564);
and UO_243 (O_243,N_2601,N_2329);
nor UO_244 (O_244,N_2862,N_2123);
and UO_245 (O_245,N_2433,N_2915);
and UO_246 (O_246,N_2415,N_2985);
and UO_247 (O_247,N_2852,N_2476);
nor UO_248 (O_248,N_2158,N_2382);
xnor UO_249 (O_249,N_2290,N_2948);
nand UO_250 (O_250,N_2402,N_2277);
or UO_251 (O_251,N_2753,N_2554);
or UO_252 (O_252,N_2085,N_2261);
nor UO_253 (O_253,N_2483,N_2091);
or UO_254 (O_254,N_2957,N_2622);
nand UO_255 (O_255,N_2062,N_2327);
and UO_256 (O_256,N_2710,N_2097);
nor UO_257 (O_257,N_2259,N_2592);
nor UO_258 (O_258,N_2162,N_2970);
and UO_259 (O_259,N_2170,N_2076);
nand UO_260 (O_260,N_2584,N_2149);
nor UO_261 (O_261,N_2611,N_2738);
nand UO_262 (O_262,N_2562,N_2917);
or UO_263 (O_263,N_2456,N_2228);
nor UO_264 (O_264,N_2727,N_2821);
xnor UO_265 (O_265,N_2011,N_2328);
or UO_266 (O_266,N_2792,N_2971);
and UO_267 (O_267,N_2626,N_2060);
nand UO_268 (O_268,N_2982,N_2040);
nor UO_269 (O_269,N_2089,N_2959);
nor UO_270 (O_270,N_2477,N_2777);
and UO_271 (O_271,N_2200,N_2620);
nand UO_272 (O_272,N_2901,N_2178);
or UO_273 (O_273,N_2169,N_2992);
nor UO_274 (O_274,N_2924,N_2820);
and UO_275 (O_275,N_2219,N_2067);
nor UO_276 (O_276,N_2514,N_2686);
or UO_277 (O_277,N_2125,N_2680);
and UO_278 (O_278,N_2816,N_2467);
nor UO_279 (O_279,N_2676,N_2107);
nor UO_280 (O_280,N_2377,N_2364);
and UO_281 (O_281,N_2489,N_2265);
nor UO_282 (O_282,N_2442,N_2585);
nor UO_283 (O_283,N_2373,N_2598);
nand UO_284 (O_284,N_2201,N_2650);
nor UO_285 (O_285,N_2270,N_2472);
or UO_286 (O_286,N_2233,N_2231);
or UO_287 (O_287,N_2444,N_2495);
nor UO_288 (O_288,N_2152,N_2184);
nand UO_289 (O_289,N_2151,N_2405);
or UO_290 (O_290,N_2481,N_2056);
and UO_291 (O_291,N_2627,N_2368);
and UO_292 (O_292,N_2931,N_2523);
nor UO_293 (O_293,N_2848,N_2203);
and UO_294 (O_294,N_2291,N_2351);
or UO_295 (O_295,N_2347,N_2098);
and UO_296 (O_296,N_2133,N_2413);
or UO_297 (O_297,N_2438,N_2432);
and UO_298 (O_298,N_2721,N_2927);
nand UO_299 (O_299,N_2312,N_2733);
or UO_300 (O_300,N_2311,N_2551);
or UO_301 (O_301,N_2761,N_2346);
or UO_302 (O_302,N_2563,N_2418);
and UO_303 (O_303,N_2878,N_2336);
nor UO_304 (O_304,N_2535,N_2379);
nor UO_305 (O_305,N_2365,N_2930);
nand UO_306 (O_306,N_2372,N_2403);
and UO_307 (O_307,N_2310,N_2582);
and UO_308 (O_308,N_2210,N_2013);
or UO_309 (O_309,N_2700,N_2645);
nor UO_310 (O_310,N_2247,N_2333);
or UO_311 (O_311,N_2825,N_2355);
or UO_312 (O_312,N_2829,N_2395);
nand UO_313 (O_313,N_2009,N_2609);
or UO_314 (O_314,N_2897,N_2160);
and UO_315 (O_315,N_2589,N_2239);
and UO_316 (O_316,N_2480,N_2422);
and UO_317 (O_317,N_2744,N_2809);
and UO_318 (O_318,N_2061,N_2946);
nor UO_319 (O_319,N_2130,N_2604);
and UO_320 (O_320,N_2243,N_2534);
and UO_321 (O_321,N_2579,N_2787);
nor UO_322 (O_322,N_2596,N_2667);
and UO_323 (O_323,N_2021,N_2177);
and UO_324 (O_324,N_2723,N_2148);
and UO_325 (O_325,N_2494,N_2498);
or UO_326 (O_326,N_2649,N_2092);
nand UO_327 (O_327,N_2995,N_2754);
and UO_328 (O_328,N_2902,N_2644);
nand UO_329 (O_329,N_2546,N_2478);
nor UO_330 (O_330,N_2190,N_2353);
nand UO_331 (O_331,N_2068,N_2670);
nand UO_332 (O_332,N_2701,N_2176);
nand UO_333 (O_333,N_2008,N_2428);
and UO_334 (O_334,N_2220,N_2425);
nor UO_335 (O_335,N_2784,N_2204);
nor UO_336 (O_336,N_2704,N_2468);
nor UO_337 (O_337,N_2115,N_2859);
and UO_338 (O_338,N_2656,N_2286);
nor UO_339 (O_339,N_2163,N_2454);
or UO_340 (O_340,N_2928,N_2459);
nor UO_341 (O_341,N_2318,N_2317);
nand UO_342 (O_342,N_2029,N_2506);
nand UO_343 (O_343,N_2880,N_2140);
nand UO_344 (O_344,N_2215,N_2875);
nor UO_345 (O_345,N_2629,N_2225);
and UO_346 (O_346,N_2421,N_2752);
nor UO_347 (O_347,N_2999,N_2702);
nand UO_348 (O_348,N_2502,N_2101);
or UO_349 (O_349,N_2445,N_2054);
or UO_350 (O_350,N_2886,N_2625);
nand UO_351 (O_351,N_2764,N_2250);
and UO_352 (O_352,N_2387,N_2526);
nand UO_353 (O_353,N_2046,N_2646);
and UO_354 (O_354,N_2631,N_2861);
and UO_355 (O_355,N_2024,N_2262);
nand UO_356 (O_356,N_2543,N_2197);
or UO_357 (O_357,N_2361,N_2131);
or UO_358 (O_358,N_2157,N_2189);
nand UO_359 (O_359,N_2866,N_2096);
nand UO_360 (O_360,N_2689,N_2832);
nor UO_361 (O_361,N_2899,N_2836);
nor UO_362 (O_362,N_2192,N_2457);
and UO_363 (O_363,N_2461,N_2801);
or UO_364 (O_364,N_2703,N_2034);
nor UO_365 (O_365,N_2014,N_2463);
nand UO_366 (O_366,N_2980,N_2396);
xor UO_367 (O_367,N_2607,N_2557);
nor UO_368 (O_368,N_2295,N_2274);
nor UO_369 (O_369,N_2026,N_2323);
nor UO_370 (O_370,N_2450,N_2117);
nor UO_371 (O_371,N_2864,N_2288);
and UO_372 (O_372,N_2530,N_2865);
nand UO_373 (O_373,N_2750,N_2573);
nand UO_374 (O_374,N_2978,N_2696);
nand UO_375 (O_375,N_2516,N_2560);
nand UO_376 (O_376,N_2652,N_2882);
nand UO_377 (O_377,N_2487,N_2474);
nor UO_378 (O_378,N_2256,N_2552);
nand UO_379 (O_379,N_2171,N_2743);
or UO_380 (O_380,N_2313,N_2033);
nor UO_381 (O_381,N_2218,N_2616);
nor UO_382 (O_382,N_2236,N_2229);
nand UO_383 (O_383,N_2118,N_2244);
nor UO_384 (O_384,N_2932,N_2536);
and UO_385 (O_385,N_2606,N_2810);
or UO_386 (O_386,N_2388,N_2823);
xor UO_387 (O_387,N_2691,N_2143);
nor UO_388 (O_388,N_2893,N_2742);
nand UO_389 (O_389,N_2179,N_2797);
nor UO_390 (O_390,N_2683,N_2449);
or UO_391 (O_391,N_2796,N_2283);
nor UO_392 (O_392,N_2342,N_2591);
nand UO_393 (O_393,N_2063,N_2105);
nand UO_394 (O_394,N_2570,N_2847);
or UO_395 (O_395,N_2298,N_2941);
or UO_396 (O_396,N_2567,N_2653);
nor UO_397 (O_397,N_2363,N_2509);
and UO_398 (O_398,N_2111,N_2776);
nor UO_399 (O_399,N_2540,N_2504);
and UO_400 (O_400,N_2803,N_2974);
nor UO_401 (O_401,N_2255,N_2791);
or UO_402 (O_402,N_2408,N_2938);
or UO_403 (O_403,N_2779,N_2898);
and UO_404 (O_404,N_2497,N_2359);
and UO_405 (O_405,N_2001,N_2617);
nand UO_406 (O_406,N_2052,N_2141);
and UO_407 (O_407,N_2669,N_2690);
nor UO_408 (O_408,N_2116,N_2624);
nand UO_409 (O_409,N_2951,N_2881);
nor UO_410 (O_410,N_2224,N_2077);
and UO_411 (O_411,N_2272,N_2760);
or UO_412 (O_412,N_2958,N_2969);
or UO_413 (O_413,N_2639,N_2769);
and UO_414 (O_414,N_2709,N_2887);
nor UO_415 (O_415,N_2424,N_2712);
and UO_416 (O_416,N_2448,N_2774);
nor UO_417 (O_417,N_2252,N_2569);
nor UO_418 (O_418,N_2041,N_2147);
or UO_419 (O_419,N_2075,N_2059);
nor UO_420 (O_420,N_2018,N_2455);
nand UO_421 (O_421,N_2267,N_2049);
or UO_422 (O_422,N_2292,N_2343);
xnor UO_423 (O_423,N_2747,N_2994);
and UO_424 (O_424,N_2349,N_2023);
nand UO_425 (O_425,N_2549,N_2548);
nand UO_426 (O_426,N_2850,N_2071);
nand UO_427 (O_427,N_2094,N_2734);
or UO_428 (O_428,N_2635,N_2989);
and UO_429 (O_429,N_2237,N_2521);
or UO_430 (O_430,N_2186,N_2871);
nand UO_431 (O_431,N_2175,N_2763);
nand UO_432 (O_432,N_2873,N_2127);
or UO_433 (O_433,N_2699,N_2294);
or UO_434 (O_434,N_2486,N_2207);
nor UO_435 (O_435,N_2370,N_2674);
nor UO_436 (O_436,N_2114,N_2035);
nand UO_437 (O_437,N_2198,N_2638);
and UO_438 (O_438,N_2458,N_2000);
nand UO_439 (O_439,N_2507,N_2087);
and UO_440 (O_440,N_2446,N_2641);
xnor UO_441 (O_441,N_2488,N_2022);
or UO_442 (O_442,N_2524,N_2386);
nand UO_443 (O_443,N_2838,N_2953);
nand UO_444 (O_444,N_2600,N_2221);
and UO_445 (O_445,N_2817,N_2692);
and UO_446 (O_446,N_2441,N_2757);
nand UO_447 (O_447,N_2044,N_2912);
nor UO_448 (O_448,N_2966,N_2853);
or UO_449 (O_449,N_2460,N_2248);
nor UO_450 (O_450,N_2997,N_2634);
and UO_451 (O_451,N_2375,N_2322);
and UO_452 (O_452,N_2735,N_2357);
or UO_453 (O_453,N_2245,N_2412);
nor UO_454 (O_454,N_2484,N_2341);
or UO_455 (O_455,N_2043,N_2937);
or UO_456 (O_456,N_2501,N_2705);
or UO_457 (O_457,N_2780,N_2340);
nor UO_458 (O_458,N_2707,N_2654);
nand UO_459 (O_459,N_2217,N_2975);
nor UO_460 (O_460,N_2773,N_2529);
nand UO_461 (O_461,N_2214,N_2222);
nor UO_462 (O_462,N_2662,N_2648);
nor UO_463 (O_463,N_2296,N_2651);
or UO_464 (O_464,N_2391,N_2520);
and UO_465 (O_465,N_2508,N_2914);
and UO_466 (O_466,N_2693,N_2533);
and UO_467 (O_467,N_2923,N_2819);
or UO_468 (O_468,N_2831,N_2708);
nor UO_469 (O_469,N_2719,N_2199);
and UO_470 (O_470,N_2661,N_2666);
or UO_471 (O_471,N_2749,N_2406);
xor UO_472 (O_472,N_2384,N_2165);
nand UO_473 (O_473,N_2376,N_2392);
and UO_474 (O_474,N_2216,N_2473);
nand UO_475 (O_475,N_2775,N_2505);
nand UO_476 (O_476,N_2150,N_2660);
nand UO_477 (O_477,N_2802,N_2321);
or UO_478 (O_478,N_2050,N_2003);
and UO_479 (O_479,N_2048,N_2212);
nand UO_480 (O_480,N_2299,N_2793);
nor UO_481 (O_481,N_2965,N_2103);
nand UO_482 (O_482,N_2427,N_2423);
nor UO_483 (O_483,N_2972,N_2610);
or UO_484 (O_484,N_2729,N_2164);
nor UO_485 (O_485,N_2174,N_2471);
nor UO_486 (O_486,N_2154,N_2845);
or UO_487 (O_487,N_2736,N_2943);
nor UO_488 (O_488,N_2435,N_2851);
nand UO_489 (O_489,N_2808,N_2998);
or UO_490 (O_490,N_2134,N_2720);
or UO_491 (O_491,N_2144,N_2672);
or UO_492 (O_492,N_2142,N_2400);
or UO_493 (O_493,N_2883,N_2302);
and UO_494 (O_494,N_2316,N_2211);
nor UO_495 (O_495,N_2037,N_2748);
nand UO_496 (O_496,N_2751,N_2800);
nand UO_497 (O_497,N_2826,N_2786);
nand UO_498 (O_498,N_2339,N_2135);
and UO_499 (O_499,N_2280,N_2136);
endmodule