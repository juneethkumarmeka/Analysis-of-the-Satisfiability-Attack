module basic_2500_25000_3000_25_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1466,In_978);
and U1 (N_1,In_364,In_183);
xnor U2 (N_2,In_1632,In_475);
nand U3 (N_3,In_2108,In_1526);
or U4 (N_4,In_1273,In_1087);
nor U5 (N_5,In_1563,In_1177);
nor U6 (N_6,In_1763,In_1794);
and U7 (N_7,In_506,In_2249);
nand U8 (N_8,In_1703,In_1025);
nand U9 (N_9,In_335,In_739);
and U10 (N_10,In_1646,In_431);
or U11 (N_11,In_1109,In_2089);
xor U12 (N_12,In_2184,In_1508);
and U13 (N_13,In_1651,In_10);
and U14 (N_14,In_2119,In_835);
and U15 (N_15,In_952,In_1486);
or U16 (N_16,In_1394,In_484);
or U17 (N_17,In_1501,In_729);
or U18 (N_18,In_2407,In_2278);
nand U19 (N_19,In_512,In_1185);
nor U20 (N_20,In_1635,In_2176);
nand U21 (N_21,In_1275,In_55);
and U22 (N_22,In_1941,In_2167);
nand U23 (N_23,In_1708,In_1055);
nor U24 (N_24,In_1931,In_683);
xor U25 (N_25,In_360,In_1731);
nor U26 (N_26,In_947,In_1347);
or U27 (N_27,In_1599,In_1584);
nand U28 (N_28,In_949,In_2396);
xor U29 (N_29,In_1863,In_1869);
and U30 (N_30,In_912,In_375);
nand U31 (N_31,In_922,In_1135);
xnor U32 (N_32,In_444,In_2145);
or U33 (N_33,In_1764,In_2292);
nand U34 (N_34,In_1525,In_1193);
or U35 (N_35,In_1441,In_118);
and U36 (N_36,In_2406,In_1798);
nand U37 (N_37,In_1366,In_871);
and U38 (N_38,In_1982,In_1494);
nor U39 (N_39,In_2455,In_1044);
nand U40 (N_40,In_1701,In_2281);
and U41 (N_41,In_1289,In_1858);
nor U42 (N_42,In_268,In_2231);
and U43 (N_43,In_388,In_1290);
nand U44 (N_44,In_1677,In_779);
xnor U45 (N_45,In_1180,In_1113);
or U46 (N_46,In_393,In_325);
and U47 (N_47,In_796,In_2188);
nor U48 (N_48,In_1740,In_322);
nand U49 (N_49,In_1242,In_942);
and U50 (N_50,In_896,In_414);
nand U51 (N_51,In_321,In_2456);
and U52 (N_52,In_792,In_1224);
nand U53 (N_53,In_1880,In_427);
and U54 (N_54,In_873,In_1364);
and U55 (N_55,In_1000,In_409);
nor U56 (N_56,In_305,In_878);
and U57 (N_57,In_361,In_1700);
or U58 (N_58,In_1848,In_1970);
or U59 (N_59,In_1483,In_433);
xor U60 (N_60,In_1714,In_1755);
or U61 (N_61,In_446,In_1234);
nor U62 (N_62,In_2172,In_869);
or U63 (N_63,In_395,In_892);
or U64 (N_64,In_2158,In_521);
or U65 (N_65,In_279,In_2387);
nand U66 (N_66,In_522,In_1996);
or U67 (N_67,In_1168,In_139);
nor U68 (N_68,In_254,In_1213);
or U69 (N_69,In_738,In_1747);
nor U70 (N_70,In_1205,In_1784);
nor U71 (N_71,In_2354,In_2006);
or U72 (N_72,In_1326,In_2484);
nor U73 (N_73,In_591,In_790);
nand U74 (N_74,In_938,In_1121);
nor U75 (N_75,In_752,In_0);
and U76 (N_76,In_1175,In_1925);
and U77 (N_77,In_1521,In_543);
xor U78 (N_78,In_1450,In_1407);
nand U79 (N_79,In_732,In_2225);
nand U80 (N_80,In_2326,In_1081);
and U81 (N_81,In_1595,In_718);
nor U82 (N_82,In_158,In_1197);
or U83 (N_83,In_1690,In_596);
and U84 (N_84,In_1116,In_2129);
xnor U85 (N_85,In_92,In_552);
xnor U86 (N_86,In_316,In_1742);
nand U87 (N_87,In_2029,In_1128);
nand U88 (N_88,In_1155,In_1598);
or U89 (N_89,In_163,In_728);
xnor U90 (N_90,In_1955,In_178);
and U91 (N_91,In_2319,In_1828);
nand U92 (N_92,In_2171,In_228);
nand U93 (N_93,In_1164,In_2163);
xnor U94 (N_94,In_888,In_1459);
and U95 (N_95,In_1513,In_2223);
nand U96 (N_96,In_197,In_2051);
nor U97 (N_97,In_966,In_2136);
or U98 (N_98,In_2007,In_905);
and U99 (N_99,In_781,In_22);
xor U100 (N_100,In_571,In_2018);
and U101 (N_101,In_1382,In_2327);
or U102 (N_102,In_598,In_109);
nand U103 (N_103,In_944,In_1829);
xor U104 (N_104,In_317,In_2118);
and U105 (N_105,In_667,In_2203);
nor U106 (N_106,In_1593,In_644);
xor U107 (N_107,In_1178,In_222);
nor U108 (N_108,In_1043,In_483);
nor U109 (N_109,In_631,In_273);
and U110 (N_110,In_945,In_1069);
nor U111 (N_111,In_899,In_1360);
nor U112 (N_112,In_25,In_362);
and U113 (N_113,In_1605,In_894);
nor U114 (N_114,In_2426,In_685);
and U115 (N_115,In_1088,In_1604);
nand U116 (N_116,In_1047,In_73);
nor U117 (N_117,In_2181,In_62);
nor U118 (N_118,In_380,In_2344);
or U119 (N_119,In_1801,In_1937);
nor U120 (N_120,In_489,In_1367);
nand U121 (N_121,In_1356,In_2028);
nor U122 (N_122,In_2334,In_255);
and U123 (N_123,In_1301,In_1350);
xnor U124 (N_124,In_374,In_2341);
nor U125 (N_125,In_2222,In_987);
or U126 (N_126,In_1916,In_150);
and U127 (N_127,In_840,In_2097);
nor U128 (N_128,In_2338,In_177);
and U129 (N_129,In_2421,In_516);
nor U130 (N_130,In_459,In_89);
nor U131 (N_131,In_784,In_1500);
or U132 (N_132,In_440,In_580);
nand U133 (N_133,In_960,In_159);
or U134 (N_134,In_384,In_555);
nand U135 (N_135,In_624,In_1669);
nor U136 (N_136,In_1706,In_2275);
xor U137 (N_137,In_2415,In_138);
nor U138 (N_138,In_2348,In_2293);
and U139 (N_139,In_1137,In_519);
or U140 (N_140,In_2159,In_1219);
nor U141 (N_141,In_520,In_579);
nor U142 (N_142,In_885,In_272);
xor U143 (N_143,In_324,In_2068);
xnor U144 (N_144,In_697,In_2198);
nand U145 (N_145,In_1733,In_303);
or U146 (N_146,In_1998,In_2195);
nor U147 (N_147,In_1924,In_396);
and U148 (N_148,In_1940,In_2112);
nor U149 (N_149,In_1556,In_1420);
nand U150 (N_150,In_2322,In_1934);
and U151 (N_151,In_680,In_494);
nor U152 (N_152,In_2234,In_2059);
xor U153 (N_153,In_1533,In_1215);
or U154 (N_154,In_1893,In_2049);
nor U155 (N_155,In_929,In_400);
and U156 (N_156,In_548,In_1030);
nand U157 (N_157,In_2117,In_1165);
nand U158 (N_158,In_2185,In_654);
or U159 (N_159,In_907,In_1460);
nor U160 (N_160,In_1298,In_1307);
or U161 (N_161,In_1012,In_2120);
nor U162 (N_162,In_2080,In_1082);
nand U163 (N_163,In_1552,In_202);
nor U164 (N_164,In_1102,In_587);
or U165 (N_165,In_973,In_2194);
nor U166 (N_166,In_2017,In_932);
or U167 (N_167,In_712,In_1850);
and U168 (N_168,In_788,In_1833);
nor U169 (N_169,In_1663,In_1373);
nand U170 (N_170,In_2309,In_830);
xnor U171 (N_171,In_1418,In_1033);
and U172 (N_172,In_1188,In_2303);
or U173 (N_173,In_3,In_1217);
or U174 (N_174,In_79,In_1448);
nor U175 (N_175,In_801,In_1603);
and U176 (N_176,In_775,In_1260);
nor U177 (N_177,In_1439,In_1281);
nor U178 (N_178,In_2485,In_1687);
nor U179 (N_179,In_2459,In_346);
nor U180 (N_180,In_2445,In_2076);
and U181 (N_181,In_1527,In_611);
xnor U182 (N_182,In_1323,In_382);
and U183 (N_183,In_2091,In_1691);
and U184 (N_184,In_946,In_2457);
nand U185 (N_185,In_120,In_1008);
nor U186 (N_186,In_1238,In_1617);
xor U187 (N_187,In_1067,In_1843);
and U188 (N_188,In_1093,In_1990);
or U189 (N_189,In_1585,In_1419);
nor U190 (N_190,In_852,In_2140);
xnor U191 (N_191,In_1567,In_1574);
or U192 (N_192,In_1952,In_2229);
nor U193 (N_193,In_241,In_258);
nor U194 (N_194,In_1997,In_803);
or U195 (N_195,In_1389,In_167);
and U196 (N_196,In_799,In_1206);
nand U197 (N_197,In_2173,In_2226);
and U198 (N_198,In_143,In_307);
or U199 (N_199,In_570,In_630);
xor U200 (N_200,In_940,In_621);
xor U201 (N_201,In_1543,In_1974);
xnor U202 (N_202,In_471,In_1465);
nand U203 (N_203,In_2467,In_606);
xnor U204 (N_204,In_146,In_556);
xor U205 (N_205,In_2472,In_2067);
nand U206 (N_206,In_403,In_2128);
or U207 (N_207,In_91,In_2113);
xnor U208 (N_208,In_701,In_1888);
or U209 (N_209,In_2332,In_1812);
or U210 (N_210,In_1068,In_2402);
nand U211 (N_211,In_1904,In_2151);
and U212 (N_212,In_2130,In_1813);
nor U213 (N_213,In_842,In_2257);
nor U214 (N_214,In_21,In_247);
xnor U215 (N_215,In_2462,In_339);
and U216 (N_216,In_1370,In_887);
xor U217 (N_217,In_1250,In_562);
xor U218 (N_218,In_1424,In_578);
nor U219 (N_219,In_1929,In_2283);
or U220 (N_220,In_1229,In_1317);
or U221 (N_221,In_2149,In_2066);
and U222 (N_222,In_1826,In_702);
xor U223 (N_223,In_2214,In_1625);
nor U224 (N_224,In_864,In_98);
and U225 (N_225,In_2252,In_2215);
nand U226 (N_226,In_1862,In_1771);
or U227 (N_227,In_963,In_1122);
or U228 (N_228,In_2266,In_1930);
xor U229 (N_229,In_190,In_2202);
or U230 (N_230,In_2191,In_48);
nor U231 (N_231,In_379,In_1944);
nand U232 (N_232,In_693,In_1616);
nor U233 (N_233,In_1098,In_1919);
nand U234 (N_234,In_481,In_2430);
and U235 (N_235,In_2123,In_2133);
nor U236 (N_236,In_1245,In_1276);
xor U237 (N_237,In_643,In_2349);
nand U238 (N_238,In_208,In_24);
or U239 (N_239,In_2463,In_6);
nor U240 (N_240,In_584,In_2137);
or U241 (N_241,In_1545,In_2132);
nor U242 (N_242,In_2383,In_833);
and U243 (N_243,In_2451,In_1657);
nor U244 (N_244,In_1633,In_184);
nand U245 (N_245,In_876,In_2147);
nand U246 (N_246,In_1387,In_2318);
nand U247 (N_247,In_2106,In_2247);
nor U248 (N_248,In_476,In_504);
or U249 (N_249,In_174,In_1753);
xnor U250 (N_250,In_2009,In_2262);
or U251 (N_251,In_882,In_1207);
nand U252 (N_252,In_1570,In_545);
and U253 (N_253,In_2282,In_2127);
and U254 (N_254,In_449,In_1950);
nand U255 (N_255,In_1073,In_677);
nor U256 (N_256,In_1036,In_329);
or U257 (N_257,In_1348,In_2015);
or U258 (N_258,In_1279,In_1672);
nor U259 (N_259,In_1475,In_20);
xnor U260 (N_260,In_612,In_744);
or U261 (N_261,In_1184,In_1300);
and U262 (N_262,In_837,In_2458);
nand U263 (N_263,In_1860,In_539);
and U264 (N_264,In_345,In_972);
xnor U265 (N_265,In_161,In_893);
nand U266 (N_266,In_1741,In_1163);
xnor U267 (N_267,In_1954,In_671);
or U268 (N_268,In_154,In_1306);
nor U269 (N_269,In_187,In_884);
nand U270 (N_270,In_11,In_558);
or U271 (N_271,In_897,In_1096);
nand U272 (N_272,In_1776,In_2267);
nand U273 (N_273,In_1660,In_1381);
nand U274 (N_274,In_2032,In_1597);
xnor U275 (N_275,In_1414,In_815);
xor U276 (N_276,In_687,In_500);
or U277 (N_277,In_1901,In_715);
nor U278 (N_278,In_848,In_1399);
or U279 (N_279,In_1992,In_2239);
nor U280 (N_280,In_1255,In_2312);
nor U281 (N_281,In_2232,In_1618);
and U282 (N_282,In_1835,In_1572);
nand U283 (N_283,In_1811,In_1469);
nor U284 (N_284,In_356,In_771);
xor U285 (N_285,In_2288,In_1);
xnor U286 (N_286,In_485,In_943);
and U287 (N_287,In_1423,In_1138);
nor U288 (N_288,In_550,In_1961);
and U289 (N_289,In_1372,In_2041);
xor U290 (N_290,In_1792,In_337);
xnor U291 (N_291,In_982,In_517);
xnor U292 (N_292,In_955,In_1917);
and U293 (N_293,In_1949,In_132);
or U294 (N_294,In_827,In_213);
nor U295 (N_295,In_1891,In_2493);
nor U296 (N_296,In_536,In_248);
and U297 (N_297,In_1696,In_1397);
xnor U298 (N_298,In_1340,In_941);
or U299 (N_299,In_1683,In_1876);
nor U300 (N_300,In_2175,In_1898);
and U301 (N_301,In_2122,In_1359);
and U302 (N_302,In_1885,In_300);
xnor U303 (N_303,In_1231,In_1673);
and U304 (N_304,In_88,In_1671);
nor U305 (N_305,In_270,In_1558);
xnor U306 (N_306,In_736,In_1684);
and U307 (N_307,In_2487,In_645);
nand U308 (N_308,In_891,In_1951);
nand U309 (N_309,In_2005,In_1622);
and U310 (N_310,In_1254,In_336);
and U311 (N_311,In_394,In_2496);
or U312 (N_312,In_2255,In_2138);
xnor U313 (N_313,In_1962,In_2263);
nor U314 (N_314,In_1571,In_2298);
nor U315 (N_315,In_181,In_917);
nor U316 (N_316,In_257,In_147);
and U317 (N_317,In_2310,In_1693);
nand U318 (N_318,In_2216,In_144);
xnor U319 (N_319,In_1640,In_625);
and U320 (N_320,In_1540,In_2448);
or U321 (N_321,In_937,In_793);
xnor U322 (N_322,In_535,In_2228);
or U323 (N_323,In_1661,In_726);
or U324 (N_324,In_287,In_130);
and U325 (N_325,In_1445,In_2135);
nand U326 (N_326,In_225,In_1564);
xnor U327 (N_327,In_108,In_817);
xor U328 (N_328,In_1544,In_2044);
or U329 (N_329,In_2331,In_496);
xor U330 (N_330,In_1587,In_2208);
xor U331 (N_331,In_1208,In_2377);
and U332 (N_332,In_385,In_1987);
nand U333 (N_333,In_925,In_2082);
nand U334 (N_334,In_2224,In_1549);
and U335 (N_335,In_2393,In_1436);
xor U336 (N_336,In_84,In_39);
and U337 (N_337,In_999,In_200);
and U338 (N_338,In_455,In_1678);
and U339 (N_339,In_662,In_2146);
nor U340 (N_340,In_920,In_1235);
or U341 (N_341,In_1831,In_975);
or U342 (N_342,In_610,In_2299);
nand U343 (N_343,In_452,In_474);
nor U344 (N_344,In_1647,In_398);
xnor U345 (N_345,In_1395,In_2466);
or U346 (N_346,In_1022,In_2302);
xor U347 (N_347,In_954,In_1286);
xnor U348 (N_348,In_1396,In_289);
nor U349 (N_349,In_710,In_1849);
nand U350 (N_350,In_1228,In_1325);
and U351 (N_351,In_785,In_1680);
or U352 (N_352,In_838,In_657);
xor U353 (N_353,In_266,In_1482);
nor U354 (N_354,In_1936,In_274);
nor U355 (N_355,In_1718,In_28);
nand U356 (N_356,In_1516,In_74);
nand U357 (N_357,In_1243,In_549);
nor U358 (N_358,In_958,In_2423);
or U359 (N_359,In_1730,In_2227);
nor U360 (N_360,In_622,In_1713);
nor U361 (N_361,In_1455,In_1251);
nor U362 (N_362,In_44,In_1409);
or U363 (N_363,In_1195,In_904);
xnor U364 (N_364,In_985,In_1903);
or U365 (N_365,In_761,In_900);
nor U366 (N_366,In_1422,In_1311);
nor U367 (N_367,In_1644,In_1592);
nor U368 (N_368,In_1086,In_767);
or U369 (N_369,In_655,In_542);
xor U370 (N_370,In_2367,In_419);
xor U371 (N_371,In_1559,In_821);
and U372 (N_372,In_1141,In_378);
nor U373 (N_373,In_212,In_1530);
xnor U374 (N_374,In_1791,In_77);
and U375 (N_375,In_443,In_1149);
xor U376 (N_376,In_2265,In_2000);
xor U377 (N_377,In_1337,In_636);
xnor U378 (N_378,In_2102,In_249);
and U379 (N_379,In_1130,In_2324);
nand U380 (N_380,In_1112,In_2022);
nand U381 (N_381,In_2026,In_2110);
xnor U382 (N_382,In_2183,In_660);
nand U383 (N_383,In_711,In_195);
and U384 (N_384,In_1006,In_1715);
xnor U385 (N_385,In_173,In_1575);
xnor U386 (N_386,In_1773,In_351);
nand U387 (N_387,In_428,In_2376);
nor U388 (N_388,In_1449,In_2362);
and U389 (N_389,In_2143,In_1821);
xnor U390 (N_390,In_2219,In_1472);
nor U391 (N_391,In_1166,In_1814);
or U392 (N_392,In_164,In_1435);
xor U393 (N_393,In_2473,In_389);
or U394 (N_394,In_642,In_970);
xor U395 (N_395,In_2052,In_466);
nand U396 (N_396,In_1415,In_753);
nor U397 (N_397,In_2072,In_172);
nor U398 (N_398,In_959,In_2301);
xor U399 (N_399,In_2142,In_581);
or U400 (N_400,In_513,In_2497);
and U401 (N_401,In_2340,In_2078);
and U402 (N_402,In_607,In_1621);
and U403 (N_403,In_1503,In_2033);
xnor U404 (N_404,In_1342,In_2204);
nor U405 (N_405,In_1031,In_2373);
or U406 (N_406,In_901,In_1859);
or U407 (N_407,In_2404,In_782);
and U408 (N_408,In_1519,In_1493);
or U409 (N_409,In_210,In_421);
nand U410 (N_410,In_1787,In_706);
nand U411 (N_411,In_1774,In_341);
xor U412 (N_412,In_1498,In_1187);
nand U413 (N_413,In_1202,In_1975);
nand U414 (N_414,In_1169,In_1820);
and U415 (N_415,In_1349,In_2398);
nand U416 (N_416,In_1977,In_755);
or U417 (N_417,In_2279,In_1304);
and U418 (N_418,In_1142,In_1352);
nor U419 (N_419,In_35,In_1745);
nand U420 (N_420,In_2372,In_217);
xnor U421 (N_421,In_2468,In_1309);
nor U422 (N_422,In_1344,In_2256);
or U423 (N_423,In_1106,In_628);
nand U424 (N_424,In_750,In_1957);
xor U425 (N_425,In_1650,In_209);
xnor U426 (N_426,In_1538,In_1895);
nor U427 (N_427,In_2246,In_1953);
or U428 (N_428,In_2011,In_340);
xor U429 (N_429,In_2307,In_686);
or U430 (N_430,In_634,In_1172);
nor U431 (N_431,In_2154,In_1171);
nor U432 (N_432,In_391,In_2399);
and U433 (N_433,In_730,In_935);
nor U434 (N_434,In_1872,In_2287);
or U435 (N_435,In_76,In_2141);
or U436 (N_436,In_2424,In_281);
and U437 (N_437,In_1629,In_2358);
xnor U438 (N_438,In_479,In_1425);
nor U439 (N_439,In_90,In_1158);
or U440 (N_440,In_1796,In_1518);
xor U441 (N_441,In_1722,In_679);
nand U442 (N_442,In_743,In_843);
or U443 (N_443,In_1882,In_991);
and U444 (N_444,In_103,In_1837);
xnor U445 (N_445,In_1426,In_523);
xor U446 (N_446,In_2054,In_1261);
or U447 (N_447,In_501,In_383);
and U448 (N_448,In_405,In_1702);
nor U449 (N_449,In_713,In_1041);
or U450 (N_450,In_65,In_1161);
or U451 (N_451,In_1314,In_1681);
xnor U452 (N_452,In_1099,In_1623);
nand U453 (N_453,In_1795,In_87);
and U454 (N_454,In_215,In_2251);
nor U455 (N_455,In_1886,In_1014);
nand U456 (N_456,In_390,In_23);
nor U457 (N_457,In_1053,In_1117);
xor U458 (N_458,In_1897,In_1676);
or U459 (N_459,In_2476,In_2408);
nand U460 (N_460,In_1966,In_2308);
or U461 (N_461,In_1001,In_1413);
xnor U462 (N_462,In_2260,In_80);
or U463 (N_463,In_1119,In_708);
and U464 (N_464,In_617,In_1920);
or U465 (N_465,In_1939,In_1284);
nand U466 (N_466,In_1363,In_198);
nand U467 (N_467,In_866,In_1579);
nand U468 (N_468,In_850,In_141);
nor U469 (N_469,In_1266,In_1505);
nand U470 (N_470,In_2134,In_1327);
and U471 (N_471,In_1489,In_1412);
nand U472 (N_472,In_2414,In_1120);
nand U473 (N_473,In_787,In_1993);
nand U474 (N_474,In_2045,In_134);
and U475 (N_475,In_1942,In_957);
and U476 (N_476,In_1656,In_1442);
nor U477 (N_477,In_196,In_2094);
nand U478 (N_478,In_2355,In_1908);
nor U479 (N_479,In_1089,In_564);
or U480 (N_480,In_983,In_277);
or U481 (N_481,In_1865,In_1510);
nand U482 (N_482,In_619,In_29);
nand U483 (N_483,In_2063,In_1697);
nor U484 (N_484,In_1437,In_694);
and U485 (N_485,In_350,In_2002);
nor U486 (N_486,In_1790,In_2410);
or U487 (N_487,In_807,In_2025);
nor U488 (N_488,In_155,In_1887);
or U489 (N_489,In_2035,In_2156);
and U490 (N_490,In_819,In_1819);
xor U491 (N_491,In_742,In_2306);
xnor U492 (N_492,In_1154,In_124);
nor U493 (N_493,In_207,In_2317);
nor U494 (N_494,In_1923,In_235);
nor U495 (N_495,In_465,In_1626);
and U496 (N_496,In_1287,In_2380);
xor U497 (N_497,In_377,In_1692);
and U498 (N_498,In_302,In_1512);
or U499 (N_499,In_699,In_1383);
xor U500 (N_500,In_1338,In_1852);
xor U501 (N_501,In_2481,In_1405);
or U502 (N_502,In_936,In_386);
nor U503 (N_503,In_822,In_1114);
or U504 (N_504,In_717,In_1578);
nand U505 (N_505,In_2197,In_633);
or U506 (N_506,In_353,In_1052);
and U507 (N_507,In_762,In_2370);
nand U508 (N_508,In_1294,In_1902);
or U509 (N_509,In_1240,In_2359);
xnor U510 (N_510,In_681,In_293);
nor U511 (N_511,In_608,In_1491);
and U512 (N_512,In_1956,In_2374);
and U513 (N_513,In_2357,In_7);
and U514 (N_514,In_49,In_1270);
xnor U515 (N_515,In_725,In_2498);
xor U516 (N_516,In_1331,In_2489);
or U517 (N_517,In_113,In_1203);
and U518 (N_518,In_2217,In_704);
nand U519 (N_519,In_1589,In_1938);
or U520 (N_520,In_2409,In_2401);
nor U521 (N_521,In_1967,In_2434);
and U522 (N_522,In_2452,In_1806);
xor U523 (N_523,In_1760,In_1265);
and U524 (N_524,In_2360,In_355);
nor U525 (N_525,In_415,In_908);
nor U526 (N_526,In_2274,In_45);
nand U527 (N_527,In_600,In_566);
or U528 (N_528,In_637,In_1816);
nand U529 (N_529,In_967,In_2253);
nand U530 (N_530,In_93,In_1480);
and U531 (N_531,In_2039,In_2100);
or U532 (N_532,In_851,In_1914);
nand U533 (N_533,In_805,In_498);
nor U534 (N_534,In_540,In_1147);
and U535 (N_535,In_369,In_142);
nand U536 (N_536,In_2148,In_370);
nor U537 (N_537,In_632,In_1464);
and U538 (N_538,In_1355,In_1293);
or U539 (N_539,In_129,In_402);
or U540 (N_540,In_392,In_658);
xnor U541 (N_541,In_2124,In_359);
xor U542 (N_542,In_1754,In_261);
nor U543 (N_543,In_2037,In_1871);
nor U544 (N_544,In_1104,In_1100);
xor U545 (N_545,In_1272,In_2034);
xnor U546 (N_546,In_703,In_853);
or U547 (N_547,In_2353,In_1018);
or U548 (N_548,In_1627,In_1057);
nand U549 (N_549,In_2162,In_748);
nand U550 (N_550,In_1076,In_716);
and U551 (N_551,In_2057,In_747);
and U552 (N_552,In_1462,In_363);
or U553 (N_553,In_906,In_839);
nor U554 (N_554,In_690,In_1484);
nor U555 (N_555,In_1196,In_916);
nor U556 (N_556,In_1485,In_656);
nor U557 (N_557,In_81,In_1761);
xnor U558 (N_558,In_810,In_1945);
and U559 (N_559,In_1262,In_204);
and U560 (N_560,In_1874,In_2092);
nor U561 (N_561,In_2389,In_1851);
xor U562 (N_562,In_1354,In_889);
nor U563 (N_563,In_844,In_376);
xnor U564 (N_564,In_514,In_956);
and U565 (N_565,In_727,In_2342);
and U566 (N_566,In_275,In_1159);
nor U567 (N_567,In_37,In_758);
nand U568 (N_568,In_1277,In_2261);
xor U569 (N_569,In_26,In_499);
xnor U570 (N_570,In_1429,In_1576);
nand U571 (N_571,In_1620,In_2179);
xor U572 (N_572,In_1810,In_43);
nand U573 (N_573,In_1928,In_2413);
or U574 (N_574,In_1151,In_586);
or U575 (N_575,In_1911,In_794);
nand U576 (N_576,In_326,In_2065);
nor U577 (N_577,In_649,In_1186);
and U578 (N_578,In_19,In_2454);
and U579 (N_579,In_698,In_676);
nor U580 (N_580,In_2335,In_1507);
nor U581 (N_581,In_1035,In_605);
and U582 (N_582,In_604,In_176);
xnor U583 (N_583,In_100,In_437);
and U584 (N_584,In_1376,In_1247);
xnor U585 (N_585,In_1230,In_1162);
or U586 (N_586,In_162,In_1094);
xor U587 (N_587,In_1638,In_1844);
and U588 (N_588,In_1440,In_734);
nor U589 (N_589,In_609,In_1658);
xor U590 (N_590,In_2276,In_594);
and U591 (N_591,In_977,In_1769);
nand U592 (N_592,In_1619,In_2230);
and U593 (N_593,In_2200,In_537);
nand U594 (N_594,In_2412,In_984);
xnor U595 (N_595,In_665,In_2323);
and U596 (N_596,In_544,In_1028);
and U597 (N_597,In_1222,In_1080);
nor U598 (N_598,In_448,In_695);
xnor U599 (N_599,In_1973,In_467);
nand U600 (N_600,In_1274,In_1979);
xnor U601 (N_601,In_572,In_1699);
or U602 (N_602,In_1038,In_1118);
and U603 (N_603,In_1529,In_436);
and U604 (N_604,In_1698,In_574);
nor U605 (N_605,In_898,In_2447);
xnor U606 (N_606,In_2220,In_1583);
nor U607 (N_607,In_487,In_774);
nor U608 (N_608,In_2321,In_236);
or U609 (N_609,In_924,In_1781);
and U610 (N_610,In_1918,In_2474);
nand U611 (N_611,In_1467,In_211);
nand U612 (N_612,In_816,In_1246);
or U613 (N_613,In_462,In_1268);
and U614 (N_614,In_282,In_1392);
xnor U615 (N_615,In_1910,In_2294);
nand U616 (N_616,In_1659,In_441);
nor U617 (N_617,In_1906,In_751);
or U618 (N_618,In_2040,In_528);
and U619 (N_619,In_1050,In_41);
xnor U620 (N_620,In_2060,In_2236);
nor U621 (N_621,In_243,In_1825);
nor U622 (N_622,In_524,In_192);
nand U623 (N_623,In_2030,In_251);
nor U624 (N_624,In_12,In_1756);
xnor U625 (N_625,In_1894,In_2075);
or U626 (N_626,In_2095,In_620);
and U627 (N_627,In_18,In_1074);
xnor U628 (N_628,In_664,In_2205);
nand U629 (N_629,In_1111,In_101);
and U630 (N_630,In_13,In_425);
or U631 (N_631,In_1841,In_447);
nor U632 (N_632,In_714,In_2088);
nand U633 (N_633,In_1269,In_175);
nand U634 (N_634,In_253,In_234);
and U635 (N_635,In_2086,In_1316);
and U636 (N_636,In_719,In_323);
xnor U637 (N_637,In_1818,In_1506);
or U638 (N_638,In_2397,In_1244);
xor U639 (N_639,In_961,In_1907);
nor U640 (N_640,In_2285,In_250);
and U641 (N_641,In_468,In_1532);
nor U642 (N_642,In_678,In_1248);
or U643 (N_643,In_618,In_1573);
nand U644 (N_644,In_1432,In_2289);
nor U645 (N_645,In_1668,In_709);
xor U646 (N_646,In_2313,In_832);
nand U647 (N_647,In_1896,In_2442);
and U648 (N_648,In_1299,In_429);
or U649 (N_649,In_691,In_372);
and U650 (N_650,In_2482,In_2004);
nor U651 (N_651,In_547,In_1146);
or U652 (N_652,In_114,In_295);
nor U653 (N_653,In_746,In_1042);
xnor U654 (N_654,In_919,In_2428);
or U655 (N_655,In_1194,In_193);
nor U656 (N_656,In_1318,In_507);
nor U657 (N_657,In_1378,In_278);
or U658 (N_658,In_2478,In_1749);
nor U659 (N_659,In_1783,In_2345);
nor U660 (N_660,In_1446,In_1181);
and U661 (N_661,In_182,In_921);
and U662 (N_662,In_2170,In_804);
nor U663 (N_663,In_2077,In_283);
xnor U664 (N_664,In_1384,In_308);
nand U665 (N_665,In_276,In_230);
nor U666 (N_666,In_623,In_2061);
nor U667 (N_667,In_52,In_849);
or U668 (N_668,In_1978,In_1972);
or U669 (N_669,In_2375,In_1115);
xnor U670 (N_670,In_1648,In_599);
nand U671 (N_671,In_352,In_541);
or U672 (N_672,In_1406,In_1964);
nand U673 (N_673,In_457,In_614);
or U674 (N_674,In_1915,In_1332);
nor U675 (N_675,In_1212,In_1034);
nor U676 (N_676,In_318,In_2019);
nor U677 (N_677,In_1569,In_588);
or U678 (N_678,In_1602,In_1346);
xor U679 (N_679,In_860,In_2411);
nand U680 (N_680,In_417,In_1649);
or U681 (N_681,In_1379,In_776);
nand U682 (N_682,In_1330,In_140);
and U683 (N_683,In_237,In_256);
nor U684 (N_684,In_2168,In_1471);
and U685 (N_685,In_149,In_214);
and U686 (N_686,In_1926,In_1836);
nand U687 (N_687,In_823,In_82);
nor U688 (N_688,In_777,In_962);
or U689 (N_689,In_526,In_15);
or U690 (N_690,In_239,In_765);
xnor U691 (N_691,In_1241,In_1322);
xnor U692 (N_692,In_2386,In_1428);
xor U693 (N_693,In_2427,In_2099);
and U694 (N_694,In_2071,In_1881);
and U695 (N_695,In_246,In_472);
nor U696 (N_696,In_2432,In_1064);
or U697 (N_697,In_31,In_2098);
and U698 (N_698,In_1523,In_1665);
or U699 (N_699,In_1478,In_1252);
nand U700 (N_700,In_684,In_357);
or U701 (N_701,In_1736,In_1751);
or U702 (N_702,In_1199,In_2101);
xor U703 (N_703,In_1766,In_1724);
nor U704 (N_704,In_188,In_226);
xor U705 (N_705,In_1534,In_9);
nor U706 (N_706,In_288,In_1292);
nor U707 (N_707,In_2405,In_1875);
nand U708 (N_708,In_661,In_2196);
nand U709 (N_709,In_56,In_2115);
nor U710 (N_710,In_1504,In_280);
and U711 (N_711,In_42,In_121);
nor U712 (N_712,In_1721,In_1225);
and U713 (N_713,In_2081,In_4);
nand U714 (N_714,In_733,In_2480);
xor U715 (N_715,In_435,In_119);
nand U716 (N_716,In_373,In_2058);
nor U717 (N_717,In_1002,In_1390);
nand U718 (N_718,In_1808,In_331);
nand U719 (N_719,In_1899,In_1971);
nand U720 (N_720,In_422,In_1126);
xor U721 (N_721,In_338,In_546);
or U722 (N_722,In_2300,In_934);
or U723 (N_723,In_227,In_1447);
xnor U724 (N_724,In_1965,In_939);
nor U725 (N_725,In_2254,In_769);
nand U726 (N_726,In_583,In_1565);
nor U727 (N_727,In_83,In_296);
nor U728 (N_728,In_64,In_616);
nand U729 (N_729,In_802,In_1707);
nor U730 (N_730,In_1652,In_123);
xor U731 (N_731,In_59,In_2337);
or U732 (N_732,In_2440,In_1223);
xnor U733 (N_733,In_1958,In_700);
nand U734 (N_734,In_1417,In_590);
nand U735 (N_735,In_450,In_1328);
nand U736 (N_736,In_2368,In_1889);
xor U737 (N_737,In_2431,In_2053);
nand U738 (N_738,In_36,In_1989);
xor U739 (N_739,In_1308,In_627);
or U740 (N_740,In_291,In_1487);
nor U741 (N_741,In_950,In_180);
and U742 (N_742,In_224,In_1800);
nand U743 (N_743,In_1960,In_1935);
and U744 (N_744,In_2272,In_868);
nand U745 (N_745,In_754,In_199);
nand U746 (N_746,In_259,In_1048);
xnor U747 (N_747,In_1335,In_861);
nor U748 (N_748,In_1148,In_1078);
xnor U749 (N_749,In_1596,In_2439);
or U750 (N_750,In_371,In_416);
nor U751 (N_751,In_151,In_1434);
nand U752 (N_752,In_2150,In_160);
xor U753 (N_753,In_2381,In_989);
nor U754 (N_754,In_58,In_495);
and U755 (N_755,In_721,In_1980);
nand U756 (N_756,In_1024,In_1675);
xor U757 (N_757,In_1900,In_1190);
xnor U758 (N_758,In_763,In_231);
xnor U759 (N_759,In_2244,In_1291);
nand U760 (N_760,In_63,In_615);
or U761 (N_761,In_576,In_46);
or U762 (N_762,In_67,In_1092);
nor U763 (N_763,In_1077,In_116);
or U764 (N_764,In_1568,In_458);
xnor U765 (N_765,In_909,In_1431);
xor U766 (N_766,In_2139,In_825);
xnor U767 (N_767,In_1430,In_2491);
and U768 (N_768,In_86,In_1010);
xor U769 (N_769,In_1461,In_722);
xor U770 (N_770,In_988,In_1134);
nor U771 (N_771,In_560,In_1438);
or U772 (N_772,In_1444,In_47);
nand U773 (N_773,In_994,In_2436);
nand U774 (N_774,In_2245,In_1357);
nor U775 (N_775,In_301,In_757);
nand U776 (N_776,In_32,In_759);
xor U777 (N_777,In_2085,In_1535);
xnor U778 (N_778,In_515,In_2259);
nor U779 (N_779,In_2010,In_647);
xor U780 (N_780,In_2036,In_503);
xnor U781 (N_781,In_1537,In_1705);
or U782 (N_782,In_668,In_1524);
nor U783 (N_783,In_1631,In_423);
nand U784 (N_784,In_927,In_315);
nand U785 (N_785,In_669,In_460);
or U786 (N_786,In_2237,In_563);
and U787 (N_787,In_601,In_189);
nor U788 (N_788,In_1016,In_1765);
and U789 (N_789,In_1288,In_1662);
or U790 (N_790,In_27,In_1492);
and U791 (N_791,In_2116,In_131);
nand U792 (N_792,In_1890,In_1866);
and U793 (N_793,In_1725,In_463);
and U794 (N_794,In_1913,In_1679);
and U795 (N_795,In_1539,In_2425);
nor U796 (N_796,In_1511,In_299);
or U797 (N_797,In_2258,In_71);
and U798 (N_798,In_2361,In_2316);
and U799 (N_799,In_1674,In_38);
and U800 (N_800,In_1375,In_327);
nand U801 (N_801,In_157,In_85);
or U802 (N_802,In_1767,In_1232);
nor U803 (N_803,In_2460,In_911);
nand U804 (N_804,In_1458,In_2048);
or U805 (N_805,In_201,In_1071);
and U806 (N_806,In_16,In_1054);
or U807 (N_807,In_1838,In_1797);
or U808 (N_808,In_2209,In_1066);
or U809 (N_809,In_1606,In_1214);
and U810 (N_810,In_1009,In_104);
xor U811 (N_811,In_1296,In_2001);
nor U812 (N_812,In_1799,In_1007);
xnor U813 (N_813,In_1912,In_979);
xnor U814 (N_814,In_406,In_1772);
xnor U815 (N_815,In_1809,In_2450);
xor U816 (N_816,In_2166,In_976);
nor U817 (N_817,In_1200,In_834);
xnor U818 (N_818,In_986,In_1667);
and U819 (N_819,In_1943,In_1404);
nor U820 (N_820,In_442,In_910);
nor U821 (N_821,In_672,In_2021);
nor U822 (N_822,In_1451,In_2042);
xnor U823 (N_823,In_1361,In_2379);
xor U824 (N_824,In_1173,In_745);
or U825 (N_825,In_2221,In_2031);
nand U826 (N_826,In_2271,In_1827);
or U827 (N_827,In_69,In_1994);
nor U828 (N_828,In_1156,In_2180);
or U829 (N_829,In_2270,In_2144);
xnor U830 (N_830,In_1345,In_70);
and U831 (N_831,In_918,In_232);
xor U832 (N_832,In_1802,In_1793);
nand U833 (N_833,In_559,In_1488);
nand U834 (N_834,In_1723,In_1611);
and U835 (N_835,In_1443,In_1476);
nand U836 (N_836,In_1748,In_244);
or U837 (N_837,In_846,In_1339);
and U838 (N_838,In_1610,In_1310);
nand U839 (N_839,In_1221,In_2240);
nor U840 (N_840,In_1546,In_117);
and U841 (N_841,In_223,In_855);
or U842 (N_842,In_1051,In_1867);
xnor U843 (N_843,In_2074,In_862);
and U844 (N_844,In_368,In_530);
or U845 (N_845,In_2248,In_1522);
and U846 (N_846,In_1013,In_1297);
and U847 (N_847,In_128,In_2284);
nand U848 (N_848,In_675,In_66);
or U849 (N_849,In_2218,In_1191);
xnor U850 (N_850,In_1209,In_858);
or U851 (N_851,In_1358,In_854);
or U852 (N_852,In_2003,In_133);
or U853 (N_853,In_1752,In_692);
or U854 (N_854,In_569,In_1877);
xnor U855 (N_855,In_1271,In_1143);
nor U856 (N_856,In_1883,In_492);
or U857 (N_857,In_1557,In_97);
xor U858 (N_858,In_2210,In_2494);
or U859 (N_859,In_2416,In_2297);
and U860 (N_860,In_51,In_1520);
and U861 (N_861,In_1732,In_313);
and U862 (N_862,In_2320,In_1032);
xor U863 (N_863,In_968,In_1682);
and U864 (N_864,In_347,In_1371);
and U865 (N_865,In_1541,In_1933);
nand U866 (N_866,In_2351,In_789);
and U867 (N_867,In_2273,In_2417);
xor U868 (N_868,In_2164,In_126);
and U869 (N_869,In_847,In_1063);
nand U870 (N_870,In_240,In_723);
xor U871 (N_871,In_168,In_990);
and U872 (N_872,In_874,In_33);
and U873 (N_873,In_365,In_2093);
nor U874 (N_874,In_1070,In_407);
xnor U875 (N_875,In_404,In_1670);
and U876 (N_876,In_1746,In_292);
nand U877 (N_877,In_57,In_348);
and U878 (N_878,In_795,In_1334);
nand U879 (N_879,In_2178,In_2385);
xor U880 (N_880,In_1388,In_2418);
nand U881 (N_881,In_1319,In_2486);
nor U882 (N_882,In_881,In_533);
nor U883 (N_883,In_527,In_298);
nand U884 (N_884,In_2464,In_14);
or U885 (N_885,In_1239,In_964);
nand U886 (N_886,In_1312,In_791);
nand U887 (N_887,In_1739,In_2212);
or U888 (N_888,In_797,In_863);
and U889 (N_889,In_216,In_1110);
xor U890 (N_890,In_1531,In_424);
nor U891 (N_891,In_2190,In_439);
xnor U892 (N_892,In_40,In_2056);
nand U893 (N_893,In_809,In_800);
and U894 (N_894,In_557,In_659);
or U895 (N_895,In_595,In_931);
nor U896 (N_896,In_1879,In_1216);
or U897 (N_897,In_1785,In_96);
and U898 (N_898,In_1295,In_1985);
xnor U899 (N_899,In_367,In_1710);
xnor U900 (N_900,In_1969,In_1468);
xor U901 (N_901,In_813,In_2437);
nand U902 (N_902,In_2403,In_870);
xnor U903 (N_903,In_1641,In_867);
and U904 (N_904,In_2155,In_2161);
nand U905 (N_905,In_2008,In_2475);
xor U906 (N_906,In_1738,In_1999);
nor U907 (N_907,In_1481,In_2121);
nand U908 (N_908,In_818,In_1257);
nand U909 (N_909,In_1129,In_772);
and U910 (N_910,In_1582,In_1321);
nor U911 (N_911,In_8,In_469);
nand U912 (N_912,In_1003,In_1720);
nor U913 (N_913,In_229,In_1803);
nand U914 (N_914,In_1233,In_2187);
nor U915 (N_915,In_1474,In_220);
nor U916 (N_916,In_2174,In_1921);
or U917 (N_917,In_2420,In_509);
and U918 (N_918,In_1770,In_1991);
nor U919 (N_919,In_420,In_879);
nand U920 (N_920,In_2055,In_72);
and U921 (N_921,In_886,In_1685);
nand U922 (N_922,In_1744,In_1857);
nand U923 (N_923,In_2073,In_1452);
or U924 (N_924,In_1182,In_1303);
or U925 (N_925,In_1150,In_2333);
or U926 (N_926,In_948,In_565);
nand U927 (N_927,In_2020,In_486);
nor U928 (N_928,In_34,In_538);
nor U929 (N_929,In_1735,In_1873);
or U930 (N_930,In_811,In_2495);
xor U931 (N_931,In_1084,In_1758);
and U932 (N_932,In_205,In_1634);
xnor U933 (N_933,In_2062,In_812);
or U934 (N_934,In_269,In_366);
nor U935 (N_935,In_2157,In_1393);
nand U936 (N_936,In_829,In_145);
nand U937 (N_937,In_342,In_1427);
or U938 (N_938,In_2160,In_1020);
nand U939 (N_939,In_1932,In_271);
or U940 (N_940,In_2369,In_2339);
nand U941 (N_941,In_505,In_95);
nand U942 (N_942,In_1624,In_1666);
nor U943 (N_943,In_2365,In_1562);
or U944 (N_944,In_1830,In_992);
or U945 (N_945,In_597,In_883);
xor U946 (N_946,In_1653,In_252);
nor U947 (N_947,In_635,In_165);
xnor U948 (N_948,In_1983,In_1267);
xor U949 (N_949,In_1011,In_105);
nand U950 (N_950,In_156,In_1189);
xor U951 (N_951,In_1136,In_262);
and U952 (N_952,In_413,In_2043);
xnor U953 (N_953,In_1283,In_333);
nand U954 (N_954,In_902,In_1017);
or U955 (N_955,In_473,In_2356);
xor U956 (N_956,In_445,In_304);
nand U957 (N_957,In_2314,In_1817);
and U958 (N_958,In_1400,In_593);
or U959 (N_959,In_267,In_930);
xnor U960 (N_960,In_2499,In_1095);
xnor U961 (N_961,In_2366,In_1853);
nand U962 (N_962,In_682,In_1847);
and U963 (N_963,In_1759,In_1547);
or U964 (N_964,In_1386,In_1023);
nand U965 (N_965,In_1591,In_1369);
and U966 (N_966,In_112,In_1613);
nand U967 (N_967,In_1410,In_1686);
and U968 (N_968,In_2291,In_1968);
and U969 (N_969,In_953,In_1160);
or U970 (N_970,In_1842,In_2169);
nor U971 (N_971,In_1768,In_1152);
xnor U972 (N_972,In_2391,In_1210);
nor U973 (N_973,In_865,In_1324);
xnor U974 (N_974,In_2296,In_349);
nor U975 (N_975,In_2211,In_242);
nand U976 (N_976,In_1855,In_314);
and U977 (N_977,In_773,In_2083);
nand U978 (N_978,In_981,In_1085);
nor U979 (N_979,In_2069,In_2107);
nand U980 (N_980,In_2264,In_641);
and U981 (N_981,In_778,In_1391);
nor U982 (N_982,In_2346,In_638);
nand U983 (N_983,In_1497,In_1249);
and U984 (N_984,In_1976,In_1514);
and U985 (N_985,In_995,In_1743);
xor U986 (N_986,In_2096,In_238);
nand U987 (N_987,In_1839,In_756);
or U988 (N_988,In_1780,In_1026);
xnor U989 (N_989,In_312,In_328);
and U990 (N_990,In_806,In_53);
xor U991 (N_991,In_491,In_2492);
or U992 (N_992,In_1709,In_332);
nand U993 (N_993,In_798,In_1108);
nor U994 (N_994,In_2350,In_2105);
or U995 (N_995,In_2378,In_786);
nor U996 (N_996,In_2165,In_1664);
nand U997 (N_997,In_1502,In_1218);
xor U998 (N_998,In_529,In_1615);
or U999 (N_999,In_2311,In_344);
nand U1000 (N_1000,In_880,In_1101);
xnor U1001 (N_1001,In_1351,N_355);
nand U1002 (N_1002,N_867,In_171);
or U1003 (N_1003,N_565,In_2186);
or U1004 (N_1004,N_872,N_134);
or U1005 (N_1005,N_396,N_442);
nand U1006 (N_1006,N_633,N_360);
xor U1007 (N_1007,N_521,N_743);
or U1008 (N_1008,N_845,N_590);
xor U1009 (N_1009,In_2014,In_1822);
and U1010 (N_1010,In_2305,N_152);
and U1011 (N_1011,N_77,N_991);
nand U1012 (N_1012,In_1864,N_446);
xnor U1013 (N_1013,N_671,N_35);
or U1014 (N_1014,N_197,In_915);
nand U1015 (N_1015,N_185,N_365);
nand U1016 (N_1016,In_453,N_174);
and U1017 (N_1017,In_652,In_1204);
nand U1018 (N_1018,N_315,In_760);
or U1019 (N_1019,N_748,N_933);
xnor U1020 (N_1020,N_645,N_286);
xor U1021 (N_1021,N_544,N_250);
and U1022 (N_1022,In_2103,N_987);
or U1023 (N_1023,N_443,N_841);
nand U1024 (N_1024,N_689,N_503);
or U1025 (N_1025,N_901,In_2109);
nand U1026 (N_1026,N_102,N_228);
and U1027 (N_1027,N_898,N_701);
and U1028 (N_1028,N_0,N_183);
and U1029 (N_1029,N_419,In_1551);
or U1030 (N_1030,N_206,N_612);
nand U1031 (N_1031,N_15,In_783);
nand U1032 (N_1032,N_575,In_1072);
nand U1033 (N_1033,In_1645,In_1909);
nand U1034 (N_1034,N_267,N_636);
or U1035 (N_1035,N_430,N_478);
xor U1036 (N_1036,In_1402,N_566);
nor U1037 (N_1037,In_1336,In_1854);
nor U1038 (N_1038,N_230,N_136);
and U1039 (N_1039,N_802,In_1091);
nand U1040 (N_1040,N_540,N_19);
or U1041 (N_1041,In_1553,N_460);
nand U1042 (N_1042,N_952,N_18);
or U1043 (N_1043,In_1884,In_411);
xor U1044 (N_1044,N_232,N_208);
nor U1045 (N_1045,N_795,In_845);
xnor U1046 (N_1046,N_275,In_426);
or U1047 (N_1047,N_877,N_660);
and U1048 (N_1048,N_614,N_104);
and U1049 (N_1049,N_382,N_855);
xor U1050 (N_1050,N_379,N_215);
or U1051 (N_1051,N_741,In_1132);
nand U1052 (N_1052,In_1103,N_860);
nand U1053 (N_1053,N_347,N_695);
nand U1054 (N_1054,N_945,N_781);
xnor U1055 (N_1055,N_370,In_820);
nand U1056 (N_1056,In_2400,N_941);
nand U1057 (N_1057,N_746,N_432);
nor U1058 (N_1058,N_148,N_497);
xor U1059 (N_1059,N_857,In_913);
nand U1060 (N_1060,In_2443,N_803);
or U1061 (N_1061,In_343,In_2);
or U1062 (N_1062,In_735,In_1636);
and U1063 (N_1063,N_637,N_667);
or U1064 (N_1064,N_218,In_1856);
nor U1065 (N_1065,In_1861,In_1315);
xnor U1066 (N_1066,In_1840,In_115);
xnor U1067 (N_1067,N_425,N_17);
and U1068 (N_1068,N_766,N_962);
or U1069 (N_1069,In_1594,In_1892);
or U1070 (N_1070,N_135,N_10);
or U1071 (N_1071,In_824,N_221);
or U1072 (N_1072,N_253,N_349);
nor U1073 (N_1073,N_725,In_169);
and U1074 (N_1074,N_778,In_1046);
nand U1075 (N_1075,N_479,N_783);
and U1076 (N_1076,N_367,N_893);
nor U1077 (N_1077,In_294,In_1341);
xor U1078 (N_1078,N_592,N_681);
nand U1079 (N_1079,N_717,N_486);
and U1080 (N_1080,N_976,N_536);
nor U1081 (N_1081,N_356,N_761);
nor U1082 (N_1082,N_62,In_577);
xor U1083 (N_1083,In_974,N_244);
nand U1084 (N_1084,In_490,N_294);
nor U1085 (N_1085,N_552,N_281);
nand U1086 (N_1086,N_409,N_490);
nand U1087 (N_1087,N_448,N_696);
nor U1088 (N_1088,N_325,N_368);
xnor U1089 (N_1089,N_533,N_115);
xor U1090 (N_1090,In_2090,N_639);
and U1091 (N_1091,N_713,N_441);
nand U1092 (N_1092,N_685,N_143);
nand U1093 (N_1093,In_68,N_792);
or U1094 (N_1094,N_679,N_264);
and U1095 (N_1095,N_587,N_881);
or U1096 (N_1096,In_770,N_57);
nand U1097 (N_1097,N_784,In_1695);
nand U1098 (N_1098,N_74,N_970);
or U1099 (N_1099,N_509,N_205);
nand U1100 (N_1100,N_394,In_99);
nand U1101 (N_1101,In_511,N_241);
or U1102 (N_1102,In_432,N_238);
xor U1103 (N_1103,N_887,N_602);
and U1104 (N_1104,N_472,N_144);
xnor U1105 (N_1105,N_388,N_569);
or U1106 (N_1106,In_971,N_630);
nand U1107 (N_1107,N_395,N_272);
or U1108 (N_1108,In_705,N_276);
xor U1109 (N_1109,In_1719,N_735);
or U1110 (N_1110,In_1157,N_782);
nor U1111 (N_1111,In_508,In_78);
nand U1112 (N_1112,N_744,In_1561);
and U1113 (N_1113,N_178,N_336);
and U1114 (N_1114,N_437,In_2104);
nand U1115 (N_1115,N_576,N_723);
xnor U1116 (N_1116,N_688,In_218);
nor U1117 (N_1117,N_538,In_914);
xor U1118 (N_1118,In_2419,In_1654);
xor U1119 (N_1119,In_1548,N_374);
xnor U1120 (N_1120,N_714,N_27);
xor U1121 (N_1121,In_2280,N_971);
xnor U1122 (N_1122,N_429,N_982);
and U1123 (N_1123,N_462,N_186);
or U1124 (N_1124,N_285,In_185);
nand U1125 (N_1125,N_234,N_157);
nor U1126 (N_1126,N_574,N_983);
xor U1127 (N_1127,N_369,N_291);
and U1128 (N_1128,N_304,In_648);
and U1129 (N_1129,N_22,In_381);
and U1130 (N_1130,N_495,N_458);
nor U1131 (N_1131,In_980,In_534);
nor U1132 (N_1132,In_245,N_164);
nor U1133 (N_1133,N_648,In_603);
nand U1134 (N_1134,N_523,In_497);
nor U1135 (N_1135,N_481,N_597);
or U1136 (N_1136,In_1905,In_319);
or U1137 (N_1137,N_141,N_635);
and U1138 (N_1138,N_620,N_457);
and U1139 (N_1139,In_2329,In_320);
and U1140 (N_1140,In_1343,N_835);
xnor U1141 (N_1141,N_311,N_44);
nand U1142 (N_1142,N_563,N_762);
nand U1143 (N_1143,In_1560,N_900);
nor U1144 (N_1144,N_665,N_939);
xnor U1145 (N_1145,In_1786,In_1083);
or U1146 (N_1146,N_345,N_979);
or U1147 (N_1147,N_879,N_322);
xnor U1148 (N_1148,N_522,In_1015);
xor U1149 (N_1149,In_780,N_306);
and U1150 (N_1150,N_265,N_530);
and U1151 (N_1151,N_651,N_615);
and U1152 (N_1152,N_116,In_106);
and U1153 (N_1153,In_1927,N_505);
nor U1154 (N_1154,N_280,N_268);
nand U1155 (N_1155,N_85,N_925);
xor U1156 (N_1156,In_1823,N_547);
or U1157 (N_1157,N_142,N_791);
xor U1158 (N_1158,N_596,N_416);
nand U1159 (N_1159,N_626,N_916);
xor U1160 (N_1160,In_740,N_708);
nor U1161 (N_1161,In_75,In_1385);
nor U1162 (N_1162,N_213,N_191);
or U1163 (N_1163,In_2330,N_156);
xor U1164 (N_1164,In_1550,N_926);
nor U1165 (N_1165,N_707,N_202);
or U1166 (N_1166,N_124,N_196);
nand U1167 (N_1167,In_2114,In_1045);
and U1168 (N_1168,N_578,N_757);
or U1169 (N_1169,N_76,N_32);
and U1170 (N_1170,N_649,N_537);
nor U1171 (N_1171,N_471,N_433);
nand U1172 (N_1172,N_715,In_306);
nand U1173 (N_1173,N_95,N_903);
nand U1174 (N_1174,N_956,N_384);
and U1175 (N_1175,N_730,N_912);
or U1176 (N_1176,N_502,N_525);
nand U1177 (N_1177,N_683,N_131);
xnor U1178 (N_1178,N_924,N_387);
nand U1179 (N_1179,In_688,In_1227);
nand U1180 (N_1180,N_172,N_112);
and U1181 (N_1181,N_830,N_98);
or U1182 (N_1182,In_2286,N_928);
or U1183 (N_1183,N_121,N_81);
xor U1184 (N_1184,In_2070,N_729);
nor U1185 (N_1185,N_591,N_151);
and U1186 (N_1186,N_63,N_198);
or U1187 (N_1187,N_390,N_201);
or U1188 (N_1188,In_2444,In_2295);
and U1189 (N_1189,N_261,In_1922);
nor U1190 (N_1190,N_884,N_105);
xor U1191 (N_1191,In_1729,In_1253);
and U1192 (N_1192,N_663,N_348);
and U1193 (N_1193,N_828,N_461);
nand U1194 (N_1194,In_2363,N_786);
nor U1195 (N_1195,In_1131,N_73);
nand U1196 (N_1196,N_551,N_814);
nor U1197 (N_1197,N_439,N_45);
nand U1198 (N_1198,N_175,N_519);
nor U1199 (N_1199,N_499,N_277);
or U1200 (N_1200,N_31,N_966);
and U1201 (N_1201,In_1058,In_1600);
nor U1202 (N_1202,N_634,N_132);
xor U1203 (N_1203,N_611,N_904);
xnor U1204 (N_1204,N_246,N_262);
and U1205 (N_1205,N_158,In_2023);
nand U1206 (N_1206,In_859,N_64);
nor U1207 (N_1207,In_749,In_1263);
xnor U1208 (N_1208,N_988,N_414);
or U1209 (N_1209,N_739,N_682);
xor U1210 (N_1210,N_313,In_1456);
and U1211 (N_1211,N_531,N_108);
nand U1212 (N_1212,In_1127,In_179);
xnor U1213 (N_1213,In_219,N_412);
or U1214 (N_1214,In_1037,N_847);
nand U1215 (N_1215,N_541,N_692);
nand U1216 (N_1216,In_330,N_29);
nand U1217 (N_1217,N_470,In_1258);
or U1218 (N_1218,N_364,N_245);
or U1219 (N_1219,N_948,N_829);
and U1220 (N_1220,N_34,N_361);
nor U1221 (N_1221,In_17,N_298);
nor U1222 (N_1222,N_40,N_317);
or U1223 (N_1223,N_475,N_968);
nor U1224 (N_1224,N_710,N_978);
or U1225 (N_1225,N_511,N_84);
and U1226 (N_1226,N_326,N_21);
or U1227 (N_1227,N_709,N_8);
nor U1228 (N_1228,N_669,N_582);
nand U1229 (N_1229,In_1555,In_650);
xor U1230 (N_1230,N_160,N_375);
xor U1231 (N_1231,In_965,In_1061);
xnor U1232 (N_1232,In_857,In_573);
and U1233 (N_1233,N_957,N_719);
nor U1234 (N_1234,N_78,N_699);
or U1235 (N_1235,N_314,In_152);
nor U1236 (N_1236,N_96,N_515);
xor U1237 (N_1237,N_343,N_127);
xnor U1238 (N_1238,In_613,N_866);
nor U1239 (N_1239,N_122,N_53);
nand U1240 (N_1240,N_929,N_55);
xor U1241 (N_1241,N_890,N_779);
or U1242 (N_1242,In_1988,N_999);
xor U1243 (N_1243,N_737,In_387);
nor U1244 (N_1244,N_48,In_1614);
nor U1245 (N_1245,N_166,N_826);
or U1246 (N_1246,N_207,N_92);
nor U1247 (N_1247,N_346,N_184);
or U1248 (N_1248,N_177,In_2024);
or U1249 (N_1249,In_1586,N_477);
or U1250 (N_1250,In_720,N_869);
or U1251 (N_1251,N_821,N_173);
nand U1252 (N_1252,N_642,In_438);
and U1253 (N_1253,N_498,In_1815);
xor U1254 (N_1254,N_953,In_2364);
xor U1255 (N_1255,N_581,N_810);
or U1256 (N_1256,In_2433,N_755);
xor U1257 (N_1257,N_372,N_65);
or U1258 (N_1258,In_2336,N_686);
and U1259 (N_1259,N_86,In_2193);
nand U1260 (N_1260,N_146,N_1);
xor U1261 (N_1261,In_410,In_531);
nor U1262 (N_1262,In_567,In_284);
or U1263 (N_1263,In_1509,N_50);
nor U1264 (N_1264,N_456,In_731);
xnor U1265 (N_1265,N_756,N_212);
and U1266 (N_1266,N_722,N_180);
nand U1267 (N_1267,N_955,N_570);
nand U1268 (N_1268,N_380,N_561);
nor U1269 (N_1269,In_933,N_584);
xnor U1270 (N_1270,In_1183,In_1333);
nand U1271 (N_1271,N_249,In_309);
nor U1272 (N_1272,N_320,In_1124);
or U1273 (N_1273,In_1580,N_450);
xnor U1274 (N_1274,N_483,N_444);
or U1275 (N_1275,N_913,N_248);
or U1276 (N_1276,N_557,N_405);
xor U1277 (N_1277,In_877,N_381);
nand U1278 (N_1278,In_464,In_674);
nor U1279 (N_1279,N_295,In_2435);
or U1280 (N_1280,N_423,In_1789);
nand U1281 (N_1281,N_885,In_1868);
and U1282 (N_1282,N_449,N_931);
xnor U1283 (N_1283,In_2206,In_1757);
nor U1284 (N_1284,N_676,N_777);
or U1285 (N_1285,N_908,In_1479);
xnor U1286 (N_1286,In_1716,In_575);
nor U1287 (N_1287,N_817,N_126);
or U1288 (N_1288,In_1170,In_2483);
nor U1289 (N_1289,In_1145,N_548);
and U1290 (N_1290,In_2269,N_59);
and U1291 (N_1291,N_106,N_629);
and U1292 (N_1292,N_12,N_338);
and U1293 (N_1293,In_166,In_1577);
nand U1294 (N_1294,In_1416,N_292);
nor U1295 (N_1295,In_50,In_875);
or U1296 (N_1296,N_188,In_1060);
nand U1297 (N_1297,N_846,In_2422);
and U1298 (N_1298,N_89,N_90);
or U1299 (N_1299,N_386,N_263);
or U1300 (N_1300,N_113,In_1090);
xnor U1301 (N_1301,In_1408,N_785);
or U1302 (N_1302,N_321,N_573);
and U1303 (N_1303,In_2441,In_2395);
and U1304 (N_1304,In_928,In_127);
or U1305 (N_1305,N_308,N_624);
and U1306 (N_1306,N_324,N_13);
nor U1307 (N_1307,In_1220,In_2046);
nand U1308 (N_1308,In_1353,N_631);
xor U1309 (N_1309,N_862,In_1517);
and U1310 (N_1310,N_693,N_327);
xor U1311 (N_1311,In_2438,In_2013);
nor U1312 (N_1312,In_707,N_51);
and U1313 (N_1313,In_408,N_974);
nand U1314 (N_1314,N_93,In_1313);
xor U1315 (N_1315,N_812,N_71);
xor U1316 (N_1316,In_2488,N_804);
and U1317 (N_1317,In_107,N_895);
xor U1318 (N_1318,N_288,In_461);
or U1319 (N_1319,In_1804,In_1499);
or U1320 (N_1320,In_923,N_410);
and U1321 (N_1321,In_2347,N_94);
nand U1322 (N_1322,N_256,N_506);
or U1323 (N_1323,N_402,N_363);
and U1324 (N_1324,N_214,In_110);
nand U1325 (N_1325,N_985,N_123);
nor U1326 (N_1326,N_816,In_764);
nand U1327 (N_1327,N_598,N_305);
or U1328 (N_1328,N_850,N_754);
xnor U1329 (N_1329,In_1832,N_674);
and U1330 (N_1330,In_2213,N_23);
nand U1331 (N_1331,In_1062,N_773);
nor U1332 (N_1332,N_351,In_1302);
xnor U1333 (N_1333,N_171,In_1566);
nor U1334 (N_1334,N_909,N_640);
or U1335 (N_1335,N_339,In_2449);
or U1336 (N_1336,N_252,N_861);
nand U1337 (N_1337,N_508,N_975);
nand U1338 (N_1338,In_1528,N_445);
nor U1339 (N_1339,N_946,N_107);
xor U1340 (N_1340,N_644,In_1065);
and U1341 (N_1341,In_1198,N_293);
nand U1342 (N_1342,N_529,N_936);
or U1343 (N_1343,N_604,In_418);
or U1344 (N_1344,N_417,In_1133);
xnor U1345 (N_1345,N_760,N_646);
or U1346 (N_1346,N_986,N_290);
xnor U1347 (N_1347,N_399,N_101);
nor U1348 (N_1348,N_964,In_592);
or U1349 (N_1349,In_895,N_532);
or U1350 (N_1350,N_467,N_476);
or U1351 (N_1351,In_2382,N_149);
nor U1352 (N_1352,N_54,N_758);
nor U1353 (N_1353,N_606,In_1457);
xor U1354 (N_1354,N_852,In_2429);
and U1355 (N_1355,N_996,N_675);
xor U1356 (N_1356,N_398,N_404);
or U1357 (N_1357,N_789,In_1039);
nor U1358 (N_1358,In_430,N_110);
nor U1359 (N_1359,N_807,N_299);
xnor U1360 (N_1360,N_874,N_535);
nand U1361 (N_1361,In_551,In_568);
nor U1362 (N_1362,N_959,In_1782);
and U1363 (N_1363,N_727,In_1995);
xnor U1364 (N_1364,N_670,In_206);
xnor U1365 (N_1365,N_79,In_2465);
xor U1366 (N_1366,N_373,N_734);
and U1367 (N_1367,N_556,In_1717);
nor U1368 (N_1368,N_41,In_2241);
nor U1369 (N_1369,N_514,N_947);
xnor U1370 (N_1370,In_1694,N_815);
nand U1371 (N_1371,N_138,N_513);
or U1372 (N_1372,In_136,N_767);
xor U1373 (N_1373,N_661,N_118);
nor U1374 (N_1374,N_678,N_740);
nor U1375 (N_1375,N_504,N_831);
xnor U1376 (N_1376,N_316,In_2250);
nand U1377 (N_1377,In_1421,N_823);
xnor U1378 (N_1378,In_1477,N_918);
nor U1379 (N_1379,In_1704,N_711);
and U1380 (N_1380,N_259,N_454);
nand U1381 (N_1381,In_1807,N_4);
and U1382 (N_1382,N_318,In_1536);
and U1383 (N_1383,In_94,In_640);
and U1384 (N_1384,N_484,In_724);
xnor U1385 (N_1385,N_849,N_463);
xnor U1386 (N_1386,In_629,N_413);
and U1387 (N_1387,N_237,N_534);
or U1388 (N_1388,N_927,N_209);
and U1389 (N_1389,N_883,N_650);
nand U1390 (N_1390,In_137,N_194);
or U1391 (N_1391,N_691,In_1004);
xor U1392 (N_1392,In_2290,N_200);
and U1393 (N_1393,N_411,In_488);
nand U1394 (N_1394,N_747,N_917);
and U1395 (N_1395,In_61,N_733);
or U1396 (N_1396,N_344,N_944);
and U1397 (N_1397,N_853,N_424);
and U1398 (N_1398,In_1264,N_824);
and U1399 (N_1399,N_28,N_383);
and U1400 (N_1400,N_937,N_447);
nand U1401 (N_1401,N_163,N_187);
or U1402 (N_1402,N_864,N_844);
nor U1403 (N_1403,N_358,N_886);
xor U1404 (N_1404,N_938,N_517);
xor U1405 (N_1405,N_422,In_1948);
nor U1406 (N_1406,N_793,N_577);
nand U1407 (N_1407,In_1453,N_528);
and U1408 (N_1408,In_1496,N_128);
nor U1409 (N_1409,N_426,In_2490);
and U1410 (N_1410,N_989,In_1542);
and U1411 (N_1411,In_1588,N_641);
or U1412 (N_1412,N_768,In_626);
and U1413 (N_1413,N_897,N_842);
or U1414 (N_1414,In_1554,In_1727);
or U1415 (N_1415,In_585,N_20);
xor U1416 (N_1416,In_1639,In_2328);
xnor U1417 (N_1417,N_67,In_1377);
xor U1418 (N_1418,In_518,N_165);
nor U1419 (N_1419,N_731,N_704);
xnor U1420 (N_1420,N_428,In_903);
and U1421 (N_1421,In_1280,In_1834);
xnor U1422 (N_1422,N_593,N_24);
or U1423 (N_1423,N_934,N_965);
and U1424 (N_1424,In_1320,In_194);
xnor U1425 (N_1425,N_623,N_453);
nor U1426 (N_1426,In_153,N_603);
nand U1427 (N_1427,In_1473,In_2394);
and U1428 (N_1428,N_455,In_1021);
or U1429 (N_1429,N_820,N_210);
or U1430 (N_1430,N_905,N_643);
and U1431 (N_1431,N_627,N_167);
and U1432 (N_1432,N_848,In_2084);
or U1433 (N_1433,In_1125,N_233);
and U1434 (N_1434,In_737,N_507);
nand U1435 (N_1435,N_858,N_66);
or U1436 (N_1436,N_972,N_408);
and U1437 (N_1437,N_545,N_677);
or U1438 (N_1438,N_68,In_2242);
nor U1439 (N_1439,N_698,N_117);
and U1440 (N_1440,In_1655,N_459);
nor U1441 (N_1441,N_610,N_619);
nand U1442 (N_1442,N_147,N_170);
nand U1443 (N_1443,N_657,N_750);
and U1444 (N_1444,In_1470,N_990);
nand U1445 (N_1445,N_806,N_951);
or U1446 (N_1446,In_1329,In_1365);
xnor U1447 (N_1447,N_876,N_851);
nor U1448 (N_1448,N_25,In_1107);
nand U1449 (N_1449,N_967,N_932);
or U1450 (N_1450,N_997,N_226);
nand U1451 (N_1451,N_618,N_752);
nor U1452 (N_1452,N_303,In_1824);
nor U1453 (N_1453,N_902,In_1778);
and U1454 (N_1454,In_856,N_921);
and U1455 (N_1455,In_2047,N_780);
nor U1456 (N_1456,N_878,N_827);
nor U1457 (N_1457,N_567,In_102);
xnor U1458 (N_1458,N_801,N_834);
xor U1459 (N_1459,N_283,N_868);
nand U1460 (N_1460,In_354,In_926);
or U1461 (N_1461,N_998,In_1612);
nor U1462 (N_1462,N_204,N_718);
nand U1463 (N_1463,In_2079,N_638);
xnor U1464 (N_1464,In_1775,In_454);
nor U1465 (N_1465,N_401,N_600);
and U1466 (N_1466,N_217,N_571);
nor U1467 (N_1467,In_510,In_1056);
nand U1468 (N_1468,N_129,In_5);
and U1469 (N_1469,In_1601,N_617);
xnor U1470 (N_1470,N_352,In_482);
nand U1471 (N_1471,In_1380,N_907);
and U1472 (N_1472,N_87,In_1689);
nor U1473 (N_1473,N_647,N_977);
xor U1474 (N_1474,N_775,N_223);
nand U1475 (N_1475,In_1123,N_607);
and U1476 (N_1476,In_1176,In_1642);
and U1477 (N_1477,N_703,In_1726);
xor U1478 (N_1478,N_697,N_473);
nand U1479 (N_1479,In_2446,In_401);
nor U1480 (N_1480,In_1278,In_2126);
or U1481 (N_1481,N_56,N_257);
and U1482 (N_1482,N_579,In_554);
nor U1483 (N_1483,N_833,In_1305);
or U1484 (N_1484,N_549,In_1981);
and U1485 (N_1485,N_616,In_766);
or U1486 (N_1486,N_341,In_1019);
nand U1487 (N_1487,N_550,N_435);
and U1488 (N_1488,N_193,N_296);
xor U1489 (N_1489,N_181,In_969);
nor U1490 (N_1490,N_880,In_493);
and U1491 (N_1491,In_1637,N_323);
xnor U1492 (N_1492,In_1590,N_625);
xnor U1493 (N_1493,In_1711,N_705);
nor U1494 (N_1494,N_894,N_46);
xnor U1495 (N_1495,N_493,In_2235);
and U1496 (N_1496,N_843,N_594);
and U1497 (N_1497,N_995,N_732);
and U1498 (N_1498,N_694,N_72);
and U1499 (N_1499,In_334,N_765);
nor U1500 (N_1500,N_583,N_192);
and U1501 (N_1501,N_609,In_434);
xnor U1502 (N_1502,N_568,N_896);
and U1503 (N_1503,In_1845,N_984);
or U1504 (N_1504,In_673,N_155);
nand U1505 (N_1505,N_496,In_1609);
and U1506 (N_1506,N_856,In_2131);
nor U1507 (N_1507,In_890,N_418);
nand U1508 (N_1508,N_328,N_109);
or U1509 (N_1509,N_482,N_7);
nor U1510 (N_1510,N_137,In_993);
and U1511 (N_1511,N_543,In_1788);
and U1512 (N_1512,In_2125,N_818);
and U1513 (N_1513,N_377,N_366);
xor U1514 (N_1514,In_186,N_702);
nand U1515 (N_1515,In_666,N_668);
and U1516 (N_1516,N_239,N_797);
xor U1517 (N_1517,In_2027,In_1140);
xnor U1518 (N_1518,In_1256,N_558);
nand U1519 (N_1519,N_813,N_666);
and U1520 (N_1520,N_763,In_264);
and U1521 (N_1521,In_2207,In_872);
nand U1522 (N_1522,N_247,N_335);
nor U1523 (N_1523,N_231,N_52);
nand U1524 (N_1524,N_220,N_488);
and U1525 (N_1525,N_287,In_1211);
nor U1526 (N_1526,N_485,N_169);
nand U1527 (N_1527,N_721,N_240);
nor U1528 (N_1528,N_251,N_33);
xnor U1529 (N_1529,In_1737,N_14);
xnor U1530 (N_1530,In_1750,In_808);
or U1531 (N_1531,In_2315,N_236);
nand U1532 (N_1532,N_736,N_700);
and U1533 (N_1533,In_286,N_431);
and U1534 (N_1534,N_599,N_133);
nor U1535 (N_1535,N_301,In_1495);
nor U1536 (N_1536,N_546,N_274);
xnor U1537 (N_1537,N_690,N_219);
xor U1538 (N_1538,N_562,In_1144);
or U1539 (N_1539,In_1777,In_2064);
xor U1540 (N_1540,N_919,N_673);
or U1541 (N_1541,N_554,In_2087);
or U1542 (N_1542,N_585,N_520);
nand U1543 (N_1543,In_111,N_451);
nor U1544 (N_1544,N_140,N_920);
nor U1545 (N_1545,N_706,In_639);
and U1546 (N_1546,N_37,N_542);
nor U1547 (N_1547,In_1947,N_510);
nor U1548 (N_1548,In_1643,N_415);
xor U1549 (N_1549,N_837,N_601);
nor U1550 (N_1550,N_342,In_2201);
nand U1551 (N_1551,N_981,N_289);
nand U1552 (N_1552,N_211,N_11);
or U1553 (N_1553,In_996,N_393);
and U1554 (N_1554,N_83,N_969);
nand U1555 (N_1555,N_553,N_873);
or U1556 (N_1556,In_1259,N_836);
xor U1557 (N_1557,In_670,In_553);
xnor U1558 (N_1558,N_330,In_1179);
xor U1559 (N_1559,In_2153,N_963);
or U1560 (N_1560,In_2352,N_595);
nor U1561 (N_1561,N_632,N_203);
and U1562 (N_1562,In_525,N_125);
and U1563 (N_1563,N_799,N_480);
or U1564 (N_1564,In_1846,In_265);
nand U1565 (N_1565,N_655,N_434);
or U1566 (N_1566,N_524,N_759);
xor U1567 (N_1567,N_353,N_684);
nand U1568 (N_1568,In_297,N_130);
nand U1569 (N_1569,In_689,In_477);
and U1570 (N_1570,N_605,N_378);
xnor U1571 (N_1571,In_125,N_279);
or U1572 (N_1572,N_466,N_464);
and U1573 (N_1573,N_589,In_1712);
or U1574 (N_1574,N_397,In_478);
nor U1575 (N_1575,In_1403,In_203);
and U1576 (N_1576,N_80,N_2);
or U1577 (N_1577,N_60,N_516);
or U1578 (N_1578,N_680,In_2243);
nand U1579 (N_1579,In_2268,N_859);
nand U1580 (N_1580,N_421,In_561);
nand U1581 (N_1581,N_870,In_1581);
or U1582 (N_1582,N_724,In_1192);
and U1583 (N_1583,N_819,In_696);
nor U1584 (N_1584,N_69,N_340);
or U1585 (N_1585,In_2233,In_1411);
and U1586 (N_1586,In_1607,N_742);
or U1587 (N_1587,In_1515,N_159);
and U1588 (N_1588,N_168,N_6);
nand U1589 (N_1589,In_1454,In_1688);
xnor U1590 (N_1590,N_656,N_284);
nand U1591 (N_1591,In_589,In_814);
nand U1592 (N_1592,N_309,In_663);
nand U1593 (N_1593,N_16,N_960);
or U1594 (N_1594,N_91,N_888);
or U1595 (N_1595,N_825,In_2152);
and U1596 (N_1596,In_263,N_329);
nor U1597 (N_1597,In_1285,N_911);
nand U1598 (N_1598,N_891,In_1805);
or U1599 (N_1599,In_841,N_229);
and U1600 (N_1600,In_2392,N_935);
and U1601 (N_1601,N_150,N_788);
xnor U1602 (N_1602,In_1959,N_222);
or U1603 (N_1603,In_2182,In_2390);
xnor U1604 (N_1604,N_822,N_474);
or U1605 (N_1605,N_749,In_741);
xor U1606 (N_1606,N_216,In_1779);
or U1607 (N_1607,N_75,N_254);
and U1608 (N_1608,N_9,N_716);
or U1609 (N_1609,In_1005,N_354);
or U1610 (N_1610,N_572,In_582);
and U1611 (N_1611,N_111,N_42);
nand U1612 (N_1612,N_728,N_664);
nor U1613 (N_1613,In_399,In_1105);
and U1614 (N_1614,N_100,In_2479);
or U1615 (N_1615,N_469,N_745);
nor U1616 (N_1616,N_243,In_998);
xnor U1617 (N_1617,N_99,In_1628);
xnor U1618 (N_1618,In_2189,In_1368);
xor U1619 (N_1619,N_297,In_2012);
nand U1620 (N_1620,N_771,In_602);
nand U1621 (N_1621,N_790,N_189);
or U1622 (N_1622,N_555,In_1374);
xnor U1623 (N_1623,N_922,In_290);
xnor U1624 (N_1624,N_942,N_266);
or U1625 (N_1625,In_502,N_539);
xnor U1626 (N_1626,In_1398,N_30);
and U1627 (N_1627,N_420,N_662);
xnor U1628 (N_1628,N_199,In_1097);
or U1629 (N_1629,N_500,N_863);
nor U1630 (N_1630,N_407,N_712);
nand U1631 (N_1631,In_2050,N_269);
xor U1632 (N_1632,N_227,N_179);
and U1633 (N_1633,In_2453,N_776);
or U1634 (N_1634,In_480,In_826);
and U1635 (N_1635,In_311,N_586);
nor U1636 (N_1636,N_726,N_564);
xnor U1637 (N_1637,N_794,N_950);
nand U1638 (N_1638,In_1728,N_333);
nor U1639 (N_1639,In_2388,N_954);
nor U1640 (N_1640,In_233,N_738);
xnor U1641 (N_1641,N_334,N_97);
nand U1642 (N_1642,In_2371,N_438);
nor U1643 (N_1643,In_54,N_350);
nand U1644 (N_1644,In_1401,In_1174);
and U1645 (N_1645,In_1059,N_452);
nand U1646 (N_1646,N_468,N_319);
nor U1647 (N_1647,N_588,In_1040);
nand U1648 (N_1648,N_832,In_135);
nand U1649 (N_1649,In_828,N_26);
nand U1650 (N_1650,N_119,N_809);
nor U1651 (N_1651,In_412,N_774);
or U1652 (N_1652,N_840,In_2384);
or U1653 (N_1653,In_1608,N_224);
nor U1654 (N_1654,In_1878,N_260);
or U1655 (N_1655,N_961,N_302);
xnor U1656 (N_1656,In_1201,In_2471);
xor U1657 (N_1657,N_337,N_494);
nor U1658 (N_1658,N_958,N_764);
or U1659 (N_1659,N_628,In_836);
xnor U1660 (N_1660,In_2470,N_36);
or U1661 (N_1661,N_653,In_646);
and U1662 (N_1662,N_103,In_285);
nor U1663 (N_1663,N_501,N_772);
nand U1664 (N_1664,N_559,N_672);
or U1665 (N_1665,In_2477,In_1029);
nand U1666 (N_1666,N_753,N_994);
nand U1667 (N_1667,N_270,N_910);
or U1668 (N_1668,N_923,In_1433);
or U1669 (N_1669,In_1167,N_839);
and U1670 (N_1670,N_892,In_170);
xnor U1671 (N_1671,N_88,N_392);
and U1672 (N_1672,N_49,N_560);
xor U1673 (N_1673,In_1226,N_371);
xor U1674 (N_1674,In_831,In_1079);
nand U1675 (N_1675,N_993,N_465);
and U1676 (N_1676,In_191,N_580);
xor U1677 (N_1677,N_258,N_875);
or U1678 (N_1678,N_980,In_310);
or U1679 (N_1679,In_456,N_278);
and U1680 (N_1680,N_436,In_2325);
xor U1681 (N_1681,N_47,In_1986);
xor U1682 (N_1682,N_654,N_808);
xnor U1683 (N_1683,N_312,N_282);
xnor U1684 (N_1684,In_2111,N_3);
xnor U1685 (N_1685,In_122,N_526);
and U1686 (N_1686,N_70,In_1236);
nor U1687 (N_1687,N_300,N_906);
or U1688 (N_1688,N_770,N_385);
and U1689 (N_1689,In_451,N_58);
nor U1690 (N_1690,N_915,In_1362);
nand U1691 (N_1691,N_440,In_651);
and U1692 (N_1692,In_2016,N_992);
nand U1693 (N_1693,In_1075,N_39);
nor U1694 (N_1694,N_114,N_273);
xor U1695 (N_1695,N_139,N_687);
and U1696 (N_1696,N_362,N_518);
nand U1697 (N_1697,N_162,N_82);
nor U1698 (N_1698,N_871,N_622);
nor U1699 (N_1699,N_235,N_608);
or U1700 (N_1700,In_1946,N_940);
xor U1701 (N_1701,N_492,In_1490);
nand U1702 (N_1702,N_331,In_1153);
and U1703 (N_1703,N_400,N_357);
nand U1704 (N_1704,N_242,N_811);
or U1705 (N_1705,N_307,In_60);
and U1706 (N_1706,N_914,In_1027);
and U1707 (N_1707,N_491,In_2177);
nor U1708 (N_1708,In_2038,N_621);
or U1709 (N_1709,N_805,N_659);
nand U1710 (N_1710,In_1870,In_2192);
nor U1711 (N_1711,N_5,N_61);
and U1712 (N_1712,N_376,N_406);
and U1713 (N_1713,N_161,In_2277);
and U1714 (N_1714,In_1762,In_148);
and U1715 (N_1715,N_613,N_798);
nor U1716 (N_1716,In_997,In_2199);
xnor U1717 (N_1717,In_653,N_195);
nand U1718 (N_1718,N_769,N_145);
xor U1719 (N_1719,N_332,N_225);
or U1720 (N_1720,N_427,N_720);
xnor U1721 (N_1721,N_176,In_470);
nor U1722 (N_1722,N_930,N_391);
or U1723 (N_1723,In_2238,N_652);
nor U1724 (N_1724,In_221,N_120);
and U1725 (N_1725,N_43,N_271);
nand U1726 (N_1726,In_1282,N_943);
and U1727 (N_1727,N_403,N_190);
xor U1728 (N_1728,N_527,In_1139);
nor U1729 (N_1729,In_2343,N_899);
nor U1730 (N_1730,N_38,N_949);
or U1731 (N_1731,N_153,In_532);
nand U1732 (N_1732,In_1630,N_487);
or U1733 (N_1733,N_882,In_951);
nor U1734 (N_1734,N_854,In_397);
nand U1735 (N_1735,In_2469,In_1984);
or U1736 (N_1736,N_359,In_2304);
nor U1737 (N_1737,N_800,N_182);
and U1738 (N_1738,In_768,N_389);
or U1739 (N_1739,In_30,N_889);
or U1740 (N_1740,N_796,N_658);
or U1741 (N_1741,N_310,In_260);
xor U1742 (N_1742,In_1463,N_865);
nor U1743 (N_1743,N_751,N_512);
and U1744 (N_1744,In_1734,In_1237);
nor U1745 (N_1745,N_973,In_358);
nor U1746 (N_1746,N_787,N_255);
xnor U1747 (N_1747,N_489,N_154);
and U1748 (N_1748,In_1963,In_2461);
and U1749 (N_1749,In_1049,N_838);
and U1750 (N_1750,N_678,In_688);
nor U1751 (N_1751,N_330,N_116);
nor U1752 (N_1752,N_894,N_315);
nor U1753 (N_1753,In_1402,N_27);
or U1754 (N_1754,N_397,N_873);
nor U1755 (N_1755,In_2422,N_470);
and U1756 (N_1756,In_179,N_942);
or U1757 (N_1757,In_1139,In_311);
and U1758 (N_1758,In_1586,N_318);
nor U1759 (N_1759,N_188,N_558);
or U1760 (N_1760,N_155,In_2186);
and U1761 (N_1761,N_739,N_851);
or U1762 (N_1762,N_497,In_2449);
nor U1763 (N_1763,In_915,N_502);
or U1764 (N_1764,N_378,In_464);
nand U1765 (N_1765,In_1717,N_103);
or U1766 (N_1766,N_206,N_122);
xnor U1767 (N_1767,In_1433,N_977);
nor U1768 (N_1768,In_1061,In_17);
and U1769 (N_1769,N_640,In_903);
nor U1770 (N_1770,In_2199,In_760);
or U1771 (N_1771,N_189,N_795);
xor U1772 (N_1772,In_17,N_193);
nor U1773 (N_1773,N_871,In_1922);
xnor U1774 (N_1774,N_35,N_218);
nor U1775 (N_1775,In_179,In_510);
nor U1776 (N_1776,N_135,N_837);
or U1777 (N_1777,N_0,N_918);
xnor U1778 (N_1778,N_958,In_2125);
xnor U1779 (N_1779,In_1636,In_1046);
and U1780 (N_1780,N_646,In_653);
and U1781 (N_1781,In_111,N_702);
or U1782 (N_1782,N_870,N_560);
or U1783 (N_1783,N_2,In_1804);
nor U1784 (N_1784,In_1145,N_70);
xnor U1785 (N_1785,In_1056,N_666);
or U1786 (N_1786,N_681,N_249);
xnor U1787 (N_1787,N_45,N_346);
nor U1788 (N_1788,In_1824,N_416);
or U1789 (N_1789,N_960,N_871);
nand U1790 (N_1790,In_1600,N_426);
nor U1791 (N_1791,N_113,In_1227);
or U1792 (N_1792,In_1107,In_1176);
xnor U1793 (N_1793,N_294,N_938);
and U1794 (N_1794,N_512,N_611);
nand U1795 (N_1795,In_1256,In_735);
or U1796 (N_1796,In_2329,In_2206);
and U1797 (N_1797,In_354,N_789);
nor U1798 (N_1798,N_879,N_523);
or U1799 (N_1799,N_286,N_453);
or U1800 (N_1800,N_655,N_366);
nor U1801 (N_1801,In_705,N_618);
nor U1802 (N_1802,In_480,N_419);
nor U1803 (N_1803,N_151,In_1892);
nand U1804 (N_1804,In_1824,N_665);
nand U1805 (N_1805,N_40,N_986);
or U1806 (N_1806,In_284,N_389);
nand U1807 (N_1807,N_144,In_110);
xor U1808 (N_1808,N_118,N_13);
nor U1809 (N_1809,In_1614,N_941);
nand U1810 (N_1810,In_696,N_242);
nor U1811 (N_1811,N_199,N_156);
nor U1812 (N_1812,In_1380,N_676);
nand U1813 (N_1813,N_589,N_363);
nand U1814 (N_1814,N_48,N_498);
and U1815 (N_1815,N_69,In_2363);
and U1816 (N_1816,N_163,N_323);
and U1817 (N_1817,N_389,N_258);
nand U1818 (N_1818,N_833,In_1496);
nor U1819 (N_1819,In_1170,N_328);
or U1820 (N_1820,N_176,In_1614);
nand U1821 (N_1821,N_903,N_500);
xnor U1822 (N_1822,In_1139,N_380);
xor U1823 (N_1823,N_705,N_340);
or U1824 (N_1824,N_837,N_699);
or U1825 (N_1825,N_36,N_831);
xor U1826 (N_1826,In_1343,In_191);
nand U1827 (N_1827,N_951,N_629);
xor U1828 (N_1828,N_325,N_703);
xnor U1829 (N_1829,N_487,N_40);
nand U1830 (N_1830,N_79,N_180);
nor U1831 (N_1831,N_323,N_200);
or U1832 (N_1832,N_555,N_405);
or U1833 (N_1833,N_783,In_203);
xor U1834 (N_1834,N_436,In_602);
nand U1835 (N_1835,N_176,In_2047);
nor U1836 (N_1836,In_2384,In_1065);
and U1837 (N_1837,In_1079,N_951);
nor U1838 (N_1838,N_478,In_1580);
or U1839 (N_1839,In_185,N_242);
and U1840 (N_1840,In_497,N_901);
and U1841 (N_1841,N_479,N_298);
xnor U1842 (N_1842,N_79,N_317);
and U1843 (N_1843,N_852,N_947);
or U1844 (N_1844,N_231,N_419);
nand U1845 (N_1845,In_264,N_747);
and U1846 (N_1846,N_609,N_109);
nand U1847 (N_1847,In_2269,In_1948);
xnor U1848 (N_1848,N_384,In_532);
nor U1849 (N_1849,In_2280,N_280);
and U1850 (N_1850,N_641,N_698);
nand U1851 (N_1851,N_869,N_427);
and U1852 (N_1852,N_982,N_786);
nand U1853 (N_1853,N_320,In_1101);
and U1854 (N_1854,In_720,N_521);
or U1855 (N_1855,N_846,In_2269);
xnor U1856 (N_1856,N_275,N_433);
nand U1857 (N_1857,N_93,N_984);
and U1858 (N_1858,In_1351,In_1577);
or U1859 (N_1859,N_6,N_579);
or U1860 (N_1860,N_387,N_62);
and U1861 (N_1861,N_686,N_137);
nand U1862 (N_1862,N_346,In_2295);
and U1863 (N_1863,N_110,In_2242);
nand U1864 (N_1864,N_419,N_215);
and U1865 (N_1865,N_377,N_605);
nor U1866 (N_1866,In_914,In_969);
nor U1867 (N_1867,In_824,In_206);
nor U1868 (N_1868,In_1845,In_148);
and U1869 (N_1869,N_87,N_37);
xor U1870 (N_1870,N_395,N_497);
or U1871 (N_1871,N_102,In_2125);
nand U1872 (N_1872,N_364,N_901);
nor U1873 (N_1873,N_966,N_476);
and U1874 (N_1874,N_219,In_1495);
or U1875 (N_1875,In_1594,In_2347);
nor U1876 (N_1876,N_784,N_398);
xor U1877 (N_1877,N_191,N_633);
xnor U1878 (N_1878,In_2490,N_465);
or U1879 (N_1879,In_1083,N_116);
and U1880 (N_1880,In_1892,In_998);
nand U1881 (N_1881,N_227,N_393);
or U1882 (N_1882,In_1694,In_629);
xnor U1883 (N_1883,N_432,In_1655);
or U1884 (N_1884,N_150,N_340);
xnor U1885 (N_1885,In_2449,N_329);
or U1886 (N_1886,N_513,In_1403);
nand U1887 (N_1887,N_587,N_112);
or U1888 (N_1888,N_950,In_1553);
xor U1889 (N_1889,In_1019,N_995);
and U1890 (N_1890,N_332,N_446);
nand U1891 (N_1891,N_973,N_468);
nand U1892 (N_1892,In_1726,N_327);
xor U1893 (N_1893,In_219,N_51);
nor U1894 (N_1894,In_1167,In_497);
xnor U1895 (N_1895,N_69,N_975);
nand U1896 (N_1896,N_31,In_68);
xor U1897 (N_1897,N_419,N_865);
and U1898 (N_1898,In_534,In_290);
nand U1899 (N_1899,N_73,In_639);
nand U1900 (N_1900,N_478,N_784);
nand U1901 (N_1901,In_1385,N_33);
or U1902 (N_1902,In_1416,N_115);
xor U1903 (N_1903,N_579,In_1421);
xor U1904 (N_1904,N_125,In_286);
xor U1905 (N_1905,In_1864,In_2443);
nand U1906 (N_1906,N_463,In_1090);
xor U1907 (N_1907,In_408,In_2290);
and U1908 (N_1908,In_1132,N_890);
or U1909 (N_1909,N_458,N_246);
nor U1910 (N_1910,In_1959,In_663);
nand U1911 (N_1911,N_987,In_1947);
and U1912 (N_1912,N_656,N_632);
and U1913 (N_1913,In_2384,N_944);
xor U1914 (N_1914,In_265,In_2269);
nand U1915 (N_1915,N_753,N_239);
xnor U1916 (N_1916,N_275,N_174);
nor U1917 (N_1917,N_748,In_2090);
or U1918 (N_1918,N_180,N_864);
nand U1919 (N_1919,N_877,In_688);
and U1920 (N_1920,N_867,N_19);
or U1921 (N_1921,N_703,In_2295);
nor U1922 (N_1922,N_828,In_397);
nor U1923 (N_1923,N_925,In_203);
and U1924 (N_1924,N_235,N_61);
xnor U1925 (N_1925,N_942,N_339);
or U1926 (N_1926,N_903,In_1453);
nor U1927 (N_1927,In_285,N_228);
xnor U1928 (N_1928,N_548,N_256);
and U1929 (N_1929,In_525,In_997);
and U1930 (N_1930,In_1343,N_881);
xnor U1931 (N_1931,In_2268,N_837);
xor U1932 (N_1932,N_676,In_233);
xnor U1933 (N_1933,N_791,N_721);
and U1934 (N_1934,In_2394,In_186);
nand U1935 (N_1935,N_831,N_405);
nand U1936 (N_1936,In_831,N_4);
nor U1937 (N_1937,N_993,N_612);
xor U1938 (N_1938,N_273,N_152);
xnor U1939 (N_1939,N_708,N_704);
xnor U1940 (N_1940,N_379,N_234);
and U1941 (N_1941,In_1065,N_652);
xor U1942 (N_1942,In_2433,N_337);
or U1943 (N_1943,In_221,N_204);
xor U1944 (N_1944,In_2488,N_163);
or U1945 (N_1945,In_1788,N_549);
or U1946 (N_1946,N_582,In_1728);
or U1947 (N_1947,N_976,N_841);
nor U1948 (N_1948,N_582,N_252);
xnor U1949 (N_1949,N_228,N_430);
and U1950 (N_1950,N_661,N_561);
or U1951 (N_1951,In_2400,N_684);
nand U1952 (N_1952,In_1655,N_412);
or U1953 (N_1953,N_473,N_349);
and U1954 (N_1954,N_755,N_397);
or U1955 (N_1955,N_598,N_786);
or U1956 (N_1956,N_367,In_646);
and U1957 (N_1957,N_201,N_341);
nor U1958 (N_1958,N_279,In_780);
nor U1959 (N_1959,N_36,N_691);
xnor U1960 (N_1960,N_915,In_310);
nor U1961 (N_1961,N_685,In_1642);
xnor U1962 (N_1962,N_604,In_2471);
nor U1963 (N_1963,In_1778,In_1719);
xor U1964 (N_1964,N_549,N_947);
nor U1965 (N_1965,N_896,In_2371);
or U1966 (N_1966,N_50,N_763);
or U1967 (N_1967,In_2046,N_490);
or U1968 (N_1968,N_95,N_362);
xnor U1969 (N_1969,N_519,In_1630);
and U1970 (N_1970,In_2277,N_40);
nand U1971 (N_1971,N_198,N_441);
nand U1972 (N_1972,In_1433,In_666);
nand U1973 (N_1973,In_1496,In_2235);
xnor U1974 (N_1974,In_1517,In_1079);
xnor U1975 (N_1975,N_778,N_166);
nor U1976 (N_1976,In_1385,N_380);
nand U1977 (N_1977,N_307,N_349);
nand U1978 (N_1978,In_2438,In_497);
or U1979 (N_1979,N_111,N_437);
nand U1980 (N_1980,N_420,In_1045);
and U1981 (N_1981,In_1554,N_623);
and U1982 (N_1982,In_1868,N_342);
or U1983 (N_1983,N_150,N_89);
and U1984 (N_1984,In_1259,N_705);
nor U1985 (N_1985,In_903,N_804);
nand U1986 (N_1986,In_2,N_610);
or U1987 (N_1987,N_962,In_923);
nor U1988 (N_1988,N_731,N_186);
nand U1989 (N_1989,N_376,N_597);
or U1990 (N_1990,N_195,N_448);
xor U1991 (N_1991,In_1139,N_728);
or U1992 (N_1992,N_411,In_2046);
nand U1993 (N_1993,N_151,N_466);
nor U1994 (N_1994,N_794,In_2470);
or U1995 (N_1995,N_547,N_466);
and U1996 (N_1996,In_2280,N_199);
or U1997 (N_1997,N_132,N_502);
xor U1998 (N_1998,N_158,N_182);
nand U1999 (N_1999,N_410,In_263);
and U2000 (N_2000,N_1344,N_1976);
xnor U2001 (N_2001,N_1933,N_1803);
nor U2002 (N_2002,N_1158,N_1365);
nor U2003 (N_2003,N_1709,N_1272);
xnor U2004 (N_2004,N_1675,N_1046);
nor U2005 (N_2005,N_1481,N_1655);
and U2006 (N_2006,N_1982,N_1128);
nor U2007 (N_2007,N_1175,N_1753);
xnor U2008 (N_2008,N_1911,N_1601);
and U2009 (N_2009,N_1864,N_1278);
xor U2010 (N_2010,N_1219,N_1463);
nand U2011 (N_2011,N_1826,N_1056);
or U2012 (N_2012,N_1673,N_1234);
nor U2013 (N_2013,N_1120,N_1904);
or U2014 (N_2014,N_1534,N_1816);
or U2015 (N_2015,N_1690,N_1104);
nor U2016 (N_2016,N_1852,N_1785);
xnor U2017 (N_2017,N_1758,N_1266);
and U2018 (N_2018,N_1943,N_1768);
nor U2019 (N_2019,N_1399,N_1134);
xor U2020 (N_2020,N_1957,N_1360);
nor U2021 (N_2021,N_1300,N_1411);
or U2022 (N_2022,N_1877,N_1420);
and U2023 (N_2023,N_1218,N_1874);
and U2024 (N_2024,N_1553,N_1710);
xnor U2025 (N_2025,N_1781,N_1107);
or U2026 (N_2026,N_1393,N_1143);
or U2027 (N_2027,N_1699,N_1116);
and U2028 (N_2028,N_1950,N_1873);
nand U2029 (N_2029,N_1189,N_1509);
and U2030 (N_2030,N_1923,N_1934);
xnor U2031 (N_2031,N_1276,N_1735);
xnor U2032 (N_2032,N_1700,N_1988);
and U2033 (N_2033,N_1053,N_1797);
and U2034 (N_2034,N_1233,N_1228);
xor U2035 (N_2035,N_1345,N_1452);
nor U2036 (N_2036,N_1722,N_1818);
nand U2037 (N_2037,N_1893,N_1497);
and U2038 (N_2038,N_1405,N_1312);
nor U2039 (N_2039,N_1440,N_1383);
nor U2040 (N_2040,N_1227,N_1930);
nand U2041 (N_2041,N_1350,N_1043);
nor U2042 (N_2042,N_1468,N_1856);
or U2043 (N_2043,N_1472,N_1010);
xnor U2044 (N_2044,N_1513,N_1188);
xor U2045 (N_2045,N_1186,N_1791);
nand U2046 (N_2046,N_1669,N_1596);
and U2047 (N_2047,N_1314,N_1038);
nor U2048 (N_2048,N_1343,N_1152);
or U2049 (N_2049,N_1646,N_1796);
or U2050 (N_2050,N_1564,N_1859);
and U2051 (N_2051,N_1938,N_1301);
and U2052 (N_2052,N_1922,N_1760);
and U2053 (N_2053,N_1090,N_1476);
nor U2054 (N_2054,N_1991,N_1321);
xor U2055 (N_2055,N_1693,N_1524);
nand U2056 (N_2056,N_1333,N_1555);
or U2057 (N_2057,N_1949,N_1133);
or U2058 (N_2058,N_1918,N_1478);
xor U2059 (N_2059,N_1637,N_1348);
nor U2060 (N_2060,N_1369,N_1725);
xor U2061 (N_2061,N_1439,N_1238);
nor U2062 (N_2062,N_1151,N_1761);
and U2063 (N_2063,N_1624,N_1719);
and U2064 (N_2064,N_1433,N_1888);
xnor U2065 (N_2065,N_1392,N_1597);
or U2066 (N_2066,N_1259,N_1800);
xnor U2067 (N_2067,N_1653,N_1883);
xor U2068 (N_2068,N_1267,N_1773);
xnor U2069 (N_2069,N_1696,N_1947);
and U2070 (N_2070,N_1268,N_1251);
xor U2071 (N_2071,N_1480,N_1215);
xnor U2072 (N_2072,N_1122,N_1082);
xor U2073 (N_2073,N_1917,N_1538);
or U2074 (N_2074,N_1762,N_1435);
nand U2075 (N_2075,N_1726,N_1823);
and U2076 (N_2076,N_1959,N_1054);
and U2077 (N_2077,N_1378,N_1491);
nor U2078 (N_2078,N_1058,N_1316);
nand U2079 (N_2079,N_1616,N_1496);
nand U2080 (N_2080,N_1289,N_1792);
nand U2081 (N_2081,N_1999,N_1181);
nand U2082 (N_2082,N_1160,N_1860);
nand U2083 (N_2083,N_1184,N_1346);
nor U2084 (N_2084,N_1121,N_1683);
and U2085 (N_2085,N_1707,N_1660);
and U2086 (N_2086,N_1114,N_1415);
or U2087 (N_2087,N_1488,N_1728);
nor U2088 (N_2088,N_1163,N_1517);
nor U2089 (N_2089,N_1937,N_1029);
or U2090 (N_2090,N_1825,N_1000);
or U2091 (N_2091,N_1750,N_1304);
or U2092 (N_2092,N_1108,N_1256);
and U2093 (N_2093,N_1337,N_1724);
xor U2094 (N_2094,N_1897,N_1093);
nand U2095 (N_2095,N_1577,N_1387);
and U2096 (N_2096,N_1824,N_1408);
nand U2097 (N_2097,N_1492,N_1389);
or U2098 (N_2098,N_1960,N_1995);
or U2099 (N_2099,N_1213,N_1868);
nor U2100 (N_2100,N_1989,N_1948);
nor U2101 (N_2101,N_1936,N_1461);
and U2102 (N_2102,N_1376,N_1772);
nand U2103 (N_2103,N_1697,N_1926);
or U2104 (N_2104,N_1559,N_1963);
xnor U2105 (N_2105,N_1743,N_1159);
and U2106 (N_2106,N_1572,N_1084);
nor U2107 (N_2107,N_1249,N_1755);
nand U2108 (N_2108,N_1741,N_1585);
and U2109 (N_2109,N_1255,N_1566);
nand U2110 (N_2110,N_1983,N_1622);
or U2111 (N_2111,N_1067,N_1263);
xnor U2112 (N_2112,N_1799,N_1171);
xnor U2113 (N_2113,N_1968,N_1017);
xnor U2114 (N_2114,N_1242,N_1554);
and U2115 (N_2115,N_1118,N_1031);
and U2116 (N_2116,N_1113,N_1739);
or U2117 (N_2117,N_1636,N_1793);
nand U2118 (N_2118,N_1662,N_1878);
nor U2119 (N_2119,N_1955,N_1150);
xor U2120 (N_2120,N_1875,N_1605);
nand U2121 (N_2121,N_1657,N_1430);
nand U2122 (N_2122,N_1055,N_1167);
nor U2123 (N_2123,N_1329,N_1672);
and U2124 (N_2124,N_1510,N_1317);
and U2125 (N_2125,N_1642,N_1581);
xor U2126 (N_2126,N_1135,N_1779);
or U2127 (N_2127,N_1362,N_1250);
xnor U2128 (N_2128,N_1196,N_1587);
nor U2129 (N_2129,N_1295,N_1907);
and U2130 (N_2130,N_1144,N_1444);
xor U2131 (N_2131,N_1115,N_1138);
and U2132 (N_2132,N_1977,N_1016);
nand U2133 (N_2133,N_1867,N_1880);
xor U2134 (N_2134,N_1347,N_1840);
nor U2135 (N_2135,N_1366,N_1375);
xnor U2136 (N_2136,N_1040,N_1521);
xnor U2137 (N_2137,N_1290,N_1361);
or U2138 (N_2138,N_1630,N_1569);
or U2139 (N_2139,N_1339,N_1821);
xor U2140 (N_2140,N_1005,N_1847);
or U2141 (N_2141,N_1179,N_1531);
and U2142 (N_2142,N_1407,N_1810);
and U2143 (N_2143,N_1428,N_1689);
and U2144 (N_2144,N_1956,N_1287);
nand U2145 (N_2145,N_1734,N_1105);
and U2146 (N_2146,N_1191,N_1216);
or U2147 (N_2147,N_1157,N_1942);
nor U2148 (N_2148,N_1532,N_1526);
nor U2149 (N_2149,N_1073,N_1895);
nand U2150 (N_2150,N_1645,N_1190);
nand U2151 (N_2151,N_1913,N_1483);
nor U2152 (N_2152,N_1342,N_1425);
or U2153 (N_2153,N_1528,N_1035);
or U2154 (N_2154,N_1098,N_1686);
nor U2155 (N_2155,N_1140,N_1633);
nor U2156 (N_2156,N_1599,N_1490);
nand U2157 (N_2157,N_1740,N_1386);
or U2158 (N_2158,N_1174,N_1853);
xor U2159 (N_2159,N_1495,N_1070);
nor U2160 (N_2160,N_1458,N_1899);
nand U2161 (N_2161,N_1870,N_1547);
and U2162 (N_2162,N_1441,N_1264);
nand U2163 (N_2163,N_1765,N_1210);
and U2164 (N_2164,N_1711,N_1909);
and U2165 (N_2165,N_1220,N_1044);
nor U2166 (N_2166,N_1431,N_1041);
or U2167 (N_2167,N_1563,N_1212);
xnor U2168 (N_2168,N_1556,N_1320);
nor U2169 (N_2169,N_1764,N_1049);
or U2170 (N_2170,N_1872,N_1901);
or U2171 (N_2171,N_1136,N_1069);
and U2172 (N_2172,N_1714,N_1292);
or U2173 (N_2173,N_1511,N_1066);
xnor U2174 (N_2174,N_1252,N_1607);
and U2175 (N_2175,N_1448,N_1668);
nor U2176 (N_2176,N_1694,N_1996);
nor U2177 (N_2177,N_1374,N_1927);
and U2178 (N_2178,N_1815,N_1450);
and U2179 (N_2179,N_1204,N_1548);
nor U2180 (N_2180,N_1195,N_1230);
nor U2181 (N_2181,N_1274,N_1822);
and U2182 (N_2182,N_1305,N_1615);
nand U2183 (N_2183,N_1703,N_1079);
or U2184 (N_2184,N_1580,N_1288);
or U2185 (N_2185,N_1368,N_1600);
xor U2186 (N_2186,N_1101,N_1447);
or U2187 (N_2187,N_1028,N_1139);
nand U2188 (N_2188,N_1454,N_1124);
nor U2189 (N_2189,N_1327,N_1299);
and U2190 (N_2190,N_1754,N_1130);
nand U2191 (N_2191,N_1200,N_1285);
or U2192 (N_2192,N_1678,N_1718);
nor U2193 (N_2193,N_1940,N_1363);
nand U2194 (N_2194,N_1892,N_1829);
nor U2195 (N_2195,N_1807,N_1153);
nor U2196 (N_2196,N_1925,N_1545);
or U2197 (N_2197,N_1030,N_1505);
nand U2198 (N_2198,N_1311,N_1391);
xnor U2199 (N_2199,N_1254,N_1384);
nand U2200 (N_2200,N_1298,N_1935);
and U2201 (N_2201,N_1328,N_1410);
or U2202 (N_2202,N_1974,N_1100);
nand U2203 (N_2203,N_1334,N_1446);
nor U2204 (N_2204,N_1089,N_1217);
and U2205 (N_2205,N_1618,N_1612);
or U2206 (N_2206,N_1059,N_1841);
or U2207 (N_2207,N_1512,N_1453);
xnor U2208 (N_2208,N_1162,N_1245);
or U2209 (N_2209,N_1687,N_1462);
and U2210 (N_2210,N_1680,N_1154);
and U2211 (N_2211,N_1381,N_1952);
and U2212 (N_2212,N_1973,N_1533);
nor U2213 (N_2213,N_1353,N_1912);
nor U2214 (N_2214,N_1225,N_1790);
nand U2215 (N_2215,N_1523,N_1352);
nor U2216 (N_2216,N_1331,N_1951);
xor U2217 (N_2217,N_1052,N_1632);
nor U2218 (N_2218,N_1103,N_1479);
xnor U2219 (N_2219,N_1315,N_1099);
nand U2220 (N_2220,N_1232,N_1241);
nor U2221 (N_2221,N_1341,N_1769);
and U2222 (N_2222,N_1731,N_1270);
xnor U2223 (N_2223,N_1804,N_1291);
nor U2224 (N_2224,N_1064,N_1306);
and U2225 (N_2225,N_1434,N_1318);
and U2226 (N_2226,N_1297,N_1654);
and U2227 (N_2227,N_1813,N_1906);
and U2228 (N_2228,N_1887,N_1080);
or U2229 (N_2229,N_1022,N_1606);
or U2230 (N_2230,N_1766,N_1953);
and U2231 (N_2231,N_1522,N_1131);
nor U2232 (N_2232,N_1309,N_1424);
and U2233 (N_2233,N_1261,N_1979);
or U2234 (N_2234,N_1487,N_1065);
and U2235 (N_2235,N_1470,N_1400);
or U2236 (N_2236,N_1507,N_1494);
nand U2237 (N_2237,N_1648,N_1187);
xor U2238 (N_2238,N_1863,N_1244);
or U2239 (N_2239,N_1096,N_1583);
xor U2240 (N_2240,N_1998,N_1565);
nor U2241 (N_2241,N_1889,N_1409);
nor U2242 (N_2242,N_1527,N_1109);
nor U2243 (N_2243,N_1861,N_1401);
or U2244 (N_2244,N_1087,N_1871);
nor U2245 (N_2245,N_1129,N_1349);
xor U2246 (N_2246,N_1777,N_1610);
xnor U2247 (N_2247,N_1598,N_1520);
nand U2248 (N_2248,N_1466,N_1223);
nand U2249 (N_2249,N_1253,N_1862);
and U2250 (N_2250,N_1783,N_1851);
nor U2251 (N_2251,N_1396,N_1809);
and U2252 (N_2252,N_1042,N_1050);
nor U2253 (N_2253,N_1727,N_1137);
and U2254 (N_2254,N_1613,N_1592);
and U2255 (N_2255,N_1033,N_1614);
nand U2256 (N_2256,N_1519,N_1504);
xor U2257 (N_2257,N_1308,N_1021);
nand U2258 (N_2258,N_1192,N_1394);
or U2259 (N_2259,N_1165,N_1723);
nor U2260 (N_2260,N_1916,N_1094);
or U2261 (N_2261,N_1670,N_1900);
nand U2262 (N_2262,N_1373,N_1202);
and U2263 (N_2263,N_1595,N_1798);
and U2264 (N_2264,N_1007,N_1385);
nand U2265 (N_2265,N_1286,N_1110);
or U2266 (N_2266,N_1656,N_1356);
nor U2267 (N_2267,N_1620,N_1965);
nand U2268 (N_2268,N_1639,N_1296);
or U2269 (N_2269,N_1627,N_1182);
xor U2270 (N_2270,N_1688,N_1229);
and U2271 (N_2271,N_1944,N_1484);
or U2272 (N_2272,N_1412,N_1908);
and U2273 (N_2273,N_1849,N_1358);
xnor U2274 (N_2274,N_1681,N_1763);
nand U2275 (N_2275,N_1106,N_1733);
xnor U2276 (N_2276,N_1771,N_1014);
or U2277 (N_2277,N_1294,N_1745);
xor U2278 (N_2278,N_1403,N_1307);
nand U2279 (N_2279,N_1265,N_1048);
nor U2280 (N_2280,N_1455,N_1177);
nand U2281 (N_2281,N_1336,N_1817);
or U2282 (N_2282,N_1176,N_1303);
or U2283 (N_2283,N_1641,N_1018);
xnor U2284 (N_2284,N_1275,N_1705);
nand U2285 (N_2285,N_1954,N_1009);
and U2286 (N_2286,N_1667,N_1183);
nor U2287 (N_2287,N_1691,N_1273);
and U2288 (N_2288,N_1661,N_1432);
xor U2289 (N_2289,N_1004,N_1617);
xnor U2290 (N_2290,N_1757,N_1149);
xor U2291 (N_2291,N_1027,N_1836);
nand U2292 (N_2292,N_1078,N_1850);
or U2293 (N_2293,N_1003,N_1964);
xor U2294 (N_2294,N_1924,N_1269);
and U2295 (N_2295,N_1537,N_1649);
xnor U2296 (N_2296,N_1015,N_1372);
and U2297 (N_2297,N_1482,N_1417);
and U2298 (N_2298,N_1514,N_1102);
and U2299 (N_2299,N_1095,N_1438);
nor U2300 (N_2300,N_1706,N_1283);
nand U2301 (N_2301,N_1736,N_1445);
nor U2302 (N_2302,N_1034,N_1051);
or U2303 (N_2303,N_1833,N_1119);
nor U2304 (N_2304,N_1846,N_1367);
or U2305 (N_2305,N_1682,N_1720);
nand U2306 (N_2306,N_1222,N_1746);
or U2307 (N_2307,N_1819,N_1919);
nor U2308 (N_2308,N_1626,N_1257);
xor U2309 (N_2309,N_1715,N_1037);
or U2310 (N_2310,N_1708,N_1418);
and U2311 (N_2311,N_1945,N_1914);
xnor U2312 (N_2312,N_1416,N_1820);
nor U2313 (N_2313,N_1932,N_1623);
nand U2314 (N_2314,N_1530,N_1025);
or U2315 (N_2315,N_1280,N_1575);
xor U2316 (N_2316,N_1588,N_1354);
or U2317 (N_2317,N_1567,N_1324);
and U2318 (N_2318,N_1885,N_1525);
and U2319 (N_2319,N_1355,N_1971);
xnor U2320 (N_2320,N_1539,N_1449);
or U2321 (N_2321,N_1414,N_1474);
nand U2322 (N_2322,N_1808,N_1744);
nand U2323 (N_2323,N_1586,N_1460);
nor U2324 (N_2324,N_1013,N_1464);
xor U2325 (N_2325,N_1075,N_1751);
nor U2326 (N_2326,N_1485,N_1894);
and U2327 (N_2327,N_1097,N_1795);
nor U2328 (N_2328,N_1112,N_1201);
xor U2329 (N_2329,N_1536,N_1881);
nor U2330 (N_2330,N_1542,N_1898);
or U2331 (N_2331,N_1207,N_1629);
nand U2332 (N_2332,N_1498,N_1582);
xor U2333 (N_2333,N_1541,N_1994);
and U2334 (N_2334,N_1173,N_1166);
xnor U2335 (N_2335,N_1060,N_1077);
nand U2336 (N_2336,N_1716,N_1986);
xor U2337 (N_2337,N_1842,N_1125);
nand U2338 (N_2338,N_1997,N_1535);
or U2339 (N_2339,N_1570,N_1621);
or U2340 (N_2340,N_1584,N_1061);
nor U2341 (N_2341,N_1117,N_1397);
xnor U2342 (N_2342,N_1008,N_1214);
nand U2343 (N_2343,N_1211,N_1987);
nand U2344 (N_2344,N_1193,N_1869);
or U2345 (N_2345,N_1395,N_1026);
nand U2346 (N_2346,N_1246,N_1156);
and U2347 (N_2347,N_1371,N_1132);
or U2348 (N_2348,N_1262,N_1359);
nand U2349 (N_2349,N_1370,N_1837);
nand U2350 (N_2350,N_1981,N_1884);
and U2351 (N_2351,N_1770,N_1155);
and U2352 (N_2352,N_1831,N_1794);
nor U2353 (N_2353,N_1429,N_1603);
xnor U2354 (N_2354,N_1910,N_1506);
nand U2355 (N_2355,N_1557,N_1260);
and U2356 (N_2356,N_1036,N_1413);
xor U2357 (N_2357,N_1208,N_1500);
nand U2358 (N_2358,N_1085,N_1774);
xnor U2359 (N_2359,N_1756,N_1659);
xor U2360 (N_2360,N_1961,N_1164);
and U2361 (N_2361,N_1062,N_1168);
xnor U2362 (N_2362,N_1471,N_1145);
or U2363 (N_2363,N_1978,N_1576);
or U2364 (N_2364,N_1185,N_1402);
xnor U2365 (N_2365,N_1692,N_1302);
or U2366 (N_2366,N_1141,N_1865);
nor U2367 (N_2367,N_1457,N_1456);
xor U2368 (N_2368,N_1380,N_1848);
nand U2369 (N_2369,N_1814,N_1839);
and U2370 (N_2370,N_1664,N_1499);
or U2371 (N_2371,N_1561,N_1489);
or U2372 (N_2372,N_1558,N_1146);
nor U2373 (N_2373,N_1560,N_1442);
nand U2374 (N_2374,N_1236,N_1473);
or U2375 (N_2375,N_1890,N_1002);
and U2376 (N_2376,N_1866,N_1406);
xor U2377 (N_2377,N_1123,N_1198);
nand U2378 (N_2378,N_1674,N_1170);
nand U2379 (N_2379,N_1398,N_1631);
and U2380 (N_2380,N_1571,N_1023);
or U2381 (N_2381,N_1088,N_1749);
nand U2382 (N_2382,N_1351,N_1006);
nor U2383 (N_2383,N_1544,N_1180);
or U2384 (N_2384,N_1501,N_1243);
or U2385 (N_2385,N_1247,N_1966);
or U2386 (N_2386,N_1992,N_1237);
nor U2387 (N_2387,N_1701,N_1529);
nand U2388 (N_2388,N_1698,N_1915);
nor U2389 (N_2389,N_1838,N_1313);
and U2390 (N_2390,N_1012,N_1747);
or U2391 (N_2391,N_1443,N_1609);
or U2392 (N_2392,N_1142,N_1666);
and U2393 (N_2393,N_1776,N_1891);
and U2394 (N_2394,N_1835,N_1011);
xor U2395 (N_2395,N_1737,N_1578);
or U2396 (N_2396,N_1967,N_1619);
or U2397 (N_2397,N_1502,N_1730);
and U2398 (N_2398,N_1282,N_1665);
or U2399 (N_2399,N_1969,N_1857);
or U2400 (N_2400,N_1604,N_1322);
or U2401 (N_2401,N_1602,N_1975);
or U2402 (N_2402,N_1568,N_1427);
xnor U2403 (N_2403,N_1319,N_1172);
xnor U2404 (N_2404,N_1608,N_1364);
and U2405 (N_2405,N_1876,N_1828);
and U2406 (N_2406,N_1235,N_1628);
and U2407 (N_2407,N_1811,N_1076);
nand U2408 (N_2408,N_1325,N_1721);
nor U2409 (N_2409,N_1467,N_1063);
and U2410 (N_2410,N_1946,N_1197);
or U2411 (N_2411,N_1640,N_1086);
xor U2412 (N_2412,N_1083,N_1832);
nor U2413 (N_2413,N_1178,N_1493);
nand U2414 (N_2414,N_1729,N_1650);
or U2415 (N_2415,N_1240,N_1310);
nand U2416 (N_2416,N_1357,N_1437);
xnor U2417 (N_2417,N_1573,N_1962);
nand U2418 (N_2418,N_1465,N_1928);
or U2419 (N_2419,N_1752,N_1068);
nor U2420 (N_2420,N_1226,N_1611);
xnor U2421 (N_2421,N_1929,N_1147);
or U2422 (N_2422,N_1993,N_1594);
xor U2423 (N_2423,N_1931,N_1845);
nor U2424 (N_2424,N_1518,N_1206);
nor U2425 (N_2425,N_1421,N_1074);
xnor U2426 (N_2426,N_1503,N_1338);
or U2427 (N_2427,N_1326,N_1419);
or U2428 (N_2428,N_1695,N_1786);
or U2429 (N_2429,N_1677,N_1844);
nand U2430 (N_2430,N_1905,N_1231);
and U2431 (N_2431,N_1676,N_1486);
xor U2432 (N_2432,N_1921,N_1647);
xor U2433 (N_2433,N_1111,N_1072);
nor U2434 (N_2434,N_1279,N_1284);
xnor U2435 (N_2435,N_1551,N_1759);
nand U2436 (N_2436,N_1780,N_1092);
xor U2437 (N_2437,N_1335,N_1091);
nand U2438 (N_2438,N_1293,N_1985);
nand U2439 (N_2439,N_1001,N_1019);
xor U2440 (N_2440,N_1330,N_1423);
nand U2441 (N_2441,N_1047,N_1020);
xnor U2442 (N_2442,N_1574,N_1939);
or U2443 (N_2443,N_1590,N_1543);
and U2444 (N_2444,N_1277,N_1045);
and U2445 (N_2445,N_1475,N_1702);
or U2446 (N_2446,N_1552,N_1802);
xnor U2447 (N_2447,N_1469,N_1209);
nor U2448 (N_2448,N_1742,N_1643);
xor U2449 (N_2449,N_1778,N_1194);
nor U2450 (N_2450,N_1591,N_1258);
and U2451 (N_2451,N_1685,N_1638);
and U2452 (N_2452,N_1958,N_1713);
xor U2453 (N_2453,N_1032,N_1775);
nor U2454 (N_2454,N_1748,N_1404);
nor U2455 (N_2455,N_1515,N_1903);
nand U2456 (N_2456,N_1858,N_1704);
and U2457 (N_2457,N_1516,N_1508);
or U2458 (N_2458,N_1579,N_1382);
and U2459 (N_2459,N_1057,N_1843);
and U2460 (N_2460,N_1071,N_1546);
nor U2461 (N_2461,N_1451,N_1199);
nor U2462 (N_2462,N_1169,N_1562);
nor U2463 (N_2463,N_1663,N_1589);
nor U2464 (N_2464,N_1281,N_1787);
or U2465 (N_2465,N_1205,N_1855);
xor U2466 (N_2466,N_1767,N_1879);
xnor U2467 (N_2467,N_1221,N_1972);
nand U2468 (N_2468,N_1024,N_1550);
and U2469 (N_2469,N_1340,N_1827);
xnor U2470 (N_2470,N_1224,N_1788);
or U2471 (N_2471,N_1377,N_1635);
nor U2472 (N_2472,N_1805,N_1127);
xnor U2473 (N_2473,N_1426,N_1920);
and U2474 (N_2474,N_1126,N_1161);
xor U2475 (N_2475,N_1801,N_1789);
xnor U2476 (N_2476,N_1738,N_1436);
nand U2477 (N_2477,N_1459,N_1712);
nand U2478 (N_2478,N_1882,N_1390);
nor U2479 (N_2479,N_1902,N_1812);
nor U2480 (N_2480,N_1239,N_1634);
xor U2481 (N_2481,N_1652,N_1684);
nand U2482 (N_2482,N_1732,N_1203);
and U2483 (N_2483,N_1984,N_1886);
and U2484 (N_2484,N_1834,N_1717);
nor U2485 (N_2485,N_1990,N_1248);
nor U2486 (N_2486,N_1970,N_1625);
or U2487 (N_2487,N_1830,N_1854);
xor U2488 (N_2488,N_1671,N_1593);
or U2489 (N_2489,N_1148,N_1081);
or U2490 (N_2490,N_1658,N_1941);
xnor U2491 (N_2491,N_1379,N_1477);
and U2492 (N_2492,N_1896,N_1782);
nand U2493 (N_2493,N_1332,N_1323);
xnor U2494 (N_2494,N_1644,N_1422);
xor U2495 (N_2495,N_1806,N_1549);
and U2496 (N_2496,N_1388,N_1784);
nor U2497 (N_2497,N_1039,N_1540);
and U2498 (N_2498,N_1271,N_1980);
nor U2499 (N_2499,N_1679,N_1651);
xor U2500 (N_2500,N_1467,N_1751);
nand U2501 (N_2501,N_1846,N_1752);
and U2502 (N_2502,N_1243,N_1099);
nor U2503 (N_2503,N_1859,N_1856);
or U2504 (N_2504,N_1271,N_1676);
xor U2505 (N_2505,N_1352,N_1118);
or U2506 (N_2506,N_1134,N_1031);
nand U2507 (N_2507,N_1296,N_1721);
and U2508 (N_2508,N_1163,N_1125);
xor U2509 (N_2509,N_1208,N_1082);
xor U2510 (N_2510,N_1780,N_1612);
nand U2511 (N_2511,N_1536,N_1665);
xnor U2512 (N_2512,N_1432,N_1493);
xnor U2513 (N_2513,N_1081,N_1546);
xnor U2514 (N_2514,N_1929,N_1854);
nand U2515 (N_2515,N_1144,N_1524);
or U2516 (N_2516,N_1583,N_1965);
and U2517 (N_2517,N_1816,N_1993);
nor U2518 (N_2518,N_1480,N_1337);
nor U2519 (N_2519,N_1112,N_1869);
nand U2520 (N_2520,N_1632,N_1660);
and U2521 (N_2521,N_1597,N_1442);
and U2522 (N_2522,N_1588,N_1383);
nor U2523 (N_2523,N_1656,N_1282);
nor U2524 (N_2524,N_1297,N_1285);
nor U2525 (N_2525,N_1692,N_1864);
nand U2526 (N_2526,N_1609,N_1971);
or U2527 (N_2527,N_1397,N_1618);
nand U2528 (N_2528,N_1502,N_1900);
and U2529 (N_2529,N_1728,N_1580);
nand U2530 (N_2530,N_1401,N_1584);
xor U2531 (N_2531,N_1163,N_1106);
or U2532 (N_2532,N_1002,N_1780);
nor U2533 (N_2533,N_1567,N_1223);
nor U2534 (N_2534,N_1518,N_1731);
and U2535 (N_2535,N_1205,N_1861);
or U2536 (N_2536,N_1339,N_1920);
or U2537 (N_2537,N_1837,N_1446);
nand U2538 (N_2538,N_1573,N_1293);
or U2539 (N_2539,N_1210,N_1868);
nor U2540 (N_2540,N_1933,N_1907);
xor U2541 (N_2541,N_1534,N_1654);
nand U2542 (N_2542,N_1718,N_1068);
xnor U2543 (N_2543,N_1623,N_1515);
nor U2544 (N_2544,N_1078,N_1491);
and U2545 (N_2545,N_1840,N_1471);
and U2546 (N_2546,N_1089,N_1056);
xor U2547 (N_2547,N_1066,N_1256);
xnor U2548 (N_2548,N_1285,N_1957);
nor U2549 (N_2549,N_1561,N_1818);
or U2550 (N_2550,N_1860,N_1897);
xor U2551 (N_2551,N_1984,N_1211);
nand U2552 (N_2552,N_1441,N_1652);
or U2553 (N_2553,N_1224,N_1750);
or U2554 (N_2554,N_1905,N_1243);
and U2555 (N_2555,N_1546,N_1102);
nand U2556 (N_2556,N_1575,N_1742);
and U2557 (N_2557,N_1087,N_1138);
and U2558 (N_2558,N_1606,N_1678);
nand U2559 (N_2559,N_1566,N_1477);
xor U2560 (N_2560,N_1075,N_1683);
or U2561 (N_2561,N_1416,N_1791);
and U2562 (N_2562,N_1842,N_1264);
and U2563 (N_2563,N_1197,N_1886);
or U2564 (N_2564,N_1752,N_1147);
nor U2565 (N_2565,N_1546,N_1164);
xnor U2566 (N_2566,N_1363,N_1938);
and U2567 (N_2567,N_1560,N_1028);
nor U2568 (N_2568,N_1860,N_1411);
xor U2569 (N_2569,N_1853,N_1571);
xor U2570 (N_2570,N_1030,N_1862);
nor U2571 (N_2571,N_1641,N_1734);
nand U2572 (N_2572,N_1060,N_1891);
nor U2573 (N_2573,N_1123,N_1839);
nor U2574 (N_2574,N_1791,N_1423);
xnor U2575 (N_2575,N_1687,N_1264);
nand U2576 (N_2576,N_1692,N_1531);
xor U2577 (N_2577,N_1963,N_1192);
nor U2578 (N_2578,N_1721,N_1469);
nand U2579 (N_2579,N_1972,N_1741);
nor U2580 (N_2580,N_1697,N_1207);
xnor U2581 (N_2581,N_1934,N_1183);
nor U2582 (N_2582,N_1570,N_1173);
and U2583 (N_2583,N_1657,N_1984);
nand U2584 (N_2584,N_1328,N_1074);
or U2585 (N_2585,N_1076,N_1019);
nand U2586 (N_2586,N_1455,N_1137);
and U2587 (N_2587,N_1616,N_1268);
or U2588 (N_2588,N_1108,N_1067);
nor U2589 (N_2589,N_1464,N_1155);
nor U2590 (N_2590,N_1492,N_1467);
or U2591 (N_2591,N_1859,N_1369);
nand U2592 (N_2592,N_1420,N_1323);
and U2593 (N_2593,N_1138,N_1797);
and U2594 (N_2594,N_1209,N_1142);
and U2595 (N_2595,N_1361,N_1233);
nor U2596 (N_2596,N_1933,N_1683);
nor U2597 (N_2597,N_1995,N_1324);
and U2598 (N_2598,N_1027,N_1026);
or U2599 (N_2599,N_1321,N_1410);
nand U2600 (N_2600,N_1817,N_1255);
nand U2601 (N_2601,N_1255,N_1132);
and U2602 (N_2602,N_1781,N_1134);
and U2603 (N_2603,N_1234,N_1064);
or U2604 (N_2604,N_1365,N_1915);
xor U2605 (N_2605,N_1822,N_1574);
nor U2606 (N_2606,N_1540,N_1542);
nand U2607 (N_2607,N_1049,N_1246);
nor U2608 (N_2608,N_1528,N_1884);
nand U2609 (N_2609,N_1474,N_1406);
nor U2610 (N_2610,N_1279,N_1572);
and U2611 (N_2611,N_1921,N_1844);
or U2612 (N_2612,N_1555,N_1550);
nand U2613 (N_2613,N_1364,N_1786);
or U2614 (N_2614,N_1249,N_1373);
or U2615 (N_2615,N_1614,N_1687);
and U2616 (N_2616,N_1015,N_1633);
or U2617 (N_2617,N_1256,N_1934);
and U2618 (N_2618,N_1210,N_1783);
nor U2619 (N_2619,N_1744,N_1975);
or U2620 (N_2620,N_1721,N_1034);
nor U2621 (N_2621,N_1659,N_1216);
or U2622 (N_2622,N_1872,N_1721);
nor U2623 (N_2623,N_1886,N_1741);
or U2624 (N_2624,N_1943,N_1744);
nand U2625 (N_2625,N_1580,N_1388);
and U2626 (N_2626,N_1685,N_1051);
nor U2627 (N_2627,N_1100,N_1802);
xor U2628 (N_2628,N_1592,N_1753);
or U2629 (N_2629,N_1837,N_1220);
xor U2630 (N_2630,N_1973,N_1340);
and U2631 (N_2631,N_1501,N_1803);
xor U2632 (N_2632,N_1284,N_1505);
nand U2633 (N_2633,N_1715,N_1847);
nand U2634 (N_2634,N_1785,N_1576);
or U2635 (N_2635,N_1430,N_1982);
xnor U2636 (N_2636,N_1915,N_1758);
or U2637 (N_2637,N_1465,N_1152);
and U2638 (N_2638,N_1964,N_1830);
and U2639 (N_2639,N_1065,N_1312);
xor U2640 (N_2640,N_1281,N_1558);
nand U2641 (N_2641,N_1207,N_1337);
xor U2642 (N_2642,N_1205,N_1601);
xnor U2643 (N_2643,N_1157,N_1172);
nand U2644 (N_2644,N_1801,N_1846);
and U2645 (N_2645,N_1863,N_1631);
and U2646 (N_2646,N_1396,N_1191);
nor U2647 (N_2647,N_1106,N_1289);
nor U2648 (N_2648,N_1228,N_1769);
or U2649 (N_2649,N_1660,N_1555);
nand U2650 (N_2650,N_1353,N_1103);
or U2651 (N_2651,N_1288,N_1013);
or U2652 (N_2652,N_1966,N_1867);
and U2653 (N_2653,N_1153,N_1192);
and U2654 (N_2654,N_1026,N_1998);
or U2655 (N_2655,N_1078,N_1275);
nand U2656 (N_2656,N_1870,N_1238);
nand U2657 (N_2657,N_1656,N_1755);
nand U2658 (N_2658,N_1961,N_1877);
nand U2659 (N_2659,N_1690,N_1059);
and U2660 (N_2660,N_1823,N_1119);
nand U2661 (N_2661,N_1194,N_1542);
and U2662 (N_2662,N_1184,N_1013);
nand U2663 (N_2663,N_1543,N_1678);
nor U2664 (N_2664,N_1332,N_1426);
xor U2665 (N_2665,N_1238,N_1268);
xor U2666 (N_2666,N_1322,N_1463);
or U2667 (N_2667,N_1843,N_1867);
nand U2668 (N_2668,N_1692,N_1890);
xor U2669 (N_2669,N_1943,N_1692);
xor U2670 (N_2670,N_1668,N_1785);
nand U2671 (N_2671,N_1221,N_1252);
and U2672 (N_2672,N_1235,N_1922);
or U2673 (N_2673,N_1293,N_1061);
xor U2674 (N_2674,N_1127,N_1232);
and U2675 (N_2675,N_1009,N_1912);
nor U2676 (N_2676,N_1210,N_1615);
xor U2677 (N_2677,N_1981,N_1637);
nor U2678 (N_2678,N_1492,N_1311);
nor U2679 (N_2679,N_1009,N_1901);
or U2680 (N_2680,N_1280,N_1232);
and U2681 (N_2681,N_1286,N_1088);
xor U2682 (N_2682,N_1884,N_1934);
or U2683 (N_2683,N_1119,N_1934);
nand U2684 (N_2684,N_1682,N_1809);
or U2685 (N_2685,N_1670,N_1630);
nand U2686 (N_2686,N_1509,N_1029);
nor U2687 (N_2687,N_1684,N_1479);
xnor U2688 (N_2688,N_1307,N_1366);
and U2689 (N_2689,N_1123,N_1210);
nand U2690 (N_2690,N_1587,N_1984);
or U2691 (N_2691,N_1866,N_1772);
nand U2692 (N_2692,N_1041,N_1999);
nand U2693 (N_2693,N_1338,N_1045);
and U2694 (N_2694,N_1217,N_1383);
xor U2695 (N_2695,N_1356,N_1497);
nor U2696 (N_2696,N_1169,N_1699);
xor U2697 (N_2697,N_1068,N_1018);
and U2698 (N_2698,N_1347,N_1759);
xnor U2699 (N_2699,N_1107,N_1486);
nor U2700 (N_2700,N_1496,N_1609);
xnor U2701 (N_2701,N_1731,N_1074);
xor U2702 (N_2702,N_1892,N_1926);
xnor U2703 (N_2703,N_1897,N_1495);
xnor U2704 (N_2704,N_1065,N_1169);
nor U2705 (N_2705,N_1833,N_1431);
nand U2706 (N_2706,N_1812,N_1958);
xor U2707 (N_2707,N_1314,N_1843);
or U2708 (N_2708,N_1914,N_1703);
and U2709 (N_2709,N_1406,N_1175);
nor U2710 (N_2710,N_1164,N_1875);
nor U2711 (N_2711,N_1955,N_1044);
nor U2712 (N_2712,N_1718,N_1927);
nor U2713 (N_2713,N_1237,N_1986);
or U2714 (N_2714,N_1204,N_1215);
nor U2715 (N_2715,N_1851,N_1747);
or U2716 (N_2716,N_1195,N_1031);
and U2717 (N_2717,N_1311,N_1738);
or U2718 (N_2718,N_1423,N_1675);
and U2719 (N_2719,N_1699,N_1484);
or U2720 (N_2720,N_1135,N_1987);
or U2721 (N_2721,N_1842,N_1249);
xnor U2722 (N_2722,N_1717,N_1132);
xnor U2723 (N_2723,N_1423,N_1070);
or U2724 (N_2724,N_1716,N_1383);
nor U2725 (N_2725,N_1600,N_1808);
nand U2726 (N_2726,N_1636,N_1257);
and U2727 (N_2727,N_1403,N_1106);
nand U2728 (N_2728,N_1923,N_1485);
nor U2729 (N_2729,N_1376,N_1293);
nor U2730 (N_2730,N_1823,N_1106);
xor U2731 (N_2731,N_1826,N_1770);
nand U2732 (N_2732,N_1669,N_1355);
nand U2733 (N_2733,N_1864,N_1785);
or U2734 (N_2734,N_1604,N_1481);
xnor U2735 (N_2735,N_1919,N_1081);
nand U2736 (N_2736,N_1553,N_1432);
nor U2737 (N_2737,N_1122,N_1964);
xor U2738 (N_2738,N_1626,N_1571);
nand U2739 (N_2739,N_1555,N_1198);
nor U2740 (N_2740,N_1100,N_1855);
and U2741 (N_2741,N_1813,N_1073);
nand U2742 (N_2742,N_1728,N_1586);
xor U2743 (N_2743,N_1683,N_1446);
or U2744 (N_2744,N_1666,N_1108);
or U2745 (N_2745,N_1717,N_1424);
nand U2746 (N_2746,N_1816,N_1411);
xnor U2747 (N_2747,N_1755,N_1032);
or U2748 (N_2748,N_1166,N_1466);
nand U2749 (N_2749,N_1241,N_1201);
or U2750 (N_2750,N_1137,N_1900);
or U2751 (N_2751,N_1630,N_1788);
and U2752 (N_2752,N_1943,N_1135);
and U2753 (N_2753,N_1327,N_1339);
nand U2754 (N_2754,N_1524,N_1163);
nor U2755 (N_2755,N_1929,N_1830);
nor U2756 (N_2756,N_1296,N_1356);
and U2757 (N_2757,N_1711,N_1317);
xnor U2758 (N_2758,N_1425,N_1682);
nor U2759 (N_2759,N_1238,N_1349);
and U2760 (N_2760,N_1980,N_1687);
nand U2761 (N_2761,N_1295,N_1298);
and U2762 (N_2762,N_1958,N_1472);
xnor U2763 (N_2763,N_1181,N_1241);
or U2764 (N_2764,N_1988,N_1963);
nand U2765 (N_2765,N_1276,N_1921);
nor U2766 (N_2766,N_1931,N_1974);
xnor U2767 (N_2767,N_1473,N_1491);
nor U2768 (N_2768,N_1542,N_1791);
nand U2769 (N_2769,N_1730,N_1252);
and U2770 (N_2770,N_1735,N_1450);
and U2771 (N_2771,N_1889,N_1290);
xor U2772 (N_2772,N_1443,N_1887);
nor U2773 (N_2773,N_1758,N_1557);
or U2774 (N_2774,N_1004,N_1510);
or U2775 (N_2775,N_1528,N_1473);
xnor U2776 (N_2776,N_1518,N_1336);
and U2777 (N_2777,N_1052,N_1174);
nand U2778 (N_2778,N_1666,N_1020);
nand U2779 (N_2779,N_1638,N_1981);
and U2780 (N_2780,N_1244,N_1782);
nand U2781 (N_2781,N_1443,N_1783);
and U2782 (N_2782,N_1096,N_1519);
nor U2783 (N_2783,N_1532,N_1359);
or U2784 (N_2784,N_1765,N_1315);
and U2785 (N_2785,N_1419,N_1435);
and U2786 (N_2786,N_1904,N_1790);
or U2787 (N_2787,N_1755,N_1818);
nand U2788 (N_2788,N_1917,N_1054);
or U2789 (N_2789,N_1502,N_1249);
and U2790 (N_2790,N_1890,N_1034);
nor U2791 (N_2791,N_1311,N_1560);
nor U2792 (N_2792,N_1099,N_1646);
nor U2793 (N_2793,N_1036,N_1476);
nand U2794 (N_2794,N_1448,N_1813);
xnor U2795 (N_2795,N_1518,N_1611);
xnor U2796 (N_2796,N_1691,N_1544);
xnor U2797 (N_2797,N_1312,N_1225);
xor U2798 (N_2798,N_1249,N_1616);
xor U2799 (N_2799,N_1602,N_1022);
or U2800 (N_2800,N_1774,N_1292);
nand U2801 (N_2801,N_1454,N_1018);
or U2802 (N_2802,N_1464,N_1150);
nand U2803 (N_2803,N_1701,N_1559);
nand U2804 (N_2804,N_1131,N_1518);
nor U2805 (N_2805,N_1786,N_1613);
and U2806 (N_2806,N_1009,N_1871);
nor U2807 (N_2807,N_1801,N_1061);
nand U2808 (N_2808,N_1525,N_1364);
nand U2809 (N_2809,N_1846,N_1580);
nor U2810 (N_2810,N_1824,N_1362);
and U2811 (N_2811,N_1723,N_1031);
xor U2812 (N_2812,N_1535,N_1251);
or U2813 (N_2813,N_1137,N_1431);
xnor U2814 (N_2814,N_1298,N_1367);
nor U2815 (N_2815,N_1301,N_1611);
nor U2816 (N_2816,N_1121,N_1188);
nand U2817 (N_2817,N_1876,N_1423);
xnor U2818 (N_2818,N_1411,N_1397);
xor U2819 (N_2819,N_1898,N_1679);
xor U2820 (N_2820,N_1874,N_1756);
nand U2821 (N_2821,N_1284,N_1830);
nand U2822 (N_2822,N_1214,N_1532);
nor U2823 (N_2823,N_1985,N_1420);
nand U2824 (N_2824,N_1990,N_1140);
nand U2825 (N_2825,N_1445,N_1772);
nand U2826 (N_2826,N_1403,N_1777);
and U2827 (N_2827,N_1598,N_1414);
and U2828 (N_2828,N_1253,N_1107);
and U2829 (N_2829,N_1127,N_1064);
or U2830 (N_2830,N_1697,N_1874);
nor U2831 (N_2831,N_1587,N_1582);
or U2832 (N_2832,N_1477,N_1228);
nor U2833 (N_2833,N_1004,N_1020);
xnor U2834 (N_2834,N_1232,N_1636);
xnor U2835 (N_2835,N_1176,N_1108);
nand U2836 (N_2836,N_1579,N_1585);
nor U2837 (N_2837,N_1782,N_1488);
nor U2838 (N_2838,N_1868,N_1422);
and U2839 (N_2839,N_1555,N_1549);
nor U2840 (N_2840,N_1686,N_1572);
xnor U2841 (N_2841,N_1977,N_1995);
or U2842 (N_2842,N_1829,N_1778);
or U2843 (N_2843,N_1693,N_1487);
nor U2844 (N_2844,N_1550,N_1314);
and U2845 (N_2845,N_1229,N_1875);
and U2846 (N_2846,N_1712,N_1697);
xnor U2847 (N_2847,N_1670,N_1935);
nor U2848 (N_2848,N_1814,N_1524);
nor U2849 (N_2849,N_1620,N_1240);
and U2850 (N_2850,N_1199,N_1996);
or U2851 (N_2851,N_1749,N_1725);
xnor U2852 (N_2852,N_1084,N_1739);
nor U2853 (N_2853,N_1598,N_1232);
nor U2854 (N_2854,N_1899,N_1363);
or U2855 (N_2855,N_1389,N_1552);
and U2856 (N_2856,N_1218,N_1258);
xnor U2857 (N_2857,N_1595,N_1219);
and U2858 (N_2858,N_1839,N_1421);
and U2859 (N_2859,N_1530,N_1952);
xor U2860 (N_2860,N_1129,N_1517);
and U2861 (N_2861,N_1971,N_1186);
nand U2862 (N_2862,N_1530,N_1975);
xor U2863 (N_2863,N_1141,N_1845);
or U2864 (N_2864,N_1604,N_1221);
and U2865 (N_2865,N_1847,N_1652);
xor U2866 (N_2866,N_1753,N_1657);
nand U2867 (N_2867,N_1988,N_1697);
xnor U2868 (N_2868,N_1506,N_1452);
and U2869 (N_2869,N_1621,N_1401);
xnor U2870 (N_2870,N_1957,N_1154);
and U2871 (N_2871,N_1863,N_1781);
or U2872 (N_2872,N_1018,N_1523);
or U2873 (N_2873,N_1264,N_1412);
nor U2874 (N_2874,N_1780,N_1063);
or U2875 (N_2875,N_1480,N_1726);
nand U2876 (N_2876,N_1916,N_1514);
xor U2877 (N_2877,N_1276,N_1085);
xnor U2878 (N_2878,N_1526,N_1071);
nor U2879 (N_2879,N_1674,N_1254);
nand U2880 (N_2880,N_1515,N_1668);
and U2881 (N_2881,N_1040,N_1630);
xor U2882 (N_2882,N_1007,N_1164);
nand U2883 (N_2883,N_1942,N_1465);
and U2884 (N_2884,N_1326,N_1619);
xnor U2885 (N_2885,N_1195,N_1457);
xor U2886 (N_2886,N_1461,N_1915);
xnor U2887 (N_2887,N_1589,N_1983);
nor U2888 (N_2888,N_1410,N_1167);
nand U2889 (N_2889,N_1514,N_1399);
nand U2890 (N_2890,N_1979,N_1963);
nand U2891 (N_2891,N_1428,N_1783);
xnor U2892 (N_2892,N_1440,N_1572);
xnor U2893 (N_2893,N_1473,N_1251);
and U2894 (N_2894,N_1612,N_1697);
nand U2895 (N_2895,N_1907,N_1843);
xnor U2896 (N_2896,N_1287,N_1118);
and U2897 (N_2897,N_1391,N_1565);
and U2898 (N_2898,N_1257,N_1069);
xnor U2899 (N_2899,N_1405,N_1325);
xor U2900 (N_2900,N_1344,N_1718);
and U2901 (N_2901,N_1025,N_1422);
xnor U2902 (N_2902,N_1399,N_1312);
or U2903 (N_2903,N_1856,N_1849);
and U2904 (N_2904,N_1262,N_1350);
or U2905 (N_2905,N_1664,N_1300);
nor U2906 (N_2906,N_1968,N_1978);
nor U2907 (N_2907,N_1762,N_1642);
xor U2908 (N_2908,N_1083,N_1188);
nand U2909 (N_2909,N_1997,N_1368);
or U2910 (N_2910,N_1026,N_1318);
and U2911 (N_2911,N_1397,N_1142);
or U2912 (N_2912,N_1792,N_1425);
xnor U2913 (N_2913,N_1201,N_1861);
xor U2914 (N_2914,N_1118,N_1422);
nand U2915 (N_2915,N_1681,N_1654);
and U2916 (N_2916,N_1178,N_1649);
xor U2917 (N_2917,N_1809,N_1218);
and U2918 (N_2918,N_1991,N_1004);
or U2919 (N_2919,N_1223,N_1749);
xnor U2920 (N_2920,N_1034,N_1089);
or U2921 (N_2921,N_1330,N_1827);
nor U2922 (N_2922,N_1736,N_1129);
xor U2923 (N_2923,N_1191,N_1572);
and U2924 (N_2924,N_1632,N_1497);
and U2925 (N_2925,N_1851,N_1734);
or U2926 (N_2926,N_1206,N_1052);
xnor U2927 (N_2927,N_1885,N_1483);
xor U2928 (N_2928,N_1271,N_1907);
nor U2929 (N_2929,N_1678,N_1760);
xor U2930 (N_2930,N_1722,N_1158);
and U2931 (N_2931,N_1676,N_1633);
nor U2932 (N_2932,N_1270,N_1389);
nor U2933 (N_2933,N_1169,N_1971);
nand U2934 (N_2934,N_1240,N_1723);
xor U2935 (N_2935,N_1546,N_1879);
nand U2936 (N_2936,N_1818,N_1118);
xnor U2937 (N_2937,N_1643,N_1104);
or U2938 (N_2938,N_1756,N_1748);
nor U2939 (N_2939,N_1453,N_1367);
xor U2940 (N_2940,N_1820,N_1381);
xor U2941 (N_2941,N_1865,N_1034);
nand U2942 (N_2942,N_1248,N_1079);
nand U2943 (N_2943,N_1156,N_1185);
and U2944 (N_2944,N_1494,N_1969);
nor U2945 (N_2945,N_1397,N_1954);
or U2946 (N_2946,N_1546,N_1287);
and U2947 (N_2947,N_1429,N_1512);
xnor U2948 (N_2948,N_1788,N_1884);
and U2949 (N_2949,N_1647,N_1175);
nand U2950 (N_2950,N_1263,N_1191);
and U2951 (N_2951,N_1756,N_1961);
nand U2952 (N_2952,N_1065,N_1951);
and U2953 (N_2953,N_1118,N_1650);
xor U2954 (N_2954,N_1903,N_1795);
xnor U2955 (N_2955,N_1815,N_1666);
nor U2956 (N_2956,N_1249,N_1122);
nand U2957 (N_2957,N_1303,N_1927);
xnor U2958 (N_2958,N_1992,N_1031);
xnor U2959 (N_2959,N_1249,N_1846);
nand U2960 (N_2960,N_1233,N_1380);
and U2961 (N_2961,N_1236,N_1826);
or U2962 (N_2962,N_1307,N_1966);
and U2963 (N_2963,N_1871,N_1890);
nor U2964 (N_2964,N_1979,N_1531);
xnor U2965 (N_2965,N_1855,N_1351);
xnor U2966 (N_2966,N_1190,N_1713);
xnor U2967 (N_2967,N_1440,N_1372);
xnor U2968 (N_2968,N_1269,N_1157);
and U2969 (N_2969,N_1770,N_1108);
xor U2970 (N_2970,N_1473,N_1415);
xnor U2971 (N_2971,N_1698,N_1822);
nand U2972 (N_2972,N_1606,N_1220);
and U2973 (N_2973,N_1421,N_1080);
nand U2974 (N_2974,N_1622,N_1781);
xor U2975 (N_2975,N_1678,N_1097);
xor U2976 (N_2976,N_1818,N_1687);
xnor U2977 (N_2977,N_1493,N_1014);
or U2978 (N_2978,N_1345,N_1047);
nand U2979 (N_2979,N_1023,N_1373);
xnor U2980 (N_2980,N_1350,N_1606);
nor U2981 (N_2981,N_1974,N_1653);
nor U2982 (N_2982,N_1876,N_1569);
nand U2983 (N_2983,N_1153,N_1534);
nor U2984 (N_2984,N_1252,N_1362);
nand U2985 (N_2985,N_1002,N_1063);
or U2986 (N_2986,N_1674,N_1669);
or U2987 (N_2987,N_1379,N_1037);
nor U2988 (N_2988,N_1665,N_1505);
nand U2989 (N_2989,N_1016,N_1543);
nor U2990 (N_2990,N_1933,N_1230);
and U2991 (N_2991,N_1950,N_1625);
or U2992 (N_2992,N_1802,N_1090);
or U2993 (N_2993,N_1870,N_1869);
xnor U2994 (N_2994,N_1949,N_1435);
or U2995 (N_2995,N_1791,N_1248);
xor U2996 (N_2996,N_1423,N_1005);
and U2997 (N_2997,N_1324,N_1811);
or U2998 (N_2998,N_1675,N_1997);
or U2999 (N_2999,N_1287,N_1569);
or U3000 (N_3000,N_2533,N_2855);
nand U3001 (N_3001,N_2199,N_2066);
or U3002 (N_3002,N_2041,N_2654);
and U3003 (N_3003,N_2682,N_2017);
or U3004 (N_3004,N_2352,N_2860);
xnor U3005 (N_3005,N_2646,N_2627);
or U3006 (N_3006,N_2923,N_2902);
and U3007 (N_3007,N_2973,N_2703);
nor U3008 (N_3008,N_2406,N_2160);
nand U3009 (N_3009,N_2382,N_2541);
and U3010 (N_3010,N_2222,N_2848);
xnor U3011 (N_3011,N_2413,N_2617);
or U3012 (N_3012,N_2478,N_2274);
xor U3013 (N_3013,N_2729,N_2584);
xor U3014 (N_3014,N_2064,N_2633);
nor U3015 (N_3015,N_2803,N_2326);
nand U3016 (N_3016,N_2576,N_2538);
nor U3017 (N_3017,N_2891,N_2163);
or U3018 (N_3018,N_2909,N_2386);
or U3019 (N_3019,N_2589,N_2399);
nor U3020 (N_3020,N_2798,N_2827);
nand U3021 (N_3021,N_2700,N_2295);
and U3022 (N_3022,N_2691,N_2348);
xnor U3023 (N_3023,N_2812,N_2258);
nand U3024 (N_3024,N_2126,N_2828);
or U3025 (N_3025,N_2928,N_2648);
or U3026 (N_3026,N_2886,N_2514);
and U3027 (N_3027,N_2754,N_2345);
xnor U3028 (N_3028,N_2238,N_2084);
or U3029 (N_3029,N_2692,N_2520);
or U3030 (N_3030,N_2546,N_2138);
xnor U3031 (N_3031,N_2402,N_2869);
or U3032 (N_3032,N_2235,N_2961);
nand U3033 (N_3033,N_2036,N_2650);
nand U3034 (N_3034,N_2548,N_2793);
nand U3035 (N_3035,N_2251,N_2733);
or U3036 (N_3036,N_2338,N_2534);
nor U3037 (N_3037,N_2963,N_2366);
nor U3038 (N_3038,N_2010,N_2512);
or U3039 (N_3039,N_2015,N_2144);
or U3040 (N_3040,N_2592,N_2822);
or U3041 (N_3041,N_2535,N_2740);
and U3042 (N_3042,N_2959,N_2350);
xnor U3043 (N_3043,N_2711,N_2819);
and U3044 (N_3044,N_2442,N_2695);
or U3045 (N_3045,N_2552,N_2025);
or U3046 (N_3046,N_2502,N_2341);
nor U3047 (N_3047,N_2018,N_2906);
or U3048 (N_3048,N_2408,N_2626);
xnor U3049 (N_3049,N_2008,N_2878);
and U3050 (N_3050,N_2192,N_2198);
and U3051 (N_3051,N_2715,N_2519);
and U3052 (N_3052,N_2521,N_2884);
nor U3053 (N_3053,N_2777,N_2311);
or U3054 (N_3054,N_2532,N_2839);
and U3055 (N_3055,N_2287,N_2965);
and U3056 (N_3056,N_2681,N_2383);
and U3057 (N_3057,N_2517,N_2489);
xnor U3058 (N_3058,N_2448,N_2292);
and U3059 (N_3059,N_2834,N_2852);
xor U3060 (N_3060,N_2438,N_2717);
and U3061 (N_3061,N_2629,N_2103);
nor U3062 (N_3062,N_2614,N_2876);
or U3063 (N_3063,N_2559,N_2677);
nor U3064 (N_3064,N_2987,N_2186);
nand U3065 (N_3065,N_2062,N_2114);
or U3066 (N_3066,N_2483,N_2527);
nor U3067 (N_3067,N_2659,N_2686);
nand U3068 (N_3068,N_2397,N_2865);
nand U3069 (N_3069,N_2652,N_2092);
nand U3070 (N_3070,N_2376,N_2197);
or U3071 (N_3071,N_2925,N_2912);
or U3072 (N_3072,N_2917,N_2095);
xnor U3073 (N_3073,N_2286,N_2823);
xnor U3074 (N_3074,N_2737,N_2093);
or U3075 (N_3075,N_2298,N_2042);
xnor U3076 (N_3076,N_2760,N_2970);
or U3077 (N_3077,N_2262,N_2571);
nand U3078 (N_3078,N_2168,N_2680);
nor U3079 (N_3079,N_2272,N_2403);
xnor U3080 (N_3080,N_2927,N_2370);
or U3081 (N_3081,N_2687,N_2841);
and U3082 (N_3082,N_2710,N_2306);
nand U3083 (N_3083,N_2797,N_2121);
nor U3084 (N_3084,N_2440,N_2599);
nand U3085 (N_3085,N_2031,N_2537);
or U3086 (N_3086,N_2707,N_2836);
nor U3087 (N_3087,N_2303,N_2786);
and U3088 (N_3088,N_2026,N_2986);
xnor U3089 (N_3089,N_2282,N_2154);
xor U3090 (N_3090,N_2771,N_2573);
and U3091 (N_3091,N_2435,N_2889);
nand U3092 (N_3092,N_2128,N_2888);
and U3093 (N_3093,N_2398,N_2916);
xnor U3094 (N_3094,N_2380,N_2935);
nand U3095 (N_3095,N_2057,N_2781);
xor U3096 (N_3096,N_2763,N_2953);
nor U3097 (N_3097,N_2053,N_2494);
or U3098 (N_3098,N_2861,N_2709);
nand U3099 (N_3099,N_2835,N_2788);
nand U3100 (N_3100,N_2701,N_2117);
nand U3101 (N_3101,N_2716,N_2216);
or U3102 (N_3102,N_2784,N_2208);
and U3103 (N_3103,N_2943,N_2881);
nor U3104 (N_3104,N_2038,N_2934);
and U3105 (N_3105,N_2672,N_2275);
and U3106 (N_3106,N_2582,N_2979);
nand U3107 (N_3107,N_2228,N_2832);
nand U3108 (N_3108,N_2211,N_2074);
nand U3109 (N_3109,N_2491,N_2735);
xnor U3110 (N_3110,N_2310,N_2866);
xnor U3111 (N_3111,N_2291,N_2256);
and U3112 (N_3112,N_2011,N_2096);
and U3113 (N_3113,N_2615,N_2391);
or U3114 (N_3114,N_2401,N_2429);
or U3115 (N_3115,N_2224,N_2164);
xor U3116 (N_3116,N_2795,N_2642);
or U3117 (N_3117,N_2213,N_2625);
xor U3118 (N_3118,N_2565,N_2296);
nor U3119 (N_3119,N_2536,N_2577);
nor U3120 (N_3120,N_2904,N_2759);
nand U3121 (N_3121,N_2858,N_2524);
xnor U3122 (N_3122,N_2436,N_2462);
xnor U3123 (N_3123,N_2469,N_2315);
and U3124 (N_3124,N_2787,N_2496);
or U3125 (N_3125,N_2032,N_2492);
or U3126 (N_3126,N_2127,N_2465);
nand U3127 (N_3127,N_2293,N_2708);
nand U3128 (N_3128,N_2568,N_2467);
or U3129 (N_3129,N_2557,N_2416);
nor U3130 (N_3130,N_2829,N_2971);
nor U3131 (N_3131,N_2149,N_2774);
xor U3132 (N_3132,N_2765,N_2265);
and U3133 (N_3133,N_2554,N_2161);
nor U3134 (N_3134,N_2574,N_2696);
nor U3135 (N_3135,N_2992,N_2718);
or U3136 (N_3136,N_2294,N_2081);
nor U3137 (N_3137,N_2993,N_2365);
or U3138 (N_3138,N_2236,N_2664);
and U3139 (N_3139,N_2638,N_2207);
nand U3140 (N_3140,N_2241,N_2896);
and U3141 (N_3141,N_2346,N_2407);
nand U3142 (N_3142,N_2751,N_2499);
nor U3143 (N_3143,N_2458,N_2676);
xor U3144 (N_3144,N_2591,N_2752);
or U3145 (N_3145,N_2052,N_2586);
or U3146 (N_3146,N_2731,N_2390);
or U3147 (N_3147,N_2741,N_2206);
nor U3148 (N_3148,N_2468,N_2892);
xnor U3149 (N_3149,N_2480,N_2049);
nor U3150 (N_3150,N_2264,N_2507);
nor U3151 (N_3151,N_2850,N_2840);
xor U3152 (N_3152,N_2649,N_2842);
nand U3153 (N_3153,N_2393,N_2178);
nor U3154 (N_3154,N_2898,N_2780);
and U3155 (N_3155,N_2673,N_2688);
xnor U3156 (N_3156,N_2485,N_2028);
xor U3157 (N_3157,N_2745,N_2431);
nand U3158 (N_3158,N_2001,N_2821);
nand U3159 (N_3159,N_2301,N_2794);
xnor U3160 (N_3160,N_2976,N_2622);
or U3161 (N_3161,N_2378,N_2080);
nor U3162 (N_3162,N_2704,N_2281);
nor U3163 (N_3163,N_2307,N_2964);
or U3164 (N_3164,N_2194,N_2563);
xnor U3165 (N_3165,N_2863,N_2356);
or U3166 (N_3166,N_2675,N_2982);
or U3167 (N_3167,N_2810,N_2868);
nor U3168 (N_3168,N_2609,N_2067);
nor U3169 (N_3169,N_2190,N_2175);
nor U3170 (N_3170,N_2856,N_2805);
or U3171 (N_3171,N_2072,N_2883);
nor U3172 (N_3172,N_2471,N_2604);
or U3173 (N_3173,N_2908,N_2547);
and U3174 (N_3174,N_2678,N_2105);
nand U3175 (N_3175,N_2369,N_2639);
nand U3176 (N_3176,N_2091,N_2619);
and U3177 (N_3177,N_2809,N_2220);
and U3178 (N_3178,N_2410,N_2593);
or U3179 (N_3179,N_2176,N_2414);
nand U3180 (N_3180,N_2088,N_2804);
nor U3181 (N_3181,N_2600,N_2359);
nor U3182 (N_3182,N_2411,N_2937);
xor U3183 (N_3183,N_2285,N_2263);
xor U3184 (N_3184,N_2044,N_2544);
xnor U3185 (N_3185,N_2513,N_2705);
xnor U3186 (N_3186,N_2820,N_2226);
and U3187 (N_3187,N_2612,N_2498);
or U3188 (N_3188,N_2252,N_2324);
nand U3189 (N_3189,N_2488,N_2231);
and U3190 (N_3190,N_2060,N_2762);
and U3191 (N_3191,N_2702,N_2583);
or U3192 (N_3192,N_2666,N_2166);
nor U3193 (N_3193,N_2463,N_2184);
xnor U3194 (N_3194,N_2016,N_2770);
and U3195 (N_3195,N_2721,N_2255);
nor U3196 (N_3196,N_2815,N_2364);
nor U3197 (N_3197,N_2969,N_2392);
and U3198 (N_3198,N_2087,N_2657);
xnor U3199 (N_3199,N_2335,N_2948);
xnor U3200 (N_3200,N_2831,N_2556);
xor U3201 (N_3201,N_2921,N_2746);
or U3202 (N_3202,N_2845,N_2297);
and U3203 (N_3203,N_2753,N_2981);
xnor U3204 (N_3204,N_2801,N_2806);
xnor U3205 (N_3205,N_2189,N_2951);
nor U3206 (N_3206,N_2219,N_2693);
nand U3207 (N_3207,N_2147,N_2640);
or U3208 (N_3208,N_2999,N_2656);
or U3209 (N_3209,N_2069,N_2165);
nand U3210 (N_3210,N_2223,N_2115);
nand U3211 (N_3211,N_2268,N_2864);
and U3212 (N_3212,N_2641,N_2671);
and U3213 (N_3213,N_2086,N_2142);
and U3214 (N_3214,N_2284,N_2932);
nor U3215 (N_3215,N_2769,N_2922);
xor U3216 (N_3216,N_2620,N_2040);
nor U3217 (N_3217,N_2441,N_2029);
nor U3218 (N_3218,N_2975,N_2791);
or U3219 (N_3219,N_2580,N_2632);
nor U3220 (N_3220,N_2336,N_2277);
or U3221 (N_3221,N_2151,N_2813);
xor U3222 (N_3222,N_2148,N_2320);
nor U3223 (N_3223,N_2385,N_2111);
nor U3224 (N_3224,N_2956,N_2954);
xnor U3225 (N_3225,N_2726,N_2977);
and U3226 (N_3226,N_2995,N_2558);
nor U3227 (N_3227,N_2260,N_2046);
or U3228 (N_3228,N_2388,N_2877);
nor U3229 (N_3229,N_2955,N_2249);
xor U3230 (N_3230,N_2332,N_2679);
nand U3231 (N_3231,N_2867,N_2423);
and U3232 (N_3232,N_2313,N_2267);
nand U3233 (N_3233,N_2108,N_2880);
xor U3234 (N_3234,N_2621,N_2996);
xnor U3235 (N_3235,N_2461,N_2553);
or U3236 (N_3236,N_2012,N_2280);
nand U3237 (N_3237,N_2177,N_2317);
nand U3238 (N_3238,N_2734,N_2572);
nand U3239 (N_3239,N_2994,N_2288);
nand U3240 (N_3240,N_2761,N_2985);
nand U3241 (N_3241,N_2050,N_2233);
or U3242 (N_3242,N_2644,N_2802);
nand U3243 (N_3243,N_2257,N_2706);
nor U3244 (N_3244,N_2434,N_2907);
nand U3245 (N_3245,N_2421,N_2611);
nor U3246 (N_3246,N_2974,N_2897);
nand U3247 (N_3247,N_2048,N_2655);
xor U3248 (N_3248,N_2594,N_2690);
nand U3249 (N_3249,N_2875,N_2487);
nand U3250 (N_3250,N_2445,N_2002);
or U3251 (N_3251,N_2045,N_2564);
or U3252 (N_3252,N_2588,N_2651);
nand U3253 (N_3253,N_2244,N_2719);
nand U3254 (N_3254,N_2919,N_2505);
xnor U3255 (N_3255,N_2417,N_2019);
and U3256 (N_3256,N_2495,N_2685);
or U3257 (N_3257,N_2635,N_2330);
nand U3258 (N_3258,N_2684,N_2446);
and U3259 (N_3259,N_2415,N_2145);
and U3260 (N_3260,N_2000,N_2089);
nand U3261 (N_3261,N_2140,N_2305);
or U3262 (N_3262,N_2323,N_2689);
or U3263 (N_3263,N_2456,N_2523);
xnor U3264 (N_3264,N_2851,N_2545);
nor U3265 (N_3265,N_2624,N_2479);
nand U3266 (N_3266,N_2887,N_2529);
xor U3267 (N_3267,N_2669,N_2585);
and U3268 (N_3268,N_2808,N_2377);
nor U3269 (N_3269,N_2811,N_2063);
nand U3270 (N_3270,N_2510,N_2363);
xnor U3271 (N_3271,N_2481,N_2447);
nand U3272 (N_3272,N_2998,N_2183);
xor U3273 (N_3273,N_2182,N_2484);
xnor U3274 (N_3274,N_2234,N_2237);
xor U3275 (N_3275,N_2670,N_2200);
nand U3276 (N_3276,N_2764,N_2490);
nor U3277 (N_3277,N_2539,N_2598);
and U3278 (N_3278,N_2373,N_2874);
nand U3279 (N_3279,N_2153,N_2312);
and U3280 (N_3280,N_2113,N_2567);
xor U3281 (N_3281,N_2561,N_2525);
xor U3282 (N_3282,N_2230,N_2605);
or U3283 (N_3283,N_2240,N_2540);
and U3284 (N_3284,N_2783,N_2090);
or U3285 (N_3285,N_2070,N_2102);
nor U3286 (N_3286,N_2404,N_2778);
nand U3287 (N_3287,N_2195,N_2185);
nand U3288 (N_3288,N_2920,N_2697);
and U3289 (N_3289,N_2844,N_2543);
xor U3290 (N_3290,N_2033,N_2453);
and U3291 (N_3291,N_2083,N_2130);
xnor U3292 (N_3292,N_2354,N_2466);
and U3293 (N_3293,N_2229,N_2039);
and U3294 (N_3294,N_2022,N_2193);
nor U3295 (N_3295,N_2261,N_2030);
nor U3296 (N_3296,N_2966,N_2618);
nand U3297 (N_3297,N_2997,N_2188);
nand U3298 (N_3298,N_2119,N_2124);
and U3299 (N_3299,N_2243,N_2381);
nand U3300 (N_3300,N_2290,N_2123);
or U3301 (N_3301,N_2169,N_2135);
nand U3302 (N_3302,N_2283,N_2125);
xnor U3303 (N_3303,N_2939,N_2530);
xnor U3304 (N_3304,N_2924,N_2551);
nor U3305 (N_3305,N_2662,N_2014);
or U3306 (N_3306,N_2172,N_2750);
xor U3307 (N_3307,N_2698,N_2503);
or U3308 (N_3308,N_2071,N_2562);
or U3309 (N_3309,N_2515,N_2419);
nand U3310 (N_3310,N_2132,N_2962);
and U3311 (N_3311,N_2930,N_2913);
nor U3312 (N_3312,N_2056,N_2796);
nor U3313 (N_3313,N_2122,N_2065);
and U3314 (N_3314,N_2949,N_2203);
or U3315 (N_3315,N_2221,N_2871);
and U3316 (N_3316,N_2107,N_2300);
nand U3317 (N_3317,N_2988,N_2329);
nor U3318 (N_3318,N_2299,N_2361);
nand U3319 (N_3319,N_2343,N_2104);
or U3320 (N_3320,N_2853,N_2816);
xor U3321 (N_3321,N_2003,N_2316);
nand U3322 (N_3322,N_2201,N_2428);
nor U3323 (N_3323,N_2109,N_2587);
xor U3324 (N_3324,N_2174,N_2073);
or U3325 (N_3325,N_2914,N_2653);
xor U3326 (N_3326,N_2351,N_2742);
xnor U3327 (N_3327,N_2023,N_2890);
nand U3328 (N_3328,N_2116,N_2007);
nor U3329 (N_3329,N_2758,N_2136);
and U3330 (N_3330,N_2824,N_2645);
nor U3331 (N_3331,N_2825,N_2162);
nand U3332 (N_3332,N_2773,N_2768);
nor U3333 (N_3333,N_2772,N_2464);
or U3334 (N_3334,N_2325,N_2205);
nor U3335 (N_3335,N_2204,N_2663);
or U3336 (N_3336,N_2344,N_2412);
xor U3337 (N_3337,N_2106,N_2833);
and U3338 (N_3338,N_2739,N_2024);
nand U3339 (N_3339,N_2112,N_2736);
nand U3340 (N_3340,N_2110,N_2933);
nor U3341 (N_3341,N_2980,N_2098);
and U3342 (N_3342,N_2712,N_2630);
or U3343 (N_3343,N_2400,N_2634);
nand U3344 (N_3344,N_2422,N_2725);
xnor U3345 (N_3345,N_2334,N_2661);
or U3346 (N_3346,N_2457,N_2699);
and U3347 (N_3347,N_2396,N_2643);
xor U3348 (N_3348,N_2035,N_2800);
and U3349 (N_3349,N_2566,N_2952);
nor U3350 (N_3350,N_2156,N_2146);
and U3351 (N_3351,N_2239,N_2387);
and U3352 (N_3352,N_2209,N_2133);
and U3353 (N_3353,N_2100,N_2202);
xnor U3354 (N_3354,N_2134,N_2054);
xnor U3355 (N_3355,N_2910,N_2347);
xnor U3356 (N_3356,N_2506,N_2027);
and U3357 (N_3357,N_2141,N_2929);
or U3358 (N_3358,N_2608,N_2248);
xor U3359 (N_3359,N_2560,N_2516);
xor U3360 (N_3360,N_2926,N_2476);
xor U3361 (N_3361,N_2418,N_2227);
or U3362 (N_3362,N_2882,N_2150);
and U3363 (N_3363,N_2501,N_2579);
nand U3364 (N_3364,N_2665,N_2047);
and U3365 (N_3365,N_2322,N_2266);
nand U3366 (N_3366,N_2006,N_2217);
nor U3367 (N_3367,N_2170,N_2606);
and U3368 (N_3368,N_2817,N_2250);
xor U3369 (N_3369,N_2938,N_2601);
and U3370 (N_3370,N_2246,N_2159);
and U3371 (N_3371,N_2319,N_2518);
or U3372 (N_3372,N_2357,N_2785);
or U3373 (N_3373,N_2021,N_2531);
and U3374 (N_3374,N_2854,N_2340);
and U3375 (N_3375,N_2394,N_2327);
or U3376 (N_3376,N_2444,N_2061);
and U3377 (N_3377,N_2637,N_2569);
xor U3378 (N_3378,N_2879,N_2972);
nand U3379 (N_3379,N_2945,N_2610);
nand U3380 (N_3380,N_2331,N_2894);
or U3381 (N_3381,N_2790,N_2129);
xor U3382 (N_3382,N_2355,N_2068);
xnor U3383 (N_3383,N_2757,N_2474);
or U3384 (N_3384,N_2254,N_2253);
xnor U3385 (N_3385,N_2658,N_2232);
nand U3386 (N_3386,N_2372,N_2732);
nand U3387 (N_3387,N_2597,N_2473);
or U3388 (N_3388,N_2748,N_2859);
nor U3389 (N_3389,N_2099,N_2968);
or U3390 (N_3390,N_2775,N_2779);
nand U3391 (N_3391,N_2034,N_2814);
nand U3392 (N_3392,N_2549,N_2171);
xor U3393 (N_3393,N_2509,N_2215);
or U3394 (N_3394,N_2602,N_2289);
and U3395 (N_3395,N_2967,N_2570);
or U3396 (N_3396,N_2747,N_2210);
or U3397 (N_3397,N_2931,N_2433);
nand U3398 (N_3398,N_2944,N_2724);
xor U3399 (N_3399,N_2857,N_2118);
or U3400 (N_3400,N_2885,N_2631);
nor U3401 (N_3401,N_2101,N_2371);
or U3402 (N_3402,N_2846,N_2075);
nand U3403 (N_3403,N_2578,N_2155);
and U3404 (N_3404,N_2694,N_2603);
xor U3405 (N_3405,N_2259,N_2475);
nand U3406 (N_3406,N_2799,N_2838);
nor U3407 (N_3407,N_2674,N_2756);
xor U3408 (N_3408,N_2903,N_2900);
or U3409 (N_3409,N_2899,N_2078);
xor U3410 (N_3410,N_2849,N_2862);
or U3411 (N_3411,N_2668,N_2905);
xor U3412 (N_3412,N_2581,N_2683);
or U3413 (N_3413,N_2451,N_2978);
xor U3414 (N_3414,N_2328,N_2942);
nor U3415 (N_3415,N_2767,N_2616);
nand U3416 (N_3416,N_2792,N_2893);
xor U3417 (N_3417,N_2379,N_2157);
nand U3418 (N_3418,N_2196,N_2308);
or U3419 (N_3419,N_2037,N_2807);
or U3420 (N_3420,N_2278,N_2660);
xnor U3421 (N_3421,N_2983,N_2728);
and U3422 (N_3422,N_2714,N_2242);
nand U3423 (N_3423,N_2059,N_2004);
or U3424 (N_3424,N_2730,N_2333);
and U3425 (N_3425,N_2443,N_2960);
xnor U3426 (N_3426,N_2437,N_2167);
or U3427 (N_3427,N_2424,N_2337);
xor U3428 (N_3428,N_2500,N_2555);
nor U3429 (N_3429,N_2782,N_2309);
or U3430 (N_3430,N_2137,N_2139);
xnor U3431 (N_3431,N_2097,N_2918);
xnor U3432 (N_3432,N_2452,N_2958);
nor U3433 (N_3433,N_2872,N_2508);
xor U3434 (N_3434,N_2304,N_2079);
nand U3435 (N_3435,N_2367,N_2940);
nor U3436 (N_3436,N_2432,N_2427);
and U3437 (N_3437,N_2218,N_2430);
or U3438 (N_3438,N_2384,N_2950);
nand U3439 (N_3439,N_2575,N_2847);
nand U3440 (N_3440,N_2405,N_2826);
or U3441 (N_3441,N_2990,N_2225);
or U3442 (N_3442,N_2339,N_2245);
xor U3443 (N_3443,N_2722,N_2276);
nand U3444 (N_3444,N_2043,N_2915);
xor U3445 (N_3445,N_2957,N_2395);
nor U3446 (N_3446,N_2449,N_2766);
nor U3447 (N_3447,N_2720,N_2450);
nor U3448 (N_3448,N_2528,N_2191);
nor U3449 (N_3449,N_2058,N_2497);
nor U3450 (N_3450,N_2459,N_2470);
or U3451 (N_3451,N_2318,N_2526);
or U3452 (N_3452,N_2991,N_2613);
and U3453 (N_3453,N_2947,N_2738);
nor U3454 (N_3454,N_2180,N_2179);
or U3455 (N_3455,N_2279,N_2187);
and U3456 (N_3456,N_2837,N_2989);
or U3457 (N_3457,N_2454,N_2085);
nand U3458 (N_3458,N_2051,N_2946);
nor U3459 (N_3459,N_2302,N_2321);
nor U3460 (N_3460,N_2830,N_2271);
and U3461 (N_3461,N_2628,N_2420);
xor U3462 (N_3462,N_2055,N_2152);
xor U3463 (N_3463,N_2486,N_2477);
xnor U3464 (N_3464,N_2212,N_2870);
xnor U3465 (N_3465,N_2789,N_2076);
nor U3466 (N_3466,N_2755,N_2723);
xor U3467 (N_3467,N_2901,N_2936);
nor U3468 (N_3468,N_2158,N_2247);
or U3469 (N_3469,N_2273,N_2460);
or U3470 (N_3470,N_2409,N_2504);
nand U3471 (N_3471,N_2360,N_2713);
and U3472 (N_3472,N_2181,N_2362);
and U3473 (N_3473,N_2143,N_2349);
xnor U3474 (N_3474,N_2120,N_2522);
or U3475 (N_3475,N_2727,N_2082);
xor U3476 (N_3476,N_2472,N_2013);
nand U3477 (N_3477,N_2873,N_2607);
xor U3478 (N_3478,N_2550,N_2776);
or U3479 (N_3479,N_2425,N_2482);
and U3480 (N_3480,N_2094,N_2077);
or U3481 (N_3481,N_2173,N_2009);
nor U3482 (N_3482,N_2426,N_2542);
nand U3483 (N_3483,N_2596,N_2667);
xor U3484 (N_3484,N_2984,N_2342);
nand U3485 (N_3485,N_2818,N_2214);
and U3486 (N_3486,N_2493,N_2744);
nor U3487 (N_3487,N_2353,N_2020);
nor U3488 (N_3488,N_2455,N_2439);
nor U3489 (N_3489,N_2595,N_2374);
or U3490 (N_3490,N_2375,N_2269);
nand U3491 (N_3491,N_2314,N_2358);
and U3492 (N_3492,N_2131,N_2005);
xor U3493 (N_3493,N_2743,N_2647);
or U3494 (N_3494,N_2511,N_2941);
and U3495 (N_3495,N_2895,N_2623);
and U3496 (N_3496,N_2636,N_2749);
or U3497 (N_3497,N_2911,N_2389);
xor U3498 (N_3498,N_2270,N_2368);
or U3499 (N_3499,N_2590,N_2843);
nand U3500 (N_3500,N_2784,N_2845);
xnor U3501 (N_3501,N_2692,N_2370);
nor U3502 (N_3502,N_2234,N_2858);
xnor U3503 (N_3503,N_2429,N_2010);
nor U3504 (N_3504,N_2439,N_2780);
nor U3505 (N_3505,N_2549,N_2965);
or U3506 (N_3506,N_2634,N_2229);
xnor U3507 (N_3507,N_2915,N_2757);
nor U3508 (N_3508,N_2442,N_2012);
nor U3509 (N_3509,N_2723,N_2528);
or U3510 (N_3510,N_2964,N_2683);
nor U3511 (N_3511,N_2621,N_2782);
or U3512 (N_3512,N_2451,N_2527);
and U3513 (N_3513,N_2786,N_2374);
nand U3514 (N_3514,N_2513,N_2018);
or U3515 (N_3515,N_2027,N_2501);
xnor U3516 (N_3516,N_2646,N_2083);
and U3517 (N_3517,N_2356,N_2899);
nor U3518 (N_3518,N_2564,N_2384);
or U3519 (N_3519,N_2581,N_2386);
and U3520 (N_3520,N_2991,N_2499);
nor U3521 (N_3521,N_2606,N_2442);
xor U3522 (N_3522,N_2692,N_2656);
nand U3523 (N_3523,N_2780,N_2563);
nor U3524 (N_3524,N_2531,N_2749);
nor U3525 (N_3525,N_2094,N_2832);
and U3526 (N_3526,N_2142,N_2087);
xor U3527 (N_3527,N_2504,N_2408);
nor U3528 (N_3528,N_2500,N_2971);
xnor U3529 (N_3529,N_2168,N_2102);
nand U3530 (N_3530,N_2229,N_2479);
or U3531 (N_3531,N_2186,N_2606);
xor U3532 (N_3532,N_2653,N_2671);
or U3533 (N_3533,N_2238,N_2741);
xnor U3534 (N_3534,N_2136,N_2518);
nor U3535 (N_3535,N_2604,N_2537);
xor U3536 (N_3536,N_2296,N_2275);
nand U3537 (N_3537,N_2225,N_2319);
or U3538 (N_3538,N_2641,N_2768);
nor U3539 (N_3539,N_2807,N_2715);
and U3540 (N_3540,N_2157,N_2947);
nand U3541 (N_3541,N_2155,N_2347);
nor U3542 (N_3542,N_2124,N_2732);
xnor U3543 (N_3543,N_2715,N_2732);
nand U3544 (N_3544,N_2731,N_2381);
nand U3545 (N_3545,N_2510,N_2654);
or U3546 (N_3546,N_2051,N_2818);
and U3547 (N_3547,N_2326,N_2152);
and U3548 (N_3548,N_2250,N_2429);
or U3549 (N_3549,N_2024,N_2084);
xor U3550 (N_3550,N_2322,N_2669);
nand U3551 (N_3551,N_2361,N_2874);
nor U3552 (N_3552,N_2273,N_2257);
and U3553 (N_3553,N_2836,N_2731);
and U3554 (N_3554,N_2111,N_2150);
or U3555 (N_3555,N_2696,N_2338);
and U3556 (N_3556,N_2663,N_2149);
nor U3557 (N_3557,N_2888,N_2777);
and U3558 (N_3558,N_2383,N_2962);
nor U3559 (N_3559,N_2188,N_2032);
nor U3560 (N_3560,N_2000,N_2525);
xnor U3561 (N_3561,N_2534,N_2675);
nand U3562 (N_3562,N_2589,N_2926);
or U3563 (N_3563,N_2918,N_2145);
or U3564 (N_3564,N_2665,N_2671);
nand U3565 (N_3565,N_2782,N_2170);
xor U3566 (N_3566,N_2342,N_2238);
nor U3567 (N_3567,N_2845,N_2880);
nand U3568 (N_3568,N_2928,N_2216);
or U3569 (N_3569,N_2437,N_2965);
and U3570 (N_3570,N_2155,N_2424);
xnor U3571 (N_3571,N_2515,N_2607);
nand U3572 (N_3572,N_2650,N_2516);
xor U3573 (N_3573,N_2353,N_2983);
nand U3574 (N_3574,N_2258,N_2435);
or U3575 (N_3575,N_2034,N_2022);
nand U3576 (N_3576,N_2173,N_2616);
or U3577 (N_3577,N_2049,N_2179);
nor U3578 (N_3578,N_2996,N_2025);
and U3579 (N_3579,N_2509,N_2494);
and U3580 (N_3580,N_2802,N_2027);
nand U3581 (N_3581,N_2065,N_2173);
nand U3582 (N_3582,N_2893,N_2363);
nand U3583 (N_3583,N_2495,N_2236);
xnor U3584 (N_3584,N_2614,N_2111);
xor U3585 (N_3585,N_2724,N_2528);
and U3586 (N_3586,N_2974,N_2357);
and U3587 (N_3587,N_2634,N_2331);
and U3588 (N_3588,N_2600,N_2272);
and U3589 (N_3589,N_2960,N_2071);
nor U3590 (N_3590,N_2361,N_2163);
nor U3591 (N_3591,N_2773,N_2191);
nand U3592 (N_3592,N_2257,N_2410);
or U3593 (N_3593,N_2997,N_2430);
nor U3594 (N_3594,N_2497,N_2826);
and U3595 (N_3595,N_2857,N_2526);
xor U3596 (N_3596,N_2254,N_2136);
nand U3597 (N_3597,N_2817,N_2450);
and U3598 (N_3598,N_2889,N_2377);
or U3599 (N_3599,N_2384,N_2160);
or U3600 (N_3600,N_2495,N_2545);
xor U3601 (N_3601,N_2063,N_2240);
and U3602 (N_3602,N_2673,N_2317);
or U3603 (N_3603,N_2839,N_2563);
nor U3604 (N_3604,N_2009,N_2957);
and U3605 (N_3605,N_2647,N_2887);
nand U3606 (N_3606,N_2462,N_2767);
or U3607 (N_3607,N_2500,N_2286);
nand U3608 (N_3608,N_2789,N_2783);
and U3609 (N_3609,N_2745,N_2901);
and U3610 (N_3610,N_2596,N_2958);
xor U3611 (N_3611,N_2770,N_2046);
nand U3612 (N_3612,N_2803,N_2505);
nor U3613 (N_3613,N_2110,N_2543);
xnor U3614 (N_3614,N_2324,N_2494);
nor U3615 (N_3615,N_2211,N_2646);
nand U3616 (N_3616,N_2262,N_2764);
xnor U3617 (N_3617,N_2930,N_2830);
xnor U3618 (N_3618,N_2740,N_2715);
nor U3619 (N_3619,N_2322,N_2593);
xor U3620 (N_3620,N_2394,N_2727);
nor U3621 (N_3621,N_2624,N_2385);
or U3622 (N_3622,N_2145,N_2512);
nand U3623 (N_3623,N_2642,N_2503);
and U3624 (N_3624,N_2920,N_2746);
xor U3625 (N_3625,N_2267,N_2359);
or U3626 (N_3626,N_2442,N_2736);
or U3627 (N_3627,N_2281,N_2921);
nand U3628 (N_3628,N_2337,N_2437);
and U3629 (N_3629,N_2217,N_2501);
or U3630 (N_3630,N_2450,N_2841);
nor U3631 (N_3631,N_2235,N_2206);
nor U3632 (N_3632,N_2678,N_2485);
nand U3633 (N_3633,N_2930,N_2792);
or U3634 (N_3634,N_2385,N_2121);
nor U3635 (N_3635,N_2444,N_2016);
or U3636 (N_3636,N_2011,N_2998);
xnor U3637 (N_3637,N_2599,N_2918);
nor U3638 (N_3638,N_2577,N_2065);
and U3639 (N_3639,N_2405,N_2720);
nand U3640 (N_3640,N_2102,N_2596);
xor U3641 (N_3641,N_2951,N_2746);
nand U3642 (N_3642,N_2070,N_2527);
or U3643 (N_3643,N_2264,N_2307);
nor U3644 (N_3644,N_2576,N_2202);
nor U3645 (N_3645,N_2149,N_2038);
nand U3646 (N_3646,N_2371,N_2402);
or U3647 (N_3647,N_2908,N_2830);
or U3648 (N_3648,N_2371,N_2123);
or U3649 (N_3649,N_2864,N_2948);
nor U3650 (N_3650,N_2015,N_2342);
xor U3651 (N_3651,N_2057,N_2808);
and U3652 (N_3652,N_2876,N_2465);
xnor U3653 (N_3653,N_2246,N_2069);
or U3654 (N_3654,N_2107,N_2696);
nor U3655 (N_3655,N_2971,N_2912);
or U3656 (N_3656,N_2425,N_2114);
nor U3657 (N_3657,N_2828,N_2169);
and U3658 (N_3658,N_2208,N_2440);
and U3659 (N_3659,N_2133,N_2360);
or U3660 (N_3660,N_2046,N_2273);
or U3661 (N_3661,N_2519,N_2009);
xor U3662 (N_3662,N_2305,N_2243);
or U3663 (N_3663,N_2948,N_2961);
nand U3664 (N_3664,N_2075,N_2886);
xor U3665 (N_3665,N_2226,N_2845);
nand U3666 (N_3666,N_2660,N_2934);
nand U3667 (N_3667,N_2787,N_2802);
or U3668 (N_3668,N_2517,N_2116);
or U3669 (N_3669,N_2980,N_2876);
and U3670 (N_3670,N_2206,N_2241);
or U3671 (N_3671,N_2275,N_2526);
nand U3672 (N_3672,N_2846,N_2597);
nand U3673 (N_3673,N_2219,N_2083);
xor U3674 (N_3674,N_2786,N_2119);
nor U3675 (N_3675,N_2017,N_2188);
nand U3676 (N_3676,N_2746,N_2396);
or U3677 (N_3677,N_2438,N_2121);
and U3678 (N_3678,N_2611,N_2620);
or U3679 (N_3679,N_2503,N_2697);
xor U3680 (N_3680,N_2477,N_2766);
nand U3681 (N_3681,N_2578,N_2546);
nand U3682 (N_3682,N_2367,N_2765);
and U3683 (N_3683,N_2025,N_2148);
nand U3684 (N_3684,N_2901,N_2502);
nor U3685 (N_3685,N_2325,N_2849);
xnor U3686 (N_3686,N_2514,N_2496);
nor U3687 (N_3687,N_2052,N_2924);
or U3688 (N_3688,N_2678,N_2189);
nor U3689 (N_3689,N_2097,N_2987);
and U3690 (N_3690,N_2498,N_2247);
or U3691 (N_3691,N_2592,N_2572);
and U3692 (N_3692,N_2171,N_2800);
and U3693 (N_3693,N_2986,N_2500);
nand U3694 (N_3694,N_2314,N_2865);
nand U3695 (N_3695,N_2377,N_2960);
xnor U3696 (N_3696,N_2874,N_2578);
nor U3697 (N_3697,N_2680,N_2074);
nand U3698 (N_3698,N_2808,N_2011);
and U3699 (N_3699,N_2543,N_2172);
or U3700 (N_3700,N_2762,N_2117);
xnor U3701 (N_3701,N_2711,N_2881);
nand U3702 (N_3702,N_2056,N_2859);
or U3703 (N_3703,N_2586,N_2141);
or U3704 (N_3704,N_2672,N_2500);
and U3705 (N_3705,N_2404,N_2465);
nor U3706 (N_3706,N_2566,N_2932);
or U3707 (N_3707,N_2181,N_2513);
xor U3708 (N_3708,N_2188,N_2673);
nand U3709 (N_3709,N_2216,N_2665);
or U3710 (N_3710,N_2272,N_2371);
and U3711 (N_3711,N_2985,N_2098);
xor U3712 (N_3712,N_2688,N_2603);
and U3713 (N_3713,N_2145,N_2519);
nand U3714 (N_3714,N_2532,N_2043);
nor U3715 (N_3715,N_2129,N_2654);
nor U3716 (N_3716,N_2915,N_2834);
nand U3717 (N_3717,N_2815,N_2570);
or U3718 (N_3718,N_2958,N_2384);
xnor U3719 (N_3719,N_2921,N_2003);
nor U3720 (N_3720,N_2360,N_2549);
nor U3721 (N_3721,N_2521,N_2122);
xor U3722 (N_3722,N_2547,N_2106);
nor U3723 (N_3723,N_2046,N_2367);
nor U3724 (N_3724,N_2013,N_2233);
nand U3725 (N_3725,N_2666,N_2270);
xnor U3726 (N_3726,N_2871,N_2792);
nand U3727 (N_3727,N_2067,N_2605);
nor U3728 (N_3728,N_2442,N_2615);
nor U3729 (N_3729,N_2817,N_2015);
nand U3730 (N_3730,N_2881,N_2453);
or U3731 (N_3731,N_2641,N_2145);
and U3732 (N_3732,N_2909,N_2318);
nand U3733 (N_3733,N_2663,N_2526);
xnor U3734 (N_3734,N_2264,N_2227);
nor U3735 (N_3735,N_2833,N_2204);
and U3736 (N_3736,N_2281,N_2000);
xnor U3737 (N_3737,N_2775,N_2026);
xnor U3738 (N_3738,N_2224,N_2061);
nor U3739 (N_3739,N_2364,N_2676);
and U3740 (N_3740,N_2281,N_2252);
or U3741 (N_3741,N_2024,N_2595);
nor U3742 (N_3742,N_2098,N_2622);
nor U3743 (N_3743,N_2290,N_2373);
nand U3744 (N_3744,N_2676,N_2928);
and U3745 (N_3745,N_2824,N_2533);
xnor U3746 (N_3746,N_2598,N_2904);
nor U3747 (N_3747,N_2870,N_2446);
and U3748 (N_3748,N_2662,N_2913);
and U3749 (N_3749,N_2424,N_2745);
or U3750 (N_3750,N_2348,N_2341);
or U3751 (N_3751,N_2627,N_2817);
nor U3752 (N_3752,N_2472,N_2952);
and U3753 (N_3753,N_2174,N_2488);
or U3754 (N_3754,N_2566,N_2798);
or U3755 (N_3755,N_2413,N_2012);
nor U3756 (N_3756,N_2369,N_2757);
nor U3757 (N_3757,N_2731,N_2780);
nand U3758 (N_3758,N_2159,N_2132);
nand U3759 (N_3759,N_2974,N_2444);
and U3760 (N_3760,N_2894,N_2054);
nand U3761 (N_3761,N_2038,N_2751);
nor U3762 (N_3762,N_2078,N_2723);
nand U3763 (N_3763,N_2516,N_2803);
nand U3764 (N_3764,N_2561,N_2624);
or U3765 (N_3765,N_2002,N_2831);
nor U3766 (N_3766,N_2209,N_2508);
or U3767 (N_3767,N_2945,N_2637);
and U3768 (N_3768,N_2374,N_2511);
xor U3769 (N_3769,N_2690,N_2783);
xnor U3770 (N_3770,N_2587,N_2416);
and U3771 (N_3771,N_2767,N_2208);
xnor U3772 (N_3772,N_2988,N_2422);
xor U3773 (N_3773,N_2714,N_2708);
or U3774 (N_3774,N_2336,N_2434);
xnor U3775 (N_3775,N_2656,N_2986);
and U3776 (N_3776,N_2983,N_2567);
or U3777 (N_3777,N_2747,N_2693);
or U3778 (N_3778,N_2989,N_2293);
nor U3779 (N_3779,N_2843,N_2739);
xnor U3780 (N_3780,N_2001,N_2304);
nand U3781 (N_3781,N_2533,N_2358);
or U3782 (N_3782,N_2228,N_2624);
or U3783 (N_3783,N_2187,N_2363);
or U3784 (N_3784,N_2246,N_2893);
nand U3785 (N_3785,N_2218,N_2844);
nor U3786 (N_3786,N_2254,N_2422);
xnor U3787 (N_3787,N_2858,N_2428);
nor U3788 (N_3788,N_2657,N_2587);
and U3789 (N_3789,N_2197,N_2097);
nor U3790 (N_3790,N_2221,N_2900);
or U3791 (N_3791,N_2488,N_2736);
nand U3792 (N_3792,N_2272,N_2395);
or U3793 (N_3793,N_2754,N_2784);
or U3794 (N_3794,N_2524,N_2737);
xor U3795 (N_3795,N_2521,N_2525);
nand U3796 (N_3796,N_2175,N_2614);
nand U3797 (N_3797,N_2298,N_2224);
or U3798 (N_3798,N_2417,N_2127);
xor U3799 (N_3799,N_2610,N_2302);
nand U3800 (N_3800,N_2212,N_2056);
or U3801 (N_3801,N_2974,N_2873);
and U3802 (N_3802,N_2954,N_2424);
xor U3803 (N_3803,N_2118,N_2416);
nand U3804 (N_3804,N_2732,N_2878);
xor U3805 (N_3805,N_2510,N_2653);
xnor U3806 (N_3806,N_2510,N_2417);
nor U3807 (N_3807,N_2027,N_2469);
nand U3808 (N_3808,N_2054,N_2468);
or U3809 (N_3809,N_2059,N_2575);
nor U3810 (N_3810,N_2516,N_2985);
or U3811 (N_3811,N_2735,N_2612);
or U3812 (N_3812,N_2675,N_2199);
nor U3813 (N_3813,N_2681,N_2649);
or U3814 (N_3814,N_2936,N_2068);
nor U3815 (N_3815,N_2738,N_2366);
or U3816 (N_3816,N_2219,N_2618);
or U3817 (N_3817,N_2602,N_2160);
and U3818 (N_3818,N_2881,N_2221);
or U3819 (N_3819,N_2450,N_2496);
nand U3820 (N_3820,N_2747,N_2897);
xnor U3821 (N_3821,N_2081,N_2893);
nand U3822 (N_3822,N_2104,N_2022);
and U3823 (N_3823,N_2108,N_2884);
and U3824 (N_3824,N_2703,N_2492);
or U3825 (N_3825,N_2739,N_2341);
nor U3826 (N_3826,N_2718,N_2812);
and U3827 (N_3827,N_2967,N_2686);
or U3828 (N_3828,N_2340,N_2188);
and U3829 (N_3829,N_2859,N_2244);
nand U3830 (N_3830,N_2794,N_2323);
or U3831 (N_3831,N_2817,N_2340);
nor U3832 (N_3832,N_2897,N_2364);
and U3833 (N_3833,N_2557,N_2881);
or U3834 (N_3834,N_2382,N_2946);
and U3835 (N_3835,N_2401,N_2071);
xnor U3836 (N_3836,N_2721,N_2919);
nor U3837 (N_3837,N_2154,N_2184);
nand U3838 (N_3838,N_2404,N_2599);
or U3839 (N_3839,N_2479,N_2776);
nand U3840 (N_3840,N_2787,N_2651);
or U3841 (N_3841,N_2047,N_2527);
nand U3842 (N_3842,N_2796,N_2680);
and U3843 (N_3843,N_2132,N_2636);
nor U3844 (N_3844,N_2335,N_2391);
xor U3845 (N_3845,N_2678,N_2607);
and U3846 (N_3846,N_2577,N_2409);
or U3847 (N_3847,N_2212,N_2309);
nand U3848 (N_3848,N_2513,N_2832);
nand U3849 (N_3849,N_2400,N_2478);
xnor U3850 (N_3850,N_2058,N_2099);
nor U3851 (N_3851,N_2352,N_2551);
and U3852 (N_3852,N_2410,N_2567);
and U3853 (N_3853,N_2789,N_2744);
or U3854 (N_3854,N_2348,N_2105);
nand U3855 (N_3855,N_2760,N_2094);
nand U3856 (N_3856,N_2590,N_2723);
nor U3857 (N_3857,N_2653,N_2647);
xnor U3858 (N_3858,N_2777,N_2588);
or U3859 (N_3859,N_2671,N_2069);
nand U3860 (N_3860,N_2016,N_2382);
xnor U3861 (N_3861,N_2427,N_2728);
or U3862 (N_3862,N_2018,N_2700);
nor U3863 (N_3863,N_2832,N_2624);
or U3864 (N_3864,N_2745,N_2900);
nand U3865 (N_3865,N_2537,N_2417);
and U3866 (N_3866,N_2169,N_2590);
nor U3867 (N_3867,N_2995,N_2296);
or U3868 (N_3868,N_2044,N_2499);
xor U3869 (N_3869,N_2335,N_2991);
xor U3870 (N_3870,N_2375,N_2718);
or U3871 (N_3871,N_2764,N_2642);
and U3872 (N_3872,N_2302,N_2438);
xnor U3873 (N_3873,N_2654,N_2979);
nand U3874 (N_3874,N_2869,N_2761);
nor U3875 (N_3875,N_2827,N_2547);
or U3876 (N_3876,N_2475,N_2434);
xnor U3877 (N_3877,N_2105,N_2622);
nand U3878 (N_3878,N_2780,N_2047);
xor U3879 (N_3879,N_2009,N_2824);
xor U3880 (N_3880,N_2935,N_2809);
nand U3881 (N_3881,N_2408,N_2477);
and U3882 (N_3882,N_2731,N_2038);
or U3883 (N_3883,N_2937,N_2932);
nand U3884 (N_3884,N_2538,N_2542);
and U3885 (N_3885,N_2853,N_2450);
and U3886 (N_3886,N_2563,N_2498);
and U3887 (N_3887,N_2003,N_2125);
nand U3888 (N_3888,N_2421,N_2014);
nand U3889 (N_3889,N_2616,N_2938);
xnor U3890 (N_3890,N_2054,N_2343);
nand U3891 (N_3891,N_2561,N_2908);
and U3892 (N_3892,N_2682,N_2214);
and U3893 (N_3893,N_2399,N_2831);
nor U3894 (N_3894,N_2000,N_2317);
nor U3895 (N_3895,N_2850,N_2234);
or U3896 (N_3896,N_2311,N_2956);
xor U3897 (N_3897,N_2568,N_2822);
xor U3898 (N_3898,N_2317,N_2962);
nand U3899 (N_3899,N_2341,N_2295);
nand U3900 (N_3900,N_2366,N_2112);
or U3901 (N_3901,N_2337,N_2134);
nand U3902 (N_3902,N_2241,N_2455);
and U3903 (N_3903,N_2709,N_2612);
nor U3904 (N_3904,N_2301,N_2360);
or U3905 (N_3905,N_2437,N_2459);
or U3906 (N_3906,N_2603,N_2683);
and U3907 (N_3907,N_2539,N_2495);
and U3908 (N_3908,N_2856,N_2579);
xor U3909 (N_3909,N_2238,N_2748);
xnor U3910 (N_3910,N_2516,N_2370);
and U3911 (N_3911,N_2154,N_2556);
and U3912 (N_3912,N_2474,N_2503);
nor U3913 (N_3913,N_2765,N_2910);
and U3914 (N_3914,N_2743,N_2223);
or U3915 (N_3915,N_2035,N_2669);
xnor U3916 (N_3916,N_2674,N_2416);
nor U3917 (N_3917,N_2458,N_2441);
or U3918 (N_3918,N_2896,N_2589);
xnor U3919 (N_3919,N_2189,N_2169);
or U3920 (N_3920,N_2667,N_2274);
and U3921 (N_3921,N_2645,N_2698);
and U3922 (N_3922,N_2218,N_2018);
and U3923 (N_3923,N_2821,N_2328);
xor U3924 (N_3924,N_2115,N_2228);
xnor U3925 (N_3925,N_2905,N_2556);
or U3926 (N_3926,N_2788,N_2401);
and U3927 (N_3927,N_2643,N_2481);
or U3928 (N_3928,N_2274,N_2781);
nand U3929 (N_3929,N_2421,N_2758);
and U3930 (N_3930,N_2620,N_2410);
xnor U3931 (N_3931,N_2963,N_2704);
xor U3932 (N_3932,N_2181,N_2306);
nand U3933 (N_3933,N_2469,N_2373);
nor U3934 (N_3934,N_2769,N_2197);
and U3935 (N_3935,N_2419,N_2281);
nand U3936 (N_3936,N_2642,N_2602);
nor U3937 (N_3937,N_2897,N_2771);
and U3938 (N_3938,N_2310,N_2239);
or U3939 (N_3939,N_2301,N_2363);
and U3940 (N_3940,N_2969,N_2224);
xnor U3941 (N_3941,N_2992,N_2876);
nand U3942 (N_3942,N_2274,N_2109);
nand U3943 (N_3943,N_2659,N_2472);
or U3944 (N_3944,N_2195,N_2929);
nor U3945 (N_3945,N_2938,N_2611);
or U3946 (N_3946,N_2039,N_2271);
or U3947 (N_3947,N_2608,N_2366);
nor U3948 (N_3948,N_2643,N_2129);
xnor U3949 (N_3949,N_2948,N_2698);
xor U3950 (N_3950,N_2522,N_2551);
xor U3951 (N_3951,N_2656,N_2599);
xor U3952 (N_3952,N_2780,N_2296);
nor U3953 (N_3953,N_2958,N_2643);
and U3954 (N_3954,N_2391,N_2306);
and U3955 (N_3955,N_2438,N_2948);
and U3956 (N_3956,N_2239,N_2649);
and U3957 (N_3957,N_2256,N_2722);
and U3958 (N_3958,N_2342,N_2018);
and U3959 (N_3959,N_2336,N_2150);
and U3960 (N_3960,N_2536,N_2262);
nand U3961 (N_3961,N_2049,N_2280);
nand U3962 (N_3962,N_2916,N_2956);
and U3963 (N_3963,N_2970,N_2009);
nor U3964 (N_3964,N_2982,N_2928);
xor U3965 (N_3965,N_2569,N_2789);
or U3966 (N_3966,N_2711,N_2478);
xor U3967 (N_3967,N_2130,N_2647);
and U3968 (N_3968,N_2205,N_2491);
xnor U3969 (N_3969,N_2835,N_2449);
xor U3970 (N_3970,N_2368,N_2187);
xor U3971 (N_3971,N_2730,N_2359);
xnor U3972 (N_3972,N_2889,N_2789);
and U3973 (N_3973,N_2107,N_2080);
or U3974 (N_3974,N_2442,N_2273);
nand U3975 (N_3975,N_2417,N_2051);
xor U3976 (N_3976,N_2947,N_2829);
nand U3977 (N_3977,N_2579,N_2382);
and U3978 (N_3978,N_2186,N_2998);
or U3979 (N_3979,N_2498,N_2315);
nor U3980 (N_3980,N_2211,N_2432);
nor U3981 (N_3981,N_2162,N_2909);
nand U3982 (N_3982,N_2196,N_2704);
xor U3983 (N_3983,N_2272,N_2629);
and U3984 (N_3984,N_2402,N_2901);
xnor U3985 (N_3985,N_2138,N_2334);
nand U3986 (N_3986,N_2087,N_2347);
xor U3987 (N_3987,N_2612,N_2515);
nand U3988 (N_3988,N_2483,N_2339);
xnor U3989 (N_3989,N_2387,N_2254);
xnor U3990 (N_3990,N_2066,N_2979);
xnor U3991 (N_3991,N_2512,N_2227);
or U3992 (N_3992,N_2777,N_2098);
nand U3993 (N_3993,N_2290,N_2707);
nor U3994 (N_3994,N_2842,N_2081);
nand U3995 (N_3995,N_2010,N_2671);
and U3996 (N_3996,N_2572,N_2466);
or U3997 (N_3997,N_2190,N_2271);
or U3998 (N_3998,N_2433,N_2932);
nand U3999 (N_3999,N_2178,N_2072);
xnor U4000 (N_4000,N_3714,N_3668);
or U4001 (N_4001,N_3495,N_3035);
nand U4002 (N_4002,N_3034,N_3690);
or U4003 (N_4003,N_3582,N_3775);
nor U4004 (N_4004,N_3733,N_3386);
and U4005 (N_4005,N_3122,N_3240);
nand U4006 (N_4006,N_3095,N_3967);
and U4007 (N_4007,N_3290,N_3719);
and U4008 (N_4008,N_3219,N_3633);
nand U4009 (N_4009,N_3667,N_3257);
or U4010 (N_4010,N_3760,N_3361);
xnor U4011 (N_4011,N_3119,N_3744);
nand U4012 (N_4012,N_3698,N_3265);
nand U4013 (N_4013,N_3634,N_3111);
xor U4014 (N_4014,N_3412,N_3162);
and U4015 (N_4015,N_3338,N_3716);
or U4016 (N_4016,N_3399,N_3340);
or U4017 (N_4017,N_3296,N_3453);
nor U4018 (N_4018,N_3170,N_3364);
and U4019 (N_4019,N_3770,N_3393);
or U4020 (N_4020,N_3443,N_3266);
or U4021 (N_4021,N_3485,N_3025);
xnor U4022 (N_4022,N_3596,N_3743);
nand U4023 (N_4023,N_3748,N_3853);
nor U4024 (N_4024,N_3534,N_3109);
and U4025 (N_4025,N_3751,N_3492);
xnor U4026 (N_4026,N_3304,N_3339);
nor U4027 (N_4027,N_3342,N_3628);
xnor U4028 (N_4028,N_3206,N_3632);
xnor U4029 (N_4029,N_3530,N_3823);
xor U4030 (N_4030,N_3283,N_3809);
xnor U4031 (N_4031,N_3933,N_3442);
nor U4032 (N_4032,N_3981,N_3145);
nand U4033 (N_4033,N_3850,N_3523);
and U4034 (N_4034,N_3227,N_3235);
nor U4035 (N_4035,N_3237,N_3648);
and U4036 (N_4036,N_3631,N_3303);
xor U4037 (N_4037,N_3154,N_3677);
xor U4038 (N_4038,N_3645,N_3194);
nor U4039 (N_4039,N_3647,N_3644);
nand U4040 (N_4040,N_3594,N_3216);
or U4041 (N_4041,N_3384,N_3617);
nand U4042 (N_4042,N_3790,N_3620);
nor U4043 (N_4043,N_3651,N_3357);
xor U4044 (N_4044,N_3861,N_3787);
or U4045 (N_4045,N_3293,N_3316);
xnor U4046 (N_4046,N_3599,N_3333);
xnor U4047 (N_4047,N_3778,N_3993);
xor U4048 (N_4048,N_3942,N_3734);
nand U4049 (N_4049,N_3371,N_3121);
and U4050 (N_4050,N_3230,N_3687);
and U4051 (N_4051,N_3782,N_3321);
nand U4052 (N_4052,N_3066,N_3385);
nor U4053 (N_4053,N_3045,N_3053);
and U4054 (N_4054,N_3692,N_3000);
xnor U4055 (N_4055,N_3577,N_3073);
nor U4056 (N_4056,N_3909,N_3921);
xor U4057 (N_4057,N_3973,N_3642);
nor U4058 (N_4058,N_3837,N_3991);
or U4059 (N_4059,N_3876,N_3014);
or U4060 (N_4060,N_3722,N_3448);
and U4061 (N_4061,N_3426,N_3427);
or U4062 (N_4062,N_3750,N_3246);
nor U4063 (N_4063,N_3055,N_3831);
and U4064 (N_4064,N_3047,N_3626);
or U4065 (N_4065,N_3226,N_3430);
xor U4066 (N_4066,N_3297,N_3665);
nand U4067 (N_4067,N_3182,N_3406);
nand U4068 (N_4068,N_3982,N_3950);
or U4069 (N_4069,N_3558,N_3540);
and U4070 (N_4070,N_3440,N_3560);
nand U4071 (N_4071,N_3731,N_3769);
nand U4072 (N_4072,N_3354,N_3874);
nor U4073 (N_4073,N_3317,N_3204);
and U4074 (N_4074,N_3435,N_3675);
nor U4075 (N_4075,N_3187,N_3547);
and U4076 (N_4076,N_3525,N_3327);
or U4077 (N_4077,N_3489,N_3139);
nand U4078 (N_4078,N_3067,N_3539);
nor U4079 (N_4079,N_3796,N_3922);
xor U4080 (N_4080,N_3330,N_3925);
and U4081 (N_4081,N_3134,N_3264);
and U4082 (N_4082,N_3696,N_3137);
nand U4083 (N_4083,N_3421,N_3510);
nand U4084 (N_4084,N_3177,N_3612);
or U4085 (N_4085,N_3484,N_3031);
nor U4086 (N_4086,N_3012,N_3326);
and U4087 (N_4087,N_3693,N_3019);
nand U4088 (N_4088,N_3550,N_3509);
xnor U4089 (N_4089,N_3449,N_3715);
xor U4090 (N_4090,N_3927,N_3171);
and U4091 (N_4091,N_3411,N_3070);
nor U4092 (N_4092,N_3001,N_3306);
or U4093 (N_4093,N_3507,N_3807);
and U4094 (N_4094,N_3115,N_3179);
or U4095 (N_4095,N_3475,N_3476);
nand U4096 (N_4096,N_3280,N_3195);
and U4097 (N_4097,N_3463,N_3785);
or U4098 (N_4098,N_3803,N_3926);
or U4099 (N_4099,N_3752,N_3804);
xnor U4100 (N_4100,N_3720,N_3331);
nand U4101 (N_4101,N_3941,N_3199);
or U4102 (N_4102,N_3639,N_3900);
or U4103 (N_4103,N_3346,N_3858);
nand U4104 (N_4104,N_3906,N_3867);
xor U4105 (N_4105,N_3027,N_3986);
nor U4106 (N_4106,N_3875,N_3060);
and U4107 (N_4107,N_3834,N_3018);
nand U4108 (N_4108,N_3529,N_3072);
nor U4109 (N_4109,N_3201,N_3205);
nand U4110 (N_4110,N_3358,N_3937);
and U4111 (N_4111,N_3746,N_3781);
and U4112 (N_4112,N_3629,N_3441);
and U4113 (N_4113,N_3911,N_3854);
and U4114 (N_4114,N_3533,N_3113);
nor U4115 (N_4115,N_3994,N_3640);
and U4116 (N_4116,N_3190,N_3168);
nor U4117 (N_4117,N_3310,N_3949);
nand U4118 (N_4118,N_3849,N_3603);
and U4119 (N_4119,N_3857,N_3673);
xnor U4120 (N_4120,N_3975,N_3391);
xor U4121 (N_4121,N_3284,N_3488);
nor U4122 (N_4122,N_3299,N_3256);
xnor U4123 (N_4123,N_3880,N_3706);
nor U4124 (N_4124,N_3788,N_3436);
or U4125 (N_4125,N_3118,N_3897);
xor U4126 (N_4126,N_3583,N_3173);
and U4127 (N_4127,N_3983,N_3958);
or U4128 (N_4128,N_3151,N_3092);
xor U4129 (N_4129,N_3120,N_3050);
xnor U4130 (N_4130,N_3262,N_3380);
or U4131 (N_4131,N_3253,N_3097);
nor U4132 (N_4132,N_3052,N_3150);
xor U4133 (N_4133,N_3791,N_3281);
nand U4134 (N_4134,N_3381,N_3130);
or U4135 (N_4135,N_3520,N_3784);
or U4136 (N_4136,N_3254,N_3434);
and U4137 (N_4137,N_3474,N_3270);
or U4138 (N_4138,N_3812,N_3454);
nor U4139 (N_4139,N_3901,N_3353);
and U4140 (N_4140,N_3163,N_3564);
xnor U4141 (N_4141,N_3833,N_3565);
or U4142 (N_4142,N_3329,N_3079);
nor U4143 (N_4143,N_3061,N_3010);
nand U4144 (N_4144,N_3102,N_3222);
nand U4145 (N_4145,N_3239,N_3409);
and U4146 (N_4146,N_3541,N_3836);
nand U4147 (N_4147,N_3248,N_3548);
and U4148 (N_4148,N_3932,N_3532);
xor U4149 (N_4149,N_3585,N_3657);
nor U4150 (N_4150,N_3065,N_3242);
nor U4151 (N_4151,N_3478,N_3114);
or U4152 (N_4152,N_3980,N_3368);
nand U4153 (N_4153,N_3502,N_3255);
nand U4154 (N_4154,N_3158,N_3403);
nor U4155 (N_4155,N_3268,N_3100);
nor U4156 (N_4156,N_3700,N_3398);
nor U4157 (N_4157,N_3608,N_3269);
or U4158 (N_4158,N_3439,N_3649);
xor U4159 (N_4159,N_3997,N_3924);
nand U4160 (N_4160,N_3383,N_3519);
and U4161 (N_4161,N_3496,N_3389);
xnor U4162 (N_4162,N_3486,N_3159);
nor U4163 (N_4163,N_3483,N_3210);
nor U4164 (N_4164,N_3978,N_3652);
nand U4165 (N_4165,N_3049,N_3545);
or U4166 (N_4166,N_3869,N_3930);
or U4167 (N_4167,N_3062,N_3007);
nor U4168 (N_4168,N_3511,N_3522);
and U4169 (N_4169,N_3919,N_3780);
xnor U4170 (N_4170,N_3971,N_3311);
nand U4171 (N_4171,N_3712,N_3605);
nand U4172 (N_4172,N_3660,N_3963);
or U4173 (N_4173,N_3043,N_3749);
xnor U4174 (N_4174,N_3462,N_3078);
xnor U4175 (N_4175,N_3764,N_3797);
xnor U4176 (N_4176,N_3955,N_3684);
xnor U4177 (N_4177,N_3029,N_3970);
or U4178 (N_4178,N_3531,N_3838);
nand U4179 (N_4179,N_3241,N_3249);
xor U4180 (N_4180,N_3794,N_3087);
nand U4181 (N_4181,N_3378,N_3360);
nor U4182 (N_4182,N_3951,N_3597);
nor U4183 (N_4183,N_3590,N_3627);
or U4184 (N_4184,N_3192,N_3345);
and U4185 (N_4185,N_3929,N_3776);
xnor U4186 (N_4186,N_3777,N_3789);
nand U4187 (N_4187,N_3745,N_3625);
or U4188 (N_4188,N_3505,N_3370);
nor U4189 (N_4189,N_3455,N_3064);
nor U4190 (N_4190,N_3783,N_3862);
nor U4191 (N_4191,N_3977,N_3197);
or U4192 (N_4192,N_3814,N_3252);
nor U4193 (N_4193,N_3232,N_3428);
or U4194 (N_4194,N_3236,N_3431);
xor U4195 (N_4195,N_3414,N_3902);
or U4196 (N_4196,N_3215,N_3481);
nand U4197 (N_4197,N_3573,N_3717);
xor U4198 (N_4198,N_3878,N_3362);
nand U4199 (N_4199,N_3852,N_3891);
xnor U4200 (N_4200,N_3148,N_3135);
or U4201 (N_4201,N_3524,N_3294);
nor U4202 (N_4202,N_3388,N_3437);
and U4203 (N_4203,N_3143,N_3348);
nand U4204 (N_4204,N_3905,N_3843);
and U4205 (N_4205,N_3356,N_3013);
nand U4206 (N_4206,N_3416,N_3638);
xor U4207 (N_4207,N_3363,N_3664);
nor U4208 (N_4208,N_3469,N_3438);
xnor U4209 (N_4209,N_3466,N_3309);
nor U4210 (N_4210,N_3107,N_3198);
nand U4211 (N_4211,N_3518,N_3561);
xor U4212 (N_4212,N_3133,N_3557);
nand U4213 (N_4213,N_3952,N_3445);
nand U4214 (N_4214,N_3225,N_3334);
and U4215 (N_4215,N_3395,N_3737);
and U4216 (N_4216,N_3429,N_3322);
and U4217 (N_4217,N_3931,N_3813);
and U4218 (N_4218,N_3514,N_3709);
nor U4219 (N_4219,N_3732,N_3680);
or U4220 (N_4220,N_3887,N_3772);
and U4221 (N_4221,N_3726,N_3576);
and U4222 (N_4222,N_3131,N_3451);
nor U4223 (N_4223,N_3944,N_3915);
nor U4224 (N_4224,N_3003,N_3051);
nand U4225 (N_4225,N_3404,N_3761);
or U4226 (N_4226,N_3465,N_3160);
or U4227 (N_4227,N_3422,N_3279);
nand U4228 (N_4228,N_3609,N_3471);
or U4229 (N_4229,N_3824,N_3801);
and U4230 (N_4230,N_3058,N_3593);
or U4231 (N_4231,N_3352,N_3896);
and U4232 (N_4232,N_3636,N_3152);
nor U4233 (N_4233,N_3702,N_3817);
and U4234 (N_4234,N_3211,N_3196);
xnor U4235 (N_4235,N_3260,N_3417);
or U4236 (N_4236,N_3341,N_3820);
and U4237 (N_4237,N_3077,N_3332);
xor U4238 (N_4238,N_3105,N_3735);
nand U4239 (N_4239,N_3841,N_3730);
nor U4240 (N_4240,N_3851,N_3091);
or U4241 (N_4241,N_3659,N_3366);
xnor U4242 (N_4242,N_3763,N_3859);
and U4243 (N_4243,N_3866,N_3899);
nor U4244 (N_4244,N_3459,N_3798);
and U4245 (N_4245,N_3602,N_3826);
or U4246 (N_4246,N_3569,N_3579);
or U4247 (N_4247,N_3877,N_3572);
nand U4248 (N_4248,N_3074,N_3960);
and U4249 (N_4249,N_3935,N_3491);
or U4250 (N_4250,N_3450,N_3616);
xor U4251 (N_4251,N_3089,N_3699);
xor U4252 (N_4252,N_3116,N_3995);
and U4253 (N_4253,N_3099,N_3968);
or U4254 (N_4254,N_3598,N_3879);
xor U4255 (N_4255,N_3164,N_3390);
nor U4256 (N_4256,N_3372,N_3203);
xnor U4257 (N_4257,N_3493,N_3516);
xor U4258 (N_4258,N_3703,N_3992);
xor U4259 (N_4259,N_3166,N_3032);
or U4260 (N_4260,N_3976,N_3231);
nor U4261 (N_4261,N_3661,N_3167);
nand U4262 (N_4262,N_3953,N_3882);
and U4263 (N_4263,N_3856,N_3697);
nand U4264 (N_4264,N_3085,N_3132);
nor U4265 (N_4265,N_3607,N_3956);
or U4266 (N_4266,N_3587,N_3604);
and U4267 (N_4267,N_3456,N_3815);
and U4268 (N_4268,N_3056,N_3172);
and U4269 (N_4269,N_3267,N_3433);
xnor U4270 (N_4270,N_3217,N_3189);
xor U4271 (N_4271,N_3979,N_3282);
and U4272 (N_4272,N_3526,N_3020);
or U4273 (N_4273,N_3939,N_3917);
nor U4274 (N_4274,N_3839,N_3562);
or U4275 (N_4275,N_3611,N_3324);
and U4276 (N_4276,N_3552,N_3914);
nand U4277 (N_4277,N_3903,N_3487);
and U4278 (N_4278,N_3081,N_3397);
and U4279 (N_4279,N_3832,N_3128);
or U4280 (N_4280,N_3300,N_3946);
nand U4281 (N_4281,N_3767,N_3676);
or U4282 (N_4282,N_3972,N_3894);
xnor U4283 (N_4283,N_3947,N_3402);
or U4284 (N_4284,N_3098,N_3344);
or U4285 (N_4285,N_3872,N_3575);
nand U4286 (N_4286,N_3373,N_3457);
nor U4287 (N_4287,N_3472,N_3110);
and U4288 (N_4288,N_3512,N_3305);
nor U4289 (N_4289,N_3686,N_3985);
and U4290 (N_4290,N_3473,N_3806);
or U4291 (N_4291,N_3885,N_3041);
nor U4292 (N_4292,N_3606,N_3551);
and U4293 (N_4293,N_3654,N_3563);
nor U4294 (N_4294,N_3556,N_3347);
and U4295 (N_4295,N_3298,N_3084);
and U4296 (N_4296,N_3191,N_3238);
and U4297 (N_4297,N_3635,N_3846);
and U4298 (N_4298,N_3538,N_3088);
or U4299 (N_4299,N_3233,N_3940);
xnor U4300 (N_4300,N_3508,N_3889);
nor U4301 (N_4301,N_3016,N_3028);
or U4302 (N_4302,N_3277,N_3181);
nand U4303 (N_4303,N_3689,N_3499);
and U4304 (N_4304,N_3873,N_3679);
xor U4305 (N_4305,N_3106,N_3033);
or U4306 (N_4306,N_3276,N_3234);
nor U4307 (N_4307,N_3096,N_3643);
xnor U4308 (N_4308,N_3786,N_3452);
nor U4309 (N_4309,N_3537,N_3581);
and U4310 (N_4310,N_3666,N_3374);
nor U4311 (N_4311,N_3757,N_3646);
nor U4312 (N_4312,N_3498,N_3365);
and U4313 (N_4313,N_3319,N_3723);
or U4314 (N_4314,N_3708,N_3559);
and U4315 (N_4315,N_3678,N_3669);
nand U4316 (N_4316,N_3998,N_3916);
nor U4317 (N_4317,N_3740,N_3890);
and U4318 (N_4318,N_3822,N_3721);
xor U4319 (N_4319,N_3432,N_3580);
xnor U4320 (N_4320,N_3287,N_3934);
or U4321 (N_4321,N_3711,N_3251);
xnor U4322 (N_4322,N_3136,N_3910);
nor U4323 (N_4323,N_3584,N_3595);
nor U4324 (N_4324,N_3323,N_3747);
xor U4325 (N_4325,N_3273,N_3213);
and U4326 (N_4326,N_3835,N_3288);
or U4327 (N_4327,N_3355,N_3513);
xnor U4328 (N_4328,N_3036,N_3156);
nor U4329 (N_4329,N_3369,N_3774);
nand U4330 (N_4330,N_3765,N_3407);
or U4331 (N_4331,N_3614,N_3157);
or U4332 (N_4332,N_3844,N_3069);
xnor U4333 (N_4333,N_3707,N_3908);
xor U4334 (N_4334,N_3898,N_3637);
nand U4335 (N_4335,N_3695,N_3479);
nor U4336 (N_4336,N_3379,N_3554);
nor U4337 (N_4337,N_3185,N_3229);
and U4338 (N_4338,N_3688,N_3672);
nand U4339 (N_4339,N_3082,N_3123);
and U4340 (N_4340,N_3682,N_3691);
or U4341 (N_4341,N_3101,N_3694);
or U4342 (N_4342,N_3002,N_3913);
nor U4343 (N_4343,N_3223,N_3104);
xor U4344 (N_4344,N_3758,N_3653);
and U4345 (N_4345,N_3615,N_3202);
and U4346 (N_4346,N_3176,N_3742);
nor U4347 (N_4347,N_3004,N_3009);
xnor U4348 (N_4348,N_3655,N_3870);
nor U4349 (N_4349,N_3613,N_3893);
or U4350 (N_4350,N_3186,N_3650);
or U4351 (N_4351,N_3816,N_3965);
nand U4352 (N_4352,N_3588,N_3800);
xnor U4353 (N_4353,N_3161,N_3146);
xnor U4354 (N_4354,N_3313,N_3762);
nand U4355 (N_4355,N_3291,N_3943);
xnor U4356 (N_4356,N_3302,N_3753);
nand U4357 (N_4357,N_3671,N_3243);
and U4358 (N_4358,N_3567,N_3108);
or U4359 (N_4359,N_3022,N_3601);
xnor U4360 (N_4360,N_3871,N_3005);
xor U4361 (N_4361,N_3656,N_3335);
nor U4362 (N_4362,N_3336,N_3208);
xor U4363 (N_4363,N_3006,N_3802);
or U4364 (N_4364,N_3739,N_3506);
or U4365 (N_4365,N_3536,N_3521);
nand U4366 (N_4366,N_3966,N_3497);
and U4367 (N_4367,N_3895,N_3883);
nor U4368 (N_4368,N_3553,N_3470);
and U4369 (N_4369,N_3017,N_3881);
and U4370 (N_4370,N_3945,N_3415);
nand U4371 (N_4371,N_3458,N_3125);
and U4372 (N_4372,N_3250,N_3845);
nand U4373 (N_4373,N_3984,N_3461);
or U4374 (N_4374,N_3912,N_3888);
and U4375 (N_4375,N_3543,N_3054);
xnor U4376 (N_4376,N_3075,N_3500);
xnor U4377 (N_4377,N_3670,N_3544);
and U4378 (N_4378,N_3863,N_3408);
and U4379 (N_4379,N_3295,N_3535);
xnor U4380 (N_4380,N_3375,N_3907);
nand U4381 (N_4381,N_3989,N_3987);
or U4382 (N_4382,N_3755,N_3261);
nor U4383 (N_4383,N_3424,N_3188);
xor U4384 (N_4384,N_3771,N_3701);
nor U4385 (N_4385,N_3400,N_3566);
and U4386 (N_4386,N_3738,N_3418);
nand U4387 (N_4387,N_3200,N_3258);
nand U4388 (N_4388,N_3938,N_3289);
nor U4389 (N_4389,N_3312,N_3224);
nor U4390 (N_4390,N_3142,N_3271);
nor U4391 (N_4391,N_3278,N_3865);
or U4392 (N_4392,N_3343,N_3377);
nor U4393 (N_4393,N_3884,N_3828);
nor U4394 (N_4394,N_3517,N_3090);
xnor U4395 (N_4395,N_3259,N_3528);
nor U4396 (N_4396,N_3568,N_3570);
nor U4397 (N_4397,N_3207,N_3503);
nor U4398 (N_4398,N_3795,N_3964);
nor U4399 (N_4399,N_3674,N_3359);
nand U4400 (N_4400,N_3328,N_3600);
nand U4401 (N_4401,N_3076,N_3209);
nor U4402 (N_4402,N_3808,N_3821);
or U4403 (N_4403,N_3094,N_3630);
and U4404 (N_4404,N_3292,N_3245);
xor U4405 (N_4405,N_3504,N_3117);
nor U4406 (N_4406,N_3464,N_3923);
xnor U4407 (N_4407,N_3999,N_3044);
nor U4408 (N_4408,N_3126,N_3768);
xnor U4409 (N_4409,N_3658,N_3578);
xor U4410 (N_4410,N_3141,N_3446);
xnor U4411 (N_4411,N_3618,N_3165);
xor U4412 (N_4412,N_3480,N_3015);
nor U4413 (N_4413,N_3683,N_3904);
nand U4414 (N_4414,N_3546,N_3641);
nor U4415 (N_4415,N_3829,N_3990);
nand U4416 (N_4416,N_3286,N_3112);
nor U4417 (N_4417,N_3855,N_3527);
and U4418 (N_4418,N_3405,N_3827);
nand U4419 (N_4419,N_3024,N_3221);
or U4420 (N_4420,N_3713,N_3140);
and U4421 (N_4421,N_3149,N_3124);
nor U4422 (N_4422,N_3961,N_3685);
nand U4423 (N_4423,N_3218,N_3811);
xnor U4424 (N_4424,N_3423,N_3467);
or U4425 (N_4425,N_3792,N_3367);
nand U4426 (N_4426,N_3799,N_3663);
nand U4427 (N_4427,N_3093,N_3301);
nand U4428 (N_4428,N_3220,N_3460);
xnor U4429 (N_4429,N_3840,N_3392);
nand U4430 (N_4430,N_3969,N_3482);
and U4431 (N_4431,N_3325,N_3957);
or U4432 (N_4432,N_3996,N_3830);
or U4433 (N_4433,N_3728,N_3574);
and U4434 (N_4434,N_3621,N_3350);
or U4435 (N_4435,N_3244,N_3619);
or U4436 (N_4436,N_3959,N_3030);
xnor U4437 (N_4437,N_3810,N_3410);
nand U4438 (N_4438,N_3586,N_3842);
xor U4439 (N_4439,N_3623,N_3180);
nand U4440 (N_4440,N_3401,N_3039);
and U4441 (N_4441,N_3736,N_3228);
nand U4442 (N_4442,N_3184,N_3396);
nand U4443 (N_4443,N_3274,N_3129);
nand U4444 (N_4444,N_3962,N_3549);
and U4445 (N_4445,N_3420,N_3083);
or U4446 (N_4446,N_3555,N_3936);
or U4447 (N_4447,N_3718,N_3622);
xnor U4448 (N_4448,N_3494,N_3848);
xnor U4449 (N_4449,N_3754,N_3477);
and U4450 (N_4450,N_3272,N_3805);
or U4451 (N_4451,N_3175,N_3868);
nand U4452 (N_4452,N_3954,N_3023);
or U4453 (N_4453,N_3918,N_3021);
or U4454 (N_4454,N_3928,N_3610);
and U4455 (N_4455,N_3727,N_3103);
nand U4456 (N_4456,N_3042,N_3263);
and U4457 (N_4457,N_3068,N_3756);
xnor U4458 (N_4458,N_3040,N_3307);
and U4459 (N_4459,N_3444,N_3315);
or U4460 (N_4460,N_3193,N_3046);
nor U4461 (N_4461,N_3948,N_3773);
and U4462 (N_4462,N_3178,N_3860);
nor U4463 (N_4463,N_3825,N_3725);
and U4464 (N_4464,N_3155,N_3988);
nor U4465 (N_4465,N_3886,N_3144);
nor U4466 (N_4466,N_3490,N_3394);
xor U4467 (N_4467,N_3864,N_3314);
xnor U4468 (N_4468,N_3382,N_3501);
nor U4469 (N_4469,N_3447,N_3153);
nor U4470 (N_4470,N_3212,N_3071);
nor U4471 (N_4471,N_3413,N_3705);
nor U4472 (N_4472,N_3320,N_3425);
xnor U4473 (N_4473,N_3086,N_3308);
or U4474 (N_4474,N_3169,N_3847);
and U4475 (N_4475,N_3048,N_3147);
nor U4476 (N_4476,N_3275,N_3337);
or U4477 (N_4477,N_3419,N_3920);
or U4478 (N_4478,N_3892,N_3351);
and U4479 (N_4479,N_3080,N_3681);
and U4480 (N_4480,N_3008,N_3247);
xor U4481 (N_4481,N_3724,N_3038);
or U4482 (N_4482,N_3138,N_3349);
xor U4483 (N_4483,N_3729,N_3057);
nor U4484 (N_4484,N_3571,N_3174);
nand U4485 (N_4485,N_3387,N_3037);
nor U4486 (N_4486,N_3376,N_3059);
nand U4487 (N_4487,N_3819,N_3624);
nor U4488 (N_4488,N_3127,N_3741);
xor U4489 (N_4489,N_3592,N_3759);
xor U4490 (N_4490,N_3766,N_3214);
nand U4491 (N_4491,N_3662,N_3818);
xor U4492 (N_4492,N_3318,N_3710);
nand U4493 (N_4493,N_3285,N_3704);
nand U4494 (N_4494,N_3974,N_3515);
xor U4495 (N_4495,N_3591,N_3468);
or U4496 (N_4496,N_3183,N_3589);
and U4497 (N_4497,N_3011,N_3026);
nor U4498 (N_4498,N_3793,N_3779);
nand U4499 (N_4499,N_3542,N_3063);
nand U4500 (N_4500,N_3834,N_3210);
or U4501 (N_4501,N_3757,N_3082);
and U4502 (N_4502,N_3781,N_3760);
and U4503 (N_4503,N_3208,N_3409);
nand U4504 (N_4504,N_3115,N_3877);
or U4505 (N_4505,N_3145,N_3757);
nor U4506 (N_4506,N_3913,N_3729);
nand U4507 (N_4507,N_3822,N_3814);
and U4508 (N_4508,N_3938,N_3043);
nor U4509 (N_4509,N_3045,N_3886);
and U4510 (N_4510,N_3876,N_3611);
nand U4511 (N_4511,N_3269,N_3171);
nand U4512 (N_4512,N_3821,N_3757);
and U4513 (N_4513,N_3520,N_3267);
or U4514 (N_4514,N_3854,N_3617);
nand U4515 (N_4515,N_3192,N_3692);
and U4516 (N_4516,N_3783,N_3242);
xor U4517 (N_4517,N_3785,N_3843);
or U4518 (N_4518,N_3131,N_3860);
nor U4519 (N_4519,N_3422,N_3812);
nand U4520 (N_4520,N_3118,N_3159);
and U4521 (N_4521,N_3014,N_3833);
xnor U4522 (N_4522,N_3630,N_3973);
and U4523 (N_4523,N_3436,N_3353);
or U4524 (N_4524,N_3018,N_3246);
xor U4525 (N_4525,N_3243,N_3673);
nor U4526 (N_4526,N_3872,N_3356);
xnor U4527 (N_4527,N_3652,N_3558);
nand U4528 (N_4528,N_3659,N_3564);
nand U4529 (N_4529,N_3659,N_3729);
xor U4530 (N_4530,N_3854,N_3130);
or U4531 (N_4531,N_3987,N_3391);
xnor U4532 (N_4532,N_3765,N_3369);
and U4533 (N_4533,N_3495,N_3281);
and U4534 (N_4534,N_3643,N_3204);
and U4535 (N_4535,N_3819,N_3470);
nand U4536 (N_4536,N_3852,N_3698);
nor U4537 (N_4537,N_3201,N_3923);
nand U4538 (N_4538,N_3772,N_3347);
xor U4539 (N_4539,N_3005,N_3478);
or U4540 (N_4540,N_3807,N_3351);
nor U4541 (N_4541,N_3905,N_3305);
or U4542 (N_4542,N_3879,N_3090);
nand U4543 (N_4543,N_3464,N_3903);
xor U4544 (N_4544,N_3182,N_3108);
nand U4545 (N_4545,N_3017,N_3031);
and U4546 (N_4546,N_3251,N_3584);
nand U4547 (N_4547,N_3210,N_3787);
xor U4548 (N_4548,N_3217,N_3486);
or U4549 (N_4549,N_3484,N_3449);
nand U4550 (N_4550,N_3868,N_3769);
nor U4551 (N_4551,N_3585,N_3038);
nand U4552 (N_4552,N_3206,N_3720);
or U4553 (N_4553,N_3674,N_3239);
and U4554 (N_4554,N_3488,N_3640);
or U4555 (N_4555,N_3419,N_3264);
or U4556 (N_4556,N_3792,N_3188);
nor U4557 (N_4557,N_3217,N_3251);
or U4558 (N_4558,N_3174,N_3757);
nor U4559 (N_4559,N_3442,N_3181);
nand U4560 (N_4560,N_3072,N_3379);
or U4561 (N_4561,N_3014,N_3228);
nand U4562 (N_4562,N_3753,N_3047);
nand U4563 (N_4563,N_3777,N_3371);
xor U4564 (N_4564,N_3800,N_3794);
nor U4565 (N_4565,N_3080,N_3358);
nor U4566 (N_4566,N_3194,N_3460);
nor U4567 (N_4567,N_3912,N_3734);
or U4568 (N_4568,N_3128,N_3066);
nor U4569 (N_4569,N_3570,N_3046);
nand U4570 (N_4570,N_3557,N_3900);
and U4571 (N_4571,N_3226,N_3722);
or U4572 (N_4572,N_3282,N_3581);
and U4573 (N_4573,N_3679,N_3782);
and U4574 (N_4574,N_3390,N_3007);
and U4575 (N_4575,N_3345,N_3483);
nand U4576 (N_4576,N_3584,N_3751);
nor U4577 (N_4577,N_3407,N_3218);
or U4578 (N_4578,N_3704,N_3465);
and U4579 (N_4579,N_3541,N_3648);
nor U4580 (N_4580,N_3065,N_3417);
or U4581 (N_4581,N_3832,N_3106);
nand U4582 (N_4582,N_3372,N_3003);
xnor U4583 (N_4583,N_3351,N_3091);
nor U4584 (N_4584,N_3653,N_3429);
nand U4585 (N_4585,N_3594,N_3441);
nor U4586 (N_4586,N_3087,N_3549);
or U4587 (N_4587,N_3386,N_3392);
or U4588 (N_4588,N_3068,N_3292);
xnor U4589 (N_4589,N_3343,N_3419);
xor U4590 (N_4590,N_3718,N_3299);
xor U4591 (N_4591,N_3803,N_3244);
nand U4592 (N_4592,N_3327,N_3228);
or U4593 (N_4593,N_3096,N_3724);
and U4594 (N_4594,N_3699,N_3480);
nand U4595 (N_4595,N_3548,N_3037);
nor U4596 (N_4596,N_3071,N_3439);
xor U4597 (N_4597,N_3492,N_3408);
xnor U4598 (N_4598,N_3439,N_3011);
nor U4599 (N_4599,N_3966,N_3624);
and U4600 (N_4600,N_3749,N_3951);
xnor U4601 (N_4601,N_3816,N_3406);
nor U4602 (N_4602,N_3850,N_3592);
xnor U4603 (N_4603,N_3291,N_3605);
nand U4604 (N_4604,N_3717,N_3292);
xnor U4605 (N_4605,N_3557,N_3111);
or U4606 (N_4606,N_3785,N_3751);
or U4607 (N_4607,N_3256,N_3977);
xnor U4608 (N_4608,N_3415,N_3446);
and U4609 (N_4609,N_3012,N_3243);
xor U4610 (N_4610,N_3864,N_3319);
nor U4611 (N_4611,N_3134,N_3216);
nor U4612 (N_4612,N_3922,N_3378);
or U4613 (N_4613,N_3596,N_3783);
xor U4614 (N_4614,N_3442,N_3825);
nand U4615 (N_4615,N_3781,N_3355);
nand U4616 (N_4616,N_3082,N_3693);
nor U4617 (N_4617,N_3212,N_3181);
nor U4618 (N_4618,N_3872,N_3134);
or U4619 (N_4619,N_3408,N_3452);
xor U4620 (N_4620,N_3791,N_3018);
nor U4621 (N_4621,N_3253,N_3350);
nand U4622 (N_4622,N_3296,N_3614);
xnor U4623 (N_4623,N_3710,N_3449);
and U4624 (N_4624,N_3251,N_3068);
and U4625 (N_4625,N_3478,N_3705);
xor U4626 (N_4626,N_3853,N_3429);
xor U4627 (N_4627,N_3151,N_3141);
nor U4628 (N_4628,N_3524,N_3056);
nand U4629 (N_4629,N_3552,N_3403);
xor U4630 (N_4630,N_3521,N_3993);
or U4631 (N_4631,N_3096,N_3481);
nor U4632 (N_4632,N_3574,N_3520);
xor U4633 (N_4633,N_3529,N_3141);
and U4634 (N_4634,N_3254,N_3695);
xor U4635 (N_4635,N_3205,N_3663);
and U4636 (N_4636,N_3651,N_3391);
and U4637 (N_4637,N_3492,N_3949);
xnor U4638 (N_4638,N_3141,N_3423);
xor U4639 (N_4639,N_3116,N_3772);
and U4640 (N_4640,N_3151,N_3928);
xnor U4641 (N_4641,N_3604,N_3043);
xnor U4642 (N_4642,N_3847,N_3266);
xnor U4643 (N_4643,N_3396,N_3809);
xor U4644 (N_4644,N_3634,N_3221);
or U4645 (N_4645,N_3928,N_3916);
and U4646 (N_4646,N_3740,N_3504);
or U4647 (N_4647,N_3282,N_3744);
xnor U4648 (N_4648,N_3570,N_3644);
nand U4649 (N_4649,N_3285,N_3542);
xnor U4650 (N_4650,N_3804,N_3237);
nand U4651 (N_4651,N_3023,N_3693);
nor U4652 (N_4652,N_3047,N_3137);
nor U4653 (N_4653,N_3596,N_3588);
xnor U4654 (N_4654,N_3117,N_3973);
or U4655 (N_4655,N_3490,N_3150);
and U4656 (N_4656,N_3737,N_3814);
xor U4657 (N_4657,N_3169,N_3734);
nor U4658 (N_4658,N_3451,N_3216);
nand U4659 (N_4659,N_3305,N_3711);
and U4660 (N_4660,N_3069,N_3753);
xor U4661 (N_4661,N_3535,N_3651);
nand U4662 (N_4662,N_3485,N_3796);
nand U4663 (N_4663,N_3828,N_3626);
nand U4664 (N_4664,N_3015,N_3808);
or U4665 (N_4665,N_3459,N_3052);
and U4666 (N_4666,N_3867,N_3584);
nor U4667 (N_4667,N_3706,N_3980);
or U4668 (N_4668,N_3820,N_3347);
nor U4669 (N_4669,N_3923,N_3128);
nor U4670 (N_4670,N_3678,N_3253);
and U4671 (N_4671,N_3092,N_3691);
xor U4672 (N_4672,N_3441,N_3690);
or U4673 (N_4673,N_3419,N_3510);
or U4674 (N_4674,N_3705,N_3668);
or U4675 (N_4675,N_3259,N_3246);
xnor U4676 (N_4676,N_3549,N_3454);
xnor U4677 (N_4677,N_3658,N_3773);
or U4678 (N_4678,N_3513,N_3112);
or U4679 (N_4679,N_3685,N_3051);
xnor U4680 (N_4680,N_3450,N_3702);
nor U4681 (N_4681,N_3506,N_3959);
or U4682 (N_4682,N_3174,N_3904);
or U4683 (N_4683,N_3628,N_3613);
nor U4684 (N_4684,N_3225,N_3570);
xnor U4685 (N_4685,N_3074,N_3064);
or U4686 (N_4686,N_3253,N_3407);
nand U4687 (N_4687,N_3347,N_3264);
nor U4688 (N_4688,N_3808,N_3992);
nand U4689 (N_4689,N_3643,N_3172);
or U4690 (N_4690,N_3852,N_3325);
and U4691 (N_4691,N_3109,N_3914);
and U4692 (N_4692,N_3887,N_3241);
and U4693 (N_4693,N_3124,N_3257);
nand U4694 (N_4694,N_3113,N_3650);
nor U4695 (N_4695,N_3472,N_3481);
or U4696 (N_4696,N_3000,N_3079);
xnor U4697 (N_4697,N_3391,N_3152);
or U4698 (N_4698,N_3090,N_3558);
and U4699 (N_4699,N_3661,N_3277);
and U4700 (N_4700,N_3744,N_3103);
and U4701 (N_4701,N_3066,N_3171);
and U4702 (N_4702,N_3270,N_3835);
nand U4703 (N_4703,N_3268,N_3732);
or U4704 (N_4704,N_3776,N_3594);
nand U4705 (N_4705,N_3787,N_3811);
and U4706 (N_4706,N_3445,N_3591);
nor U4707 (N_4707,N_3009,N_3132);
nor U4708 (N_4708,N_3438,N_3288);
xor U4709 (N_4709,N_3556,N_3696);
nand U4710 (N_4710,N_3373,N_3604);
nor U4711 (N_4711,N_3697,N_3428);
nand U4712 (N_4712,N_3652,N_3746);
and U4713 (N_4713,N_3968,N_3620);
xor U4714 (N_4714,N_3151,N_3153);
nand U4715 (N_4715,N_3661,N_3563);
xnor U4716 (N_4716,N_3298,N_3258);
nor U4717 (N_4717,N_3987,N_3333);
xor U4718 (N_4718,N_3343,N_3696);
nand U4719 (N_4719,N_3704,N_3141);
nand U4720 (N_4720,N_3033,N_3790);
or U4721 (N_4721,N_3548,N_3522);
or U4722 (N_4722,N_3085,N_3198);
nand U4723 (N_4723,N_3238,N_3660);
nand U4724 (N_4724,N_3641,N_3367);
or U4725 (N_4725,N_3286,N_3103);
or U4726 (N_4726,N_3511,N_3240);
nand U4727 (N_4727,N_3406,N_3598);
nor U4728 (N_4728,N_3052,N_3852);
nor U4729 (N_4729,N_3907,N_3920);
nor U4730 (N_4730,N_3649,N_3657);
nand U4731 (N_4731,N_3902,N_3862);
or U4732 (N_4732,N_3116,N_3518);
and U4733 (N_4733,N_3653,N_3618);
and U4734 (N_4734,N_3361,N_3283);
and U4735 (N_4735,N_3563,N_3505);
nand U4736 (N_4736,N_3324,N_3235);
and U4737 (N_4737,N_3622,N_3985);
nand U4738 (N_4738,N_3973,N_3963);
and U4739 (N_4739,N_3523,N_3165);
nand U4740 (N_4740,N_3630,N_3146);
or U4741 (N_4741,N_3638,N_3256);
nor U4742 (N_4742,N_3438,N_3730);
xnor U4743 (N_4743,N_3309,N_3031);
and U4744 (N_4744,N_3948,N_3359);
and U4745 (N_4745,N_3498,N_3368);
or U4746 (N_4746,N_3732,N_3041);
or U4747 (N_4747,N_3245,N_3056);
nand U4748 (N_4748,N_3413,N_3180);
and U4749 (N_4749,N_3380,N_3287);
nand U4750 (N_4750,N_3326,N_3493);
and U4751 (N_4751,N_3662,N_3446);
nor U4752 (N_4752,N_3159,N_3748);
and U4753 (N_4753,N_3373,N_3121);
and U4754 (N_4754,N_3968,N_3248);
xor U4755 (N_4755,N_3025,N_3882);
and U4756 (N_4756,N_3167,N_3623);
and U4757 (N_4757,N_3475,N_3023);
and U4758 (N_4758,N_3799,N_3810);
nor U4759 (N_4759,N_3074,N_3609);
and U4760 (N_4760,N_3411,N_3133);
nor U4761 (N_4761,N_3120,N_3269);
nor U4762 (N_4762,N_3643,N_3763);
xnor U4763 (N_4763,N_3594,N_3921);
or U4764 (N_4764,N_3224,N_3397);
and U4765 (N_4765,N_3174,N_3557);
and U4766 (N_4766,N_3811,N_3082);
nand U4767 (N_4767,N_3102,N_3518);
and U4768 (N_4768,N_3323,N_3181);
and U4769 (N_4769,N_3328,N_3014);
nor U4770 (N_4770,N_3227,N_3136);
xor U4771 (N_4771,N_3822,N_3405);
and U4772 (N_4772,N_3341,N_3024);
and U4773 (N_4773,N_3274,N_3102);
and U4774 (N_4774,N_3977,N_3786);
and U4775 (N_4775,N_3042,N_3029);
and U4776 (N_4776,N_3106,N_3696);
xnor U4777 (N_4777,N_3879,N_3296);
or U4778 (N_4778,N_3762,N_3969);
nor U4779 (N_4779,N_3535,N_3588);
and U4780 (N_4780,N_3881,N_3948);
nor U4781 (N_4781,N_3466,N_3948);
nor U4782 (N_4782,N_3615,N_3801);
xnor U4783 (N_4783,N_3783,N_3034);
or U4784 (N_4784,N_3968,N_3726);
nand U4785 (N_4785,N_3182,N_3118);
and U4786 (N_4786,N_3584,N_3892);
nand U4787 (N_4787,N_3557,N_3408);
or U4788 (N_4788,N_3112,N_3268);
xor U4789 (N_4789,N_3329,N_3250);
or U4790 (N_4790,N_3177,N_3856);
nor U4791 (N_4791,N_3959,N_3317);
nand U4792 (N_4792,N_3864,N_3006);
or U4793 (N_4793,N_3761,N_3693);
nor U4794 (N_4794,N_3561,N_3109);
and U4795 (N_4795,N_3077,N_3473);
nor U4796 (N_4796,N_3245,N_3725);
or U4797 (N_4797,N_3670,N_3389);
and U4798 (N_4798,N_3554,N_3064);
xor U4799 (N_4799,N_3491,N_3029);
xor U4800 (N_4800,N_3687,N_3345);
nor U4801 (N_4801,N_3348,N_3281);
xnor U4802 (N_4802,N_3163,N_3344);
nand U4803 (N_4803,N_3277,N_3871);
xnor U4804 (N_4804,N_3156,N_3139);
or U4805 (N_4805,N_3309,N_3808);
nand U4806 (N_4806,N_3983,N_3876);
nor U4807 (N_4807,N_3097,N_3255);
and U4808 (N_4808,N_3111,N_3681);
xor U4809 (N_4809,N_3763,N_3389);
nor U4810 (N_4810,N_3333,N_3057);
or U4811 (N_4811,N_3476,N_3870);
or U4812 (N_4812,N_3504,N_3515);
and U4813 (N_4813,N_3027,N_3740);
nand U4814 (N_4814,N_3770,N_3624);
or U4815 (N_4815,N_3584,N_3192);
and U4816 (N_4816,N_3060,N_3750);
xnor U4817 (N_4817,N_3982,N_3615);
nor U4818 (N_4818,N_3658,N_3331);
xor U4819 (N_4819,N_3191,N_3711);
nand U4820 (N_4820,N_3893,N_3248);
or U4821 (N_4821,N_3312,N_3212);
nand U4822 (N_4822,N_3348,N_3245);
or U4823 (N_4823,N_3091,N_3678);
and U4824 (N_4824,N_3420,N_3540);
xnor U4825 (N_4825,N_3244,N_3334);
or U4826 (N_4826,N_3686,N_3472);
and U4827 (N_4827,N_3409,N_3415);
nor U4828 (N_4828,N_3719,N_3412);
xnor U4829 (N_4829,N_3828,N_3125);
or U4830 (N_4830,N_3970,N_3210);
or U4831 (N_4831,N_3851,N_3896);
nor U4832 (N_4832,N_3440,N_3952);
nor U4833 (N_4833,N_3876,N_3759);
nor U4834 (N_4834,N_3384,N_3534);
and U4835 (N_4835,N_3569,N_3025);
nor U4836 (N_4836,N_3591,N_3237);
xnor U4837 (N_4837,N_3185,N_3431);
and U4838 (N_4838,N_3608,N_3717);
nor U4839 (N_4839,N_3762,N_3019);
and U4840 (N_4840,N_3280,N_3119);
nand U4841 (N_4841,N_3559,N_3891);
nor U4842 (N_4842,N_3771,N_3766);
xnor U4843 (N_4843,N_3825,N_3038);
nor U4844 (N_4844,N_3079,N_3950);
or U4845 (N_4845,N_3459,N_3448);
and U4846 (N_4846,N_3180,N_3785);
xor U4847 (N_4847,N_3052,N_3373);
nand U4848 (N_4848,N_3087,N_3415);
or U4849 (N_4849,N_3189,N_3759);
or U4850 (N_4850,N_3761,N_3890);
or U4851 (N_4851,N_3126,N_3564);
and U4852 (N_4852,N_3011,N_3477);
nand U4853 (N_4853,N_3560,N_3129);
nor U4854 (N_4854,N_3732,N_3696);
or U4855 (N_4855,N_3209,N_3579);
and U4856 (N_4856,N_3171,N_3850);
xnor U4857 (N_4857,N_3529,N_3264);
or U4858 (N_4858,N_3187,N_3433);
xnor U4859 (N_4859,N_3080,N_3914);
and U4860 (N_4860,N_3036,N_3003);
xor U4861 (N_4861,N_3170,N_3003);
and U4862 (N_4862,N_3156,N_3881);
or U4863 (N_4863,N_3012,N_3374);
or U4864 (N_4864,N_3624,N_3836);
and U4865 (N_4865,N_3559,N_3927);
or U4866 (N_4866,N_3664,N_3991);
xor U4867 (N_4867,N_3025,N_3126);
and U4868 (N_4868,N_3022,N_3227);
or U4869 (N_4869,N_3873,N_3189);
or U4870 (N_4870,N_3551,N_3492);
and U4871 (N_4871,N_3264,N_3708);
nor U4872 (N_4872,N_3044,N_3630);
nand U4873 (N_4873,N_3283,N_3428);
or U4874 (N_4874,N_3920,N_3445);
nand U4875 (N_4875,N_3821,N_3129);
nor U4876 (N_4876,N_3558,N_3996);
nor U4877 (N_4877,N_3354,N_3014);
or U4878 (N_4878,N_3704,N_3606);
nand U4879 (N_4879,N_3640,N_3779);
nor U4880 (N_4880,N_3605,N_3824);
or U4881 (N_4881,N_3746,N_3138);
and U4882 (N_4882,N_3987,N_3269);
nand U4883 (N_4883,N_3757,N_3500);
or U4884 (N_4884,N_3172,N_3341);
nand U4885 (N_4885,N_3850,N_3490);
xnor U4886 (N_4886,N_3101,N_3536);
nand U4887 (N_4887,N_3684,N_3210);
or U4888 (N_4888,N_3857,N_3084);
xnor U4889 (N_4889,N_3975,N_3367);
and U4890 (N_4890,N_3440,N_3349);
nand U4891 (N_4891,N_3475,N_3829);
xor U4892 (N_4892,N_3400,N_3707);
and U4893 (N_4893,N_3035,N_3750);
nor U4894 (N_4894,N_3423,N_3347);
xor U4895 (N_4895,N_3449,N_3577);
xnor U4896 (N_4896,N_3118,N_3486);
nor U4897 (N_4897,N_3685,N_3983);
xnor U4898 (N_4898,N_3589,N_3708);
xnor U4899 (N_4899,N_3899,N_3782);
or U4900 (N_4900,N_3639,N_3558);
nor U4901 (N_4901,N_3546,N_3233);
nor U4902 (N_4902,N_3447,N_3361);
and U4903 (N_4903,N_3248,N_3554);
or U4904 (N_4904,N_3374,N_3720);
and U4905 (N_4905,N_3371,N_3948);
xnor U4906 (N_4906,N_3598,N_3195);
and U4907 (N_4907,N_3381,N_3062);
or U4908 (N_4908,N_3028,N_3667);
nand U4909 (N_4909,N_3500,N_3666);
and U4910 (N_4910,N_3369,N_3326);
and U4911 (N_4911,N_3896,N_3377);
and U4912 (N_4912,N_3273,N_3084);
and U4913 (N_4913,N_3749,N_3918);
nand U4914 (N_4914,N_3709,N_3973);
and U4915 (N_4915,N_3258,N_3389);
and U4916 (N_4916,N_3267,N_3401);
xnor U4917 (N_4917,N_3963,N_3353);
and U4918 (N_4918,N_3593,N_3489);
and U4919 (N_4919,N_3111,N_3370);
xnor U4920 (N_4920,N_3104,N_3356);
nand U4921 (N_4921,N_3664,N_3149);
xnor U4922 (N_4922,N_3168,N_3373);
or U4923 (N_4923,N_3911,N_3181);
or U4924 (N_4924,N_3015,N_3001);
nand U4925 (N_4925,N_3949,N_3179);
and U4926 (N_4926,N_3958,N_3943);
nand U4927 (N_4927,N_3101,N_3064);
and U4928 (N_4928,N_3261,N_3584);
or U4929 (N_4929,N_3429,N_3870);
xor U4930 (N_4930,N_3969,N_3467);
nand U4931 (N_4931,N_3884,N_3780);
nor U4932 (N_4932,N_3360,N_3012);
xnor U4933 (N_4933,N_3762,N_3715);
or U4934 (N_4934,N_3733,N_3581);
nand U4935 (N_4935,N_3559,N_3897);
xnor U4936 (N_4936,N_3837,N_3929);
nor U4937 (N_4937,N_3849,N_3979);
or U4938 (N_4938,N_3995,N_3592);
nand U4939 (N_4939,N_3904,N_3513);
and U4940 (N_4940,N_3000,N_3108);
or U4941 (N_4941,N_3768,N_3094);
and U4942 (N_4942,N_3780,N_3910);
and U4943 (N_4943,N_3992,N_3701);
nor U4944 (N_4944,N_3466,N_3997);
nand U4945 (N_4945,N_3402,N_3877);
or U4946 (N_4946,N_3125,N_3777);
and U4947 (N_4947,N_3049,N_3866);
or U4948 (N_4948,N_3205,N_3947);
and U4949 (N_4949,N_3822,N_3490);
nor U4950 (N_4950,N_3933,N_3795);
and U4951 (N_4951,N_3812,N_3789);
or U4952 (N_4952,N_3736,N_3436);
nand U4953 (N_4953,N_3909,N_3824);
nor U4954 (N_4954,N_3093,N_3355);
nand U4955 (N_4955,N_3602,N_3849);
nor U4956 (N_4956,N_3120,N_3252);
xor U4957 (N_4957,N_3479,N_3033);
and U4958 (N_4958,N_3179,N_3902);
and U4959 (N_4959,N_3088,N_3033);
and U4960 (N_4960,N_3890,N_3936);
nor U4961 (N_4961,N_3975,N_3229);
nand U4962 (N_4962,N_3128,N_3807);
and U4963 (N_4963,N_3665,N_3980);
nand U4964 (N_4964,N_3906,N_3367);
or U4965 (N_4965,N_3476,N_3497);
xnor U4966 (N_4966,N_3038,N_3899);
nand U4967 (N_4967,N_3577,N_3470);
nand U4968 (N_4968,N_3513,N_3564);
nor U4969 (N_4969,N_3692,N_3037);
or U4970 (N_4970,N_3769,N_3554);
xnor U4971 (N_4971,N_3581,N_3403);
xor U4972 (N_4972,N_3925,N_3845);
xnor U4973 (N_4973,N_3126,N_3477);
xor U4974 (N_4974,N_3794,N_3722);
nand U4975 (N_4975,N_3206,N_3607);
and U4976 (N_4976,N_3532,N_3221);
nor U4977 (N_4977,N_3682,N_3352);
xor U4978 (N_4978,N_3153,N_3885);
and U4979 (N_4979,N_3081,N_3858);
nor U4980 (N_4980,N_3742,N_3443);
xnor U4981 (N_4981,N_3583,N_3194);
xor U4982 (N_4982,N_3721,N_3731);
nor U4983 (N_4983,N_3536,N_3179);
xnor U4984 (N_4984,N_3810,N_3803);
nor U4985 (N_4985,N_3727,N_3865);
and U4986 (N_4986,N_3889,N_3305);
and U4987 (N_4987,N_3626,N_3405);
or U4988 (N_4988,N_3493,N_3171);
or U4989 (N_4989,N_3863,N_3832);
nand U4990 (N_4990,N_3951,N_3948);
or U4991 (N_4991,N_3956,N_3844);
and U4992 (N_4992,N_3061,N_3877);
xnor U4993 (N_4993,N_3387,N_3888);
nor U4994 (N_4994,N_3266,N_3325);
or U4995 (N_4995,N_3187,N_3559);
nor U4996 (N_4996,N_3748,N_3590);
xnor U4997 (N_4997,N_3404,N_3636);
nand U4998 (N_4998,N_3435,N_3406);
nand U4999 (N_4999,N_3153,N_3611);
nand U5000 (N_5000,N_4784,N_4845);
and U5001 (N_5001,N_4677,N_4967);
nand U5002 (N_5002,N_4119,N_4616);
xnor U5003 (N_5003,N_4620,N_4462);
nand U5004 (N_5004,N_4068,N_4155);
nand U5005 (N_5005,N_4292,N_4198);
xor U5006 (N_5006,N_4955,N_4093);
nand U5007 (N_5007,N_4558,N_4126);
nor U5008 (N_5008,N_4702,N_4442);
xor U5009 (N_5009,N_4939,N_4515);
xor U5010 (N_5010,N_4688,N_4820);
or U5011 (N_5011,N_4831,N_4072);
nor U5012 (N_5012,N_4221,N_4559);
nor U5013 (N_5013,N_4195,N_4511);
xnor U5014 (N_5014,N_4672,N_4798);
and U5015 (N_5015,N_4656,N_4226);
or U5016 (N_5016,N_4641,N_4086);
or U5017 (N_5017,N_4942,N_4239);
xnor U5018 (N_5018,N_4051,N_4583);
xnor U5019 (N_5019,N_4213,N_4461);
nor U5020 (N_5020,N_4017,N_4897);
or U5021 (N_5021,N_4855,N_4290);
xor U5022 (N_5022,N_4116,N_4458);
and U5023 (N_5023,N_4993,N_4351);
nand U5024 (N_5024,N_4959,N_4542);
and U5025 (N_5025,N_4539,N_4666);
xnor U5026 (N_5026,N_4143,N_4994);
or U5027 (N_5027,N_4886,N_4124);
and U5028 (N_5028,N_4541,N_4575);
xnor U5029 (N_5029,N_4907,N_4841);
or U5030 (N_5030,N_4060,N_4451);
and U5031 (N_5031,N_4110,N_4170);
and U5032 (N_5032,N_4070,N_4052);
or U5033 (N_5033,N_4495,N_4755);
nor U5034 (N_5034,N_4840,N_4503);
and U5035 (N_5035,N_4890,N_4626);
and U5036 (N_5036,N_4349,N_4333);
xor U5037 (N_5037,N_4745,N_4824);
xor U5038 (N_5038,N_4567,N_4737);
xnor U5039 (N_5039,N_4122,N_4336);
nand U5040 (N_5040,N_4781,N_4319);
nand U5041 (N_5041,N_4083,N_4001);
and U5042 (N_5042,N_4906,N_4700);
nor U5043 (N_5043,N_4506,N_4173);
and U5044 (N_5044,N_4657,N_4299);
nand U5045 (N_5045,N_4443,N_4302);
or U5046 (N_5046,N_4652,N_4777);
or U5047 (N_5047,N_4976,N_4312);
nand U5048 (N_5048,N_4560,N_4115);
and U5049 (N_5049,N_4960,N_4147);
and U5050 (N_5050,N_4929,N_4637);
nor U5051 (N_5051,N_4731,N_4538);
or U5052 (N_5052,N_4785,N_4827);
nor U5053 (N_5053,N_4973,N_4923);
nand U5054 (N_5054,N_4026,N_4609);
nand U5055 (N_5055,N_4732,N_4882);
nand U5056 (N_5056,N_4535,N_4928);
and U5057 (N_5057,N_4747,N_4184);
and U5058 (N_5058,N_4012,N_4801);
or U5059 (N_5059,N_4870,N_4985);
xor U5060 (N_5060,N_4377,N_4573);
nand U5061 (N_5061,N_4338,N_4386);
or U5062 (N_5062,N_4169,N_4261);
xnor U5063 (N_5063,N_4197,N_4715);
or U5064 (N_5064,N_4596,N_4681);
xor U5065 (N_5065,N_4662,N_4859);
or U5066 (N_5066,N_4809,N_4724);
nor U5067 (N_5067,N_4521,N_4281);
or U5068 (N_5068,N_4876,N_4120);
nand U5069 (N_5069,N_4076,N_4146);
or U5070 (N_5070,N_4056,N_4621);
and U5071 (N_5071,N_4565,N_4502);
xor U5072 (N_5072,N_4211,N_4977);
nor U5073 (N_5073,N_4329,N_4933);
and U5074 (N_5074,N_4316,N_4220);
nor U5075 (N_5075,N_4986,N_4125);
xor U5076 (N_5076,N_4199,N_4912);
xnor U5077 (N_5077,N_4729,N_4137);
nor U5078 (N_5078,N_4383,N_4874);
xor U5079 (N_5079,N_4382,N_4414);
nor U5080 (N_5080,N_4748,N_4074);
and U5081 (N_5081,N_4758,N_4266);
nand U5082 (N_5082,N_4008,N_4712);
or U5083 (N_5083,N_4649,N_4309);
nor U5084 (N_5084,N_4645,N_4523);
nand U5085 (N_5085,N_4154,N_4482);
nor U5086 (N_5086,N_4634,N_4029);
or U5087 (N_5087,N_4839,N_4471);
nor U5088 (N_5088,N_4133,N_4448);
nor U5089 (N_5089,N_4038,N_4200);
xnor U5090 (N_5090,N_4454,N_4420);
or U5091 (N_5091,N_4332,N_4011);
xor U5092 (N_5092,N_4648,N_4061);
nor U5093 (N_5093,N_4048,N_4815);
nor U5094 (N_5094,N_4172,N_4880);
xnor U5095 (N_5095,N_4171,N_4524);
nand U5096 (N_5096,N_4167,N_4370);
xnor U5097 (N_5097,N_4468,N_4948);
and U5098 (N_5098,N_4527,N_4698);
nand U5099 (N_5099,N_4162,N_4690);
nand U5100 (N_5100,N_4837,N_4530);
nor U5101 (N_5101,N_4188,N_4556);
nand U5102 (N_5102,N_4186,N_4362);
or U5103 (N_5103,N_4087,N_4988);
nor U5104 (N_5104,N_4278,N_4099);
nand U5105 (N_5105,N_4297,N_4310);
xor U5106 (N_5106,N_4821,N_4224);
or U5107 (N_5107,N_4668,N_4078);
nand U5108 (N_5108,N_4926,N_4418);
and U5109 (N_5109,N_4619,N_4847);
nor U5110 (N_5110,N_4036,N_4954);
nor U5111 (N_5111,N_4103,N_4006);
and U5112 (N_5112,N_4699,N_4135);
or U5113 (N_5113,N_4991,N_4021);
or U5114 (N_5114,N_4400,N_4091);
and U5115 (N_5115,N_4630,N_4434);
or U5116 (N_5116,N_4673,N_4982);
and U5117 (N_5117,N_4315,N_4084);
nand U5118 (N_5118,N_4148,N_4919);
or U5119 (N_5119,N_4459,N_4854);
xor U5120 (N_5120,N_4202,N_4944);
and U5121 (N_5121,N_4417,N_4764);
nor U5122 (N_5122,N_4812,N_4075);
nor U5123 (N_5123,N_4819,N_4168);
or U5124 (N_5124,N_4520,N_4872);
xor U5125 (N_5125,N_4331,N_4144);
and U5126 (N_5126,N_4768,N_4488);
or U5127 (N_5127,N_4212,N_4437);
and U5128 (N_5128,N_4532,N_4646);
xor U5129 (N_5129,N_4958,N_4256);
nand U5130 (N_5130,N_4943,N_4592);
xor U5131 (N_5131,N_4574,N_4658);
nand U5132 (N_5132,N_4746,N_4406);
nand U5133 (N_5133,N_4893,N_4483);
nand U5134 (N_5134,N_4273,N_4194);
nor U5135 (N_5135,N_4725,N_4177);
or U5136 (N_5136,N_4306,N_4741);
nor U5137 (N_5137,N_4247,N_4989);
or U5138 (N_5138,N_4275,N_4693);
nand U5139 (N_5139,N_4572,N_4248);
and U5140 (N_5140,N_4174,N_4582);
xnor U5141 (N_5141,N_4618,N_4342);
nor U5142 (N_5142,N_4891,N_4394);
or U5143 (N_5143,N_4723,N_4262);
nand U5144 (N_5144,N_4384,N_4296);
nand U5145 (N_5145,N_4347,N_4799);
and U5146 (N_5146,N_4487,N_4667);
xor U5147 (N_5147,N_4114,N_4294);
nor U5148 (N_5148,N_4424,N_4516);
or U5149 (N_5149,N_4337,N_4661);
nor U5150 (N_5150,N_4217,N_4271);
and U5151 (N_5151,N_4356,N_4354);
nor U5152 (N_5152,N_4480,N_4403);
and U5153 (N_5153,N_4361,N_4359);
nor U5154 (N_5154,N_4773,N_4762);
nand U5155 (N_5155,N_4033,N_4323);
nand U5156 (N_5156,N_4774,N_4178);
or U5157 (N_5157,N_4749,N_4372);
nand U5158 (N_5158,N_4863,N_4376);
or U5159 (N_5159,N_4025,N_4612);
and U5160 (N_5160,N_4833,N_4796);
or U5161 (N_5161,N_4655,N_4554);
and U5162 (N_5162,N_4816,N_4380);
xor U5163 (N_5163,N_4234,N_4166);
and U5164 (N_5164,N_4628,N_4090);
xnor U5165 (N_5165,N_4650,N_4623);
nand U5166 (N_5166,N_4015,N_4852);
or U5167 (N_5167,N_4259,N_4439);
and U5168 (N_5168,N_4606,N_4498);
and U5169 (N_5169,N_4335,N_4563);
nor U5170 (N_5170,N_4676,N_4340);
nor U5171 (N_5171,N_4037,N_4407);
nand U5172 (N_5172,N_4549,N_4627);
nor U5173 (N_5173,N_4836,N_4811);
nor U5174 (N_5174,N_4536,N_4499);
xnor U5175 (N_5175,N_4846,N_4111);
xor U5176 (N_5176,N_4694,N_4586);
and U5177 (N_5177,N_4832,N_4871);
nand U5178 (N_5178,N_4569,N_4776);
or U5179 (N_5179,N_4921,N_4447);
xnor U5180 (N_5180,N_4924,N_4002);
nand U5181 (N_5181,N_4020,N_4877);
nor U5182 (N_5182,N_4121,N_4899);
xor U5183 (N_5183,N_4970,N_4622);
and U5184 (N_5184,N_4587,N_4671);
nor U5185 (N_5185,N_4601,N_4106);
and U5186 (N_5186,N_4455,N_4940);
nor U5187 (N_5187,N_4716,N_4851);
and U5188 (N_5188,N_4714,N_4428);
and U5189 (N_5189,N_4004,N_4644);
xnor U5190 (N_5190,N_4624,N_4964);
nand U5191 (N_5191,N_4486,N_4680);
xor U5192 (N_5192,N_4632,N_4467);
or U5193 (N_5193,N_4794,N_4157);
xor U5194 (N_5194,N_4440,N_4100);
xor U5195 (N_5195,N_4733,N_4274);
xor U5196 (N_5196,N_4128,N_4325);
nand U5197 (N_5197,N_4810,N_4346);
nor U5198 (N_5198,N_4317,N_4311);
nand U5199 (N_5199,N_4485,N_4260);
nand U5200 (N_5200,N_4436,N_4223);
and U5201 (N_5201,N_4508,N_4584);
or U5202 (N_5202,N_4856,N_4295);
or U5203 (N_5203,N_4105,N_4463);
and U5204 (N_5204,N_4429,N_4005);
nor U5205 (N_5205,N_4949,N_4608);
xor U5206 (N_5206,N_4279,N_4250);
and U5207 (N_5207,N_4088,N_4931);
nand U5208 (N_5208,N_4210,N_4547);
xnor U5209 (N_5209,N_4718,N_4687);
or U5210 (N_5210,N_4510,N_4113);
or U5211 (N_5211,N_4981,N_4425);
and U5212 (N_5212,N_4790,N_4187);
or U5213 (N_5213,N_4564,N_4579);
or U5214 (N_5214,N_4862,N_4719);
nor U5215 (N_5215,N_4829,N_4185);
nand U5216 (N_5216,N_4997,N_4441);
nor U5217 (N_5217,N_4932,N_4334);
xnor U5218 (N_5218,N_4016,N_4358);
and U5219 (N_5219,N_4066,N_4770);
nor U5220 (N_5220,N_4058,N_4481);
and U5221 (N_5221,N_4270,N_4867);
xnor U5222 (N_5222,N_4085,N_4158);
and U5223 (N_5223,N_4800,N_4956);
nand U5224 (N_5224,N_4385,N_4357);
nand U5225 (N_5225,N_4904,N_4965);
nor U5226 (N_5226,N_4971,N_4484);
nor U5227 (N_5227,N_4720,N_4922);
nand U5228 (N_5228,N_4686,N_4684);
xor U5229 (N_5229,N_4426,N_4995);
nand U5230 (N_5230,N_4389,N_4938);
or U5231 (N_5231,N_4138,N_4947);
and U5232 (N_5232,N_4098,N_4313);
xor U5233 (N_5233,N_4452,N_4046);
xnor U5234 (N_5234,N_4284,N_4276);
nor U5235 (N_5235,N_4685,N_4464);
nor U5236 (N_5236,N_4553,N_4397);
and U5237 (N_5237,N_4507,N_4878);
xnor U5238 (N_5238,N_4307,N_4934);
xor U5239 (N_5239,N_4175,N_4813);
xor U5240 (N_5240,N_4423,N_4303);
or U5241 (N_5241,N_4513,N_4225);
and U5242 (N_5242,N_4314,N_4818);
xor U5243 (N_5243,N_4682,N_4610);
nor U5244 (N_5244,N_4388,N_4551);
and U5245 (N_5245,N_4022,N_4301);
xnor U5246 (N_5246,N_4850,N_4433);
nand U5247 (N_5247,N_4230,N_4916);
xnor U5248 (N_5248,N_4229,N_4902);
nand U5249 (N_5249,N_4208,N_4219);
and U5250 (N_5250,N_4660,N_4131);
xnor U5251 (N_5251,N_4324,N_4364);
nor U5252 (N_5252,N_4793,N_4501);
nor U5253 (N_5253,N_4097,N_4438);
nand U5254 (N_5254,N_4884,N_4915);
nand U5255 (N_5255,N_4979,N_4760);
or U5256 (N_5256,N_4548,N_4101);
xnor U5257 (N_5257,N_4288,N_4010);
nand U5258 (N_5258,N_4864,N_4478);
nor U5259 (N_5259,N_4024,N_4589);
nand U5260 (N_5260,N_4898,N_4014);
or U5261 (N_5261,N_4722,N_4743);
and U5262 (N_5262,N_4390,N_4215);
nor U5263 (N_5263,N_4865,N_4123);
nand U5264 (N_5264,N_4003,N_4925);
or U5265 (N_5265,N_4348,N_4889);
nor U5266 (N_5266,N_4639,N_4398);
nand U5267 (N_5267,N_4327,N_4590);
xnor U5268 (N_5268,N_4164,N_4431);
nor U5269 (N_5269,N_4607,N_4849);
and U5270 (N_5270,N_4065,N_4079);
nand U5271 (N_5271,N_4231,N_4092);
or U5272 (N_5272,N_4300,N_4251);
nor U5273 (N_5273,N_4952,N_4265);
nor U5274 (N_5274,N_4858,N_4792);
or U5275 (N_5275,N_4375,N_4756);
nor U5276 (N_5276,N_4726,N_4242);
xor U5277 (N_5277,N_4528,N_4405);
or U5278 (N_5278,N_4509,N_4069);
nor U5279 (N_5279,N_4214,N_4449);
xor U5280 (N_5280,N_4780,N_4435);
or U5281 (N_5281,N_4363,N_4419);
nor U5282 (N_5282,N_4089,N_4585);
xnor U5283 (N_5283,N_4761,N_4857);
or U5284 (N_5284,N_4096,N_4318);
nand U5285 (N_5285,N_4228,N_4129);
xor U5286 (N_5286,N_4765,N_4491);
and U5287 (N_5287,N_4190,N_4692);
or U5288 (N_5288,N_4603,N_4055);
or U5289 (N_5289,N_4489,N_4593);
and U5290 (N_5290,N_4401,N_4514);
nor U5291 (N_5291,N_4206,N_4717);
xnor U5292 (N_5292,N_4980,N_4803);
xnor U5293 (N_5293,N_4411,N_4936);
nor U5294 (N_5294,N_4704,N_4064);
and U5295 (N_5295,N_4267,N_4320);
nand U5296 (N_5296,N_4328,N_4496);
nor U5297 (N_5297,N_4151,N_4413);
and U5298 (N_5298,N_4191,N_4469);
or U5299 (N_5299,N_4580,N_4544);
nor U5300 (N_5300,N_4935,N_4653);
or U5301 (N_5301,N_4689,N_4475);
nand U5302 (N_5302,N_4222,N_4396);
and U5303 (N_5303,N_4152,N_4629);
xnor U5304 (N_5304,N_4028,N_4599);
nand U5305 (N_5305,N_4734,N_4561);
nand U5306 (N_5306,N_4611,N_4600);
nor U5307 (N_5307,N_4412,N_4557);
xor U5308 (N_5308,N_4473,N_4830);
nand U5309 (N_5309,N_4393,N_4264);
xnor U5310 (N_5310,N_4032,N_4246);
nor U5311 (N_5311,N_4059,N_4373);
nor U5312 (N_5312,N_4102,N_4588);
and U5313 (N_5313,N_4041,N_4255);
nor U5314 (N_5314,N_4848,N_4945);
nand U5315 (N_5315,N_4139,N_4866);
nand U5316 (N_5316,N_4404,N_4263);
and U5317 (N_5317,N_4027,N_4752);
xnor U5318 (N_5318,N_4444,N_4035);
nor U5319 (N_5319,N_4067,N_4739);
nor U5320 (N_5320,N_4062,N_4695);
xnor U5321 (N_5321,N_4636,N_4176);
or U5322 (N_5322,N_4504,N_4132);
or U5323 (N_5323,N_4237,N_4408);
xnor U5324 (N_5324,N_4531,N_4806);
and U5325 (N_5325,N_4550,N_4127);
xnor U5326 (N_5326,N_4961,N_4844);
nand U5327 (N_5327,N_4422,N_4713);
nand U5328 (N_5328,N_4141,N_4345);
and U5329 (N_5329,N_4142,N_4512);
or U5330 (N_5330,N_4783,N_4570);
xor U5331 (N_5331,N_4631,N_4642);
or U5332 (N_5332,N_4159,N_4181);
and U5333 (N_5333,N_4838,N_4571);
nor U5334 (N_5334,N_4913,N_4814);
and U5335 (N_5335,N_4771,N_4000);
xor U5336 (N_5336,N_4978,N_4663);
nand U5337 (N_5337,N_4670,N_4227);
nor U5338 (N_5338,N_4081,N_4283);
nor U5339 (N_5339,N_4826,N_4387);
or U5340 (N_5340,N_4243,N_4875);
and U5341 (N_5341,N_4497,N_4740);
nand U5342 (N_5342,N_4769,N_4465);
or U5343 (N_5343,N_4707,N_4145);
nand U5344 (N_5344,N_4754,N_4709);
or U5345 (N_5345,N_4355,N_4410);
nor U5346 (N_5346,N_4823,N_4804);
nand U5347 (N_5347,N_4339,N_4697);
nor U5348 (N_5348,N_4703,N_4957);
nor U5349 (N_5349,N_4946,N_4282);
xnor U5350 (N_5350,N_4492,N_4134);
or U5351 (N_5351,N_4277,N_4753);
nor U5352 (N_5352,N_4540,N_4216);
nor U5353 (N_5353,N_4604,N_4537);
nor U5354 (N_5354,N_4992,N_4107);
and U5355 (N_5355,N_4330,N_4232);
and U5356 (N_5356,N_4039,N_4007);
and U5357 (N_5357,N_4533,N_4254);
or U5358 (N_5358,N_4990,N_4920);
nand U5359 (N_5359,N_4892,N_4050);
and U5360 (N_5360,N_4043,N_4552);
or U5361 (N_5361,N_4885,N_4253);
or U5362 (N_5362,N_4708,N_4545);
xnor U5363 (N_5363,N_4817,N_4183);
or U5364 (N_5364,N_4706,N_4835);
and U5365 (N_5365,N_4470,N_4625);
or U5366 (N_5366,N_4711,N_4918);
xnor U5367 (N_5367,N_4368,N_4117);
or U5368 (N_5368,N_4034,N_4257);
and U5369 (N_5369,N_4189,N_4427);
xor U5370 (N_5370,N_4019,N_4280);
and U5371 (N_5371,N_4905,N_4675);
xor U5372 (N_5372,N_4238,N_4853);
nand U5373 (N_5373,N_4365,N_4192);
nand U5374 (N_5374,N_4472,N_4252);
nor U5375 (N_5375,N_4900,N_4615);
xor U5376 (N_5376,N_4937,N_4416);
nor U5377 (N_5377,N_4710,N_4240);
or U5378 (N_5378,N_4291,N_4054);
and U5379 (N_5379,N_4391,N_4647);
nor U5380 (N_5380,N_4374,N_4903);
xnor U5381 (N_5381,N_4179,N_4304);
xor U5382 (N_5382,N_4529,N_4289);
nand U5383 (N_5383,N_4379,N_4298);
or U5384 (N_5384,N_4972,N_4366);
and U5385 (N_5385,N_4788,N_4999);
or U5386 (N_5386,N_4352,N_4402);
nor U5387 (N_5387,N_4742,N_4236);
xor U5388 (N_5388,N_4802,N_4705);
nor U5389 (N_5389,N_4235,N_4165);
nor U5390 (N_5390,N_4479,N_4969);
and U5391 (N_5391,N_4910,N_4805);
nand U5392 (N_5392,N_4578,N_4888);
and U5393 (N_5393,N_4577,N_4868);
nor U5394 (N_5394,N_4305,N_4456);
or U5395 (N_5395,N_4104,N_4901);
and U5396 (N_5396,N_4828,N_4778);
or U5397 (N_5397,N_4927,N_4595);
and U5398 (N_5398,N_4998,N_4180);
nor U5399 (N_5399,N_4911,N_4322);
or U5400 (N_5400,N_4450,N_4679);
nor U5401 (N_5401,N_4633,N_4562);
nor U5402 (N_5402,N_4951,N_4082);
nor U5403 (N_5403,N_4201,N_4343);
and U5404 (N_5404,N_4047,N_4094);
nor U5405 (N_5405,N_4518,N_4205);
or U5406 (N_5406,N_4797,N_4669);
nor U5407 (N_5407,N_4160,N_4080);
nand U5408 (N_5408,N_4807,N_4635);
nand U5409 (N_5409,N_4842,N_4156);
nand U5410 (N_5410,N_4987,N_4466);
nand U5411 (N_5411,N_4258,N_4738);
and U5412 (N_5412,N_4789,N_4775);
xnor U5413 (N_5413,N_4244,N_4204);
nor U5414 (N_5414,N_4203,N_4245);
nor U5415 (N_5415,N_4353,N_4963);
nor U5416 (N_5416,N_4526,N_4566);
nor U5417 (N_5417,N_4009,N_4453);
nor U5418 (N_5418,N_4367,N_4654);
or U5419 (N_5419,N_4730,N_4045);
or U5420 (N_5420,N_4728,N_4822);
nor U5421 (N_5421,N_4053,N_4108);
or U5422 (N_5422,N_4869,N_4984);
nand U5423 (N_5423,N_4207,N_4895);
xor U5424 (N_5424,N_4941,N_4744);
xor U5425 (N_5425,N_4613,N_4140);
xor U5426 (N_5426,N_4446,N_4750);
nand U5427 (N_5427,N_4568,N_4136);
nor U5428 (N_5428,N_4791,N_4782);
or U5429 (N_5429,N_4130,N_4371);
or U5430 (N_5430,N_4721,N_4505);
and U5431 (N_5431,N_4163,N_4182);
nor U5432 (N_5432,N_4736,N_4534);
xor U5433 (N_5433,N_4474,N_4786);
xor U5434 (N_5434,N_4759,N_4643);
nand U5435 (N_5435,N_4543,N_4665);
or U5436 (N_5436,N_4308,N_4879);
nand U5437 (N_5437,N_4696,N_4883);
nor U5438 (N_5438,N_4861,N_4241);
xnor U5439 (N_5439,N_4896,N_4153);
xnor U5440 (N_5440,N_4095,N_4691);
xnor U5441 (N_5441,N_4968,N_4350);
and U5442 (N_5442,N_4909,N_4285);
nor U5443 (N_5443,N_4873,N_4779);
nand U5444 (N_5444,N_4787,N_4651);
xnor U5445 (N_5445,N_4602,N_4605);
nor U5446 (N_5446,N_4218,N_4576);
and U5447 (N_5447,N_4966,N_4767);
xor U5448 (N_5448,N_4494,N_4326);
xor U5449 (N_5449,N_4042,N_4555);
nand U5450 (N_5450,N_4040,N_4983);
and U5451 (N_5451,N_4415,N_4023);
xnor U5452 (N_5452,N_4766,N_4460);
or U5453 (N_5453,N_4678,N_4445);
nor U5454 (N_5454,N_4378,N_4735);
or U5455 (N_5455,N_4757,N_4617);
xor U5456 (N_5456,N_4293,N_4057);
xor U5457 (N_5457,N_4477,N_4953);
nand U5458 (N_5458,N_4522,N_4395);
xor U5459 (N_5459,N_4917,N_4430);
nor U5460 (N_5460,N_4109,N_4392);
xor U5461 (N_5461,N_4598,N_4887);
xnor U5462 (N_5462,N_4196,N_4268);
nor U5463 (N_5463,N_4381,N_4112);
nor U5464 (N_5464,N_4150,N_4272);
or U5465 (N_5465,N_4763,N_4808);
nor U5466 (N_5466,N_4881,N_4664);
nor U5467 (N_5467,N_4825,N_4674);
xnor U5468 (N_5468,N_4209,N_4233);
nand U5469 (N_5469,N_4500,N_4344);
or U5470 (N_5470,N_4049,N_4269);
nor U5471 (N_5471,N_4597,N_4341);
nor U5472 (N_5472,N_4950,N_4287);
xor U5473 (N_5473,N_4421,N_4581);
and U5474 (N_5474,N_4894,N_4683);
nor U5475 (N_5475,N_4594,N_4321);
xnor U5476 (N_5476,N_4432,N_4795);
xnor U5477 (N_5477,N_4161,N_4525);
xnor U5478 (N_5478,N_4399,N_4930);
or U5479 (N_5479,N_4073,N_4030);
and U5480 (N_5480,N_4772,N_4409);
or U5481 (N_5481,N_4476,N_4490);
nor U5482 (N_5482,N_4974,N_4638);
and U5483 (N_5483,N_4360,N_4457);
or U5484 (N_5484,N_4013,N_4908);
or U5485 (N_5485,N_4071,N_4834);
and U5486 (N_5486,N_4751,N_4914);
and U5487 (N_5487,N_4063,N_4149);
and U5488 (N_5488,N_4546,N_4493);
or U5489 (N_5489,N_4193,N_4860);
nor U5490 (N_5490,N_4591,N_4018);
nor U5491 (N_5491,N_4996,N_4369);
and U5492 (N_5492,N_4519,N_4659);
and U5493 (N_5493,N_4640,N_4031);
and U5494 (N_5494,N_4843,N_4517);
xor U5495 (N_5495,N_4962,N_4118);
nor U5496 (N_5496,N_4975,N_4614);
nand U5497 (N_5497,N_4727,N_4249);
nor U5498 (N_5498,N_4044,N_4701);
xnor U5499 (N_5499,N_4077,N_4286);
xor U5500 (N_5500,N_4972,N_4092);
and U5501 (N_5501,N_4298,N_4552);
or U5502 (N_5502,N_4759,N_4733);
xnor U5503 (N_5503,N_4470,N_4705);
nand U5504 (N_5504,N_4724,N_4951);
xnor U5505 (N_5505,N_4962,N_4894);
and U5506 (N_5506,N_4397,N_4043);
xnor U5507 (N_5507,N_4404,N_4322);
xor U5508 (N_5508,N_4540,N_4730);
nand U5509 (N_5509,N_4991,N_4848);
and U5510 (N_5510,N_4845,N_4871);
xnor U5511 (N_5511,N_4632,N_4548);
or U5512 (N_5512,N_4389,N_4978);
and U5513 (N_5513,N_4035,N_4711);
or U5514 (N_5514,N_4434,N_4101);
or U5515 (N_5515,N_4723,N_4869);
nor U5516 (N_5516,N_4092,N_4331);
or U5517 (N_5517,N_4400,N_4255);
and U5518 (N_5518,N_4724,N_4390);
and U5519 (N_5519,N_4750,N_4905);
or U5520 (N_5520,N_4334,N_4160);
or U5521 (N_5521,N_4800,N_4770);
nand U5522 (N_5522,N_4264,N_4158);
xor U5523 (N_5523,N_4770,N_4728);
xor U5524 (N_5524,N_4059,N_4170);
nor U5525 (N_5525,N_4927,N_4413);
and U5526 (N_5526,N_4421,N_4593);
and U5527 (N_5527,N_4357,N_4121);
or U5528 (N_5528,N_4276,N_4838);
nand U5529 (N_5529,N_4281,N_4113);
nand U5530 (N_5530,N_4534,N_4957);
and U5531 (N_5531,N_4610,N_4384);
xor U5532 (N_5532,N_4857,N_4907);
xor U5533 (N_5533,N_4741,N_4876);
nand U5534 (N_5534,N_4565,N_4300);
nand U5535 (N_5535,N_4524,N_4056);
nor U5536 (N_5536,N_4522,N_4565);
and U5537 (N_5537,N_4127,N_4312);
nand U5538 (N_5538,N_4927,N_4196);
or U5539 (N_5539,N_4187,N_4200);
xor U5540 (N_5540,N_4588,N_4221);
xnor U5541 (N_5541,N_4709,N_4214);
xnor U5542 (N_5542,N_4226,N_4091);
or U5543 (N_5543,N_4525,N_4173);
and U5544 (N_5544,N_4920,N_4413);
xor U5545 (N_5545,N_4639,N_4219);
and U5546 (N_5546,N_4120,N_4950);
xnor U5547 (N_5547,N_4888,N_4091);
nand U5548 (N_5548,N_4662,N_4235);
nor U5549 (N_5549,N_4142,N_4544);
xor U5550 (N_5550,N_4751,N_4947);
nand U5551 (N_5551,N_4598,N_4198);
and U5552 (N_5552,N_4479,N_4231);
xnor U5553 (N_5553,N_4152,N_4649);
nand U5554 (N_5554,N_4505,N_4922);
nand U5555 (N_5555,N_4081,N_4433);
nor U5556 (N_5556,N_4109,N_4485);
nor U5557 (N_5557,N_4339,N_4869);
xor U5558 (N_5558,N_4244,N_4078);
or U5559 (N_5559,N_4981,N_4189);
and U5560 (N_5560,N_4712,N_4453);
xnor U5561 (N_5561,N_4129,N_4981);
xnor U5562 (N_5562,N_4189,N_4111);
nand U5563 (N_5563,N_4307,N_4763);
or U5564 (N_5564,N_4206,N_4165);
and U5565 (N_5565,N_4323,N_4094);
nand U5566 (N_5566,N_4821,N_4151);
nand U5567 (N_5567,N_4965,N_4001);
or U5568 (N_5568,N_4076,N_4215);
xor U5569 (N_5569,N_4103,N_4118);
or U5570 (N_5570,N_4607,N_4080);
nand U5571 (N_5571,N_4094,N_4449);
nor U5572 (N_5572,N_4228,N_4577);
and U5573 (N_5573,N_4648,N_4224);
and U5574 (N_5574,N_4028,N_4023);
nand U5575 (N_5575,N_4915,N_4323);
or U5576 (N_5576,N_4189,N_4018);
xor U5577 (N_5577,N_4708,N_4269);
and U5578 (N_5578,N_4422,N_4861);
xnor U5579 (N_5579,N_4540,N_4009);
nor U5580 (N_5580,N_4793,N_4564);
and U5581 (N_5581,N_4704,N_4530);
nor U5582 (N_5582,N_4424,N_4968);
xor U5583 (N_5583,N_4815,N_4037);
nor U5584 (N_5584,N_4107,N_4605);
nand U5585 (N_5585,N_4628,N_4827);
xnor U5586 (N_5586,N_4445,N_4937);
and U5587 (N_5587,N_4663,N_4388);
or U5588 (N_5588,N_4983,N_4584);
or U5589 (N_5589,N_4221,N_4314);
and U5590 (N_5590,N_4621,N_4007);
nand U5591 (N_5591,N_4292,N_4908);
nor U5592 (N_5592,N_4690,N_4285);
and U5593 (N_5593,N_4817,N_4772);
nor U5594 (N_5594,N_4078,N_4233);
nand U5595 (N_5595,N_4474,N_4196);
and U5596 (N_5596,N_4453,N_4005);
xor U5597 (N_5597,N_4250,N_4069);
or U5598 (N_5598,N_4910,N_4376);
nand U5599 (N_5599,N_4981,N_4898);
and U5600 (N_5600,N_4426,N_4120);
xor U5601 (N_5601,N_4418,N_4468);
xor U5602 (N_5602,N_4192,N_4391);
nor U5603 (N_5603,N_4649,N_4504);
nand U5604 (N_5604,N_4090,N_4975);
xnor U5605 (N_5605,N_4259,N_4045);
nand U5606 (N_5606,N_4317,N_4851);
xor U5607 (N_5607,N_4714,N_4004);
xor U5608 (N_5608,N_4577,N_4451);
and U5609 (N_5609,N_4888,N_4436);
nor U5610 (N_5610,N_4495,N_4076);
and U5611 (N_5611,N_4746,N_4876);
nor U5612 (N_5612,N_4627,N_4822);
nor U5613 (N_5613,N_4516,N_4528);
nand U5614 (N_5614,N_4297,N_4412);
nor U5615 (N_5615,N_4550,N_4410);
xor U5616 (N_5616,N_4233,N_4800);
xor U5617 (N_5617,N_4803,N_4848);
nand U5618 (N_5618,N_4019,N_4068);
or U5619 (N_5619,N_4054,N_4780);
and U5620 (N_5620,N_4495,N_4135);
and U5621 (N_5621,N_4629,N_4021);
and U5622 (N_5622,N_4543,N_4917);
and U5623 (N_5623,N_4150,N_4256);
xnor U5624 (N_5624,N_4303,N_4688);
nor U5625 (N_5625,N_4261,N_4697);
or U5626 (N_5626,N_4474,N_4894);
xor U5627 (N_5627,N_4169,N_4564);
xor U5628 (N_5628,N_4716,N_4126);
nand U5629 (N_5629,N_4652,N_4771);
nor U5630 (N_5630,N_4750,N_4483);
or U5631 (N_5631,N_4742,N_4819);
or U5632 (N_5632,N_4155,N_4417);
nand U5633 (N_5633,N_4665,N_4383);
and U5634 (N_5634,N_4707,N_4384);
and U5635 (N_5635,N_4394,N_4276);
and U5636 (N_5636,N_4694,N_4010);
nor U5637 (N_5637,N_4423,N_4417);
nand U5638 (N_5638,N_4791,N_4270);
and U5639 (N_5639,N_4516,N_4552);
or U5640 (N_5640,N_4175,N_4063);
and U5641 (N_5641,N_4115,N_4752);
or U5642 (N_5642,N_4611,N_4136);
and U5643 (N_5643,N_4528,N_4751);
or U5644 (N_5644,N_4881,N_4832);
nor U5645 (N_5645,N_4267,N_4941);
and U5646 (N_5646,N_4262,N_4635);
nand U5647 (N_5647,N_4586,N_4457);
and U5648 (N_5648,N_4468,N_4745);
and U5649 (N_5649,N_4834,N_4387);
nand U5650 (N_5650,N_4707,N_4447);
nand U5651 (N_5651,N_4188,N_4056);
or U5652 (N_5652,N_4581,N_4624);
or U5653 (N_5653,N_4128,N_4764);
or U5654 (N_5654,N_4497,N_4219);
nor U5655 (N_5655,N_4019,N_4294);
nand U5656 (N_5656,N_4957,N_4411);
and U5657 (N_5657,N_4852,N_4434);
nor U5658 (N_5658,N_4055,N_4156);
and U5659 (N_5659,N_4228,N_4413);
and U5660 (N_5660,N_4614,N_4304);
and U5661 (N_5661,N_4825,N_4800);
nor U5662 (N_5662,N_4192,N_4755);
nor U5663 (N_5663,N_4011,N_4931);
nand U5664 (N_5664,N_4164,N_4790);
or U5665 (N_5665,N_4941,N_4988);
nand U5666 (N_5666,N_4104,N_4688);
nor U5667 (N_5667,N_4942,N_4784);
nand U5668 (N_5668,N_4371,N_4362);
or U5669 (N_5669,N_4641,N_4229);
and U5670 (N_5670,N_4932,N_4985);
and U5671 (N_5671,N_4729,N_4448);
xnor U5672 (N_5672,N_4461,N_4102);
nor U5673 (N_5673,N_4166,N_4868);
nor U5674 (N_5674,N_4617,N_4813);
or U5675 (N_5675,N_4344,N_4939);
or U5676 (N_5676,N_4895,N_4476);
nand U5677 (N_5677,N_4009,N_4623);
xor U5678 (N_5678,N_4507,N_4437);
nand U5679 (N_5679,N_4704,N_4413);
or U5680 (N_5680,N_4425,N_4620);
and U5681 (N_5681,N_4484,N_4388);
nor U5682 (N_5682,N_4074,N_4529);
xnor U5683 (N_5683,N_4170,N_4749);
or U5684 (N_5684,N_4247,N_4543);
and U5685 (N_5685,N_4446,N_4605);
nand U5686 (N_5686,N_4040,N_4945);
or U5687 (N_5687,N_4192,N_4280);
and U5688 (N_5688,N_4749,N_4712);
nand U5689 (N_5689,N_4070,N_4207);
xnor U5690 (N_5690,N_4880,N_4013);
and U5691 (N_5691,N_4431,N_4011);
nor U5692 (N_5692,N_4115,N_4464);
nor U5693 (N_5693,N_4781,N_4987);
xnor U5694 (N_5694,N_4058,N_4827);
nand U5695 (N_5695,N_4166,N_4593);
nand U5696 (N_5696,N_4259,N_4310);
and U5697 (N_5697,N_4197,N_4776);
nor U5698 (N_5698,N_4051,N_4303);
nor U5699 (N_5699,N_4755,N_4942);
or U5700 (N_5700,N_4480,N_4538);
nand U5701 (N_5701,N_4248,N_4894);
nor U5702 (N_5702,N_4517,N_4408);
or U5703 (N_5703,N_4368,N_4503);
or U5704 (N_5704,N_4224,N_4922);
nand U5705 (N_5705,N_4648,N_4726);
nor U5706 (N_5706,N_4881,N_4628);
xor U5707 (N_5707,N_4320,N_4362);
or U5708 (N_5708,N_4124,N_4535);
nand U5709 (N_5709,N_4314,N_4300);
or U5710 (N_5710,N_4967,N_4635);
xnor U5711 (N_5711,N_4983,N_4765);
and U5712 (N_5712,N_4599,N_4392);
nor U5713 (N_5713,N_4513,N_4201);
nand U5714 (N_5714,N_4406,N_4688);
nand U5715 (N_5715,N_4247,N_4723);
nor U5716 (N_5716,N_4127,N_4729);
xnor U5717 (N_5717,N_4501,N_4881);
xnor U5718 (N_5718,N_4337,N_4890);
xor U5719 (N_5719,N_4388,N_4676);
nand U5720 (N_5720,N_4848,N_4572);
and U5721 (N_5721,N_4143,N_4845);
nand U5722 (N_5722,N_4148,N_4499);
xor U5723 (N_5723,N_4785,N_4341);
nand U5724 (N_5724,N_4942,N_4876);
and U5725 (N_5725,N_4492,N_4308);
or U5726 (N_5726,N_4472,N_4157);
nand U5727 (N_5727,N_4590,N_4059);
and U5728 (N_5728,N_4609,N_4325);
nand U5729 (N_5729,N_4130,N_4653);
and U5730 (N_5730,N_4096,N_4293);
or U5731 (N_5731,N_4536,N_4474);
nor U5732 (N_5732,N_4762,N_4150);
nand U5733 (N_5733,N_4463,N_4554);
or U5734 (N_5734,N_4590,N_4720);
xor U5735 (N_5735,N_4903,N_4824);
nor U5736 (N_5736,N_4081,N_4061);
xnor U5737 (N_5737,N_4532,N_4016);
xnor U5738 (N_5738,N_4785,N_4398);
and U5739 (N_5739,N_4112,N_4158);
xnor U5740 (N_5740,N_4189,N_4496);
nand U5741 (N_5741,N_4980,N_4758);
or U5742 (N_5742,N_4068,N_4627);
nor U5743 (N_5743,N_4983,N_4638);
and U5744 (N_5744,N_4799,N_4590);
xnor U5745 (N_5745,N_4242,N_4861);
or U5746 (N_5746,N_4817,N_4603);
nor U5747 (N_5747,N_4456,N_4132);
xor U5748 (N_5748,N_4270,N_4077);
xor U5749 (N_5749,N_4046,N_4134);
nand U5750 (N_5750,N_4320,N_4768);
nand U5751 (N_5751,N_4501,N_4756);
nor U5752 (N_5752,N_4277,N_4270);
xor U5753 (N_5753,N_4573,N_4714);
and U5754 (N_5754,N_4960,N_4332);
or U5755 (N_5755,N_4345,N_4734);
nor U5756 (N_5756,N_4299,N_4415);
or U5757 (N_5757,N_4375,N_4112);
or U5758 (N_5758,N_4525,N_4162);
xnor U5759 (N_5759,N_4570,N_4479);
xor U5760 (N_5760,N_4506,N_4621);
or U5761 (N_5761,N_4541,N_4516);
nor U5762 (N_5762,N_4130,N_4610);
or U5763 (N_5763,N_4685,N_4180);
or U5764 (N_5764,N_4114,N_4934);
nand U5765 (N_5765,N_4666,N_4001);
or U5766 (N_5766,N_4047,N_4621);
xor U5767 (N_5767,N_4697,N_4272);
or U5768 (N_5768,N_4931,N_4247);
nor U5769 (N_5769,N_4937,N_4825);
nand U5770 (N_5770,N_4645,N_4322);
nor U5771 (N_5771,N_4784,N_4943);
or U5772 (N_5772,N_4709,N_4397);
and U5773 (N_5773,N_4531,N_4509);
or U5774 (N_5774,N_4778,N_4932);
nand U5775 (N_5775,N_4251,N_4384);
nand U5776 (N_5776,N_4092,N_4045);
nor U5777 (N_5777,N_4719,N_4429);
xor U5778 (N_5778,N_4868,N_4881);
or U5779 (N_5779,N_4263,N_4847);
or U5780 (N_5780,N_4038,N_4125);
and U5781 (N_5781,N_4043,N_4348);
nand U5782 (N_5782,N_4649,N_4666);
nor U5783 (N_5783,N_4779,N_4436);
nor U5784 (N_5784,N_4322,N_4345);
nor U5785 (N_5785,N_4310,N_4255);
xnor U5786 (N_5786,N_4985,N_4574);
nor U5787 (N_5787,N_4458,N_4279);
or U5788 (N_5788,N_4874,N_4104);
and U5789 (N_5789,N_4740,N_4120);
and U5790 (N_5790,N_4555,N_4177);
xor U5791 (N_5791,N_4216,N_4602);
nand U5792 (N_5792,N_4821,N_4107);
xnor U5793 (N_5793,N_4407,N_4109);
xor U5794 (N_5794,N_4203,N_4897);
nand U5795 (N_5795,N_4524,N_4591);
xor U5796 (N_5796,N_4075,N_4808);
or U5797 (N_5797,N_4904,N_4024);
xor U5798 (N_5798,N_4251,N_4691);
nand U5799 (N_5799,N_4166,N_4341);
or U5800 (N_5800,N_4625,N_4913);
nand U5801 (N_5801,N_4264,N_4808);
nor U5802 (N_5802,N_4623,N_4799);
xor U5803 (N_5803,N_4549,N_4562);
and U5804 (N_5804,N_4990,N_4149);
and U5805 (N_5805,N_4288,N_4428);
and U5806 (N_5806,N_4388,N_4694);
or U5807 (N_5807,N_4146,N_4327);
or U5808 (N_5808,N_4033,N_4727);
nor U5809 (N_5809,N_4309,N_4606);
or U5810 (N_5810,N_4230,N_4999);
nand U5811 (N_5811,N_4470,N_4472);
xnor U5812 (N_5812,N_4736,N_4972);
and U5813 (N_5813,N_4864,N_4340);
and U5814 (N_5814,N_4971,N_4241);
or U5815 (N_5815,N_4114,N_4111);
and U5816 (N_5816,N_4234,N_4508);
and U5817 (N_5817,N_4532,N_4652);
nor U5818 (N_5818,N_4967,N_4697);
nor U5819 (N_5819,N_4431,N_4323);
nor U5820 (N_5820,N_4201,N_4651);
xor U5821 (N_5821,N_4236,N_4047);
and U5822 (N_5822,N_4376,N_4092);
or U5823 (N_5823,N_4497,N_4768);
or U5824 (N_5824,N_4782,N_4338);
nand U5825 (N_5825,N_4347,N_4432);
nand U5826 (N_5826,N_4569,N_4942);
nand U5827 (N_5827,N_4339,N_4757);
nor U5828 (N_5828,N_4970,N_4389);
xor U5829 (N_5829,N_4313,N_4091);
or U5830 (N_5830,N_4690,N_4268);
nor U5831 (N_5831,N_4375,N_4690);
and U5832 (N_5832,N_4044,N_4421);
nand U5833 (N_5833,N_4376,N_4482);
nor U5834 (N_5834,N_4569,N_4762);
or U5835 (N_5835,N_4381,N_4365);
or U5836 (N_5836,N_4664,N_4651);
xnor U5837 (N_5837,N_4680,N_4662);
and U5838 (N_5838,N_4369,N_4632);
nand U5839 (N_5839,N_4194,N_4396);
nand U5840 (N_5840,N_4509,N_4800);
xor U5841 (N_5841,N_4049,N_4829);
xnor U5842 (N_5842,N_4348,N_4699);
and U5843 (N_5843,N_4512,N_4468);
and U5844 (N_5844,N_4130,N_4542);
nor U5845 (N_5845,N_4560,N_4499);
nor U5846 (N_5846,N_4630,N_4657);
nor U5847 (N_5847,N_4719,N_4289);
and U5848 (N_5848,N_4060,N_4795);
nor U5849 (N_5849,N_4779,N_4327);
and U5850 (N_5850,N_4659,N_4720);
nor U5851 (N_5851,N_4185,N_4538);
xnor U5852 (N_5852,N_4257,N_4079);
nand U5853 (N_5853,N_4952,N_4724);
nor U5854 (N_5854,N_4488,N_4811);
or U5855 (N_5855,N_4303,N_4088);
nand U5856 (N_5856,N_4892,N_4829);
nor U5857 (N_5857,N_4225,N_4832);
or U5858 (N_5858,N_4777,N_4031);
or U5859 (N_5859,N_4119,N_4597);
and U5860 (N_5860,N_4782,N_4475);
xor U5861 (N_5861,N_4847,N_4001);
nand U5862 (N_5862,N_4831,N_4716);
nand U5863 (N_5863,N_4370,N_4157);
or U5864 (N_5864,N_4855,N_4497);
nand U5865 (N_5865,N_4666,N_4683);
nand U5866 (N_5866,N_4004,N_4254);
or U5867 (N_5867,N_4761,N_4672);
or U5868 (N_5868,N_4466,N_4866);
nor U5869 (N_5869,N_4929,N_4629);
or U5870 (N_5870,N_4613,N_4051);
xnor U5871 (N_5871,N_4101,N_4860);
xnor U5872 (N_5872,N_4253,N_4843);
nand U5873 (N_5873,N_4134,N_4131);
or U5874 (N_5874,N_4145,N_4630);
nand U5875 (N_5875,N_4107,N_4266);
and U5876 (N_5876,N_4054,N_4102);
and U5877 (N_5877,N_4807,N_4311);
nand U5878 (N_5878,N_4793,N_4381);
nand U5879 (N_5879,N_4252,N_4129);
and U5880 (N_5880,N_4630,N_4332);
nor U5881 (N_5881,N_4870,N_4831);
nor U5882 (N_5882,N_4858,N_4098);
and U5883 (N_5883,N_4935,N_4889);
nor U5884 (N_5884,N_4855,N_4905);
xor U5885 (N_5885,N_4390,N_4890);
and U5886 (N_5886,N_4531,N_4517);
nand U5887 (N_5887,N_4715,N_4535);
or U5888 (N_5888,N_4546,N_4558);
xor U5889 (N_5889,N_4918,N_4504);
nand U5890 (N_5890,N_4316,N_4764);
and U5891 (N_5891,N_4262,N_4284);
xor U5892 (N_5892,N_4044,N_4920);
and U5893 (N_5893,N_4831,N_4747);
nor U5894 (N_5894,N_4932,N_4434);
nor U5895 (N_5895,N_4134,N_4571);
nor U5896 (N_5896,N_4873,N_4092);
or U5897 (N_5897,N_4743,N_4634);
nand U5898 (N_5898,N_4638,N_4728);
or U5899 (N_5899,N_4257,N_4427);
nor U5900 (N_5900,N_4955,N_4568);
or U5901 (N_5901,N_4061,N_4720);
nand U5902 (N_5902,N_4782,N_4799);
or U5903 (N_5903,N_4987,N_4970);
nand U5904 (N_5904,N_4281,N_4227);
or U5905 (N_5905,N_4455,N_4604);
or U5906 (N_5906,N_4328,N_4468);
nand U5907 (N_5907,N_4621,N_4142);
nand U5908 (N_5908,N_4835,N_4982);
or U5909 (N_5909,N_4763,N_4552);
and U5910 (N_5910,N_4374,N_4623);
or U5911 (N_5911,N_4498,N_4462);
xnor U5912 (N_5912,N_4238,N_4463);
and U5913 (N_5913,N_4982,N_4517);
nor U5914 (N_5914,N_4493,N_4715);
nor U5915 (N_5915,N_4444,N_4218);
nor U5916 (N_5916,N_4837,N_4503);
xor U5917 (N_5917,N_4344,N_4430);
xor U5918 (N_5918,N_4388,N_4131);
and U5919 (N_5919,N_4239,N_4389);
and U5920 (N_5920,N_4471,N_4797);
and U5921 (N_5921,N_4651,N_4351);
or U5922 (N_5922,N_4344,N_4625);
or U5923 (N_5923,N_4092,N_4963);
or U5924 (N_5924,N_4262,N_4621);
nor U5925 (N_5925,N_4680,N_4163);
nor U5926 (N_5926,N_4024,N_4562);
nand U5927 (N_5927,N_4691,N_4831);
nor U5928 (N_5928,N_4312,N_4726);
xor U5929 (N_5929,N_4909,N_4957);
xor U5930 (N_5930,N_4483,N_4997);
xnor U5931 (N_5931,N_4029,N_4942);
nand U5932 (N_5932,N_4147,N_4433);
and U5933 (N_5933,N_4537,N_4184);
or U5934 (N_5934,N_4853,N_4211);
and U5935 (N_5935,N_4568,N_4696);
or U5936 (N_5936,N_4450,N_4302);
nand U5937 (N_5937,N_4650,N_4790);
or U5938 (N_5938,N_4323,N_4925);
and U5939 (N_5939,N_4639,N_4871);
nor U5940 (N_5940,N_4138,N_4132);
and U5941 (N_5941,N_4176,N_4341);
and U5942 (N_5942,N_4335,N_4963);
or U5943 (N_5943,N_4370,N_4553);
or U5944 (N_5944,N_4095,N_4503);
and U5945 (N_5945,N_4091,N_4628);
and U5946 (N_5946,N_4290,N_4383);
and U5947 (N_5947,N_4406,N_4863);
xor U5948 (N_5948,N_4688,N_4790);
or U5949 (N_5949,N_4147,N_4266);
nor U5950 (N_5950,N_4520,N_4009);
nand U5951 (N_5951,N_4014,N_4088);
or U5952 (N_5952,N_4906,N_4194);
nor U5953 (N_5953,N_4808,N_4686);
or U5954 (N_5954,N_4871,N_4162);
or U5955 (N_5955,N_4557,N_4007);
or U5956 (N_5956,N_4011,N_4159);
nand U5957 (N_5957,N_4793,N_4279);
xnor U5958 (N_5958,N_4507,N_4984);
nor U5959 (N_5959,N_4003,N_4882);
xnor U5960 (N_5960,N_4835,N_4179);
nor U5961 (N_5961,N_4842,N_4675);
nor U5962 (N_5962,N_4172,N_4943);
xor U5963 (N_5963,N_4741,N_4282);
xnor U5964 (N_5964,N_4662,N_4195);
nand U5965 (N_5965,N_4866,N_4972);
and U5966 (N_5966,N_4496,N_4346);
or U5967 (N_5967,N_4682,N_4461);
xnor U5968 (N_5968,N_4695,N_4685);
nand U5969 (N_5969,N_4811,N_4374);
or U5970 (N_5970,N_4139,N_4884);
nand U5971 (N_5971,N_4526,N_4984);
and U5972 (N_5972,N_4842,N_4545);
nand U5973 (N_5973,N_4027,N_4491);
nor U5974 (N_5974,N_4084,N_4108);
and U5975 (N_5975,N_4882,N_4479);
or U5976 (N_5976,N_4757,N_4288);
and U5977 (N_5977,N_4999,N_4721);
or U5978 (N_5978,N_4051,N_4900);
xor U5979 (N_5979,N_4807,N_4725);
and U5980 (N_5980,N_4149,N_4585);
xor U5981 (N_5981,N_4967,N_4498);
and U5982 (N_5982,N_4484,N_4935);
or U5983 (N_5983,N_4165,N_4255);
and U5984 (N_5984,N_4898,N_4227);
xor U5985 (N_5985,N_4014,N_4712);
nand U5986 (N_5986,N_4841,N_4162);
nor U5987 (N_5987,N_4113,N_4942);
xnor U5988 (N_5988,N_4572,N_4830);
nand U5989 (N_5989,N_4019,N_4835);
nor U5990 (N_5990,N_4374,N_4788);
nand U5991 (N_5991,N_4805,N_4719);
xor U5992 (N_5992,N_4488,N_4138);
nand U5993 (N_5993,N_4024,N_4320);
and U5994 (N_5994,N_4876,N_4098);
xnor U5995 (N_5995,N_4759,N_4922);
and U5996 (N_5996,N_4427,N_4087);
xnor U5997 (N_5997,N_4712,N_4013);
nand U5998 (N_5998,N_4954,N_4287);
nor U5999 (N_5999,N_4442,N_4701);
and U6000 (N_6000,N_5645,N_5141);
or U6001 (N_6001,N_5860,N_5493);
nor U6002 (N_6002,N_5047,N_5420);
xor U6003 (N_6003,N_5211,N_5407);
or U6004 (N_6004,N_5812,N_5589);
nand U6005 (N_6005,N_5334,N_5419);
nor U6006 (N_6006,N_5185,N_5929);
xor U6007 (N_6007,N_5956,N_5290);
nand U6008 (N_6008,N_5619,N_5488);
and U6009 (N_6009,N_5104,N_5487);
nor U6010 (N_6010,N_5457,N_5733);
or U6011 (N_6011,N_5077,N_5202);
nand U6012 (N_6012,N_5971,N_5554);
or U6013 (N_6013,N_5530,N_5118);
nor U6014 (N_6014,N_5258,N_5542);
or U6015 (N_6015,N_5351,N_5189);
nor U6016 (N_6016,N_5865,N_5361);
or U6017 (N_6017,N_5350,N_5581);
nor U6018 (N_6018,N_5596,N_5228);
and U6019 (N_6019,N_5509,N_5900);
xnor U6020 (N_6020,N_5021,N_5230);
xor U6021 (N_6021,N_5379,N_5630);
or U6022 (N_6022,N_5825,N_5239);
xnor U6023 (N_6023,N_5867,N_5483);
xor U6024 (N_6024,N_5293,N_5845);
nand U6025 (N_6025,N_5218,N_5306);
xor U6026 (N_6026,N_5615,N_5428);
nand U6027 (N_6027,N_5526,N_5832);
and U6028 (N_6028,N_5355,N_5169);
and U6029 (N_6029,N_5314,N_5690);
nor U6030 (N_6030,N_5089,N_5841);
nor U6031 (N_6031,N_5548,N_5344);
nor U6032 (N_6032,N_5943,N_5128);
and U6033 (N_6033,N_5427,N_5133);
nand U6034 (N_6034,N_5784,N_5498);
xor U6035 (N_6035,N_5363,N_5553);
nand U6036 (N_6036,N_5154,N_5013);
and U6037 (N_6037,N_5364,N_5651);
nand U6038 (N_6038,N_5280,N_5255);
nor U6039 (N_6039,N_5271,N_5269);
xnor U6040 (N_6040,N_5728,N_5816);
or U6041 (N_6041,N_5541,N_5009);
or U6042 (N_6042,N_5932,N_5330);
or U6043 (N_6043,N_5850,N_5472);
or U6044 (N_6044,N_5066,N_5984);
or U6045 (N_6045,N_5511,N_5741);
nand U6046 (N_6046,N_5224,N_5672);
and U6047 (N_6047,N_5256,N_5573);
nand U6048 (N_6048,N_5312,N_5222);
nor U6049 (N_6049,N_5149,N_5432);
nor U6050 (N_6050,N_5975,N_5112);
or U6051 (N_6051,N_5979,N_5138);
and U6052 (N_6052,N_5757,N_5952);
or U6053 (N_6053,N_5086,N_5034);
xnor U6054 (N_6054,N_5147,N_5491);
or U6055 (N_6055,N_5756,N_5729);
and U6056 (N_6056,N_5958,N_5988);
xor U6057 (N_6057,N_5715,N_5270);
nand U6058 (N_6058,N_5950,N_5263);
xnor U6059 (N_6059,N_5347,N_5685);
nor U6060 (N_6060,N_5305,N_5377);
nor U6061 (N_6061,N_5739,N_5215);
nand U6062 (N_6062,N_5699,N_5184);
xor U6063 (N_6063,N_5083,N_5074);
and U6064 (N_6064,N_5858,N_5539);
and U6065 (N_6065,N_5571,N_5521);
nor U6066 (N_6066,N_5054,N_5558);
and U6067 (N_6067,N_5041,N_5309);
xnor U6068 (N_6068,N_5423,N_5879);
or U6069 (N_6069,N_5180,N_5683);
or U6070 (N_6070,N_5694,N_5060);
xnor U6071 (N_6071,N_5899,N_5671);
or U6072 (N_6072,N_5249,N_5406);
and U6073 (N_6073,N_5643,N_5904);
nor U6074 (N_6074,N_5325,N_5183);
nor U6075 (N_6075,N_5523,N_5804);
or U6076 (N_6076,N_5079,N_5378);
xor U6077 (N_6077,N_5072,N_5916);
and U6078 (N_6078,N_5486,N_5259);
nor U6079 (N_6079,N_5278,N_5903);
xnor U6080 (N_6080,N_5459,N_5385);
and U6081 (N_6081,N_5976,N_5076);
xnor U6082 (N_6082,N_5106,N_5452);
xnor U6083 (N_6083,N_5182,N_5028);
or U6084 (N_6084,N_5122,N_5124);
or U6085 (N_6085,N_5603,N_5474);
nand U6086 (N_6086,N_5114,N_5875);
nor U6087 (N_6087,N_5982,N_5636);
xor U6088 (N_6088,N_5000,N_5084);
or U6089 (N_6089,N_5235,N_5968);
and U6090 (N_6090,N_5092,N_5658);
nand U6091 (N_6091,N_5640,N_5939);
nand U6092 (N_6092,N_5050,N_5796);
nand U6093 (N_6093,N_5856,N_5513);
and U6094 (N_6094,N_5338,N_5771);
xnor U6095 (N_6095,N_5160,N_5388);
and U6096 (N_6096,N_5605,N_5700);
nor U6097 (N_6097,N_5930,N_5425);
or U6098 (N_6098,N_5518,N_5246);
xor U6099 (N_6099,N_5620,N_5641);
or U6100 (N_6100,N_5404,N_5579);
nor U6101 (N_6101,N_5545,N_5873);
and U6102 (N_6102,N_5177,N_5460);
or U6103 (N_6103,N_5842,N_5310);
nor U6104 (N_6104,N_5260,N_5098);
or U6105 (N_6105,N_5787,N_5225);
or U6106 (N_6106,N_5667,N_5399);
nand U6107 (N_6107,N_5738,N_5265);
xor U6108 (N_6108,N_5241,N_5924);
and U6109 (N_6109,N_5445,N_5071);
nor U6110 (N_6110,N_5535,N_5159);
or U6111 (N_6111,N_5520,N_5876);
nor U6112 (N_6112,N_5957,N_5618);
or U6113 (N_6113,N_5512,N_5301);
nand U6114 (N_6114,N_5203,N_5770);
nand U6115 (N_6115,N_5067,N_5917);
or U6116 (N_6116,N_5623,N_5110);
nand U6117 (N_6117,N_5100,N_5023);
nor U6118 (N_6118,N_5552,N_5343);
or U6119 (N_6119,N_5339,N_5781);
nand U6120 (N_6120,N_5284,N_5938);
nor U6121 (N_6121,N_5393,N_5703);
nor U6122 (N_6122,N_5614,N_5172);
xnor U6123 (N_6123,N_5760,N_5580);
xnor U6124 (N_6124,N_5540,N_5257);
and U6125 (N_6125,N_5805,N_5758);
and U6126 (N_6126,N_5859,N_5161);
nor U6127 (N_6127,N_5806,N_5061);
xnor U6128 (N_6128,N_5598,N_5019);
xor U6129 (N_6129,N_5358,N_5820);
and U6130 (N_6130,N_5441,N_5735);
nor U6131 (N_6131,N_5208,N_5666);
nand U6132 (N_6132,N_5273,N_5788);
and U6133 (N_6133,N_5676,N_5148);
and U6134 (N_6134,N_5763,N_5102);
nor U6135 (N_6135,N_5800,N_5433);
and U6136 (N_6136,N_5714,N_5550);
xnor U6137 (N_6137,N_5704,N_5489);
nand U6138 (N_6138,N_5448,N_5769);
nand U6139 (N_6139,N_5582,N_5568);
nor U6140 (N_6140,N_5337,N_5267);
xor U6141 (N_6141,N_5586,N_5017);
or U6142 (N_6142,N_5707,N_5212);
xor U6143 (N_6143,N_5204,N_5368);
nor U6144 (N_6144,N_5458,N_5549);
nand U6145 (N_6145,N_5893,N_5918);
and U6146 (N_6146,N_5570,N_5990);
and U6147 (N_6147,N_5164,N_5591);
xnor U6148 (N_6148,N_5555,N_5977);
and U6149 (N_6149,N_5340,N_5109);
nor U6150 (N_6150,N_5562,N_5536);
and U6151 (N_6151,N_5751,N_5687);
and U6152 (N_6152,N_5882,N_5995);
nand U6153 (N_6153,N_5969,N_5680);
nand U6154 (N_6154,N_5702,N_5030);
and U6155 (N_6155,N_5025,N_5986);
and U6156 (N_6156,N_5219,N_5966);
nor U6157 (N_6157,N_5561,N_5413);
or U6158 (N_6158,N_5889,N_5764);
nor U6159 (N_6159,N_5798,N_5048);
nand U6160 (N_6160,N_5371,N_5035);
and U6161 (N_6161,N_5409,N_5120);
or U6162 (N_6162,N_5972,N_5888);
and U6163 (N_6163,N_5229,N_5813);
nand U6164 (N_6164,N_5892,N_5942);
and U6165 (N_6165,N_5822,N_5283);
and U6166 (N_6166,N_5901,N_5116);
and U6167 (N_6167,N_5342,N_5624);
or U6168 (N_6168,N_5998,N_5611);
nor U6169 (N_6169,N_5210,N_5227);
nor U6170 (N_6170,N_5849,N_5522);
and U6171 (N_6171,N_5890,N_5261);
or U6172 (N_6172,N_5543,N_5201);
nand U6173 (N_6173,N_5031,N_5776);
nand U6174 (N_6174,N_5115,N_5839);
xnor U6175 (N_6175,N_5983,N_5497);
and U6176 (N_6176,N_5818,N_5987);
and U6177 (N_6177,N_5723,N_5479);
xnor U6178 (N_6178,N_5237,N_5682);
and U6179 (N_6179,N_5401,N_5248);
or U6180 (N_6180,N_5777,N_5285);
nor U6181 (N_6181,N_5463,N_5477);
nand U6182 (N_6182,N_5604,N_5706);
and U6183 (N_6183,N_5473,N_5754);
or U6184 (N_6184,N_5710,N_5322);
nor U6185 (N_6185,N_5029,N_5455);
nor U6186 (N_6186,N_5327,N_5417);
nand U6187 (N_6187,N_5366,N_5236);
and U6188 (N_6188,N_5033,N_5991);
xor U6189 (N_6189,N_5563,N_5588);
or U6190 (N_6190,N_5332,N_5716);
xor U6191 (N_6191,N_5912,N_5181);
nand U6192 (N_6192,N_5302,N_5962);
and U6193 (N_6193,N_5864,N_5008);
or U6194 (N_6194,N_5557,N_5802);
and U6195 (N_6195,N_5176,N_5749);
and U6196 (N_6196,N_5386,N_5069);
nor U6197 (N_6197,N_5383,N_5575);
xnor U6198 (N_6198,N_5747,N_5357);
or U6199 (N_6199,N_5884,N_5701);
nand U6200 (N_6200,N_5855,N_5821);
nand U6201 (N_6201,N_5384,N_5346);
or U6202 (N_6202,N_5765,N_5315);
nand U6203 (N_6203,N_5251,N_5577);
xnor U6204 (N_6204,N_5380,N_5585);
nand U6205 (N_6205,N_5944,N_5226);
nor U6206 (N_6206,N_5426,N_5453);
nand U6207 (N_6207,N_5827,N_5424);
or U6208 (N_6208,N_5403,N_5913);
nand U6209 (N_6209,N_5705,N_5005);
and U6210 (N_6210,N_5398,N_5949);
nand U6211 (N_6211,N_5857,N_5602);
xnor U6212 (N_6212,N_5783,N_5768);
nand U6213 (N_6213,N_5815,N_5199);
xor U6214 (N_6214,N_5915,N_5049);
and U6215 (N_6215,N_5253,N_5797);
nor U6216 (N_6216,N_5795,N_5078);
or U6217 (N_6217,N_5119,N_5170);
and U6218 (N_6218,N_5967,N_5300);
xor U6219 (N_6219,N_5501,N_5297);
or U6220 (N_6220,N_5410,N_5039);
nand U6221 (N_6221,N_5247,N_5779);
or U6222 (N_6222,N_5252,N_5157);
nand U6223 (N_6223,N_5923,N_5447);
or U6224 (N_6224,N_5625,N_5209);
xor U6225 (N_6225,N_5935,N_5730);
or U6226 (N_6226,N_5907,N_5782);
xnor U6227 (N_6227,N_5131,N_5173);
and U6228 (N_6228,N_5608,N_5742);
xor U6229 (N_6229,N_5087,N_5055);
nor U6230 (N_6230,N_5759,N_5853);
or U6231 (N_6231,N_5767,N_5878);
and U6232 (N_6232,N_5994,N_5367);
and U6233 (N_6233,N_5593,N_5231);
nand U6234 (N_6234,N_5547,N_5153);
xnor U6235 (N_6235,N_5387,N_5809);
nor U6236 (N_6236,N_5633,N_5937);
or U6237 (N_6237,N_5877,N_5693);
xor U6238 (N_6238,N_5438,N_5725);
and U6239 (N_6239,N_5740,N_5205);
xnor U6240 (N_6240,N_5003,N_5885);
xnor U6241 (N_6241,N_5179,N_5674);
xor U6242 (N_6242,N_5372,N_5429);
and U6243 (N_6243,N_5773,N_5287);
nor U6244 (N_6244,N_5093,N_5673);
nand U6245 (N_6245,N_5369,N_5471);
and U6246 (N_6246,N_5648,N_5908);
nor U6247 (N_6247,N_5277,N_5400);
or U6248 (N_6248,N_5774,N_5635);
and U6249 (N_6249,N_5750,N_5657);
nand U6250 (N_6250,N_5799,N_5794);
or U6251 (N_6251,N_5391,N_5188);
or U6252 (N_6252,N_5838,N_5698);
nand U6253 (N_6253,N_5091,N_5217);
nand U6254 (N_6254,N_5677,N_5151);
nand U6255 (N_6255,N_5663,N_5508);
or U6256 (N_6256,N_5282,N_5684);
nor U6257 (N_6257,N_5560,N_5466);
nor U6258 (N_6258,N_5303,N_5503);
xor U6259 (N_6259,N_5175,N_5482);
and U6260 (N_6260,N_5524,N_5254);
nor U6261 (N_6261,N_5318,N_5243);
nand U6262 (N_6262,N_5960,N_5238);
or U6263 (N_6263,N_5103,N_5389);
or U6264 (N_6264,N_5519,N_5527);
nand U6265 (N_6265,N_5496,N_5475);
nor U6266 (N_6266,N_5370,N_5381);
nand U6267 (N_6267,N_5495,N_5748);
and U6268 (N_6268,N_5057,N_5360);
xor U6269 (N_6269,N_5135,N_5016);
or U6270 (N_6270,N_5947,N_5286);
nor U6271 (N_6271,N_5652,N_5439);
or U6272 (N_6272,N_5661,N_5974);
or U6273 (N_6273,N_5814,N_5861);
nor U6274 (N_6274,N_5992,N_5697);
nand U6275 (N_6275,N_5752,N_5801);
nand U6276 (N_6276,N_5090,N_5951);
and U6277 (N_6277,N_5689,N_5140);
nor U6278 (N_6278,N_5584,N_5245);
and U6279 (N_6279,N_5056,N_5022);
or U6280 (N_6280,N_5139,N_5043);
nand U6281 (N_6281,N_5727,N_5015);
or U6282 (N_6282,N_5696,N_5601);
xnor U6283 (N_6283,N_5333,N_5392);
nor U6284 (N_6284,N_5510,N_5440);
or U6285 (N_6285,N_5150,N_5376);
nand U6286 (N_6286,N_5668,N_5127);
nand U6287 (N_6287,N_5528,N_5617);
or U6288 (N_6288,N_5349,N_5365);
or U6289 (N_6289,N_5559,N_5037);
nand U6290 (N_6290,N_5088,N_5639);
xor U6291 (N_6291,N_5921,N_5772);
nand U6292 (N_6292,N_5791,N_5662);
nor U6293 (N_6293,N_5324,N_5709);
or U6294 (N_6294,N_5281,N_5665);
xnor U6295 (N_6295,N_5162,N_5163);
xnor U6296 (N_6296,N_5627,N_5394);
or U6297 (N_6297,N_5922,N_5828);
nor U6298 (N_6298,N_5085,N_5279);
or U6299 (N_6299,N_5823,N_5631);
xor U6300 (N_6300,N_5111,N_5012);
xor U6301 (N_6301,N_5020,N_5925);
nor U6302 (N_6302,N_5565,N_5691);
nand U6303 (N_6303,N_5973,N_5240);
or U6304 (N_6304,N_5027,N_5637);
xnor U6305 (N_6305,N_5656,N_5412);
nor U6306 (N_6306,N_5449,N_5762);
nand U6307 (N_6307,N_5062,N_5080);
or U6308 (N_6308,N_5946,N_5854);
xnor U6309 (N_6309,N_5775,N_5959);
and U6310 (N_6310,N_5507,N_5713);
and U6311 (N_6311,N_5026,N_5622);
or U6312 (N_6312,N_5965,N_5011);
xnor U6313 (N_6313,N_5634,N_5505);
xnor U6314 (N_6314,N_5985,N_5961);
xnor U6315 (N_6315,N_5874,N_5955);
nand U6316 (N_6316,N_5356,N_5712);
nand U6317 (N_6317,N_5166,N_5650);
and U6318 (N_6318,N_5444,N_5534);
or U6319 (N_6319,N_5107,N_5038);
and U6320 (N_6320,N_5004,N_5316);
and U6321 (N_6321,N_5953,N_5353);
or U6322 (N_6322,N_5606,N_5736);
nand U6323 (N_6323,N_5213,N_5362);
xor U6324 (N_6324,N_5233,N_5099);
nor U6325 (N_6325,N_5590,N_5051);
or U6326 (N_6326,N_5480,N_5272);
and U6327 (N_6327,N_5517,N_5044);
or U6328 (N_6328,N_5970,N_5121);
nand U6329 (N_6329,N_5108,N_5612);
xnor U6330 (N_6330,N_5328,N_5808);
and U6331 (N_6331,N_5345,N_5375);
or U6332 (N_6332,N_5920,N_5926);
xor U6333 (N_6333,N_5997,N_5834);
nand U6334 (N_6334,N_5569,N_5819);
xor U6335 (N_6335,N_5105,N_5018);
xnor U6336 (N_6336,N_5313,N_5137);
xnor U6337 (N_6337,N_5195,N_5826);
or U6338 (N_6338,N_5145,N_5533);
nand U6339 (N_6339,N_5803,N_5167);
or U6340 (N_6340,N_5894,N_5152);
and U6341 (N_6341,N_5928,N_5659);
nand U6342 (N_6342,N_5244,N_5075);
and U6343 (N_6343,N_5686,N_5556);
and U6344 (N_6344,N_5307,N_5927);
and U6345 (N_6345,N_5609,N_5616);
nand U6346 (N_6346,N_5500,N_5341);
or U6347 (N_6347,N_5352,N_5430);
and U6348 (N_6348,N_5649,N_5442);
or U6349 (N_6349,N_5531,N_5397);
nand U6350 (N_6350,N_5905,N_5276);
and U6351 (N_6351,N_5416,N_5989);
nand U6352 (N_6352,N_5792,N_5669);
nand U6353 (N_6353,N_5870,N_5024);
nand U6354 (N_6354,N_5132,N_5732);
xor U6355 (N_6355,N_5469,N_5001);
xnor U6356 (N_6356,N_5722,N_5978);
nor U6357 (N_6357,N_5123,N_5654);
nand U6358 (N_6358,N_5317,N_5296);
and U6359 (N_6359,N_5506,N_5817);
or U6360 (N_6360,N_5014,N_5436);
and U6361 (N_6361,N_5902,N_5094);
and U6362 (N_6362,N_5117,N_5156);
xor U6363 (N_6363,N_5931,N_5653);
and U6364 (N_6364,N_5097,N_5996);
or U6365 (N_6365,N_5896,N_5963);
nor U6366 (N_6366,N_5191,N_5232);
or U6367 (N_6367,N_5032,N_5871);
and U6368 (N_6368,N_5354,N_5909);
and U6369 (N_6369,N_5190,N_5600);
xor U6370 (N_6370,N_5734,N_5485);
xor U6371 (N_6371,N_5621,N_5793);
nand U6372 (N_6372,N_5846,N_5880);
nor U6373 (N_6373,N_5134,N_5451);
nor U6374 (N_6374,N_5544,N_5396);
or U6375 (N_6375,N_5036,N_5264);
nand U6376 (N_6376,N_5981,N_5664);
and U6377 (N_6377,N_5829,N_5242);
nor U6378 (N_6378,N_5359,N_5578);
nand U6379 (N_6379,N_5143,N_5298);
nor U6380 (N_6380,N_5613,N_5414);
and U6381 (N_6381,N_5868,N_5187);
nor U6382 (N_6382,N_5848,N_5844);
or U6383 (N_6383,N_5484,N_5010);
xor U6384 (N_6384,N_5395,N_5895);
nor U6385 (N_6385,N_5743,N_5638);
or U6386 (N_6386,N_5288,N_5872);
nor U6387 (N_6387,N_5766,N_5335);
or U6388 (N_6388,N_5113,N_5833);
and U6389 (N_6389,N_5807,N_5964);
or U6390 (N_6390,N_5142,N_5891);
or U6391 (N_6391,N_5655,N_5411);
nand U6392 (N_6392,N_5945,N_5897);
and U6393 (N_6393,N_5914,N_5171);
and U6394 (N_6394,N_5476,N_5464);
or U6395 (N_6395,N_5761,N_5726);
and U6396 (N_6396,N_5786,N_5869);
xnor U6397 (N_6397,N_5262,N_5144);
nor U6398 (N_6398,N_5502,N_5192);
nand U6399 (N_6399,N_5268,N_5538);
or U6400 (N_6400,N_5193,N_5745);
nor U6401 (N_6401,N_5574,N_5478);
and U6402 (N_6402,N_5980,N_5331);
xnor U6403 (N_6403,N_5717,N_5881);
xor U6404 (N_6404,N_5883,N_5940);
and U6405 (N_6405,N_5007,N_5753);
xor U6406 (N_6406,N_5678,N_5824);
xor U6407 (N_6407,N_5304,N_5168);
or U6408 (N_6408,N_5450,N_5592);
xnor U6409 (N_6409,N_5186,N_5852);
and U6410 (N_6410,N_5461,N_5642);
nand U6411 (N_6411,N_5576,N_5390);
nand U6412 (N_6412,N_5587,N_5688);
xnor U6413 (N_6413,N_5529,N_5146);
nand U6414 (N_6414,N_5468,N_5954);
xnor U6415 (N_6415,N_5059,N_5374);
and U6416 (N_6416,N_5421,N_5719);
nor U6417 (N_6417,N_5126,N_5525);
xor U6418 (N_6418,N_5681,N_5721);
nor U6419 (N_6419,N_5494,N_5125);
or U6420 (N_6420,N_5155,N_5220);
nor U6421 (N_6421,N_5632,N_5999);
or U6422 (N_6422,N_5382,N_5886);
nand U6423 (N_6423,N_5898,N_5418);
and U6424 (N_6424,N_5470,N_5647);
nor U6425 (N_6425,N_5724,N_5831);
nor U6426 (N_6426,N_5081,N_5408);
nor U6427 (N_6427,N_5197,N_5564);
nand U6428 (N_6428,N_5308,N_5311);
and U6429 (N_6429,N_5434,N_5454);
nor U6430 (N_6430,N_5910,N_5594);
or U6431 (N_6431,N_5065,N_5336);
nor U6432 (N_6432,N_5670,N_5207);
and U6433 (N_6433,N_5064,N_5446);
and U6434 (N_6434,N_5504,N_5289);
nor U6435 (N_6435,N_5790,N_5830);
or U6436 (N_6436,N_5045,N_5292);
or U6437 (N_6437,N_5068,N_5058);
and U6438 (N_6438,N_5082,N_5266);
xnor U6439 (N_6439,N_5490,N_5934);
nand U6440 (N_6440,N_5042,N_5053);
xnor U6441 (N_6441,N_5708,N_5250);
xnor U6442 (N_6442,N_5194,N_5443);
or U6443 (N_6443,N_5836,N_5415);
or U6444 (N_6444,N_5597,N_5595);
and U6445 (N_6445,N_5679,N_5435);
or U6446 (N_6446,N_5373,N_5862);
xnor U6447 (N_6447,N_5214,N_5835);
xnor U6448 (N_6448,N_5002,N_5198);
nor U6449 (N_6449,N_5348,N_5866);
nand U6450 (N_6450,N_5499,N_5936);
nand U6451 (N_6451,N_5863,N_5933);
nand U6452 (N_6452,N_5040,N_5626);
xnor U6453 (N_6453,N_5514,N_5223);
and U6454 (N_6454,N_5583,N_5063);
nand U6455 (N_6455,N_5843,N_5101);
and U6456 (N_6456,N_5158,N_5737);
xnor U6457 (N_6457,N_5274,N_5178);
nand U6458 (N_6458,N_5326,N_5811);
xor U6459 (N_6459,N_5718,N_5275);
nor U6460 (N_6460,N_5295,N_5789);
xnor U6461 (N_6461,N_5422,N_5607);
nor U6462 (N_6462,N_5206,N_5052);
nand U6463 (N_6463,N_5948,N_5129);
xnor U6464 (N_6464,N_5993,N_5216);
nand U6465 (N_6465,N_5196,N_5136);
and U6466 (N_6466,N_5840,N_5046);
nand U6467 (N_6467,N_5516,N_5644);
or U6468 (N_6468,N_5566,N_5096);
nand U6469 (N_6469,N_5746,N_5755);
nand U6470 (N_6470,N_5660,N_5646);
or U6471 (N_6471,N_5720,N_5329);
or U6472 (N_6472,N_5465,N_5405);
and U6473 (N_6473,N_5492,N_5887);
nor U6474 (N_6474,N_5291,N_5006);
nor U6475 (N_6475,N_5567,N_5321);
and U6476 (N_6476,N_5323,N_5778);
nand U6477 (N_6477,N_5851,N_5234);
and U6478 (N_6478,N_5095,N_5599);
or U6479 (N_6479,N_5174,N_5431);
or U6480 (N_6480,N_5456,N_5402);
xnor U6481 (N_6481,N_5537,N_5070);
nand U6482 (N_6482,N_5221,N_5780);
nand U6483 (N_6483,N_5299,N_5711);
xor U6484 (N_6484,N_5073,N_5810);
nand U6485 (N_6485,N_5675,N_5200);
nor U6486 (N_6486,N_5130,N_5628);
xnor U6487 (N_6487,N_5906,N_5744);
nor U6488 (N_6488,N_5695,N_5462);
nor U6489 (N_6489,N_5610,N_5546);
nand U6490 (N_6490,N_5572,N_5319);
nand U6491 (N_6491,N_5847,N_5532);
nand U6492 (N_6492,N_5941,N_5515);
nand U6493 (N_6493,N_5294,N_5551);
and U6494 (N_6494,N_5837,N_5629);
nor U6495 (N_6495,N_5785,N_5919);
or U6496 (N_6496,N_5692,N_5467);
nand U6497 (N_6497,N_5165,N_5437);
and U6498 (N_6498,N_5911,N_5320);
and U6499 (N_6499,N_5731,N_5481);
nand U6500 (N_6500,N_5415,N_5642);
or U6501 (N_6501,N_5878,N_5891);
xnor U6502 (N_6502,N_5286,N_5518);
and U6503 (N_6503,N_5509,N_5635);
nor U6504 (N_6504,N_5644,N_5359);
nor U6505 (N_6505,N_5525,N_5924);
nor U6506 (N_6506,N_5623,N_5348);
nor U6507 (N_6507,N_5076,N_5373);
nor U6508 (N_6508,N_5005,N_5350);
nand U6509 (N_6509,N_5482,N_5185);
xor U6510 (N_6510,N_5445,N_5089);
or U6511 (N_6511,N_5198,N_5098);
nor U6512 (N_6512,N_5219,N_5836);
or U6513 (N_6513,N_5399,N_5819);
nor U6514 (N_6514,N_5442,N_5712);
and U6515 (N_6515,N_5476,N_5712);
and U6516 (N_6516,N_5673,N_5903);
xnor U6517 (N_6517,N_5493,N_5940);
nor U6518 (N_6518,N_5727,N_5473);
nor U6519 (N_6519,N_5461,N_5152);
nand U6520 (N_6520,N_5892,N_5211);
and U6521 (N_6521,N_5002,N_5216);
xnor U6522 (N_6522,N_5340,N_5336);
nor U6523 (N_6523,N_5381,N_5166);
or U6524 (N_6524,N_5651,N_5418);
nor U6525 (N_6525,N_5423,N_5982);
and U6526 (N_6526,N_5574,N_5442);
or U6527 (N_6527,N_5693,N_5751);
nor U6528 (N_6528,N_5936,N_5430);
nand U6529 (N_6529,N_5005,N_5384);
and U6530 (N_6530,N_5078,N_5090);
xor U6531 (N_6531,N_5527,N_5805);
nand U6532 (N_6532,N_5484,N_5950);
nor U6533 (N_6533,N_5276,N_5033);
nor U6534 (N_6534,N_5753,N_5332);
nor U6535 (N_6535,N_5376,N_5027);
nor U6536 (N_6536,N_5070,N_5113);
and U6537 (N_6537,N_5577,N_5189);
nand U6538 (N_6538,N_5846,N_5298);
xor U6539 (N_6539,N_5655,N_5790);
or U6540 (N_6540,N_5917,N_5538);
nand U6541 (N_6541,N_5465,N_5835);
and U6542 (N_6542,N_5560,N_5404);
and U6543 (N_6543,N_5199,N_5297);
and U6544 (N_6544,N_5312,N_5688);
xnor U6545 (N_6545,N_5304,N_5990);
nand U6546 (N_6546,N_5015,N_5704);
or U6547 (N_6547,N_5684,N_5861);
or U6548 (N_6548,N_5979,N_5615);
xor U6549 (N_6549,N_5514,N_5866);
or U6550 (N_6550,N_5060,N_5944);
or U6551 (N_6551,N_5712,N_5031);
or U6552 (N_6552,N_5153,N_5724);
xnor U6553 (N_6553,N_5448,N_5272);
or U6554 (N_6554,N_5104,N_5759);
or U6555 (N_6555,N_5390,N_5809);
nor U6556 (N_6556,N_5253,N_5891);
or U6557 (N_6557,N_5823,N_5593);
or U6558 (N_6558,N_5675,N_5165);
nand U6559 (N_6559,N_5109,N_5198);
nand U6560 (N_6560,N_5156,N_5161);
and U6561 (N_6561,N_5351,N_5679);
or U6562 (N_6562,N_5429,N_5313);
nor U6563 (N_6563,N_5894,N_5183);
or U6564 (N_6564,N_5747,N_5686);
nand U6565 (N_6565,N_5061,N_5187);
and U6566 (N_6566,N_5408,N_5235);
nand U6567 (N_6567,N_5528,N_5560);
and U6568 (N_6568,N_5632,N_5394);
nor U6569 (N_6569,N_5374,N_5873);
xnor U6570 (N_6570,N_5886,N_5884);
nor U6571 (N_6571,N_5158,N_5942);
and U6572 (N_6572,N_5677,N_5033);
or U6573 (N_6573,N_5104,N_5090);
or U6574 (N_6574,N_5751,N_5859);
nand U6575 (N_6575,N_5216,N_5266);
nand U6576 (N_6576,N_5397,N_5002);
nor U6577 (N_6577,N_5875,N_5804);
and U6578 (N_6578,N_5650,N_5528);
nand U6579 (N_6579,N_5705,N_5691);
or U6580 (N_6580,N_5240,N_5278);
or U6581 (N_6581,N_5650,N_5215);
xor U6582 (N_6582,N_5811,N_5678);
nand U6583 (N_6583,N_5767,N_5806);
or U6584 (N_6584,N_5130,N_5738);
and U6585 (N_6585,N_5178,N_5561);
or U6586 (N_6586,N_5867,N_5823);
nand U6587 (N_6587,N_5103,N_5956);
nand U6588 (N_6588,N_5452,N_5082);
and U6589 (N_6589,N_5968,N_5404);
or U6590 (N_6590,N_5393,N_5405);
xor U6591 (N_6591,N_5088,N_5423);
nand U6592 (N_6592,N_5518,N_5370);
nand U6593 (N_6593,N_5599,N_5048);
and U6594 (N_6594,N_5510,N_5744);
nand U6595 (N_6595,N_5133,N_5457);
or U6596 (N_6596,N_5496,N_5939);
nor U6597 (N_6597,N_5698,N_5019);
or U6598 (N_6598,N_5840,N_5394);
xnor U6599 (N_6599,N_5047,N_5100);
or U6600 (N_6600,N_5270,N_5174);
nand U6601 (N_6601,N_5105,N_5670);
nand U6602 (N_6602,N_5106,N_5319);
nor U6603 (N_6603,N_5507,N_5684);
xor U6604 (N_6604,N_5404,N_5849);
nor U6605 (N_6605,N_5942,N_5672);
nor U6606 (N_6606,N_5952,N_5815);
nand U6607 (N_6607,N_5519,N_5900);
or U6608 (N_6608,N_5497,N_5144);
and U6609 (N_6609,N_5012,N_5144);
or U6610 (N_6610,N_5451,N_5822);
xor U6611 (N_6611,N_5041,N_5873);
xnor U6612 (N_6612,N_5832,N_5826);
and U6613 (N_6613,N_5392,N_5636);
nor U6614 (N_6614,N_5852,N_5599);
or U6615 (N_6615,N_5829,N_5389);
or U6616 (N_6616,N_5439,N_5922);
and U6617 (N_6617,N_5743,N_5765);
and U6618 (N_6618,N_5062,N_5845);
xor U6619 (N_6619,N_5439,N_5825);
and U6620 (N_6620,N_5870,N_5653);
xnor U6621 (N_6621,N_5665,N_5021);
nand U6622 (N_6622,N_5154,N_5859);
nor U6623 (N_6623,N_5539,N_5049);
nand U6624 (N_6624,N_5632,N_5551);
or U6625 (N_6625,N_5406,N_5140);
and U6626 (N_6626,N_5448,N_5444);
nand U6627 (N_6627,N_5431,N_5581);
or U6628 (N_6628,N_5356,N_5180);
nor U6629 (N_6629,N_5935,N_5819);
or U6630 (N_6630,N_5533,N_5703);
and U6631 (N_6631,N_5632,N_5650);
xnor U6632 (N_6632,N_5852,N_5822);
or U6633 (N_6633,N_5289,N_5781);
and U6634 (N_6634,N_5929,N_5649);
xor U6635 (N_6635,N_5367,N_5178);
and U6636 (N_6636,N_5190,N_5523);
xor U6637 (N_6637,N_5358,N_5832);
xor U6638 (N_6638,N_5672,N_5759);
xor U6639 (N_6639,N_5927,N_5801);
and U6640 (N_6640,N_5899,N_5698);
and U6641 (N_6641,N_5528,N_5036);
nand U6642 (N_6642,N_5195,N_5875);
or U6643 (N_6643,N_5349,N_5963);
and U6644 (N_6644,N_5011,N_5889);
nand U6645 (N_6645,N_5698,N_5286);
nor U6646 (N_6646,N_5200,N_5436);
xnor U6647 (N_6647,N_5094,N_5906);
xnor U6648 (N_6648,N_5682,N_5756);
or U6649 (N_6649,N_5083,N_5839);
or U6650 (N_6650,N_5787,N_5321);
nor U6651 (N_6651,N_5228,N_5018);
or U6652 (N_6652,N_5884,N_5142);
or U6653 (N_6653,N_5191,N_5330);
xor U6654 (N_6654,N_5919,N_5333);
nor U6655 (N_6655,N_5050,N_5884);
nand U6656 (N_6656,N_5922,N_5686);
and U6657 (N_6657,N_5908,N_5100);
and U6658 (N_6658,N_5953,N_5982);
xnor U6659 (N_6659,N_5888,N_5830);
xnor U6660 (N_6660,N_5203,N_5379);
and U6661 (N_6661,N_5062,N_5254);
nor U6662 (N_6662,N_5187,N_5210);
or U6663 (N_6663,N_5246,N_5103);
nand U6664 (N_6664,N_5408,N_5358);
nand U6665 (N_6665,N_5702,N_5447);
or U6666 (N_6666,N_5146,N_5007);
nand U6667 (N_6667,N_5924,N_5235);
or U6668 (N_6668,N_5617,N_5018);
nor U6669 (N_6669,N_5832,N_5372);
xnor U6670 (N_6670,N_5766,N_5196);
nor U6671 (N_6671,N_5065,N_5955);
or U6672 (N_6672,N_5251,N_5473);
xnor U6673 (N_6673,N_5810,N_5655);
or U6674 (N_6674,N_5683,N_5416);
xnor U6675 (N_6675,N_5700,N_5336);
or U6676 (N_6676,N_5969,N_5842);
nand U6677 (N_6677,N_5330,N_5028);
nand U6678 (N_6678,N_5868,N_5893);
and U6679 (N_6679,N_5659,N_5849);
or U6680 (N_6680,N_5519,N_5374);
or U6681 (N_6681,N_5882,N_5516);
nand U6682 (N_6682,N_5198,N_5405);
nor U6683 (N_6683,N_5813,N_5850);
and U6684 (N_6684,N_5628,N_5595);
and U6685 (N_6685,N_5501,N_5652);
or U6686 (N_6686,N_5783,N_5963);
nand U6687 (N_6687,N_5962,N_5012);
xor U6688 (N_6688,N_5440,N_5365);
and U6689 (N_6689,N_5426,N_5974);
xnor U6690 (N_6690,N_5385,N_5049);
and U6691 (N_6691,N_5817,N_5365);
nor U6692 (N_6692,N_5804,N_5393);
nor U6693 (N_6693,N_5187,N_5620);
or U6694 (N_6694,N_5961,N_5372);
and U6695 (N_6695,N_5026,N_5402);
and U6696 (N_6696,N_5603,N_5813);
nand U6697 (N_6697,N_5409,N_5440);
nand U6698 (N_6698,N_5286,N_5784);
or U6699 (N_6699,N_5826,N_5657);
nor U6700 (N_6700,N_5713,N_5946);
xnor U6701 (N_6701,N_5017,N_5846);
nor U6702 (N_6702,N_5926,N_5312);
nand U6703 (N_6703,N_5155,N_5034);
nor U6704 (N_6704,N_5343,N_5518);
nand U6705 (N_6705,N_5961,N_5258);
nand U6706 (N_6706,N_5832,N_5549);
nor U6707 (N_6707,N_5252,N_5671);
xor U6708 (N_6708,N_5126,N_5009);
nand U6709 (N_6709,N_5570,N_5606);
or U6710 (N_6710,N_5942,N_5606);
or U6711 (N_6711,N_5207,N_5609);
and U6712 (N_6712,N_5101,N_5733);
nor U6713 (N_6713,N_5870,N_5405);
nand U6714 (N_6714,N_5313,N_5757);
xor U6715 (N_6715,N_5031,N_5183);
nand U6716 (N_6716,N_5866,N_5117);
nand U6717 (N_6717,N_5212,N_5699);
or U6718 (N_6718,N_5921,N_5939);
nand U6719 (N_6719,N_5674,N_5572);
or U6720 (N_6720,N_5761,N_5793);
or U6721 (N_6721,N_5515,N_5287);
xor U6722 (N_6722,N_5300,N_5685);
xnor U6723 (N_6723,N_5555,N_5094);
xor U6724 (N_6724,N_5692,N_5610);
xor U6725 (N_6725,N_5967,N_5448);
nand U6726 (N_6726,N_5431,N_5309);
xnor U6727 (N_6727,N_5886,N_5656);
and U6728 (N_6728,N_5038,N_5908);
and U6729 (N_6729,N_5710,N_5043);
and U6730 (N_6730,N_5486,N_5852);
xor U6731 (N_6731,N_5119,N_5228);
nand U6732 (N_6732,N_5212,N_5957);
nor U6733 (N_6733,N_5490,N_5544);
nor U6734 (N_6734,N_5932,N_5880);
nand U6735 (N_6735,N_5975,N_5925);
nor U6736 (N_6736,N_5961,N_5166);
nor U6737 (N_6737,N_5567,N_5280);
or U6738 (N_6738,N_5334,N_5923);
and U6739 (N_6739,N_5591,N_5519);
or U6740 (N_6740,N_5449,N_5888);
or U6741 (N_6741,N_5918,N_5805);
or U6742 (N_6742,N_5658,N_5937);
and U6743 (N_6743,N_5238,N_5885);
nor U6744 (N_6744,N_5991,N_5937);
nor U6745 (N_6745,N_5944,N_5031);
nor U6746 (N_6746,N_5929,N_5887);
nand U6747 (N_6747,N_5075,N_5620);
nor U6748 (N_6748,N_5616,N_5640);
nand U6749 (N_6749,N_5925,N_5206);
nand U6750 (N_6750,N_5741,N_5375);
or U6751 (N_6751,N_5582,N_5385);
or U6752 (N_6752,N_5222,N_5904);
or U6753 (N_6753,N_5850,N_5174);
and U6754 (N_6754,N_5660,N_5307);
nand U6755 (N_6755,N_5068,N_5623);
nand U6756 (N_6756,N_5949,N_5339);
or U6757 (N_6757,N_5192,N_5650);
xnor U6758 (N_6758,N_5125,N_5046);
and U6759 (N_6759,N_5362,N_5294);
nand U6760 (N_6760,N_5737,N_5544);
nand U6761 (N_6761,N_5788,N_5770);
nand U6762 (N_6762,N_5387,N_5235);
or U6763 (N_6763,N_5913,N_5284);
or U6764 (N_6764,N_5627,N_5762);
nor U6765 (N_6765,N_5954,N_5448);
nand U6766 (N_6766,N_5032,N_5110);
xnor U6767 (N_6767,N_5437,N_5711);
nor U6768 (N_6768,N_5666,N_5158);
or U6769 (N_6769,N_5370,N_5664);
nand U6770 (N_6770,N_5354,N_5638);
nand U6771 (N_6771,N_5546,N_5809);
or U6772 (N_6772,N_5687,N_5590);
or U6773 (N_6773,N_5526,N_5979);
and U6774 (N_6774,N_5170,N_5881);
or U6775 (N_6775,N_5346,N_5734);
nor U6776 (N_6776,N_5412,N_5778);
nor U6777 (N_6777,N_5196,N_5571);
and U6778 (N_6778,N_5116,N_5825);
xor U6779 (N_6779,N_5298,N_5892);
xor U6780 (N_6780,N_5868,N_5724);
nor U6781 (N_6781,N_5791,N_5746);
xnor U6782 (N_6782,N_5571,N_5504);
and U6783 (N_6783,N_5182,N_5119);
and U6784 (N_6784,N_5196,N_5373);
xor U6785 (N_6785,N_5016,N_5039);
xnor U6786 (N_6786,N_5181,N_5899);
or U6787 (N_6787,N_5499,N_5538);
nand U6788 (N_6788,N_5249,N_5422);
xnor U6789 (N_6789,N_5728,N_5550);
nor U6790 (N_6790,N_5186,N_5863);
nor U6791 (N_6791,N_5823,N_5329);
xnor U6792 (N_6792,N_5598,N_5005);
and U6793 (N_6793,N_5885,N_5739);
nand U6794 (N_6794,N_5770,N_5772);
and U6795 (N_6795,N_5077,N_5837);
or U6796 (N_6796,N_5972,N_5295);
or U6797 (N_6797,N_5759,N_5842);
nor U6798 (N_6798,N_5286,N_5556);
nor U6799 (N_6799,N_5018,N_5692);
or U6800 (N_6800,N_5886,N_5345);
nor U6801 (N_6801,N_5144,N_5836);
and U6802 (N_6802,N_5436,N_5250);
or U6803 (N_6803,N_5686,N_5524);
nor U6804 (N_6804,N_5538,N_5206);
nor U6805 (N_6805,N_5419,N_5216);
and U6806 (N_6806,N_5747,N_5644);
nor U6807 (N_6807,N_5788,N_5988);
nand U6808 (N_6808,N_5942,N_5159);
nand U6809 (N_6809,N_5974,N_5563);
xnor U6810 (N_6810,N_5812,N_5336);
or U6811 (N_6811,N_5000,N_5255);
or U6812 (N_6812,N_5577,N_5751);
nand U6813 (N_6813,N_5024,N_5011);
or U6814 (N_6814,N_5732,N_5465);
and U6815 (N_6815,N_5625,N_5007);
or U6816 (N_6816,N_5151,N_5685);
nor U6817 (N_6817,N_5468,N_5885);
nor U6818 (N_6818,N_5959,N_5660);
or U6819 (N_6819,N_5474,N_5786);
or U6820 (N_6820,N_5977,N_5858);
or U6821 (N_6821,N_5956,N_5425);
and U6822 (N_6822,N_5528,N_5781);
nand U6823 (N_6823,N_5528,N_5195);
nor U6824 (N_6824,N_5041,N_5535);
or U6825 (N_6825,N_5292,N_5787);
nor U6826 (N_6826,N_5789,N_5369);
and U6827 (N_6827,N_5575,N_5243);
or U6828 (N_6828,N_5397,N_5194);
and U6829 (N_6829,N_5553,N_5325);
and U6830 (N_6830,N_5108,N_5556);
nand U6831 (N_6831,N_5399,N_5463);
or U6832 (N_6832,N_5474,N_5271);
xnor U6833 (N_6833,N_5108,N_5898);
xor U6834 (N_6834,N_5876,N_5165);
or U6835 (N_6835,N_5001,N_5577);
and U6836 (N_6836,N_5095,N_5629);
nor U6837 (N_6837,N_5816,N_5013);
nor U6838 (N_6838,N_5194,N_5286);
xor U6839 (N_6839,N_5382,N_5455);
nor U6840 (N_6840,N_5727,N_5809);
and U6841 (N_6841,N_5616,N_5503);
nand U6842 (N_6842,N_5240,N_5609);
nor U6843 (N_6843,N_5213,N_5804);
nor U6844 (N_6844,N_5458,N_5762);
and U6845 (N_6845,N_5817,N_5711);
xor U6846 (N_6846,N_5886,N_5102);
xnor U6847 (N_6847,N_5104,N_5628);
nor U6848 (N_6848,N_5068,N_5236);
nor U6849 (N_6849,N_5031,N_5170);
xor U6850 (N_6850,N_5082,N_5681);
and U6851 (N_6851,N_5771,N_5837);
nand U6852 (N_6852,N_5896,N_5164);
or U6853 (N_6853,N_5169,N_5145);
nor U6854 (N_6854,N_5345,N_5650);
or U6855 (N_6855,N_5301,N_5527);
xor U6856 (N_6856,N_5930,N_5555);
nand U6857 (N_6857,N_5151,N_5171);
nor U6858 (N_6858,N_5264,N_5835);
and U6859 (N_6859,N_5653,N_5366);
and U6860 (N_6860,N_5427,N_5547);
and U6861 (N_6861,N_5227,N_5441);
or U6862 (N_6862,N_5133,N_5094);
and U6863 (N_6863,N_5214,N_5307);
nand U6864 (N_6864,N_5809,N_5085);
nand U6865 (N_6865,N_5637,N_5968);
nand U6866 (N_6866,N_5426,N_5140);
nand U6867 (N_6867,N_5662,N_5801);
and U6868 (N_6868,N_5278,N_5803);
nor U6869 (N_6869,N_5926,N_5784);
or U6870 (N_6870,N_5146,N_5306);
and U6871 (N_6871,N_5406,N_5911);
and U6872 (N_6872,N_5352,N_5941);
nand U6873 (N_6873,N_5568,N_5488);
and U6874 (N_6874,N_5690,N_5784);
nand U6875 (N_6875,N_5001,N_5799);
nor U6876 (N_6876,N_5858,N_5642);
xor U6877 (N_6877,N_5296,N_5909);
xor U6878 (N_6878,N_5829,N_5162);
nand U6879 (N_6879,N_5763,N_5668);
and U6880 (N_6880,N_5974,N_5620);
nor U6881 (N_6881,N_5160,N_5991);
xnor U6882 (N_6882,N_5286,N_5625);
xnor U6883 (N_6883,N_5429,N_5395);
nor U6884 (N_6884,N_5129,N_5234);
and U6885 (N_6885,N_5169,N_5120);
nor U6886 (N_6886,N_5977,N_5359);
xor U6887 (N_6887,N_5255,N_5217);
nor U6888 (N_6888,N_5972,N_5393);
nand U6889 (N_6889,N_5605,N_5003);
or U6890 (N_6890,N_5411,N_5721);
nand U6891 (N_6891,N_5021,N_5810);
and U6892 (N_6892,N_5254,N_5566);
nor U6893 (N_6893,N_5064,N_5479);
or U6894 (N_6894,N_5499,N_5858);
nand U6895 (N_6895,N_5932,N_5758);
xnor U6896 (N_6896,N_5608,N_5960);
and U6897 (N_6897,N_5644,N_5776);
or U6898 (N_6898,N_5513,N_5478);
xnor U6899 (N_6899,N_5519,N_5285);
nand U6900 (N_6900,N_5316,N_5640);
xnor U6901 (N_6901,N_5944,N_5347);
xnor U6902 (N_6902,N_5224,N_5401);
xnor U6903 (N_6903,N_5999,N_5516);
and U6904 (N_6904,N_5163,N_5539);
xnor U6905 (N_6905,N_5262,N_5104);
nand U6906 (N_6906,N_5963,N_5009);
nor U6907 (N_6907,N_5401,N_5598);
xnor U6908 (N_6908,N_5427,N_5841);
nor U6909 (N_6909,N_5889,N_5776);
xor U6910 (N_6910,N_5814,N_5676);
or U6911 (N_6911,N_5296,N_5786);
xor U6912 (N_6912,N_5394,N_5323);
nand U6913 (N_6913,N_5602,N_5309);
nand U6914 (N_6914,N_5891,N_5465);
or U6915 (N_6915,N_5516,N_5817);
xnor U6916 (N_6916,N_5117,N_5867);
nor U6917 (N_6917,N_5666,N_5597);
nor U6918 (N_6918,N_5358,N_5082);
nor U6919 (N_6919,N_5395,N_5413);
and U6920 (N_6920,N_5870,N_5967);
xnor U6921 (N_6921,N_5772,N_5039);
or U6922 (N_6922,N_5663,N_5186);
xnor U6923 (N_6923,N_5410,N_5605);
and U6924 (N_6924,N_5789,N_5892);
xnor U6925 (N_6925,N_5753,N_5468);
nand U6926 (N_6926,N_5677,N_5488);
or U6927 (N_6927,N_5532,N_5977);
nor U6928 (N_6928,N_5699,N_5912);
and U6929 (N_6929,N_5658,N_5496);
nor U6930 (N_6930,N_5502,N_5140);
and U6931 (N_6931,N_5508,N_5400);
nor U6932 (N_6932,N_5620,N_5041);
nand U6933 (N_6933,N_5222,N_5121);
or U6934 (N_6934,N_5057,N_5533);
and U6935 (N_6935,N_5365,N_5205);
nor U6936 (N_6936,N_5148,N_5843);
and U6937 (N_6937,N_5786,N_5480);
nand U6938 (N_6938,N_5747,N_5071);
nand U6939 (N_6939,N_5693,N_5007);
xor U6940 (N_6940,N_5739,N_5573);
and U6941 (N_6941,N_5327,N_5899);
or U6942 (N_6942,N_5029,N_5227);
or U6943 (N_6943,N_5434,N_5681);
or U6944 (N_6944,N_5056,N_5351);
nor U6945 (N_6945,N_5213,N_5756);
and U6946 (N_6946,N_5525,N_5034);
and U6947 (N_6947,N_5918,N_5820);
and U6948 (N_6948,N_5143,N_5721);
nand U6949 (N_6949,N_5843,N_5655);
or U6950 (N_6950,N_5313,N_5560);
nor U6951 (N_6951,N_5543,N_5933);
or U6952 (N_6952,N_5300,N_5947);
nor U6953 (N_6953,N_5575,N_5747);
and U6954 (N_6954,N_5711,N_5788);
xnor U6955 (N_6955,N_5977,N_5516);
nand U6956 (N_6956,N_5868,N_5338);
or U6957 (N_6957,N_5062,N_5097);
and U6958 (N_6958,N_5899,N_5586);
nor U6959 (N_6959,N_5247,N_5242);
xor U6960 (N_6960,N_5964,N_5759);
and U6961 (N_6961,N_5512,N_5706);
nor U6962 (N_6962,N_5375,N_5390);
xnor U6963 (N_6963,N_5420,N_5306);
and U6964 (N_6964,N_5195,N_5383);
nand U6965 (N_6965,N_5251,N_5152);
and U6966 (N_6966,N_5923,N_5784);
and U6967 (N_6967,N_5403,N_5834);
nor U6968 (N_6968,N_5611,N_5823);
or U6969 (N_6969,N_5747,N_5051);
xnor U6970 (N_6970,N_5081,N_5968);
or U6971 (N_6971,N_5815,N_5251);
nand U6972 (N_6972,N_5100,N_5986);
xnor U6973 (N_6973,N_5556,N_5478);
nor U6974 (N_6974,N_5425,N_5080);
nand U6975 (N_6975,N_5114,N_5732);
and U6976 (N_6976,N_5319,N_5024);
and U6977 (N_6977,N_5894,N_5181);
and U6978 (N_6978,N_5165,N_5513);
and U6979 (N_6979,N_5569,N_5165);
nand U6980 (N_6980,N_5271,N_5030);
and U6981 (N_6981,N_5592,N_5989);
nand U6982 (N_6982,N_5508,N_5192);
nand U6983 (N_6983,N_5265,N_5725);
nand U6984 (N_6984,N_5206,N_5796);
nor U6985 (N_6985,N_5271,N_5195);
nor U6986 (N_6986,N_5849,N_5215);
and U6987 (N_6987,N_5521,N_5375);
nand U6988 (N_6988,N_5929,N_5504);
xor U6989 (N_6989,N_5924,N_5089);
xor U6990 (N_6990,N_5711,N_5204);
and U6991 (N_6991,N_5491,N_5562);
or U6992 (N_6992,N_5086,N_5380);
nand U6993 (N_6993,N_5597,N_5968);
or U6994 (N_6994,N_5587,N_5205);
or U6995 (N_6995,N_5959,N_5133);
and U6996 (N_6996,N_5266,N_5084);
and U6997 (N_6997,N_5335,N_5070);
nand U6998 (N_6998,N_5695,N_5327);
nand U6999 (N_6999,N_5430,N_5768);
xnor U7000 (N_7000,N_6385,N_6227);
nand U7001 (N_7001,N_6536,N_6180);
and U7002 (N_7002,N_6110,N_6029);
and U7003 (N_7003,N_6311,N_6562);
or U7004 (N_7004,N_6132,N_6326);
nand U7005 (N_7005,N_6465,N_6701);
and U7006 (N_7006,N_6447,N_6048);
or U7007 (N_7007,N_6964,N_6357);
and U7008 (N_7008,N_6542,N_6533);
or U7009 (N_7009,N_6984,N_6639);
nor U7010 (N_7010,N_6320,N_6990);
xnor U7011 (N_7011,N_6500,N_6787);
or U7012 (N_7012,N_6561,N_6010);
xor U7013 (N_7013,N_6345,N_6987);
and U7014 (N_7014,N_6434,N_6036);
and U7015 (N_7015,N_6379,N_6605);
and U7016 (N_7016,N_6023,N_6479);
nor U7017 (N_7017,N_6680,N_6633);
and U7018 (N_7018,N_6150,N_6917);
or U7019 (N_7019,N_6943,N_6052);
nor U7020 (N_7020,N_6902,N_6773);
or U7021 (N_7021,N_6386,N_6769);
nand U7022 (N_7022,N_6178,N_6470);
and U7023 (N_7023,N_6962,N_6521);
nand U7024 (N_7024,N_6634,N_6472);
nor U7025 (N_7025,N_6147,N_6926);
xnor U7026 (N_7026,N_6328,N_6684);
or U7027 (N_7027,N_6154,N_6976);
xor U7028 (N_7028,N_6181,N_6160);
xor U7029 (N_7029,N_6547,N_6495);
xnor U7030 (N_7030,N_6259,N_6431);
and U7031 (N_7031,N_6724,N_6486);
xor U7032 (N_7032,N_6318,N_6281);
and U7033 (N_7033,N_6493,N_6941);
or U7034 (N_7034,N_6515,N_6854);
nand U7035 (N_7035,N_6895,N_6784);
nor U7036 (N_7036,N_6645,N_6407);
or U7037 (N_7037,N_6354,N_6882);
nand U7038 (N_7038,N_6835,N_6912);
nand U7039 (N_7039,N_6372,N_6143);
nand U7040 (N_7040,N_6254,N_6793);
and U7041 (N_7041,N_6878,N_6919);
nor U7042 (N_7042,N_6842,N_6316);
or U7043 (N_7043,N_6258,N_6846);
nor U7044 (N_7044,N_6122,N_6975);
and U7045 (N_7045,N_6603,N_6828);
or U7046 (N_7046,N_6136,N_6839);
nand U7047 (N_7047,N_6346,N_6757);
and U7048 (N_7048,N_6667,N_6790);
or U7049 (N_7049,N_6806,N_6035);
nor U7050 (N_7050,N_6167,N_6678);
or U7051 (N_7051,N_6795,N_6004);
nand U7052 (N_7052,N_6657,N_6303);
and U7053 (N_7053,N_6522,N_6717);
or U7054 (N_7054,N_6060,N_6568);
and U7055 (N_7055,N_6378,N_6703);
nor U7056 (N_7056,N_6800,N_6451);
and U7057 (N_7057,N_6174,N_6428);
and U7058 (N_7058,N_6856,N_6774);
nor U7059 (N_7059,N_6400,N_6636);
nand U7060 (N_7060,N_6333,N_6435);
or U7061 (N_7061,N_6754,N_6362);
or U7062 (N_7062,N_6766,N_6598);
nor U7063 (N_7063,N_6292,N_6125);
xor U7064 (N_7064,N_6767,N_6492);
or U7065 (N_7065,N_6900,N_6991);
nand U7066 (N_7066,N_6276,N_6686);
nand U7067 (N_7067,N_6802,N_6121);
or U7068 (N_7068,N_6871,N_6692);
and U7069 (N_7069,N_6512,N_6661);
and U7070 (N_7070,N_6954,N_6865);
xor U7071 (N_7071,N_6459,N_6008);
xor U7072 (N_7072,N_6450,N_6245);
nand U7073 (N_7073,N_6716,N_6021);
and U7074 (N_7074,N_6051,N_6261);
xnor U7075 (N_7075,N_6243,N_6709);
and U7076 (N_7076,N_6045,N_6710);
or U7077 (N_7077,N_6898,N_6421);
nand U7078 (N_7078,N_6159,N_6211);
nor U7079 (N_7079,N_6437,N_6705);
xor U7080 (N_7080,N_6874,N_6376);
nand U7081 (N_7081,N_6652,N_6002);
xnor U7082 (N_7082,N_6315,N_6584);
nand U7083 (N_7083,N_6706,N_6507);
nand U7084 (N_7084,N_6455,N_6868);
nand U7085 (N_7085,N_6073,N_6758);
and U7086 (N_7086,N_6108,N_6807);
nand U7087 (N_7087,N_6711,N_6586);
nor U7088 (N_7088,N_6785,N_6949);
or U7089 (N_7089,N_6221,N_6475);
or U7090 (N_7090,N_6393,N_6195);
and U7091 (N_7091,N_6144,N_6877);
nor U7092 (N_7092,N_6454,N_6436);
nor U7093 (N_7093,N_6194,N_6031);
and U7094 (N_7094,N_6323,N_6140);
nor U7095 (N_7095,N_6582,N_6062);
or U7096 (N_7096,N_6197,N_6597);
or U7097 (N_7097,N_6755,N_6216);
xnor U7098 (N_7098,N_6775,N_6129);
nand U7099 (N_7099,N_6752,N_6067);
xnor U7100 (N_7100,N_6336,N_6145);
nor U7101 (N_7101,N_6420,N_6952);
or U7102 (N_7102,N_6084,N_6527);
xor U7103 (N_7103,N_6574,N_6047);
or U7104 (N_7104,N_6079,N_6207);
or U7105 (N_7105,N_6786,N_6370);
nand U7106 (N_7106,N_6511,N_6950);
xnor U7107 (N_7107,N_6443,N_6402);
or U7108 (N_7108,N_6738,N_6074);
or U7109 (N_7109,N_6841,N_6439);
or U7110 (N_7110,N_6630,N_6414);
xnor U7111 (N_7111,N_6904,N_6413);
nand U7112 (N_7112,N_6293,N_6018);
xor U7113 (N_7113,N_6749,N_6737);
and U7114 (N_7114,N_6165,N_6487);
xnor U7115 (N_7115,N_6498,N_6575);
and U7116 (N_7116,N_6938,N_6973);
or U7117 (N_7117,N_6816,N_6914);
nor U7118 (N_7118,N_6302,N_6005);
nor U7119 (N_7119,N_6642,N_6727);
or U7120 (N_7120,N_6388,N_6484);
nor U7121 (N_7121,N_6913,N_6212);
xor U7122 (N_7122,N_6933,N_6595);
and U7123 (N_7123,N_6128,N_6820);
nor U7124 (N_7124,N_6324,N_6344);
nand U7125 (N_7125,N_6761,N_6891);
and U7126 (N_7126,N_6556,N_6702);
nand U7127 (N_7127,N_6291,N_6055);
nor U7128 (N_7128,N_6285,N_6377);
nand U7129 (N_7129,N_6860,N_6552);
nor U7130 (N_7130,N_6011,N_6674);
nor U7131 (N_7131,N_6383,N_6741);
nor U7132 (N_7132,N_6873,N_6744);
and U7133 (N_7133,N_6267,N_6646);
xnor U7134 (N_7134,N_6200,N_6551);
and U7135 (N_7135,N_6229,N_6228);
and U7136 (N_7136,N_6412,N_6573);
or U7137 (N_7137,N_6999,N_6814);
xnor U7138 (N_7138,N_6422,N_6960);
and U7139 (N_7139,N_6763,N_6528);
or U7140 (N_7140,N_6689,N_6957);
and U7141 (N_7141,N_6248,N_6359);
and U7142 (N_7142,N_6695,N_6676);
nor U7143 (N_7143,N_6631,N_6290);
xnor U7144 (N_7144,N_6264,N_6924);
xor U7145 (N_7145,N_6054,N_6635);
and U7146 (N_7146,N_6649,N_6664);
xnor U7147 (N_7147,N_6751,N_6683);
xor U7148 (N_7148,N_6628,N_6650);
nor U7149 (N_7149,N_6825,N_6343);
and U7150 (N_7150,N_6833,N_6007);
or U7151 (N_7151,N_6813,N_6456);
and U7152 (N_7152,N_6809,N_6563);
nor U7153 (N_7153,N_6355,N_6797);
nor U7154 (N_7154,N_6287,N_6395);
nand U7155 (N_7155,N_6672,N_6148);
nand U7156 (N_7156,N_6858,N_6351);
nand U7157 (N_7157,N_6022,N_6946);
or U7158 (N_7158,N_6955,N_6837);
or U7159 (N_7159,N_6064,N_6277);
or U7160 (N_7160,N_6049,N_6843);
nor U7161 (N_7161,N_6516,N_6085);
nand U7162 (N_7162,N_6896,N_6997);
or U7163 (N_7163,N_6930,N_6374);
nor U7164 (N_7164,N_6959,N_6480);
xor U7165 (N_7165,N_6391,N_6998);
nor U7166 (N_7166,N_6546,N_6619);
and U7167 (N_7167,N_6819,N_6305);
and U7168 (N_7168,N_6732,N_6430);
or U7169 (N_7169,N_6131,N_6020);
nor U7170 (N_7170,N_6583,N_6517);
xor U7171 (N_7171,N_6932,N_6916);
and U7172 (N_7172,N_6901,N_6513);
nor U7173 (N_7173,N_6776,N_6219);
or U7174 (N_7174,N_6623,N_6381);
xnor U7175 (N_7175,N_6665,N_6215);
nand U7176 (N_7176,N_6530,N_6153);
nor U7177 (N_7177,N_6698,N_6094);
xnor U7178 (N_7178,N_6101,N_6471);
nand U7179 (N_7179,N_6273,N_6262);
xnor U7180 (N_7180,N_6840,N_6849);
or U7181 (N_7181,N_6935,N_6231);
nand U7182 (N_7182,N_6275,N_6587);
xnor U7183 (N_7183,N_6770,N_6765);
and U7184 (N_7184,N_6453,N_6659);
nand U7185 (N_7185,N_6445,N_6739);
or U7186 (N_7186,N_6030,N_6994);
nand U7187 (N_7187,N_6970,N_6821);
nand U7188 (N_7188,N_6670,N_6756);
nand U7189 (N_7189,N_6884,N_6156);
xor U7190 (N_7190,N_6588,N_6353);
nor U7191 (N_7191,N_6024,N_6832);
nor U7192 (N_7192,N_6151,N_6392);
or U7193 (N_7193,N_6410,N_6899);
nand U7194 (N_7194,N_6114,N_6466);
or U7195 (N_7195,N_6099,N_6923);
xnor U7196 (N_7196,N_6482,N_6988);
xnor U7197 (N_7197,N_6429,N_6349);
nand U7198 (N_7198,N_6585,N_6003);
or U7199 (N_7199,N_6265,N_6685);
and U7200 (N_7200,N_6815,N_6557);
xor U7201 (N_7201,N_6278,N_6523);
nand U7202 (N_7202,N_6508,N_6016);
or U7203 (N_7203,N_6968,N_6851);
nor U7204 (N_7204,N_6170,N_6647);
nand U7205 (N_7205,N_6779,N_6330);
nor U7206 (N_7206,N_6251,N_6506);
xor U7207 (N_7207,N_6071,N_6463);
or U7208 (N_7208,N_6116,N_6892);
xnor U7209 (N_7209,N_6538,N_6284);
nand U7210 (N_7210,N_6720,N_6590);
or U7211 (N_7211,N_6894,N_6643);
and U7212 (N_7212,N_6117,N_6982);
nor U7213 (N_7213,N_6554,N_6539);
xnor U7214 (N_7214,N_6066,N_6390);
xnor U7215 (N_7215,N_6087,N_6308);
and U7216 (N_7216,N_6951,N_6403);
nand U7217 (N_7217,N_6225,N_6387);
xnor U7218 (N_7218,N_6600,N_6577);
nand U7219 (N_7219,N_6166,N_6112);
nand U7220 (N_7220,N_6632,N_6548);
xnor U7221 (N_7221,N_6827,N_6502);
or U7222 (N_7222,N_6416,N_6105);
or U7223 (N_7223,N_6411,N_6995);
nand U7224 (N_7224,N_6476,N_6501);
nor U7225 (N_7225,N_6233,N_6876);
or U7226 (N_7226,N_6905,N_6130);
and U7227 (N_7227,N_6679,N_6468);
or U7228 (N_7228,N_6615,N_6721);
xnor U7229 (N_7229,N_6288,N_6038);
nand U7230 (N_7230,N_6525,N_6505);
xnor U7231 (N_7231,N_6581,N_6338);
or U7232 (N_7232,N_6193,N_6804);
xnor U7233 (N_7233,N_6304,N_6286);
and U7234 (N_7234,N_6782,N_6347);
nor U7235 (N_7235,N_6830,N_6762);
and U7236 (N_7236,N_6618,N_6172);
nor U7237 (N_7237,N_6425,N_6203);
or U7238 (N_7238,N_6253,N_6081);
nor U7239 (N_7239,N_6075,N_6341);
xnor U7240 (N_7240,N_6009,N_6715);
nor U7241 (N_7241,N_6857,N_6558);
nor U7242 (N_7242,N_6818,N_6875);
and U7243 (N_7243,N_6707,N_6969);
or U7244 (N_7244,N_6269,N_6090);
xor U7245 (N_7245,N_6179,N_6747);
nand U7246 (N_7246,N_6983,N_6714);
nand U7247 (N_7247,N_6544,N_6032);
nor U7248 (N_7248,N_6535,N_6545);
nor U7249 (N_7249,N_6423,N_6115);
nor U7250 (N_7250,N_6234,N_6396);
nor U7251 (N_7251,N_6928,N_6307);
nand U7252 (N_7252,N_6602,N_6188);
xnor U7253 (N_7253,N_6593,N_6176);
nor U7254 (N_7254,N_6161,N_6204);
and U7255 (N_7255,N_6006,N_6967);
or U7256 (N_7256,N_6244,N_6072);
nand U7257 (N_7257,N_6549,N_6576);
or U7258 (N_7258,N_6280,N_6726);
nor U7259 (N_7259,N_6268,N_6663);
or U7260 (N_7260,N_6452,N_6373);
nor U7261 (N_7261,N_6367,N_6432);
and U7262 (N_7262,N_6015,N_6838);
xnor U7263 (N_7263,N_6571,N_6137);
or U7264 (N_7264,N_6653,N_6102);
and U7265 (N_7265,N_6237,N_6929);
and U7266 (N_7266,N_6332,N_6191);
nor U7267 (N_7267,N_6164,N_6750);
nand U7268 (N_7268,N_6850,N_6731);
or U7269 (N_7269,N_6728,N_6580);
nor U7270 (N_7270,N_6440,N_6799);
or U7271 (N_7271,N_6599,N_6504);
nand U7272 (N_7272,N_6086,N_6089);
nand U7273 (N_7273,N_6158,N_6266);
nand U7274 (N_7274,N_6570,N_6283);
xnor U7275 (N_7275,N_6666,N_6978);
or U7276 (N_7276,N_6417,N_6907);
or U7277 (N_7277,N_6250,N_6648);
and U7278 (N_7278,N_6668,N_6252);
or U7279 (N_7279,N_6608,N_6339);
nor U7280 (N_7280,N_6397,N_6931);
nor U7281 (N_7281,N_6406,N_6723);
xor U7282 (N_7282,N_6327,N_6862);
or U7283 (N_7283,N_6963,N_6034);
nand U7284 (N_7284,N_6350,N_6936);
or U7285 (N_7285,N_6043,N_6001);
and U7286 (N_7286,N_6469,N_6772);
nor U7287 (N_7287,N_6944,N_6569);
xor U7288 (N_7288,N_6046,N_6342);
or U7289 (N_7289,N_6039,N_6184);
nand U7290 (N_7290,N_6553,N_6824);
or U7291 (N_7291,N_6885,N_6399);
or U7292 (N_7292,N_6753,N_6255);
nand U7293 (N_7293,N_6177,N_6694);
nor U7294 (N_7294,N_6771,N_6699);
and U7295 (N_7295,N_6325,N_6607);
and U7296 (N_7296,N_6524,N_6065);
and U7297 (N_7297,N_6922,N_6514);
or U7298 (N_7298,N_6398,N_6260);
nor U7299 (N_7299,N_6192,N_6272);
and U7300 (N_7300,N_6735,N_6889);
nand U7301 (N_7301,N_6897,N_6915);
xor U7302 (N_7302,N_6295,N_6579);
nand U7303 (N_7303,N_6477,N_6247);
nand U7304 (N_7304,N_6119,N_6503);
and U7305 (N_7305,N_6682,N_6317);
and U7306 (N_7306,N_6358,N_6687);
or U7307 (N_7307,N_6822,N_6171);
xor U7308 (N_7308,N_6314,N_6230);
nor U7309 (N_7309,N_6920,N_6778);
nor U7310 (N_7310,N_6893,N_6058);
nor U7311 (N_7311,N_6209,N_6427);
nor U7312 (N_7312,N_6489,N_6606);
or U7313 (N_7313,N_6263,N_6473);
nor U7314 (N_7314,N_6257,N_6866);
nand U7315 (N_7315,N_6675,N_6214);
nand U7316 (N_7316,N_6133,N_6961);
and U7317 (N_7317,N_6322,N_6578);
or U7318 (N_7318,N_6014,N_6852);
nand U7319 (N_7319,N_6040,N_6887);
nand U7320 (N_7320,N_6220,N_6729);
and U7321 (N_7321,N_6082,N_6104);
or U7322 (N_7322,N_6394,N_6743);
nand U7323 (N_7323,N_6491,N_6296);
nor U7324 (N_7324,N_6168,N_6310);
xnor U7325 (N_7325,N_6939,N_6791);
xor U7326 (N_7326,N_6446,N_6028);
nor U7327 (N_7327,N_6641,N_6061);
or U7328 (N_7328,N_6925,N_6053);
xnor U7329 (N_7329,N_6027,N_6056);
nor U7330 (N_7330,N_6173,N_6796);
nor U7331 (N_7331,N_6945,N_6488);
xor U7332 (N_7332,N_6369,N_6444);
nor U7333 (N_7333,N_6458,N_6077);
nor U7334 (N_7334,N_6235,N_6654);
xnor U7335 (N_7335,N_6669,N_6989);
nor U7336 (N_7336,N_6190,N_6033);
or U7337 (N_7337,N_6748,N_6518);
or U7338 (N_7338,N_6497,N_6540);
and U7339 (N_7339,N_6240,N_6224);
xnor U7340 (N_7340,N_6000,N_6134);
and U7341 (N_7341,N_6025,N_6478);
nand U7342 (N_7342,N_6927,N_6113);
xnor U7343 (N_7343,N_6911,N_6496);
xor U7344 (N_7344,N_6356,N_6213);
nor U7345 (N_7345,N_6823,N_6185);
nor U7346 (N_7346,N_6651,N_6609);
and U7347 (N_7347,N_6098,N_6270);
or U7348 (N_7348,N_6481,N_6906);
nand U7349 (N_7349,N_6050,N_6848);
nand U7350 (N_7350,N_6713,N_6965);
nor U7351 (N_7351,N_6734,N_6124);
nand U7352 (N_7352,N_6853,N_6801);
and U7353 (N_7353,N_6937,N_6910);
nand U7354 (N_7354,N_6974,N_6183);
nand U7355 (N_7355,N_6218,N_6780);
or U7356 (N_7356,N_6198,N_6543);
xnor U7357 (N_7357,N_6870,N_6106);
nor U7358 (N_7358,N_6604,N_6205);
or U7359 (N_7359,N_6629,N_6520);
nor U7360 (N_7360,N_6348,N_6861);
or U7361 (N_7361,N_6594,N_6360);
nand U7362 (N_7362,N_6375,N_6321);
nand U7363 (N_7363,N_6109,N_6120);
nor U7364 (N_7364,N_6196,N_6733);
and U7365 (N_7365,N_6187,N_6312);
xnor U7366 (N_7366,N_6746,N_6097);
xnor U7367 (N_7367,N_6693,N_6217);
or U7368 (N_7368,N_6986,N_6942);
nor U7369 (N_7369,N_6494,N_6026);
nor U7370 (N_7370,N_6810,N_6289);
or U7371 (N_7371,N_6610,N_6340);
or U7372 (N_7372,N_6621,N_6155);
nand U7373 (N_7373,N_6279,N_6844);
and U7374 (N_7374,N_6637,N_6464);
nor U7375 (N_7375,N_6163,N_6953);
nor U7376 (N_7376,N_6918,N_6335);
xor U7377 (N_7377,N_6592,N_6474);
and U7378 (N_7378,N_6088,N_6589);
or U7379 (N_7379,N_6123,N_6100);
or U7380 (N_7380,N_6169,N_6981);
xnor U7381 (N_7381,N_6834,N_6091);
or U7382 (N_7382,N_6627,N_6696);
nand U7383 (N_7383,N_6566,N_6222);
and U7384 (N_7384,N_6700,N_6798);
and U7385 (N_7385,N_6424,N_6677);
nor U7386 (N_7386,N_6712,N_6719);
and U7387 (N_7387,N_6118,N_6760);
and U7388 (N_7388,N_6940,N_6206);
nand U7389 (N_7389,N_6808,N_6111);
or U7390 (N_7390,N_6068,N_6658);
nor U7391 (N_7391,N_6811,N_6859);
or U7392 (N_7392,N_6408,N_6805);
and U7393 (N_7393,N_6282,N_6363);
nand U7394 (N_7394,N_6881,N_6980);
and U7395 (N_7395,N_6238,N_6826);
and U7396 (N_7396,N_6223,N_6688);
xnor U7397 (N_7397,N_6294,N_6236);
nor U7398 (N_7398,N_6186,N_6175);
nand U7399 (N_7399,N_6829,N_6534);
xnor U7400 (N_7400,N_6956,N_6418);
or U7401 (N_7401,N_6442,N_6368);
nor U7402 (N_7402,N_6037,N_6135);
nor U7403 (N_7403,N_6300,N_6704);
nand U7404 (N_7404,N_6781,N_6141);
or U7405 (N_7405,N_6909,N_6298);
nand U7406 (N_7406,N_6485,N_6127);
or U7407 (N_7407,N_6958,N_6382);
and U7408 (N_7408,N_6380,N_6596);
or U7409 (N_7409,N_6162,N_6948);
nor U7410 (N_7410,N_6888,N_6880);
and U7411 (N_7411,N_6626,N_6872);
or U7412 (N_7412,N_6934,N_6541);
or U7413 (N_7413,N_6438,N_6836);
and U7414 (N_7414,N_6662,N_6992);
or U7415 (N_7415,N_6070,N_6483);
or U7416 (N_7416,N_6519,N_6979);
or U7417 (N_7417,N_6625,N_6673);
xor U7418 (N_7418,N_6457,N_6655);
nand U7419 (N_7419,N_6242,N_6564);
or U7420 (N_7420,N_6297,N_6745);
xor U7421 (N_7421,N_6201,N_6966);
nand U7422 (N_7422,N_6433,N_6817);
and U7423 (N_7423,N_6057,N_6644);
or U7424 (N_7424,N_6241,N_6803);
nand U7425 (N_7425,N_6409,N_6921);
and U7426 (N_7426,N_6365,N_6789);
xor U7427 (N_7427,N_6681,N_6309);
and U7428 (N_7428,N_6908,N_6232);
or U7429 (N_7429,N_6299,N_6638);
xor U7430 (N_7430,N_6614,N_6531);
xnor U7431 (N_7431,N_6783,N_6977);
and U7432 (N_7432,N_6611,N_6301);
xor U7433 (N_7433,N_6189,N_6069);
or U7434 (N_7434,N_6691,N_6149);
or U7435 (N_7435,N_6510,N_6730);
and U7436 (N_7436,N_6017,N_6886);
nand U7437 (N_7437,N_6718,N_6864);
xor U7438 (N_7438,N_6622,N_6337);
nand U7439 (N_7439,N_6059,N_6078);
and U7440 (N_7440,N_6560,N_6426);
xnor U7441 (N_7441,N_6526,N_6690);
xor U7442 (N_7442,N_6855,N_6208);
nor U7443 (N_7443,N_6095,N_6274);
or U7444 (N_7444,N_6863,N_6624);
nand U7445 (N_7445,N_6537,N_6565);
nor U7446 (N_7446,N_6182,N_6449);
xnor U7447 (N_7447,N_6401,N_6617);
and U7448 (N_7448,N_6601,N_6740);
xnor U7449 (N_7449,N_6559,N_6334);
xnor U7450 (N_7450,N_6845,N_6139);
nand U7451 (N_7451,N_6613,N_6019);
xnor U7452 (N_7452,N_6364,N_6404);
and U7453 (N_7453,N_6329,N_6384);
xnor U7454 (N_7454,N_6371,N_6126);
xnor U7455 (N_7455,N_6319,N_6080);
and U7456 (N_7456,N_6759,N_6042);
or U7457 (N_7457,N_6768,N_6448);
nand U7458 (N_7458,N_6202,N_6499);
xnor U7459 (N_7459,N_6152,N_6640);
xnor U7460 (N_7460,N_6012,N_6529);
nor U7461 (N_7461,N_6869,N_6996);
and U7462 (N_7462,N_6947,N_6063);
xor U7463 (N_7463,N_6697,N_6722);
or U7464 (N_7464,N_6777,N_6041);
nor U7465 (N_7465,N_6331,N_6993);
nand U7466 (N_7466,N_6249,N_6550);
or U7467 (N_7467,N_6616,N_6083);
xor U7468 (N_7468,N_6157,N_6903);
xor U7469 (N_7469,N_6764,N_6146);
and U7470 (N_7470,N_6405,N_6092);
xor U7471 (N_7471,N_6794,N_6509);
xnor U7472 (N_7472,N_6013,N_6460);
or U7473 (N_7473,N_6096,N_6490);
or U7474 (N_7474,N_6532,N_6612);
nor U7475 (N_7475,N_6591,N_6142);
and U7476 (N_7476,N_6107,N_6352);
xor U7477 (N_7477,N_6441,N_6879);
xor U7478 (N_7478,N_6199,N_6419);
xor U7479 (N_7479,N_6725,N_6572);
or U7480 (N_7480,N_6792,N_6883);
and U7481 (N_7481,N_6867,N_6461);
and U7482 (N_7482,N_6742,N_6847);
or U7483 (N_7483,N_6389,N_6138);
or U7484 (N_7484,N_6708,N_6239);
nor U7485 (N_7485,N_6271,N_6306);
or U7486 (N_7486,N_6620,N_6415);
xnor U7487 (N_7487,N_6076,N_6246);
nor U7488 (N_7488,N_6366,N_6226);
nor U7489 (N_7489,N_6313,N_6812);
and U7490 (N_7490,N_6890,N_6985);
nand U7491 (N_7491,N_6103,N_6361);
and U7492 (N_7492,N_6972,N_6736);
and U7493 (N_7493,N_6660,N_6467);
xor U7494 (N_7494,N_6462,N_6093);
and U7495 (N_7495,N_6671,N_6567);
nand U7496 (N_7496,N_6971,N_6210);
xor U7497 (N_7497,N_6788,N_6555);
xor U7498 (N_7498,N_6044,N_6831);
nand U7499 (N_7499,N_6656,N_6256);
nor U7500 (N_7500,N_6402,N_6067);
nand U7501 (N_7501,N_6329,N_6453);
nand U7502 (N_7502,N_6628,N_6999);
or U7503 (N_7503,N_6011,N_6654);
nand U7504 (N_7504,N_6467,N_6183);
nor U7505 (N_7505,N_6922,N_6579);
xor U7506 (N_7506,N_6864,N_6299);
xnor U7507 (N_7507,N_6617,N_6538);
or U7508 (N_7508,N_6319,N_6950);
xor U7509 (N_7509,N_6502,N_6940);
xnor U7510 (N_7510,N_6617,N_6934);
and U7511 (N_7511,N_6535,N_6748);
nand U7512 (N_7512,N_6218,N_6554);
nor U7513 (N_7513,N_6181,N_6158);
and U7514 (N_7514,N_6168,N_6267);
nor U7515 (N_7515,N_6915,N_6653);
xor U7516 (N_7516,N_6720,N_6804);
and U7517 (N_7517,N_6548,N_6906);
nor U7518 (N_7518,N_6030,N_6960);
nor U7519 (N_7519,N_6332,N_6514);
or U7520 (N_7520,N_6124,N_6490);
or U7521 (N_7521,N_6925,N_6138);
or U7522 (N_7522,N_6178,N_6702);
or U7523 (N_7523,N_6614,N_6276);
and U7524 (N_7524,N_6775,N_6096);
or U7525 (N_7525,N_6022,N_6197);
xnor U7526 (N_7526,N_6555,N_6060);
or U7527 (N_7527,N_6669,N_6115);
nor U7528 (N_7528,N_6509,N_6086);
nand U7529 (N_7529,N_6027,N_6487);
nand U7530 (N_7530,N_6654,N_6425);
nand U7531 (N_7531,N_6397,N_6864);
nand U7532 (N_7532,N_6916,N_6383);
and U7533 (N_7533,N_6478,N_6901);
xnor U7534 (N_7534,N_6534,N_6644);
or U7535 (N_7535,N_6226,N_6655);
nand U7536 (N_7536,N_6019,N_6629);
nand U7537 (N_7537,N_6475,N_6696);
nand U7538 (N_7538,N_6311,N_6376);
nor U7539 (N_7539,N_6316,N_6472);
or U7540 (N_7540,N_6445,N_6698);
xnor U7541 (N_7541,N_6500,N_6897);
and U7542 (N_7542,N_6788,N_6626);
nand U7543 (N_7543,N_6877,N_6490);
xnor U7544 (N_7544,N_6904,N_6126);
nand U7545 (N_7545,N_6935,N_6211);
nor U7546 (N_7546,N_6398,N_6902);
nor U7547 (N_7547,N_6394,N_6609);
nand U7548 (N_7548,N_6605,N_6610);
nand U7549 (N_7549,N_6175,N_6762);
nand U7550 (N_7550,N_6941,N_6640);
xor U7551 (N_7551,N_6619,N_6106);
nand U7552 (N_7552,N_6273,N_6305);
xnor U7553 (N_7553,N_6214,N_6774);
nor U7554 (N_7554,N_6891,N_6030);
nor U7555 (N_7555,N_6472,N_6111);
or U7556 (N_7556,N_6126,N_6481);
and U7557 (N_7557,N_6082,N_6119);
nor U7558 (N_7558,N_6573,N_6959);
and U7559 (N_7559,N_6522,N_6290);
xor U7560 (N_7560,N_6728,N_6450);
or U7561 (N_7561,N_6346,N_6005);
nand U7562 (N_7562,N_6526,N_6639);
nor U7563 (N_7563,N_6791,N_6159);
xnor U7564 (N_7564,N_6309,N_6767);
xor U7565 (N_7565,N_6197,N_6674);
or U7566 (N_7566,N_6180,N_6901);
nor U7567 (N_7567,N_6750,N_6056);
xor U7568 (N_7568,N_6832,N_6319);
xnor U7569 (N_7569,N_6644,N_6116);
and U7570 (N_7570,N_6020,N_6591);
or U7571 (N_7571,N_6776,N_6237);
nand U7572 (N_7572,N_6432,N_6091);
xnor U7573 (N_7573,N_6163,N_6267);
and U7574 (N_7574,N_6388,N_6804);
nand U7575 (N_7575,N_6324,N_6896);
or U7576 (N_7576,N_6031,N_6898);
nor U7577 (N_7577,N_6127,N_6088);
xor U7578 (N_7578,N_6912,N_6942);
and U7579 (N_7579,N_6950,N_6604);
xnor U7580 (N_7580,N_6306,N_6871);
or U7581 (N_7581,N_6337,N_6850);
xor U7582 (N_7582,N_6709,N_6893);
nor U7583 (N_7583,N_6203,N_6928);
and U7584 (N_7584,N_6695,N_6866);
and U7585 (N_7585,N_6805,N_6073);
xnor U7586 (N_7586,N_6880,N_6039);
xor U7587 (N_7587,N_6730,N_6743);
nor U7588 (N_7588,N_6797,N_6038);
nor U7589 (N_7589,N_6525,N_6907);
or U7590 (N_7590,N_6479,N_6882);
xor U7591 (N_7591,N_6853,N_6835);
and U7592 (N_7592,N_6139,N_6545);
xnor U7593 (N_7593,N_6274,N_6713);
xor U7594 (N_7594,N_6990,N_6000);
nand U7595 (N_7595,N_6756,N_6298);
or U7596 (N_7596,N_6674,N_6023);
or U7597 (N_7597,N_6391,N_6360);
nor U7598 (N_7598,N_6555,N_6850);
xor U7599 (N_7599,N_6680,N_6310);
nor U7600 (N_7600,N_6741,N_6728);
nand U7601 (N_7601,N_6450,N_6950);
xnor U7602 (N_7602,N_6895,N_6311);
and U7603 (N_7603,N_6458,N_6059);
nor U7604 (N_7604,N_6743,N_6164);
nand U7605 (N_7605,N_6641,N_6070);
nand U7606 (N_7606,N_6335,N_6518);
or U7607 (N_7607,N_6527,N_6875);
xor U7608 (N_7608,N_6887,N_6914);
nand U7609 (N_7609,N_6891,N_6319);
nand U7610 (N_7610,N_6813,N_6016);
nand U7611 (N_7611,N_6376,N_6557);
nand U7612 (N_7612,N_6392,N_6388);
xnor U7613 (N_7613,N_6540,N_6656);
xnor U7614 (N_7614,N_6132,N_6054);
nand U7615 (N_7615,N_6500,N_6096);
nand U7616 (N_7616,N_6104,N_6670);
nand U7617 (N_7617,N_6182,N_6650);
and U7618 (N_7618,N_6761,N_6661);
nor U7619 (N_7619,N_6421,N_6315);
and U7620 (N_7620,N_6685,N_6872);
or U7621 (N_7621,N_6256,N_6700);
and U7622 (N_7622,N_6275,N_6115);
or U7623 (N_7623,N_6736,N_6509);
nand U7624 (N_7624,N_6542,N_6139);
and U7625 (N_7625,N_6403,N_6870);
and U7626 (N_7626,N_6905,N_6132);
xor U7627 (N_7627,N_6335,N_6070);
and U7628 (N_7628,N_6753,N_6351);
xor U7629 (N_7629,N_6711,N_6744);
nand U7630 (N_7630,N_6031,N_6766);
and U7631 (N_7631,N_6355,N_6985);
nor U7632 (N_7632,N_6876,N_6385);
nand U7633 (N_7633,N_6285,N_6077);
nor U7634 (N_7634,N_6233,N_6829);
xor U7635 (N_7635,N_6053,N_6396);
and U7636 (N_7636,N_6464,N_6937);
nor U7637 (N_7637,N_6405,N_6817);
or U7638 (N_7638,N_6278,N_6180);
nor U7639 (N_7639,N_6353,N_6938);
xnor U7640 (N_7640,N_6978,N_6572);
or U7641 (N_7641,N_6792,N_6230);
or U7642 (N_7642,N_6026,N_6529);
nor U7643 (N_7643,N_6981,N_6215);
xnor U7644 (N_7644,N_6480,N_6222);
nor U7645 (N_7645,N_6202,N_6843);
or U7646 (N_7646,N_6898,N_6306);
or U7647 (N_7647,N_6990,N_6937);
and U7648 (N_7648,N_6440,N_6876);
xor U7649 (N_7649,N_6277,N_6160);
nor U7650 (N_7650,N_6653,N_6905);
and U7651 (N_7651,N_6284,N_6700);
xor U7652 (N_7652,N_6046,N_6293);
nand U7653 (N_7653,N_6566,N_6754);
and U7654 (N_7654,N_6682,N_6560);
xnor U7655 (N_7655,N_6786,N_6808);
and U7656 (N_7656,N_6858,N_6019);
or U7657 (N_7657,N_6924,N_6913);
xnor U7658 (N_7658,N_6447,N_6947);
xor U7659 (N_7659,N_6755,N_6427);
or U7660 (N_7660,N_6243,N_6442);
xnor U7661 (N_7661,N_6560,N_6754);
or U7662 (N_7662,N_6448,N_6125);
nand U7663 (N_7663,N_6757,N_6749);
nor U7664 (N_7664,N_6107,N_6824);
nor U7665 (N_7665,N_6941,N_6080);
or U7666 (N_7666,N_6139,N_6394);
nand U7667 (N_7667,N_6894,N_6611);
nand U7668 (N_7668,N_6170,N_6438);
and U7669 (N_7669,N_6926,N_6189);
nand U7670 (N_7670,N_6097,N_6161);
nand U7671 (N_7671,N_6741,N_6431);
or U7672 (N_7672,N_6111,N_6379);
and U7673 (N_7673,N_6864,N_6471);
xnor U7674 (N_7674,N_6294,N_6692);
or U7675 (N_7675,N_6720,N_6400);
xor U7676 (N_7676,N_6439,N_6772);
and U7677 (N_7677,N_6176,N_6098);
nand U7678 (N_7678,N_6663,N_6588);
nor U7679 (N_7679,N_6607,N_6031);
or U7680 (N_7680,N_6765,N_6843);
and U7681 (N_7681,N_6919,N_6142);
nor U7682 (N_7682,N_6195,N_6093);
and U7683 (N_7683,N_6501,N_6505);
and U7684 (N_7684,N_6758,N_6913);
nor U7685 (N_7685,N_6281,N_6416);
nand U7686 (N_7686,N_6232,N_6087);
xnor U7687 (N_7687,N_6774,N_6979);
and U7688 (N_7688,N_6127,N_6836);
xnor U7689 (N_7689,N_6764,N_6715);
or U7690 (N_7690,N_6552,N_6784);
nor U7691 (N_7691,N_6051,N_6434);
nor U7692 (N_7692,N_6552,N_6937);
or U7693 (N_7693,N_6705,N_6294);
nand U7694 (N_7694,N_6053,N_6367);
or U7695 (N_7695,N_6863,N_6384);
xnor U7696 (N_7696,N_6678,N_6839);
or U7697 (N_7697,N_6901,N_6604);
nor U7698 (N_7698,N_6146,N_6306);
nand U7699 (N_7699,N_6688,N_6034);
or U7700 (N_7700,N_6547,N_6473);
nand U7701 (N_7701,N_6801,N_6245);
and U7702 (N_7702,N_6182,N_6764);
nor U7703 (N_7703,N_6484,N_6010);
or U7704 (N_7704,N_6491,N_6728);
and U7705 (N_7705,N_6423,N_6447);
or U7706 (N_7706,N_6408,N_6486);
or U7707 (N_7707,N_6518,N_6376);
nor U7708 (N_7708,N_6858,N_6123);
xor U7709 (N_7709,N_6037,N_6913);
and U7710 (N_7710,N_6971,N_6567);
xor U7711 (N_7711,N_6251,N_6885);
nand U7712 (N_7712,N_6074,N_6599);
nor U7713 (N_7713,N_6510,N_6858);
xnor U7714 (N_7714,N_6778,N_6772);
and U7715 (N_7715,N_6818,N_6456);
nor U7716 (N_7716,N_6564,N_6902);
xor U7717 (N_7717,N_6152,N_6817);
nor U7718 (N_7718,N_6909,N_6863);
and U7719 (N_7719,N_6025,N_6109);
xnor U7720 (N_7720,N_6135,N_6820);
xnor U7721 (N_7721,N_6369,N_6053);
nor U7722 (N_7722,N_6891,N_6858);
or U7723 (N_7723,N_6547,N_6656);
or U7724 (N_7724,N_6509,N_6987);
or U7725 (N_7725,N_6516,N_6426);
nand U7726 (N_7726,N_6384,N_6997);
nor U7727 (N_7727,N_6638,N_6693);
and U7728 (N_7728,N_6193,N_6082);
or U7729 (N_7729,N_6298,N_6124);
nor U7730 (N_7730,N_6209,N_6035);
xnor U7731 (N_7731,N_6091,N_6801);
nand U7732 (N_7732,N_6490,N_6541);
nor U7733 (N_7733,N_6789,N_6230);
nand U7734 (N_7734,N_6216,N_6215);
xnor U7735 (N_7735,N_6477,N_6877);
or U7736 (N_7736,N_6854,N_6473);
nor U7737 (N_7737,N_6333,N_6217);
xnor U7738 (N_7738,N_6762,N_6052);
xnor U7739 (N_7739,N_6989,N_6831);
or U7740 (N_7740,N_6710,N_6919);
nor U7741 (N_7741,N_6577,N_6114);
xor U7742 (N_7742,N_6554,N_6709);
or U7743 (N_7743,N_6290,N_6709);
nand U7744 (N_7744,N_6400,N_6875);
or U7745 (N_7745,N_6936,N_6724);
and U7746 (N_7746,N_6676,N_6721);
nand U7747 (N_7747,N_6213,N_6250);
and U7748 (N_7748,N_6228,N_6900);
nand U7749 (N_7749,N_6721,N_6270);
xnor U7750 (N_7750,N_6886,N_6749);
nand U7751 (N_7751,N_6428,N_6674);
and U7752 (N_7752,N_6915,N_6345);
nand U7753 (N_7753,N_6201,N_6345);
or U7754 (N_7754,N_6243,N_6944);
xnor U7755 (N_7755,N_6946,N_6153);
nand U7756 (N_7756,N_6165,N_6191);
nor U7757 (N_7757,N_6687,N_6772);
xnor U7758 (N_7758,N_6654,N_6212);
nand U7759 (N_7759,N_6506,N_6288);
and U7760 (N_7760,N_6170,N_6960);
nor U7761 (N_7761,N_6683,N_6167);
xor U7762 (N_7762,N_6163,N_6470);
and U7763 (N_7763,N_6476,N_6935);
nand U7764 (N_7764,N_6425,N_6532);
nand U7765 (N_7765,N_6705,N_6453);
nor U7766 (N_7766,N_6107,N_6228);
xnor U7767 (N_7767,N_6971,N_6850);
nand U7768 (N_7768,N_6305,N_6564);
xor U7769 (N_7769,N_6589,N_6850);
xnor U7770 (N_7770,N_6269,N_6623);
and U7771 (N_7771,N_6766,N_6975);
and U7772 (N_7772,N_6113,N_6526);
xor U7773 (N_7773,N_6306,N_6836);
nor U7774 (N_7774,N_6701,N_6877);
nor U7775 (N_7775,N_6445,N_6089);
xor U7776 (N_7776,N_6476,N_6560);
xnor U7777 (N_7777,N_6549,N_6490);
nor U7778 (N_7778,N_6617,N_6904);
xor U7779 (N_7779,N_6927,N_6412);
nor U7780 (N_7780,N_6314,N_6635);
nor U7781 (N_7781,N_6216,N_6203);
xnor U7782 (N_7782,N_6268,N_6509);
and U7783 (N_7783,N_6664,N_6046);
nand U7784 (N_7784,N_6284,N_6335);
or U7785 (N_7785,N_6236,N_6436);
nor U7786 (N_7786,N_6810,N_6098);
nor U7787 (N_7787,N_6920,N_6158);
or U7788 (N_7788,N_6313,N_6099);
and U7789 (N_7789,N_6271,N_6856);
nor U7790 (N_7790,N_6031,N_6717);
xnor U7791 (N_7791,N_6822,N_6008);
or U7792 (N_7792,N_6582,N_6256);
xnor U7793 (N_7793,N_6693,N_6507);
or U7794 (N_7794,N_6081,N_6781);
xnor U7795 (N_7795,N_6657,N_6202);
nor U7796 (N_7796,N_6385,N_6104);
or U7797 (N_7797,N_6228,N_6185);
and U7798 (N_7798,N_6215,N_6257);
nand U7799 (N_7799,N_6690,N_6702);
nor U7800 (N_7800,N_6856,N_6753);
or U7801 (N_7801,N_6421,N_6566);
and U7802 (N_7802,N_6800,N_6218);
or U7803 (N_7803,N_6268,N_6473);
nand U7804 (N_7804,N_6075,N_6130);
or U7805 (N_7805,N_6757,N_6173);
xor U7806 (N_7806,N_6821,N_6281);
xor U7807 (N_7807,N_6732,N_6715);
and U7808 (N_7808,N_6341,N_6736);
nor U7809 (N_7809,N_6846,N_6593);
and U7810 (N_7810,N_6222,N_6732);
nor U7811 (N_7811,N_6544,N_6945);
and U7812 (N_7812,N_6571,N_6621);
and U7813 (N_7813,N_6394,N_6536);
and U7814 (N_7814,N_6159,N_6998);
and U7815 (N_7815,N_6462,N_6169);
or U7816 (N_7816,N_6629,N_6590);
xnor U7817 (N_7817,N_6601,N_6852);
xnor U7818 (N_7818,N_6965,N_6188);
nor U7819 (N_7819,N_6528,N_6996);
and U7820 (N_7820,N_6137,N_6462);
xnor U7821 (N_7821,N_6341,N_6353);
nand U7822 (N_7822,N_6867,N_6826);
or U7823 (N_7823,N_6421,N_6857);
and U7824 (N_7824,N_6007,N_6570);
nor U7825 (N_7825,N_6972,N_6702);
and U7826 (N_7826,N_6107,N_6067);
and U7827 (N_7827,N_6058,N_6240);
and U7828 (N_7828,N_6524,N_6669);
or U7829 (N_7829,N_6425,N_6250);
xnor U7830 (N_7830,N_6682,N_6687);
or U7831 (N_7831,N_6302,N_6355);
or U7832 (N_7832,N_6977,N_6525);
xnor U7833 (N_7833,N_6194,N_6881);
nor U7834 (N_7834,N_6335,N_6094);
xnor U7835 (N_7835,N_6412,N_6899);
and U7836 (N_7836,N_6155,N_6375);
nand U7837 (N_7837,N_6550,N_6612);
nor U7838 (N_7838,N_6491,N_6502);
xor U7839 (N_7839,N_6848,N_6589);
or U7840 (N_7840,N_6107,N_6686);
nor U7841 (N_7841,N_6074,N_6183);
or U7842 (N_7842,N_6655,N_6250);
nand U7843 (N_7843,N_6196,N_6641);
or U7844 (N_7844,N_6453,N_6455);
nand U7845 (N_7845,N_6374,N_6495);
nand U7846 (N_7846,N_6303,N_6779);
or U7847 (N_7847,N_6518,N_6764);
and U7848 (N_7848,N_6385,N_6165);
nand U7849 (N_7849,N_6964,N_6832);
and U7850 (N_7850,N_6964,N_6422);
nand U7851 (N_7851,N_6807,N_6993);
or U7852 (N_7852,N_6974,N_6994);
or U7853 (N_7853,N_6449,N_6019);
xor U7854 (N_7854,N_6776,N_6497);
xnor U7855 (N_7855,N_6312,N_6398);
nand U7856 (N_7856,N_6804,N_6667);
nor U7857 (N_7857,N_6895,N_6668);
or U7858 (N_7858,N_6577,N_6688);
nor U7859 (N_7859,N_6610,N_6737);
xor U7860 (N_7860,N_6545,N_6875);
or U7861 (N_7861,N_6813,N_6632);
or U7862 (N_7862,N_6180,N_6643);
nor U7863 (N_7863,N_6703,N_6458);
or U7864 (N_7864,N_6871,N_6973);
xor U7865 (N_7865,N_6991,N_6043);
nor U7866 (N_7866,N_6270,N_6011);
nor U7867 (N_7867,N_6157,N_6867);
nor U7868 (N_7868,N_6454,N_6191);
and U7869 (N_7869,N_6983,N_6771);
nor U7870 (N_7870,N_6324,N_6863);
nor U7871 (N_7871,N_6385,N_6412);
and U7872 (N_7872,N_6571,N_6514);
and U7873 (N_7873,N_6139,N_6167);
nand U7874 (N_7874,N_6367,N_6597);
xor U7875 (N_7875,N_6634,N_6426);
xor U7876 (N_7876,N_6999,N_6066);
or U7877 (N_7877,N_6190,N_6808);
nor U7878 (N_7878,N_6007,N_6557);
nand U7879 (N_7879,N_6965,N_6729);
or U7880 (N_7880,N_6907,N_6133);
or U7881 (N_7881,N_6317,N_6647);
nor U7882 (N_7882,N_6444,N_6934);
nand U7883 (N_7883,N_6438,N_6220);
or U7884 (N_7884,N_6214,N_6816);
and U7885 (N_7885,N_6960,N_6676);
nor U7886 (N_7886,N_6333,N_6348);
and U7887 (N_7887,N_6367,N_6444);
and U7888 (N_7888,N_6108,N_6899);
xnor U7889 (N_7889,N_6854,N_6924);
nor U7890 (N_7890,N_6966,N_6328);
nor U7891 (N_7891,N_6433,N_6543);
nand U7892 (N_7892,N_6887,N_6122);
nor U7893 (N_7893,N_6429,N_6417);
nand U7894 (N_7894,N_6108,N_6630);
or U7895 (N_7895,N_6134,N_6608);
nor U7896 (N_7896,N_6147,N_6479);
nand U7897 (N_7897,N_6609,N_6896);
or U7898 (N_7898,N_6415,N_6662);
xnor U7899 (N_7899,N_6080,N_6370);
and U7900 (N_7900,N_6182,N_6260);
xor U7901 (N_7901,N_6570,N_6386);
xor U7902 (N_7902,N_6560,N_6643);
or U7903 (N_7903,N_6820,N_6464);
nor U7904 (N_7904,N_6155,N_6799);
and U7905 (N_7905,N_6542,N_6617);
nor U7906 (N_7906,N_6111,N_6273);
nor U7907 (N_7907,N_6003,N_6135);
nand U7908 (N_7908,N_6052,N_6241);
nand U7909 (N_7909,N_6696,N_6883);
and U7910 (N_7910,N_6071,N_6112);
xor U7911 (N_7911,N_6101,N_6718);
or U7912 (N_7912,N_6742,N_6961);
and U7913 (N_7913,N_6218,N_6049);
xor U7914 (N_7914,N_6681,N_6671);
or U7915 (N_7915,N_6554,N_6893);
nor U7916 (N_7916,N_6256,N_6481);
nand U7917 (N_7917,N_6191,N_6362);
nor U7918 (N_7918,N_6628,N_6885);
nand U7919 (N_7919,N_6524,N_6955);
or U7920 (N_7920,N_6183,N_6310);
nand U7921 (N_7921,N_6978,N_6103);
or U7922 (N_7922,N_6196,N_6830);
xnor U7923 (N_7923,N_6649,N_6206);
and U7924 (N_7924,N_6548,N_6011);
and U7925 (N_7925,N_6147,N_6322);
nand U7926 (N_7926,N_6520,N_6194);
or U7927 (N_7927,N_6717,N_6755);
or U7928 (N_7928,N_6054,N_6937);
xnor U7929 (N_7929,N_6337,N_6251);
and U7930 (N_7930,N_6455,N_6126);
nor U7931 (N_7931,N_6548,N_6703);
nand U7932 (N_7932,N_6383,N_6664);
nor U7933 (N_7933,N_6537,N_6825);
nand U7934 (N_7934,N_6051,N_6965);
nor U7935 (N_7935,N_6729,N_6886);
or U7936 (N_7936,N_6087,N_6660);
nor U7937 (N_7937,N_6437,N_6390);
or U7938 (N_7938,N_6479,N_6239);
nand U7939 (N_7939,N_6066,N_6982);
nor U7940 (N_7940,N_6582,N_6689);
or U7941 (N_7941,N_6596,N_6540);
or U7942 (N_7942,N_6734,N_6913);
xor U7943 (N_7943,N_6678,N_6713);
xnor U7944 (N_7944,N_6093,N_6587);
or U7945 (N_7945,N_6399,N_6019);
and U7946 (N_7946,N_6705,N_6995);
nand U7947 (N_7947,N_6495,N_6382);
xnor U7948 (N_7948,N_6617,N_6035);
xnor U7949 (N_7949,N_6578,N_6195);
and U7950 (N_7950,N_6133,N_6676);
nor U7951 (N_7951,N_6793,N_6780);
nor U7952 (N_7952,N_6817,N_6527);
nand U7953 (N_7953,N_6381,N_6118);
or U7954 (N_7954,N_6600,N_6139);
and U7955 (N_7955,N_6734,N_6121);
or U7956 (N_7956,N_6283,N_6852);
xor U7957 (N_7957,N_6987,N_6735);
xor U7958 (N_7958,N_6858,N_6686);
nand U7959 (N_7959,N_6590,N_6420);
xnor U7960 (N_7960,N_6352,N_6345);
nand U7961 (N_7961,N_6382,N_6269);
nor U7962 (N_7962,N_6906,N_6728);
and U7963 (N_7963,N_6006,N_6160);
xnor U7964 (N_7964,N_6479,N_6769);
nand U7965 (N_7965,N_6984,N_6781);
nand U7966 (N_7966,N_6354,N_6679);
and U7967 (N_7967,N_6997,N_6022);
nor U7968 (N_7968,N_6403,N_6634);
nor U7969 (N_7969,N_6715,N_6382);
nand U7970 (N_7970,N_6179,N_6257);
or U7971 (N_7971,N_6079,N_6676);
and U7972 (N_7972,N_6875,N_6946);
nor U7973 (N_7973,N_6076,N_6374);
or U7974 (N_7974,N_6633,N_6152);
nand U7975 (N_7975,N_6697,N_6996);
nor U7976 (N_7976,N_6666,N_6846);
and U7977 (N_7977,N_6018,N_6797);
xor U7978 (N_7978,N_6134,N_6449);
nand U7979 (N_7979,N_6608,N_6673);
xnor U7980 (N_7980,N_6908,N_6192);
and U7981 (N_7981,N_6482,N_6888);
xnor U7982 (N_7982,N_6005,N_6328);
nand U7983 (N_7983,N_6773,N_6295);
or U7984 (N_7984,N_6991,N_6957);
xnor U7985 (N_7985,N_6457,N_6437);
or U7986 (N_7986,N_6964,N_6149);
xor U7987 (N_7987,N_6550,N_6321);
nand U7988 (N_7988,N_6456,N_6770);
nor U7989 (N_7989,N_6786,N_6235);
and U7990 (N_7990,N_6134,N_6994);
and U7991 (N_7991,N_6817,N_6374);
nor U7992 (N_7992,N_6169,N_6837);
xor U7993 (N_7993,N_6908,N_6746);
nand U7994 (N_7994,N_6810,N_6676);
xor U7995 (N_7995,N_6911,N_6117);
or U7996 (N_7996,N_6665,N_6389);
nand U7997 (N_7997,N_6265,N_6069);
xor U7998 (N_7998,N_6671,N_6949);
nand U7999 (N_7999,N_6818,N_6257);
xnor U8000 (N_8000,N_7800,N_7311);
or U8001 (N_8001,N_7192,N_7527);
nand U8002 (N_8002,N_7920,N_7531);
nand U8003 (N_8003,N_7475,N_7607);
and U8004 (N_8004,N_7133,N_7126);
nor U8005 (N_8005,N_7547,N_7259);
nand U8006 (N_8006,N_7304,N_7706);
nand U8007 (N_8007,N_7479,N_7303);
xnor U8008 (N_8008,N_7209,N_7046);
and U8009 (N_8009,N_7541,N_7322);
xor U8010 (N_8010,N_7513,N_7953);
nor U8011 (N_8011,N_7723,N_7766);
or U8012 (N_8012,N_7592,N_7963);
xor U8013 (N_8013,N_7058,N_7077);
nand U8014 (N_8014,N_7786,N_7495);
nor U8015 (N_8015,N_7840,N_7150);
or U8016 (N_8016,N_7299,N_7526);
and U8017 (N_8017,N_7941,N_7110);
xnor U8018 (N_8018,N_7249,N_7178);
xor U8019 (N_8019,N_7960,N_7971);
and U8020 (N_8020,N_7424,N_7091);
xor U8021 (N_8021,N_7632,N_7595);
nor U8022 (N_8022,N_7198,N_7929);
or U8023 (N_8023,N_7462,N_7961);
xnor U8024 (N_8024,N_7431,N_7896);
nand U8025 (N_8025,N_7180,N_7887);
xor U8026 (N_8026,N_7845,N_7329);
xnor U8027 (N_8027,N_7289,N_7662);
xor U8028 (N_8028,N_7038,N_7269);
xnor U8029 (N_8029,N_7957,N_7990);
xnor U8030 (N_8030,N_7219,N_7707);
xnor U8031 (N_8031,N_7391,N_7035);
or U8032 (N_8032,N_7555,N_7335);
xor U8033 (N_8033,N_7827,N_7146);
nand U8034 (N_8034,N_7678,N_7710);
nand U8035 (N_8035,N_7725,N_7759);
or U8036 (N_8036,N_7429,N_7125);
nand U8037 (N_8037,N_7435,N_7208);
nor U8038 (N_8038,N_7925,N_7411);
and U8039 (N_8039,N_7293,N_7865);
xor U8040 (N_8040,N_7366,N_7212);
nor U8041 (N_8041,N_7317,N_7023);
or U8042 (N_8042,N_7296,N_7338);
nor U8043 (N_8043,N_7457,N_7735);
or U8044 (N_8044,N_7911,N_7739);
nand U8045 (N_8045,N_7380,N_7397);
xor U8046 (N_8046,N_7181,N_7994);
xor U8047 (N_8047,N_7423,N_7666);
or U8048 (N_8048,N_7367,N_7128);
xnor U8049 (N_8049,N_7717,N_7230);
nor U8050 (N_8050,N_7959,N_7202);
or U8051 (N_8051,N_7408,N_7593);
nor U8052 (N_8052,N_7647,N_7798);
nor U8053 (N_8053,N_7825,N_7747);
nor U8054 (N_8054,N_7331,N_7697);
nand U8055 (N_8055,N_7818,N_7882);
and U8056 (N_8056,N_7458,N_7363);
xnor U8057 (N_8057,N_7660,N_7403);
and U8058 (N_8058,N_7740,N_7471);
nand U8059 (N_8059,N_7797,N_7536);
xor U8060 (N_8060,N_7646,N_7453);
nand U8061 (N_8061,N_7651,N_7998);
nand U8062 (N_8062,N_7060,N_7467);
or U8063 (N_8063,N_7567,N_7654);
nor U8064 (N_8064,N_7315,N_7732);
xnor U8065 (N_8065,N_7681,N_7897);
xor U8066 (N_8066,N_7412,N_7116);
xor U8067 (N_8067,N_7179,N_7688);
or U8068 (N_8068,N_7982,N_7696);
and U8069 (N_8069,N_7078,N_7701);
or U8070 (N_8070,N_7578,N_7068);
xnor U8071 (N_8071,N_7055,N_7967);
and U8072 (N_8072,N_7835,N_7670);
and U8073 (N_8073,N_7885,N_7398);
nor U8074 (N_8074,N_7124,N_7459);
and U8075 (N_8075,N_7502,N_7040);
nor U8076 (N_8076,N_7444,N_7190);
and U8077 (N_8077,N_7045,N_7746);
xnor U8078 (N_8078,N_7251,N_7463);
nand U8079 (N_8079,N_7748,N_7067);
and U8080 (N_8080,N_7011,N_7652);
xnor U8081 (N_8081,N_7007,N_7912);
nand U8082 (N_8082,N_7501,N_7901);
nor U8083 (N_8083,N_7785,N_7553);
or U8084 (N_8084,N_7240,N_7573);
or U8085 (N_8085,N_7616,N_7935);
xnor U8086 (N_8086,N_7523,N_7884);
xnor U8087 (N_8087,N_7056,N_7191);
or U8088 (N_8088,N_7503,N_7954);
and U8089 (N_8089,N_7917,N_7194);
nand U8090 (N_8090,N_7017,N_7522);
or U8091 (N_8091,N_7724,N_7637);
nor U8092 (N_8092,N_7783,N_7628);
and U8093 (N_8093,N_7810,N_7499);
xnor U8094 (N_8094,N_7227,N_7563);
and U8095 (N_8095,N_7619,N_7385);
or U8096 (N_8096,N_7184,N_7330);
nor U8097 (N_8097,N_7610,N_7399);
nand U8098 (N_8098,N_7942,N_7348);
nor U8099 (N_8099,N_7000,N_7430);
or U8100 (N_8100,N_7490,N_7332);
or U8101 (N_8101,N_7373,N_7656);
xor U8102 (N_8102,N_7460,N_7653);
nor U8103 (N_8103,N_7505,N_7736);
or U8104 (N_8104,N_7402,N_7611);
nand U8105 (N_8105,N_7745,N_7493);
nand U8106 (N_8106,N_7864,N_7859);
nor U8107 (N_8107,N_7254,N_7873);
or U8108 (N_8108,N_7674,N_7152);
and U8109 (N_8109,N_7443,N_7438);
or U8110 (N_8110,N_7253,N_7881);
nand U8111 (N_8111,N_7708,N_7709);
or U8112 (N_8112,N_7326,N_7137);
nor U8113 (N_8113,N_7496,N_7819);
or U8114 (N_8114,N_7236,N_7115);
nand U8115 (N_8115,N_7451,N_7816);
xor U8116 (N_8116,N_7050,N_7968);
nand U8117 (N_8117,N_7649,N_7053);
or U8118 (N_8118,N_7312,N_7266);
and U8119 (N_8119,N_7980,N_7770);
nor U8120 (N_8120,N_7114,N_7988);
and U8121 (N_8121,N_7310,N_7339);
xor U8122 (N_8122,N_7158,N_7700);
or U8123 (N_8123,N_7521,N_7229);
and U8124 (N_8124,N_7323,N_7016);
or U8125 (N_8125,N_7188,N_7215);
or U8126 (N_8126,N_7083,N_7672);
and U8127 (N_8127,N_7029,N_7956);
nand U8128 (N_8128,N_7744,N_7549);
or U8129 (N_8129,N_7342,N_7716);
xnor U8130 (N_8130,N_7472,N_7528);
nand U8131 (N_8131,N_7879,N_7794);
nand U8132 (N_8132,N_7504,N_7009);
nand U8133 (N_8133,N_7066,N_7142);
and U8134 (N_8134,N_7109,N_7842);
xnor U8135 (N_8135,N_7659,N_7689);
nor U8136 (N_8136,N_7924,N_7934);
nor U8137 (N_8137,N_7583,N_7404);
nor U8138 (N_8138,N_7589,N_7914);
and U8139 (N_8139,N_7880,N_7764);
or U8140 (N_8140,N_7750,N_7564);
and U8141 (N_8141,N_7422,N_7347);
nand U8142 (N_8142,N_7006,N_7359);
and U8143 (N_8143,N_7650,N_7939);
and U8144 (N_8144,N_7540,N_7871);
xor U8145 (N_8145,N_7878,N_7407);
nor U8146 (N_8146,N_7409,N_7135);
nand U8147 (N_8147,N_7612,N_7313);
xnor U8148 (N_8148,N_7099,N_7103);
nor U8149 (N_8149,N_7532,N_7134);
xnor U8150 (N_8150,N_7774,N_7364);
nor U8151 (N_8151,N_7262,N_7480);
xnor U8152 (N_8152,N_7092,N_7233);
and U8153 (N_8153,N_7287,N_7014);
xnor U8154 (N_8154,N_7515,N_7157);
xnor U8155 (N_8155,N_7870,N_7148);
and U8156 (N_8156,N_7602,N_7594);
and U8157 (N_8157,N_7183,N_7519);
nor U8158 (N_8158,N_7591,N_7173);
and U8159 (N_8159,N_7905,N_7857);
nor U8160 (N_8160,N_7909,N_7626);
nor U8161 (N_8161,N_7343,N_7437);
or U8162 (N_8162,N_7906,N_7787);
xor U8163 (N_8163,N_7605,N_7379);
nand U8164 (N_8164,N_7966,N_7974);
nor U8165 (N_8165,N_7627,N_7383);
or U8166 (N_8166,N_7965,N_7280);
xnor U8167 (N_8167,N_7439,N_7096);
nor U8168 (N_8168,N_7769,N_7828);
and U8169 (N_8169,N_7100,N_7107);
nand U8170 (N_8170,N_7903,N_7345);
nand U8171 (N_8171,N_7111,N_7354);
xor U8172 (N_8172,N_7761,N_7288);
nor U8173 (N_8173,N_7946,N_7557);
and U8174 (N_8174,N_7441,N_7510);
nand U8175 (N_8175,N_7143,N_7071);
nor U8176 (N_8176,N_7369,N_7203);
xor U8177 (N_8177,N_7042,N_7846);
xnor U8178 (N_8178,N_7093,N_7820);
or U8179 (N_8179,N_7534,N_7639);
nor U8180 (N_8180,N_7734,N_7085);
nor U8181 (N_8181,N_7175,N_7772);
or U8182 (N_8182,N_7738,N_7763);
nor U8183 (N_8183,N_7353,N_7687);
or U8184 (N_8184,N_7168,N_7374);
xor U8185 (N_8185,N_7396,N_7350);
nand U8186 (N_8186,N_7052,N_7976);
nand U8187 (N_8187,N_7756,N_7377);
and U8188 (N_8188,N_7908,N_7705);
nand U8189 (N_8189,N_7642,N_7235);
and U8190 (N_8190,N_7730,N_7973);
nand U8191 (N_8191,N_7643,N_7415);
or U8192 (N_8192,N_7483,N_7552);
or U8193 (N_8193,N_7948,N_7144);
or U8194 (N_8194,N_7847,N_7722);
xor U8195 (N_8195,N_7788,N_7558);
nand U8196 (N_8196,N_7789,N_7599);
or U8197 (N_8197,N_7305,N_7225);
and U8198 (N_8198,N_7172,N_7655);
or U8199 (N_8199,N_7349,N_7586);
xor U8200 (N_8200,N_7623,N_7294);
nand U8201 (N_8201,N_7520,N_7970);
and U8202 (N_8202,N_7661,N_7321);
xor U8203 (N_8203,N_7962,N_7702);
nand U8204 (N_8204,N_7197,N_7488);
xnor U8205 (N_8205,N_7242,N_7665);
and U8206 (N_8206,N_7171,N_7297);
nor U8207 (N_8207,N_7693,N_7445);
xnor U8208 (N_8208,N_7365,N_7755);
xor U8209 (N_8209,N_7270,N_7476);
or U8210 (N_8210,N_7440,N_7875);
and U8211 (N_8211,N_7999,N_7153);
xnor U8212 (N_8212,N_7837,N_7683);
xnor U8213 (N_8213,N_7856,N_7267);
or U8214 (N_8214,N_7389,N_7018);
or U8215 (N_8215,N_7617,N_7587);
xnor U8216 (N_8216,N_7640,N_7664);
xor U8217 (N_8217,N_7570,N_7216);
or U8218 (N_8218,N_7778,N_7868);
xor U8219 (N_8219,N_7084,N_7596);
nor U8220 (N_8220,N_7757,N_7630);
or U8221 (N_8221,N_7600,N_7393);
and U8222 (N_8222,N_7516,N_7826);
or U8223 (N_8223,N_7069,N_7370);
or U8224 (N_8224,N_7768,N_7392);
xnor U8225 (N_8225,N_7395,N_7509);
and U8226 (N_8226,N_7104,N_7162);
nor U8227 (N_8227,N_7727,N_7484);
nand U8228 (N_8228,N_7063,N_7576);
and U8229 (N_8229,N_7613,N_7489);
or U8230 (N_8230,N_7244,N_7057);
nand U8231 (N_8231,N_7442,N_7074);
or U8232 (N_8232,N_7585,N_7200);
nor U8233 (N_8233,N_7477,N_7160);
nand U8234 (N_8234,N_7633,N_7760);
and U8235 (N_8235,N_7933,N_7079);
and U8236 (N_8236,N_7986,N_7718);
and U8237 (N_8237,N_7132,N_7138);
or U8238 (N_8238,N_7806,N_7070);
nor U8239 (N_8239,N_7386,N_7360);
xor U8240 (N_8240,N_7784,N_7316);
nor U8241 (N_8241,N_7945,N_7852);
and U8242 (N_8242,N_7106,N_7185);
and U8243 (N_8243,N_7921,N_7944);
and U8244 (N_8244,N_7765,N_7877);
xnor U8245 (N_8245,N_7663,N_7196);
nand U8246 (N_8246,N_7743,N_7276);
nand U8247 (N_8247,N_7927,N_7416);
xor U8248 (N_8248,N_7469,N_7985);
or U8249 (N_8249,N_7679,N_7898);
nor U8250 (N_8250,N_7265,N_7087);
nor U8251 (N_8251,N_7812,N_7801);
and U8252 (N_8252,N_7910,N_7170);
xor U8253 (N_8253,N_7657,N_7274);
nor U8254 (N_8254,N_7932,N_7952);
nand U8255 (N_8255,N_7686,N_7206);
and U8256 (N_8256,N_7947,N_7487);
nand U8257 (N_8257,N_7072,N_7327);
nor U8258 (N_8258,N_7560,N_7382);
nand U8259 (N_8259,N_7166,N_7533);
or U8260 (N_8260,N_7234,N_7448);
xor U8261 (N_8261,N_7538,N_7036);
nor U8262 (N_8262,N_7177,N_7543);
nand U8263 (N_8263,N_7728,N_7972);
or U8264 (N_8264,N_7086,N_7272);
nand U8265 (N_8265,N_7039,N_7207);
nand U8266 (N_8266,N_7456,N_7530);
nand U8267 (N_8267,N_7804,N_7088);
xnor U8268 (N_8268,N_7913,N_7995);
nand U8269 (N_8269,N_7983,N_7062);
xor U8270 (N_8270,N_7400,N_7454);
xnor U8271 (N_8271,N_7685,N_7928);
or U8272 (N_8272,N_7569,N_7899);
nand U8273 (N_8273,N_7387,N_7836);
nor U8274 (N_8274,N_7256,N_7518);
and U8275 (N_8275,N_7824,N_7465);
and U8276 (N_8276,N_7466,N_7277);
nor U8277 (N_8277,N_7580,N_7022);
and U8278 (N_8278,N_7893,N_7468);
nor U8279 (N_8279,N_7565,N_7830);
nor U8280 (N_8280,N_7636,N_7620);
and U8281 (N_8281,N_7449,N_7119);
nor U8282 (N_8282,N_7147,N_7224);
or U8283 (N_8283,N_7575,N_7507);
nor U8284 (N_8284,N_7482,N_7891);
xnor U8285 (N_8285,N_7300,N_7497);
nor U8286 (N_8286,N_7481,N_7869);
nor U8287 (N_8287,N_7264,N_7777);
xor U8288 (N_8288,N_7075,N_7268);
xnor U8289 (N_8289,N_7217,N_7361);
and U8290 (N_8290,N_7904,N_7714);
and U8291 (N_8291,N_7950,N_7043);
nor U8292 (N_8292,N_7936,N_7394);
xnor U8293 (N_8293,N_7559,N_7817);
nor U8294 (N_8294,N_7969,N_7426);
nor U8295 (N_8295,N_7117,N_7427);
and U8296 (N_8296,N_7260,N_7461);
xor U8297 (N_8297,N_7922,N_7434);
xnor U8298 (N_8298,N_7252,N_7711);
xor U8299 (N_8299,N_7669,N_7713);
nand U8300 (N_8300,N_7680,N_7937);
xor U8301 (N_8301,N_7888,N_7129);
xnor U8302 (N_8302,N_7691,N_7958);
and U8303 (N_8303,N_7989,N_7436);
xnor U8304 (N_8304,N_7566,N_7771);
nor U8305 (N_8305,N_7991,N_7275);
or U8306 (N_8306,N_7556,N_7250);
xor U8307 (N_8307,N_7384,N_7588);
and U8308 (N_8308,N_7841,N_7858);
and U8309 (N_8309,N_7019,N_7065);
and U8310 (N_8310,N_7892,N_7625);
nand U8311 (N_8311,N_7237,N_7694);
xnor U8312 (N_8312,N_7120,N_7273);
or U8313 (N_8313,N_7352,N_7889);
nand U8314 (N_8314,N_7163,N_7512);
or U8315 (N_8315,N_7601,N_7930);
nand U8316 (N_8316,N_7780,N_7314);
and U8317 (N_8317,N_7742,N_7608);
nor U8318 (N_8318,N_7145,N_7975);
xor U8319 (N_8319,N_7076,N_7005);
or U8320 (N_8320,N_7634,N_7306);
xor U8321 (N_8321,N_7658,N_7049);
nand U8322 (N_8322,N_7095,N_7692);
and U8323 (N_8323,N_7261,N_7285);
and U8324 (N_8324,N_7508,N_7413);
or U8325 (N_8325,N_7328,N_7378);
xor U8326 (N_8326,N_7539,N_7101);
xor U8327 (N_8327,N_7337,N_7815);
xnor U8328 (N_8328,N_7258,N_7997);
or U8329 (N_8329,N_7105,N_7517);
and U8330 (N_8330,N_7492,N_7542);
nand U8331 (N_8331,N_7803,N_7102);
nor U8332 (N_8332,N_7562,N_7161);
or U8333 (N_8333,N_7123,N_7025);
xnor U8334 (N_8334,N_7210,N_7080);
nand U8335 (N_8335,N_7853,N_7221);
or U8336 (N_8336,N_7834,N_7059);
xor U8337 (N_8337,N_7844,N_7604);
or U8338 (N_8338,N_7715,N_7420);
and U8339 (N_8339,N_7464,N_7341);
nand U8340 (N_8340,N_7176,N_7829);
or U8341 (N_8341,N_7452,N_7606);
xnor U8342 (N_8342,N_7579,N_7141);
and U8343 (N_8343,N_7703,N_7298);
xor U8344 (N_8344,N_7597,N_7895);
and U8345 (N_8345,N_7098,N_7428);
and U8346 (N_8346,N_7546,N_7598);
or U8347 (N_8347,N_7823,N_7336);
nand U8348 (N_8348,N_7618,N_7245);
or U8349 (N_8349,N_7187,N_7228);
xnor U8350 (N_8350,N_7358,N_7799);
xnor U8351 (N_8351,N_7248,N_7247);
and U8352 (N_8352,N_7561,N_7622);
or U8353 (N_8353,N_7741,N_7964);
nor U8354 (N_8354,N_7432,N_7271);
and U8355 (N_8355,N_7455,N_7406);
nor U8356 (N_8356,N_7796,N_7319);
nand U8357 (N_8357,N_7401,N_7676);
xnor U8358 (N_8358,N_7008,N_7381);
and U8359 (N_8359,N_7281,N_7189);
xor U8360 (N_8360,N_7047,N_7118);
and U8361 (N_8361,N_7218,N_7222);
nand U8362 (N_8362,N_7450,N_7726);
nor U8363 (N_8363,N_7851,N_7226);
xnor U8364 (N_8364,N_7886,N_7108);
nand U8365 (N_8365,N_7839,N_7807);
or U8366 (N_8366,N_7026,N_7902);
xnor U8367 (N_8367,N_7193,N_7849);
nor U8368 (N_8368,N_7822,N_7122);
xnor U8369 (N_8369,N_7729,N_7671);
and U8370 (N_8370,N_7165,N_7325);
xor U8371 (N_8371,N_7609,N_7243);
or U8372 (N_8372,N_7511,N_7506);
nand U8373 (N_8373,N_7791,N_7758);
nor U8374 (N_8374,N_7308,N_7500);
xnor U8375 (N_8375,N_7872,N_7677);
or U8376 (N_8376,N_7199,N_7907);
xor U8377 (N_8377,N_7376,N_7793);
and U8378 (N_8378,N_7894,N_7890);
nor U8379 (N_8379,N_7255,N_7590);
nor U8380 (N_8380,N_7213,N_7773);
xor U8381 (N_8381,N_7003,N_7239);
nand U8382 (N_8382,N_7603,N_7082);
xnor U8383 (N_8383,N_7550,N_7012);
or U8384 (N_8384,N_7195,N_7848);
nor U8385 (N_8385,N_7802,N_7446);
nand U8386 (N_8386,N_7978,N_7548);
and U8387 (N_8387,N_7667,N_7309);
xnor U8388 (N_8388,N_7641,N_7149);
nand U8389 (N_8389,N_7544,N_7916);
nand U8390 (N_8390,N_7987,N_7470);
nor U8391 (N_8391,N_7372,N_7169);
nand U8392 (N_8392,N_7535,N_7028);
and U8393 (N_8393,N_7155,N_7863);
or U8394 (N_8394,N_7231,N_7290);
nand U8395 (N_8395,N_7582,N_7673);
and U8396 (N_8396,N_7425,N_7238);
xor U8397 (N_8397,N_7151,N_7733);
or U8398 (N_8398,N_7286,N_7356);
nand U8399 (N_8399,N_7776,N_7631);
xnor U8400 (N_8400,N_7010,N_7127);
nor U8401 (N_8401,N_7719,N_7645);
and U8402 (N_8402,N_7362,N_7205);
nor U8403 (N_8403,N_7346,N_7048);
xor U8404 (N_8404,N_7615,N_7320);
or U8405 (N_8405,N_7574,N_7767);
nor U8406 (N_8406,N_7112,N_7090);
nand U8407 (N_8407,N_7644,N_7943);
and U8408 (N_8408,N_7027,N_7167);
xor U8409 (N_8409,N_7186,N_7241);
and U8410 (N_8410,N_7278,N_7751);
nand U8411 (N_8411,N_7781,N_7139);
xor U8412 (N_8412,N_7762,N_7291);
nor U8413 (N_8413,N_7821,N_7201);
or U8414 (N_8414,N_7949,N_7979);
nor U8415 (N_8415,N_7473,N_7577);
or U8416 (N_8416,N_7390,N_7081);
or U8417 (N_8417,N_7371,N_7204);
nor U8418 (N_8418,N_7182,N_7981);
nor U8419 (N_8419,N_7926,N_7737);
or U8420 (N_8420,N_7699,N_7675);
and U8421 (N_8421,N_7485,N_7993);
or U8422 (N_8422,N_7094,N_7919);
nor U8423 (N_8423,N_7813,N_7375);
or U8424 (N_8424,N_7494,N_7614);
and U8425 (N_8425,N_7690,N_7792);
nor U8426 (N_8426,N_7032,N_7862);
nor U8427 (N_8427,N_7782,N_7417);
nand U8428 (N_8428,N_7918,N_7779);
xor U8429 (N_8429,N_7355,N_7021);
and U8430 (N_8430,N_7754,N_7302);
xor U8431 (N_8431,N_7002,N_7866);
and U8432 (N_8432,N_7915,N_7140);
or U8433 (N_8433,N_7051,N_7214);
nor U8434 (N_8434,N_7638,N_7874);
or U8435 (N_8435,N_7414,N_7033);
xor U8436 (N_8436,N_7900,N_7704);
or U8437 (N_8437,N_7156,N_7113);
and U8438 (N_8438,N_7698,N_7833);
or U8439 (N_8439,N_7131,N_7838);
and U8440 (N_8440,N_7004,N_7854);
xnor U8441 (N_8441,N_7860,N_7753);
xor U8442 (N_8442,N_7572,N_7097);
nor U8443 (N_8443,N_7324,N_7537);
and U8444 (N_8444,N_7232,N_7568);
nor U8445 (N_8445,N_7292,N_7861);
or U8446 (N_8446,N_7013,N_7938);
nor U8447 (N_8447,N_7931,N_7211);
nor U8448 (N_8448,N_7174,N_7015);
nor U8449 (N_8449,N_7977,N_7037);
nand U8450 (N_8450,N_7418,N_7486);
nand U8451 (N_8451,N_7811,N_7668);
and U8452 (N_8452,N_7164,N_7447);
nor U8453 (N_8453,N_7020,N_7996);
nand U8454 (N_8454,N_7301,N_7031);
xnor U8455 (N_8455,N_7635,N_7334);
nand U8456 (N_8456,N_7581,N_7024);
xnor U8457 (N_8457,N_7344,N_7984);
nor U8458 (N_8458,N_7279,N_7629);
xor U8459 (N_8459,N_7808,N_7529);
xnor U8460 (N_8460,N_7720,N_7831);
xnor U8461 (N_8461,N_7054,N_7405);
or U8462 (N_8462,N_7089,N_7357);
or U8463 (N_8463,N_7855,N_7571);
nor U8464 (N_8464,N_7525,N_7551);
nand U8465 (N_8465,N_7041,N_7030);
xnor U8466 (N_8466,N_7621,N_7421);
xnor U8467 (N_8467,N_7712,N_7136);
or U8468 (N_8468,N_7951,N_7814);
nor U8469 (N_8469,N_7064,N_7263);
and U8470 (N_8470,N_7992,N_7001);
or U8471 (N_8471,N_7368,N_7283);
and U8472 (N_8472,N_7955,N_7775);
or U8473 (N_8473,N_7514,N_7223);
nor U8474 (N_8474,N_7795,N_7257);
or U8475 (N_8475,N_7333,N_7419);
xnor U8476 (N_8476,N_7121,N_7624);
nor U8477 (N_8477,N_7433,N_7220);
xnor U8478 (N_8478,N_7876,N_7034);
and U8479 (N_8479,N_7284,N_7923);
nand U8480 (N_8480,N_7809,N_7159);
and U8481 (N_8481,N_7478,N_7154);
nand U8482 (N_8482,N_7061,N_7351);
nor U8483 (N_8483,N_7340,N_7790);
nand U8484 (N_8484,N_7584,N_7295);
nand U8485 (N_8485,N_7307,N_7498);
nand U8486 (N_8486,N_7545,N_7130);
nor U8487 (N_8487,N_7648,N_7721);
or U8488 (N_8488,N_7282,N_7491);
xnor U8489 (N_8489,N_7752,N_7832);
or U8490 (N_8490,N_7850,N_7073);
and U8491 (N_8491,N_7246,N_7474);
and U8492 (N_8492,N_7695,N_7554);
or U8493 (N_8493,N_7044,N_7731);
xor U8494 (N_8494,N_7940,N_7805);
nor U8495 (N_8495,N_7749,N_7410);
xor U8496 (N_8496,N_7867,N_7843);
nand U8497 (N_8497,N_7318,N_7883);
and U8498 (N_8498,N_7682,N_7388);
nand U8499 (N_8499,N_7524,N_7684);
nor U8500 (N_8500,N_7961,N_7882);
nand U8501 (N_8501,N_7266,N_7754);
nand U8502 (N_8502,N_7094,N_7897);
nand U8503 (N_8503,N_7232,N_7927);
and U8504 (N_8504,N_7874,N_7813);
and U8505 (N_8505,N_7298,N_7573);
and U8506 (N_8506,N_7427,N_7120);
and U8507 (N_8507,N_7627,N_7092);
and U8508 (N_8508,N_7797,N_7150);
xnor U8509 (N_8509,N_7619,N_7426);
nor U8510 (N_8510,N_7807,N_7098);
nor U8511 (N_8511,N_7348,N_7370);
xnor U8512 (N_8512,N_7543,N_7192);
nor U8513 (N_8513,N_7247,N_7735);
and U8514 (N_8514,N_7686,N_7994);
nand U8515 (N_8515,N_7003,N_7514);
nor U8516 (N_8516,N_7279,N_7458);
nor U8517 (N_8517,N_7698,N_7376);
and U8518 (N_8518,N_7859,N_7219);
nor U8519 (N_8519,N_7560,N_7352);
and U8520 (N_8520,N_7994,N_7232);
xor U8521 (N_8521,N_7803,N_7872);
or U8522 (N_8522,N_7149,N_7798);
nor U8523 (N_8523,N_7657,N_7485);
nand U8524 (N_8524,N_7107,N_7961);
nand U8525 (N_8525,N_7432,N_7366);
nor U8526 (N_8526,N_7687,N_7096);
and U8527 (N_8527,N_7659,N_7359);
nand U8528 (N_8528,N_7104,N_7657);
nand U8529 (N_8529,N_7764,N_7219);
nor U8530 (N_8530,N_7367,N_7906);
xor U8531 (N_8531,N_7686,N_7679);
or U8532 (N_8532,N_7057,N_7549);
or U8533 (N_8533,N_7057,N_7436);
and U8534 (N_8534,N_7933,N_7075);
or U8535 (N_8535,N_7328,N_7103);
or U8536 (N_8536,N_7881,N_7527);
or U8537 (N_8537,N_7113,N_7613);
and U8538 (N_8538,N_7274,N_7016);
and U8539 (N_8539,N_7025,N_7412);
and U8540 (N_8540,N_7391,N_7098);
or U8541 (N_8541,N_7419,N_7312);
and U8542 (N_8542,N_7182,N_7786);
and U8543 (N_8543,N_7087,N_7842);
or U8544 (N_8544,N_7072,N_7222);
xnor U8545 (N_8545,N_7875,N_7990);
nor U8546 (N_8546,N_7994,N_7280);
xor U8547 (N_8547,N_7541,N_7534);
nor U8548 (N_8548,N_7628,N_7554);
or U8549 (N_8549,N_7524,N_7316);
or U8550 (N_8550,N_7389,N_7676);
and U8551 (N_8551,N_7606,N_7715);
xnor U8552 (N_8552,N_7699,N_7497);
nand U8553 (N_8553,N_7354,N_7784);
nand U8554 (N_8554,N_7575,N_7815);
and U8555 (N_8555,N_7406,N_7154);
xnor U8556 (N_8556,N_7929,N_7379);
nand U8557 (N_8557,N_7670,N_7174);
and U8558 (N_8558,N_7544,N_7733);
or U8559 (N_8559,N_7314,N_7873);
and U8560 (N_8560,N_7910,N_7960);
nand U8561 (N_8561,N_7286,N_7635);
nor U8562 (N_8562,N_7363,N_7389);
nor U8563 (N_8563,N_7602,N_7907);
nand U8564 (N_8564,N_7962,N_7242);
xnor U8565 (N_8565,N_7463,N_7315);
or U8566 (N_8566,N_7660,N_7543);
nor U8567 (N_8567,N_7450,N_7075);
and U8568 (N_8568,N_7178,N_7225);
or U8569 (N_8569,N_7900,N_7398);
and U8570 (N_8570,N_7309,N_7479);
and U8571 (N_8571,N_7260,N_7173);
nor U8572 (N_8572,N_7161,N_7151);
xor U8573 (N_8573,N_7059,N_7479);
xor U8574 (N_8574,N_7756,N_7576);
nor U8575 (N_8575,N_7090,N_7489);
nand U8576 (N_8576,N_7268,N_7897);
xor U8577 (N_8577,N_7101,N_7111);
xor U8578 (N_8578,N_7116,N_7433);
or U8579 (N_8579,N_7347,N_7672);
and U8580 (N_8580,N_7823,N_7233);
nor U8581 (N_8581,N_7659,N_7386);
xnor U8582 (N_8582,N_7724,N_7177);
nand U8583 (N_8583,N_7711,N_7417);
and U8584 (N_8584,N_7260,N_7115);
nor U8585 (N_8585,N_7232,N_7846);
and U8586 (N_8586,N_7039,N_7462);
xnor U8587 (N_8587,N_7067,N_7677);
nor U8588 (N_8588,N_7322,N_7599);
or U8589 (N_8589,N_7417,N_7991);
or U8590 (N_8590,N_7282,N_7995);
nor U8591 (N_8591,N_7714,N_7031);
nor U8592 (N_8592,N_7603,N_7668);
nand U8593 (N_8593,N_7847,N_7066);
xnor U8594 (N_8594,N_7854,N_7886);
xor U8595 (N_8595,N_7230,N_7700);
or U8596 (N_8596,N_7347,N_7269);
nor U8597 (N_8597,N_7506,N_7100);
xnor U8598 (N_8598,N_7427,N_7193);
nand U8599 (N_8599,N_7442,N_7072);
xnor U8600 (N_8600,N_7894,N_7346);
and U8601 (N_8601,N_7970,N_7488);
or U8602 (N_8602,N_7805,N_7416);
xor U8603 (N_8603,N_7775,N_7703);
nand U8604 (N_8604,N_7521,N_7624);
and U8605 (N_8605,N_7193,N_7477);
and U8606 (N_8606,N_7544,N_7224);
or U8607 (N_8607,N_7468,N_7768);
or U8608 (N_8608,N_7223,N_7359);
xor U8609 (N_8609,N_7200,N_7565);
or U8610 (N_8610,N_7527,N_7851);
xnor U8611 (N_8611,N_7834,N_7810);
and U8612 (N_8612,N_7549,N_7757);
or U8613 (N_8613,N_7523,N_7236);
and U8614 (N_8614,N_7896,N_7022);
and U8615 (N_8615,N_7617,N_7368);
nor U8616 (N_8616,N_7846,N_7618);
or U8617 (N_8617,N_7387,N_7350);
and U8618 (N_8618,N_7497,N_7619);
and U8619 (N_8619,N_7106,N_7634);
nand U8620 (N_8620,N_7544,N_7483);
and U8621 (N_8621,N_7425,N_7447);
xnor U8622 (N_8622,N_7106,N_7055);
nor U8623 (N_8623,N_7582,N_7441);
and U8624 (N_8624,N_7875,N_7475);
and U8625 (N_8625,N_7150,N_7606);
and U8626 (N_8626,N_7876,N_7029);
nand U8627 (N_8627,N_7793,N_7200);
and U8628 (N_8628,N_7086,N_7270);
and U8629 (N_8629,N_7250,N_7627);
nand U8630 (N_8630,N_7936,N_7102);
nand U8631 (N_8631,N_7412,N_7854);
or U8632 (N_8632,N_7148,N_7308);
nand U8633 (N_8633,N_7374,N_7000);
or U8634 (N_8634,N_7625,N_7797);
nor U8635 (N_8635,N_7719,N_7734);
nor U8636 (N_8636,N_7799,N_7932);
and U8637 (N_8637,N_7410,N_7091);
and U8638 (N_8638,N_7232,N_7582);
and U8639 (N_8639,N_7829,N_7828);
or U8640 (N_8640,N_7688,N_7660);
nor U8641 (N_8641,N_7217,N_7657);
nand U8642 (N_8642,N_7535,N_7684);
or U8643 (N_8643,N_7288,N_7380);
nor U8644 (N_8644,N_7216,N_7133);
and U8645 (N_8645,N_7598,N_7154);
or U8646 (N_8646,N_7011,N_7294);
and U8647 (N_8647,N_7684,N_7735);
nor U8648 (N_8648,N_7930,N_7627);
xor U8649 (N_8649,N_7322,N_7808);
xor U8650 (N_8650,N_7040,N_7207);
nand U8651 (N_8651,N_7767,N_7723);
and U8652 (N_8652,N_7864,N_7186);
nor U8653 (N_8653,N_7307,N_7778);
xnor U8654 (N_8654,N_7187,N_7548);
nand U8655 (N_8655,N_7889,N_7133);
and U8656 (N_8656,N_7715,N_7996);
nor U8657 (N_8657,N_7107,N_7583);
nor U8658 (N_8658,N_7846,N_7776);
nor U8659 (N_8659,N_7937,N_7114);
xor U8660 (N_8660,N_7360,N_7068);
xnor U8661 (N_8661,N_7995,N_7823);
nor U8662 (N_8662,N_7563,N_7692);
xor U8663 (N_8663,N_7343,N_7563);
nand U8664 (N_8664,N_7700,N_7494);
nor U8665 (N_8665,N_7514,N_7101);
nor U8666 (N_8666,N_7280,N_7258);
nor U8667 (N_8667,N_7586,N_7012);
and U8668 (N_8668,N_7351,N_7539);
nand U8669 (N_8669,N_7762,N_7629);
nor U8670 (N_8670,N_7576,N_7712);
and U8671 (N_8671,N_7542,N_7952);
nand U8672 (N_8672,N_7017,N_7045);
xnor U8673 (N_8673,N_7585,N_7494);
nand U8674 (N_8674,N_7410,N_7935);
nand U8675 (N_8675,N_7070,N_7517);
nand U8676 (N_8676,N_7054,N_7298);
nand U8677 (N_8677,N_7597,N_7871);
or U8678 (N_8678,N_7301,N_7381);
and U8679 (N_8679,N_7980,N_7087);
nand U8680 (N_8680,N_7433,N_7496);
or U8681 (N_8681,N_7028,N_7152);
nand U8682 (N_8682,N_7363,N_7443);
xnor U8683 (N_8683,N_7141,N_7685);
nor U8684 (N_8684,N_7915,N_7556);
xnor U8685 (N_8685,N_7872,N_7134);
and U8686 (N_8686,N_7566,N_7515);
nand U8687 (N_8687,N_7143,N_7190);
nand U8688 (N_8688,N_7087,N_7397);
xor U8689 (N_8689,N_7155,N_7858);
nor U8690 (N_8690,N_7406,N_7287);
or U8691 (N_8691,N_7744,N_7634);
nand U8692 (N_8692,N_7587,N_7553);
and U8693 (N_8693,N_7686,N_7197);
or U8694 (N_8694,N_7333,N_7539);
nor U8695 (N_8695,N_7769,N_7394);
xnor U8696 (N_8696,N_7872,N_7376);
nor U8697 (N_8697,N_7434,N_7983);
and U8698 (N_8698,N_7151,N_7561);
nand U8699 (N_8699,N_7812,N_7563);
nor U8700 (N_8700,N_7428,N_7968);
and U8701 (N_8701,N_7976,N_7931);
xor U8702 (N_8702,N_7189,N_7123);
or U8703 (N_8703,N_7539,N_7590);
nor U8704 (N_8704,N_7507,N_7176);
or U8705 (N_8705,N_7848,N_7835);
nor U8706 (N_8706,N_7992,N_7464);
nor U8707 (N_8707,N_7536,N_7294);
nand U8708 (N_8708,N_7963,N_7642);
nor U8709 (N_8709,N_7584,N_7145);
or U8710 (N_8710,N_7429,N_7355);
or U8711 (N_8711,N_7467,N_7977);
nor U8712 (N_8712,N_7031,N_7256);
nor U8713 (N_8713,N_7826,N_7265);
and U8714 (N_8714,N_7735,N_7678);
or U8715 (N_8715,N_7584,N_7783);
xnor U8716 (N_8716,N_7541,N_7307);
or U8717 (N_8717,N_7219,N_7724);
or U8718 (N_8718,N_7172,N_7878);
nand U8719 (N_8719,N_7810,N_7413);
xnor U8720 (N_8720,N_7870,N_7659);
nand U8721 (N_8721,N_7697,N_7104);
or U8722 (N_8722,N_7041,N_7689);
and U8723 (N_8723,N_7525,N_7415);
and U8724 (N_8724,N_7451,N_7080);
and U8725 (N_8725,N_7325,N_7218);
or U8726 (N_8726,N_7067,N_7439);
xnor U8727 (N_8727,N_7145,N_7036);
nand U8728 (N_8728,N_7558,N_7386);
nand U8729 (N_8729,N_7486,N_7742);
or U8730 (N_8730,N_7506,N_7743);
nand U8731 (N_8731,N_7919,N_7152);
or U8732 (N_8732,N_7816,N_7434);
nand U8733 (N_8733,N_7116,N_7283);
nand U8734 (N_8734,N_7712,N_7671);
nor U8735 (N_8735,N_7035,N_7287);
nand U8736 (N_8736,N_7418,N_7389);
xnor U8737 (N_8737,N_7646,N_7943);
nor U8738 (N_8738,N_7463,N_7551);
xor U8739 (N_8739,N_7345,N_7341);
nor U8740 (N_8740,N_7494,N_7274);
xor U8741 (N_8741,N_7399,N_7376);
and U8742 (N_8742,N_7918,N_7949);
nor U8743 (N_8743,N_7014,N_7987);
and U8744 (N_8744,N_7558,N_7954);
and U8745 (N_8745,N_7705,N_7152);
nor U8746 (N_8746,N_7483,N_7310);
nand U8747 (N_8747,N_7979,N_7242);
and U8748 (N_8748,N_7976,N_7155);
and U8749 (N_8749,N_7481,N_7014);
or U8750 (N_8750,N_7686,N_7644);
and U8751 (N_8751,N_7822,N_7381);
or U8752 (N_8752,N_7321,N_7624);
or U8753 (N_8753,N_7929,N_7884);
xor U8754 (N_8754,N_7373,N_7197);
and U8755 (N_8755,N_7978,N_7244);
xnor U8756 (N_8756,N_7638,N_7708);
nor U8757 (N_8757,N_7502,N_7772);
and U8758 (N_8758,N_7415,N_7368);
or U8759 (N_8759,N_7026,N_7321);
or U8760 (N_8760,N_7784,N_7905);
or U8761 (N_8761,N_7475,N_7074);
and U8762 (N_8762,N_7269,N_7818);
xor U8763 (N_8763,N_7513,N_7305);
and U8764 (N_8764,N_7318,N_7743);
or U8765 (N_8765,N_7209,N_7988);
nor U8766 (N_8766,N_7515,N_7656);
nand U8767 (N_8767,N_7949,N_7139);
nand U8768 (N_8768,N_7262,N_7044);
nand U8769 (N_8769,N_7757,N_7352);
or U8770 (N_8770,N_7840,N_7010);
xor U8771 (N_8771,N_7705,N_7715);
nor U8772 (N_8772,N_7565,N_7878);
or U8773 (N_8773,N_7211,N_7728);
or U8774 (N_8774,N_7578,N_7142);
and U8775 (N_8775,N_7252,N_7796);
and U8776 (N_8776,N_7985,N_7917);
or U8777 (N_8777,N_7415,N_7255);
nor U8778 (N_8778,N_7728,N_7115);
and U8779 (N_8779,N_7989,N_7982);
or U8780 (N_8780,N_7800,N_7636);
nor U8781 (N_8781,N_7927,N_7541);
xnor U8782 (N_8782,N_7861,N_7653);
or U8783 (N_8783,N_7860,N_7117);
and U8784 (N_8784,N_7538,N_7274);
nand U8785 (N_8785,N_7519,N_7520);
nor U8786 (N_8786,N_7446,N_7948);
nand U8787 (N_8787,N_7193,N_7214);
xor U8788 (N_8788,N_7639,N_7645);
or U8789 (N_8789,N_7701,N_7313);
and U8790 (N_8790,N_7304,N_7923);
xor U8791 (N_8791,N_7362,N_7140);
nand U8792 (N_8792,N_7300,N_7850);
nand U8793 (N_8793,N_7361,N_7236);
xor U8794 (N_8794,N_7766,N_7784);
or U8795 (N_8795,N_7173,N_7204);
and U8796 (N_8796,N_7000,N_7698);
or U8797 (N_8797,N_7837,N_7198);
nand U8798 (N_8798,N_7343,N_7611);
xor U8799 (N_8799,N_7803,N_7123);
xnor U8800 (N_8800,N_7139,N_7763);
and U8801 (N_8801,N_7028,N_7237);
and U8802 (N_8802,N_7534,N_7858);
nor U8803 (N_8803,N_7768,N_7366);
or U8804 (N_8804,N_7775,N_7841);
nand U8805 (N_8805,N_7665,N_7869);
nor U8806 (N_8806,N_7456,N_7582);
and U8807 (N_8807,N_7658,N_7301);
and U8808 (N_8808,N_7311,N_7686);
xor U8809 (N_8809,N_7467,N_7585);
and U8810 (N_8810,N_7020,N_7786);
or U8811 (N_8811,N_7896,N_7522);
nand U8812 (N_8812,N_7508,N_7556);
xnor U8813 (N_8813,N_7134,N_7141);
and U8814 (N_8814,N_7293,N_7348);
and U8815 (N_8815,N_7015,N_7919);
and U8816 (N_8816,N_7389,N_7094);
nand U8817 (N_8817,N_7790,N_7120);
or U8818 (N_8818,N_7055,N_7610);
and U8819 (N_8819,N_7280,N_7925);
or U8820 (N_8820,N_7541,N_7188);
and U8821 (N_8821,N_7450,N_7428);
or U8822 (N_8822,N_7598,N_7908);
xor U8823 (N_8823,N_7730,N_7010);
xnor U8824 (N_8824,N_7808,N_7670);
xor U8825 (N_8825,N_7948,N_7206);
xor U8826 (N_8826,N_7276,N_7422);
xnor U8827 (N_8827,N_7672,N_7341);
nor U8828 (N_8828,N_7506,N_7063);
or U8829 (N_8829,N_7609,N_7647);
or U8830 (N_8830,N_7133,N_7249);
xor U8831 (N_8831,N_7466,N_7463);
or U8832 (N_8832,N_7104,N_7836);
nor U8833 (N_8833,N_7698,N_7057);
or U8834 (N_8834,N_7149,N_7155);
xor U8835 (N_8835,N_7636,N_7698);
and U8836 (N_8836,N_7306,N_7223);
or U8837 (N_8837,N_7455,N_7283);
nor U8838 (N_8838,N_7136,N_7352);
nand U8839 (N_8839,N_7006,N_7877);
nand U8840 (N_8840,N_7741,N_7018);
xor U8841 (N_8841,N_7175,N_7669);
and U8842 (N_8842,N_7804,N_7883);
and U8843 (N_8843,N_7112,N_7539);
and U8844 (N_8844,N_7276,N_7315);
or U8845 (N_8845,N_7389,N_7133);
nand U8846 (N_8846,N_7608,N_7764);
or U8847 (N_8847,N_7081,N_7136);
or U8848 (N_8848,N_7266,N_7121);
and U8849 (N_8849,N_7181,N_7714);
nand U8850 (N_8850,N_7669,N_7856);
nand U8851 (N_8851,N_7253,N_7153);
and U8852 (N_8852,N_7188,N_7554);
or U8853 (N_8853,N_7683,N_7057);
and U8854 (N_8854,N_7935,N_7406);
or U8855 (N_8855,N_7140,N_7795);
or U8856 (N_8856,N_7115,N_7702);
nor U8857 (N_8857,N_7044,N_7148);
and U8858 (N_8858,N_7873,N_7388);
and U8859 (N_8859,N_7234,N_7809);
nand U8860 (N_8860,N_7755,N_7344);
or U8861 (N_8861,N_7785,N_7388);
xor U8862 (N_8862,N_7584,N_7192);
xor U8863 (N_8863,N_7745,N_7458);
or U8864 (N_8864,N_7139,N_7830);
nand U8865 (N_8865,N_7045,N_7056);
nor U8866 (N_8866,N_7378,N_7902);
xnor U8867 (N_8867,N_7048,N_7587);
or U8868 (N_8868,N_7570,N_7646);
nor U8869 (N_8869,N_7413,N_7202);
nor U8870 (N_8870,N_7408,N_7868);
and U8871 (N_8871,N_7267,N_7913);
and U8872 (N_8872,N_7279,N_7466);
xnor U8873 (N_8873,N_7427,N_7141);
nor U8874 (N_8874,N_7329,N_7989);
and U8875 (N_8875,N_7698,N_7239);
xor U8876 (N_8876,N_7217,N_7277);
nor U8877 (N_8877,N_7870,N_7546);
and U8878 (N_8878,N_7035,N_7676);
nor U8879 (N_8879,N_7316,N_7466);
or U8880 (N_8880,N_7322,N_7327);
xor U8881 (N_8881,N_7848,N_7139);
or U8882 (N_8882,N_7293,N_7774);
nor U8883 (N_8883,N_7837,N_7148);
and U8884 (N_8884,N_7579,N_7339);
xnor U8885 (N_8885,N_7563,N_7683);
or U8886 (N_8886,N_7263,N_7261);
and U8887 (N_8887,N_7214,N_7952);
and U8888 (N_8888,N_7369,N_7305);
nand U8889 (N_8889,N_7654,N_7262);
or U8890 (N_8890,N_7329,N_7468);
or U8891 (N_8891,N_7063,N_7879);
nand U8892 (N_8892,N_7270,N_7976);
nand U8893 (N_8893,N_7491,N_7305);
xor U8894 (N_8894,N_7079,N_7298);
nor U8895 (N_8895,N_7755,N_7421);
nand U8896 (N_8896,N_7539,N_7039);
nor U8897 (N_8897,N_7162,N_7260);
or U8898 (N_8898,N_7266,N_7802);
nor U8899 (N_8899,N_7016,N_7114);
or U8900 (N_8900,N_7551,N_7185);
or U8901 (N_8901,N_7910,N_7018);
or U8902 (N_8902,N_7495,N_7232);
xor U8903 (N_8903,N_7294,N_7568);
xnor U8904 (N_8904,N_7785,N_7702);
nand U8905 (N_8905,N_7946,N_7132);
or U8906 (N_8906,N_7545,N_7118);
or U8907 (N_8907,N_7179,N_7657);
and U8908 (N_8908,N_7322,N_7629);
xor U8909 (N_8909,N_7849,N_7854);
nand U8910 (N_8910,N_7470,N_7465);
nand U8911 (N_8911,N_7913,N_7780);
xnor U8912 (N_8912,N_7022,N_7118);
nand U8913 (N_8913,N_7675,N_7408);
nand U8914 (N_8914,N_7912,N_7503);
nand U8915 (N_8915,N_7333,N_7614);
nand U8916 (N_8916,N_7325,N_7609);
nor U8917 (N_8917,N_7477,N_7367);
and U8918 (N_8918,N_7003,N_7134);
or U8919 (N_8919,N_7845,N_7574);
xnor U8920 (N_8920,N_7864,N_7641);
nor U8921 (N_8921,N_7929,N_7145);
xnor U8922 (N_8922,N_7139,N_7874);
and U8923 (N_8923,N_7782,N_7640);
and U8924 (N_8924,N_7701,N_7458);
and U8925 (N_8925,N_7250,N_7994);
and U8926 (N_8926,N_7116,N_7953);
nor U8927 (N_8927,N_7598,N_7922);
nor U8928 (N_8928,N_7378,N_7885);
nand U8929 (N_8929,N_7839,N_7196);
nor U8930 (N_8930,N_7008,N_7452);
nor U8931 (N_8931,N_7136,N_7366);
or U8932 (N_8932,N_7586,N_7890);
nand U8933 (N_8933,N_7398,N_7010);
nor U8934 (N_8934,N_7354,N_7113);
xnor U8935 (N_8935,N_7340,N_7766);
nor U8936 (N_8936,N_7872,N_7055);
and U8937 (N_8937,N_7513,N_7821);
or U8938 (N_8938,N_7259,N_7191);
nand U8939 (N_8939,N_7467,N_7906);
nand U8940 (N_8940,N_7582,N_7170);
nor U8941 (N_8941,N_7853,N_7785);
or U8942 (N_8942,N_7100,N_7389);
xor U8943 (N_8943,N_7748,N_7515);
and U8944 (N_8944,N_7295,N_7212);
xor U8945 (N_8945,N_7064,N_7163);
nor U8946 (N_8946,N_7344,N_7149);
or U8947 (N_8947,N_7696,N_7300);
nand U8948 (N_8948,N_7260,N_7054);
or U8949 (N_8949,N_7788,N_7956);
and U8950 (N_8950,N_7064,N_7967);
nand U8951 (N_8951,N_7665,N_7615);
and U8952 (N_8952,N_7712,N_7692);
and U8953 (N_8953,N_7402,N_7800);
nand U8954 (N_8954,N_7702,N_7866);
xnor U8955 (N_8955,N_7999,N_7050);
nor U8956 (N_8956,N_7660,N_7254);
nand U8957 (N_8957,N_7938,N_7353);
nand U8958 (N_8958,N_7773,N_7448);
xnor U8959 (N_8959,N_7773,N_7073);
xnor U8960 (N_8960,N_7294,N_7256);
nor U8961 (N_8961,N_7802,N_7939);
xor U8962 (N_8962,N_7802,N_7679);
or U8963 (N_8963,N_7231,N_7717);
xnor U8964 (N_8964,N_7209,N_7159);
and U8965 (N_8965,N_7879,N_7164);
nand U8966 (N_8966,N_7049,N_7162);
and U8967 (N_8967,N_7878,N_7687);
nor U8968 (N_8968,N_7275,N_7670);
xor U8969 (N_8969,N_7977,N_7573);
nand U8970 (N_8970,N_7101,N_7832);
nor U8971 (N_8971,N_7914,N_7985);
xor U8972 (N_8972,N_7955,N_7818);
and U8973 (N_8973,N_7381,N_7097);
and U8974 (N_8974,N_7053,N_7277);
xnor U8975 (N_8975,N_7126,N_7773);
or U8976 (N_8976,N_7198,N_7159);
xor U8977 (N_8977,N_7338,N_7389);
nand U8978 (N_8978,N_7436,N_7566);
and U8979 (N_8979,N_7686,N_7701);
and U8980 (N_8980,N_7176,N_7047);
nand U8981 (N_8981,N_7177,N_7314);
and U8982 (N_8982,N_7471,N_7850);
nand U8983 (N_8983,N_7310,N_7033);
nand U8984 (N_8984,N_7177,N_7590);
and U8985 (N_8985,N_7870,N_7033);
xnor U8986 (N_8986,N_7153,N_7914);
xnor U8987 (N_8987,N_7464,N_7443);
nor U8988 (N_8988,N_7975,N_7441);
xor U8989 (N_8989,N_7770,N_7598);
and U8990 (N_8990,N_7457,N_7771);
nor U8991 (N_8991,N_7743,N_7119);
nand U8992 (N_8992,N_7657,N_7635);
or U8993 (N_8993,N_7217,N_7113);
nand U8994 (N_8994,N_7198,N_7336);
xor U8995 (N_8995,N_7244,N_7694);
and U8996 (N_8996,N_7793,N_7148);
and U8997 (N_8997,N_7218,N_7377);
nor U8998 (N_8998,N_7174,N_7034);
and U8999 (N_8999,N_7375,N_7954);
nand U9000 (N_9000,N_8318,N_8894);
and U9001 (N_9001,N_8736,N_8222);
nand U9002 (N_9002,N_8740,N_8492);
or U9003 (N_9003,N_8432,N_8677);
nand U9004 (N_9004,N_8914,N_8895);
nand U9005 (N_9005,N_8235,N_8339);
or U9006 (N_9006,N_8147,N_8421);
nand U9007 (N_9007,N_8460,N_8859);
nor U9008 (N_9008,N_8933,N_8729);
xor U9009 (N_9009,N_8756,N_8488);
and U9010 (N_9010,N_8745,N_8277);
and U9011 (N_9011,N_8387,N_8417);
or U9012 (N_9012,N_8509,N_8924);
nor U9013 (N_9013,N_8600,N_8438);
nor U9014 (N_9014,N_8798,N_8270);
and U9015 (N_9015,N_8682,N_8818);
nand U9016 (N_9016,N_8987,N_8319);
and U9017 (N_9017,N_8060,N_8086);
or U9018 (N_9018,N_8253,N_8074);
or U9019 (N_9019,N_8344,N_8370);
nand U9020 (N_9020,N_8940,N_8218);
nor U9021 (N_9021,N_8008,N_8288);
nand U9022 (N_9022,N_8955,N_8590);
xnor U9023 (N_9023,N_8063,N_8337);
and U9024 (N_9024,N_8472,N_8484);
and U9025 (N_9025,N_8949,N_8988);
and U9026 (N_9026,N_8236,N_8816);
nor U9027 (N_9027,N_8813,N_8611);
nor U9028 (N_9028,N_8331,N_8477);
and U9029 (N_9029,N_8992,N_8698);
nor U9030 (N_9030,N_8011,N_8833);
and U9031 (N_9031,N_8877,N_8025);
and U9032 (N_9032,N_8479,N_8462);
and U9033 (N_9033,N_8545,N_8657);
or U9034 (N_9034,N_8773,N_8765);
or U9035 (N_9035,N_8723,N_8350);
and U9036 (N_9036,N_8822,N_8364);
and U9037 (N_9037,N_8367,N_8125);
nor U9038 (N_9038,N_8978,N_8839);
nand U9039 (N_9039,N_8070,N_8834);
nand U9040 (N_9040,N_8827,N_8412);
or U9041 (N_9041,N_8369,N_8466);
nand U9042 (N_9042,N_8075,N_8298);
xnor U9043 (N_9043,N_8844,N_8311);
nor U9044 (N_9044,N_8631,N_8137);
nor U9045 (N_9045,N_8242,N_8216);
xnor U9046 (N_9046,N_8393,N_8644);
and U9047 (N_9047,N_8335,N_8101);
nand U9048 (N_9048,N_8416,N_8610);
or U9049 (N_9049,N_8341,N_8150);
nand U9050 (N_9050,N_8093,N_8800);
and U9051 (N_9051,N_8155,N_8574);
nand U9052 (N_9052,N_8221,N_8860);
xnor U9053 (N_9053,N_8095,N_8603);
nor U9054 (N_9054,N_8098,N_8983);
nand U9055 (N_9055,N_8120,N_8510);
or U9056 (N_9056,N_8379,N_8414);
nand U9057 (N_9057,N_8708,N_8751);
or U9058 (N_9058,N_8343,N_8871);
xnor U9059 (N_9059,N_8825,N_8501);
nand U9060 (N_9060,N_8539,N_8680);
and U9061 (N_9061,N_8009,N_8873);
nand U9062 (N_9062,N_8586,N_8964);
and U9063 (N_9063,N_8465,N_8498);
nor U9064 (N_9064,N_8205,N_8258);
or U9065 (N_9065,N_8937,N_8958);
and U9066 (N_9066,N_8374,N_8490);
nor U9067 (N_9067,N_8685,N_8872);
and U9068 (N_9068,N_8255,N_8938);
or U9069 (N_9069,N_8832,N_8826);
xnor U9070 (N_9070,N_8170,N_8007);
xnor U9071 (N_9071,N_8293,N_8476);
and U9072 (N_9072,N_8806,N_8819);
nor U9073 (N_9073,N_8925,N_8415);
or U9074 (N_9074,N_8409,N_8457);
and U9075 (N_9075,N_8923,N_8652);
nor U9076 (N_9076,N_8398,N_8783);
xnor U9077 (N_9077,N_8779,N_8139);
or U9078 (N_9078,N_8107,N_8560);
nor U9079 (N_9079,N_8148,N_8434);
and U9080 (N_9080,N_8194,N_8902);
or U9081 (N_9081,N_8252,N_8720);
xnor U9082 (N_9082,N_8089,N_8407);
nand U9083 (N_9083,N_8926,N_8525);
or U9084 (N_9084,N_8592,N_8024);
and U9085 (N_9085,N_8468,N_8100);
xnor U9086 (N_9086,N_8977,N_8061);
or U9087 (N_9087,N_8917,N_8506);
xnor U9088 (N_9088,N_8368,N_8326);
nand U9089 (N_9089,N_8947,N_8934);
and U9090 (N_9090,N_8687,N_8542);
xor U9091 (N_9091,N_8126,N_8463);
nor U9092 (N_9092,N_8874,N_8799);
nor U9093 (N_9093,N_8360,N_8559);
or U9094 (N_9094,N_8880,N_8742);
nor U9095 (N_9095,N_8608,N_8786);
nor U9096 (N_9096,N_8726,N_8516);
and U9097 (N_9097,N_8951,N_8553);
xor U9098 (N_9098,N_8596,N_8225);
and U9099 (N_9099,N_8283,N_8012);
nand U9100 (N_9100,N_8437,N_8519);
or U9101 (N_9101,N_8733,N_8342);
xor U9102 (N_9102,N_8849,N_8946);
and U9103 (N_9103,N_8156,N_8950);
or U9104 (N_9104,N_8327,N_8357);
or U9105 (N_9105,N_8200,N_8470);
nand U9106 (N_9106,N_8758,N_8634);
and U9107 (N_9107,N_8188,N_8371);
and U9108 (N_9108,N_8079,N_8239);
nand U9109 (N_9109,N_8418,N_8683);
or U9110 (N_9110,N_8062,N_8856);
xor U9111 (N_9111,N_8945,N_8588);
and U9112 (N_9112,N_8004,N_8899);
or U9113 (N_9113,N_8186,N_8980);
or U9114 (N_9114,N_8276,N_8797);
nor U9115 (N_9115,N_8931,N_8215);
and U9116 (N_9116,N_8151,N_8046);
nor U9117 (N_9117,N_8648,N_8065);
nor U9118 (N_9118,N_8246,N_8203);
nor U9119 (N_9119,N_8781,N_8010);
nand U9120 (N_9120,N_8442,N_8094);
xnor U9121 (N_9121,N_8626,N_8981);
nor U9122 (N_9122,N_8140,N_8537);
nand U9123 (N_9123,N_8660,N_8824);
xnor U9124 (N_9124,N_8124,N_8443);
and U9125 (N_9125,N_8961,N_8994);
xor U9126 (N_9126,N_8759,N_8702);
nand U9127 (N_9127,N_8535,N_8718);
and U9128 (N_9128,N_8753,N_8711);
or U9129 (N_9129,N_8295,N_8345);
xnor U9130 (N_9130,N_8482,N_8817);
nor U9131 (N_9131,N_8142,N_8640);
or U9132 (N_9132,N_8320,N_8868);
or U9133 (N_9133,N_8424,N_8068);
or U9134 (N_9134,N_8830,N_8807);
nand U9135 (N_9135,N_8309,N_8523);
or U9136 (N_9136,N_8558,N_8582);
and U9137 (N_9137,N_8738,N_8966);
or U9138 (N_9138,N_8570,N_8267);
nand U9139 (N_9139,N_8731,N_8475);
nand U9140 (N_9140,N_8069,N_8767);
nor U9141 (N_9141,N_8347,N_8426);
xnor U9142 (N_9142,N_8549,N_8885);
nor U9143 (N_9143,N_8499,N_8129);
nor U9144 (N_9144,N_8187,N_8670);
xor U9145 (N_9145,N_8245,N_8551);
nor U9146 (N_9146,N_8518,N_8845);
nand U9147 (N_9147,N_8587,N_8546);
xnor U9148 (N_9148,N_8423,N_8152);
nand U9149 (N_9149,N_8058,N_8659);
nor U9150 (N_9150,N_8021,N_8449);
nor U9151 (N_9151,N_8508,N_8392);
xnor U9152 (N_9152,N_8285,N_8281);
xnor U9153 (N_9153,N_8425,N_8990);
nor U9154 (N_9154,N_8780,N_8037);
nor U9155 (N_9155,N_8422,N_8909);
or U9156 (N_9156,N_8384,N_8540);
or U9157 (N_9157,N_8633,N_8127);
nand U9158 (N_9158,N_8183,N_8497);
nand U9159 (N_9159,N_8158,N_8473);
xnor U9160 (N_9160,N_8199,N_8308);
nand U9161 (N_9161,N_8864,N_8378);
or U9162 (N_9162,N_8340,N_8420);
or U9163 (N_9163,N_8448,N_8145);
nand U9164 (N_9164,N_8583,N_8930);
nand U9165 (N_9165,N_8777,N_8632);
and U9166 (N_9166,N_8348,N_8865);
nand U9167 (N_9167,N_8211,N_8134);
xnor U9168 (N_9168,N_8628,N_8247);
xnor U9169 (N_9169,N_8858,N_8483);
nor U9170 (N_9170,N_8645,N_8737);
and U9171 (N_9171,N_8389,N_8333);
nor U9172 (N_9172,N_8505,N_8260);
nor U9173 (N_9173,N_8787,N_8695);
or U9174 (N_9174,N_8027,N_8249);
or U9175 (N_9175,N_8122,N_8087);
xnor U9176 (N_9176,N_8898,N_8030);
or U9177 (N_9177,N_8566,N_8772);
and U9178 (N_9178,N_8679,N_8085);
and U9179 (N_9179,N_8986,N_8612);
and U9180 (N_9180,N_8663,N_8688);
nor U9181 (N_9181,N_8039,N_8793);
or U9182 (N_9182,N_8624,N_8495);
nand U9183 (N_9183,N_8848,N_8257);
nand U9184 (N_9184,N_8173,N_8213);
nor U9185 (N_9185,N_8067,N_8489);
nand U9186 (N_9186,N_8703,N_8684);
and U9187 (N_9187,N_8710,N_8905);
nor U9188 (N_9188,N_8761,N_8439);
or U9189 (N_9189,N_8664,N_8323);
xor U9190 (N_9190,N_8513,N_8804);
nand U9191 (N_9191,N_8565,N_8287);
nand U9192 (N_9192,N_8223,N_8694);
nand U9193 (N_9193,N_8176,N_8597);
xor U9194 (N_9194,N_8088,N_8296);
and U9195 (N_9195,N_8271,N_8689);
nand U9196 (N_9196,N_8890,N_8748);
nand U9197 (N_9197,N_8811,N_8328);
or U9198 (N_9198,N_8397,N_8228);
xor U9199 (N_9199,N_8055,N_8831);
and U9200 (N_9200,N_8109,N_8051);
and U9201 (N_9201,N_8855,N_8707);
xnor U9202 (N_9202,N_8942,N_8604);
nand U9203 (N_9203,N_8891,N_8517);
or U9204 (N_9204,N_8968,N_8979);
xnor U9205 (N_9205,N_8638,N_8321);
nor U9206 (N_9206,N_8447,N_8478);
xor U9207 (N_9207,N_8507,N_8214);
xor U9208 (N_9208,N_8117,N_8690);
and U9209 (N_9209,N_8362,N_8430);
and U9210 (N_9210,N_8863,N_8927);
nand U9211 (N_9211,N_8149,N_8607);
xor U9212 (N_9212,N_8274,N_8240);
nand U9213 (N_9213,N_8103,N_8036);
xor U9214 (N_9214,N_8163,N_8042);
nor U9215 (N_9215,N_8372,N_8616);
nand U9216 (N_9216,N_8629,N_8232);
xnor U9217 (N_9217,N_8269,N_8573);
nor U9218 (N_9218,N_8224,N_8052);
xnor U9219 (N_9219,N_8212,N_8165);
nand U9220 (N_9220,N_8172,N_8901);
and U9221 (N_9221,N_8835,N_8598);
and U9222 (N_9222,N_8280,N_8837);
and U9223 (N_9223,N_8536,N_8643);
xnor U9224 (N_9224,N_8303,N_8716);
xor U9225 (N_9225,N_8493,N_8119);
or U9226 (N_9226,N_8778,N_8091);
xor U9227 (N_9227,N_8918,N_8671);
nand U9228 (N_9228,N_8975,N_8678);
nor U9229 (N_9229,N_8047,N_8013);
xor U9230 (N_9230,N_8965,N_8850);
xor U9231 (N_9231,N_8291,N_8441);
xor U9232 (N_9232,N_8693,N_8001);
xnor U9233 (N_9233,N_8656,N_8529);
nor U9234 (N_9234,N_8511,N_8166);
and U9235 (N_9235,N_8615,N_8264);
nor U9236 (N_9236,N_8391,N_8076);
or U9237 (N_9237,N_8712,N_8016);
xnor U9238 (N_9238,N_8960,N_8485);
nand U9239 (N_9239,N_8233,N_8550);
or U9240 (N_9240,N_8760,N_8580);
or U9241 (N_9241,N_8408,N_8669);
or U9242 (N_9242,N_8450,N_8622);
nand U9243 (N_9243,N_8038,N_8724);
nor U9244 (N_9244,N_8658,N_8429);
and U9245 (N_9245,N_8533,N_8775);
and U9246 (N_9246,N_8512,N_8732);
nand U9247 (N_9247,N_8202,N_8851);
and U9248 (N_9248,N_8705,N_8941);
and U9249 (N_9249,N_8359,N_8044);
nor U9250 (N_9250,N_8538,N_8770);
xnor U9251 (N_9251,N_8018,N_8962);
or U9252 (N_9252,N_8217,N_8469);
and U9253 (N_9253,N_8717,N_8916);
xor U9254 (N_9254,N_8179,N_8900);
xor U9255 (N_9255,N_8358,N_8180);
xor U9256 (N_9256,N_8380,N_8821);
xor U9257 (N_9257,N_8956,N_8105);
nor U9258 (N_9258,N_8195,N_8167);
or U9259 (N_9259,N_8810,N_8351);
and U9260 (N_9260,N_8329,N_8504);
and U9261 (N_9261,N_8883,N_8735);
xnor U9262 (N_9262,N_8936,N_8790);
nor U9263 (N_9263,N_8928,N_8279);
or U9264 (N_9264,N_8268,N_8130);
or U9265 (N_9265,N_8273,N_8486);
and U9266 (N_9266,N_8118,N_8991);
or U9267 (N_9267,N_8602,N_8154);
or U9268 (N_9268,N_8569,N_8861);
or U9269 (N_9269,N_8814,N_8033);
and U9270 (N_9270,N_8520,N_8433);
and U9271 (N_9271,N_8059,N_8593);
and U9272 (N_9272,N_8647,N_8725);
nand U9273 (N_9273,N_8701,N_8576);
or U9274 (N_9274,N_8177,N_8557);
and U9275 (N_9275,N_8757,N_8887);
nand U9276 (N_9276,N_8244,N_8719);
nor U9277 (N_9277,N_8621,N_8164);
and U9278 (N_9278,N_8043,N_8266);
nor U9279 (N_9279,N_8912,N_8561);
or U9280 (N_9280,N_8932,N_8136);
or U9281 (N_9281,N_8886,N_8704);
nand U9282 (N_9282,N_8769,N_8792);
or U9283 (N_9283,N_8455,N_8275);
and U9284 (N_9284,N_8528,N_8642);
nor U9285 (N_9285,N_8714,N_8096);
and U9286 (N_9286,N_8458,N_8402);
nand U9287 (N_9287,N_8325,N_8355);
and U9288 (N_9288,N_8954,N_8383);
and U9289 (N_9289,N_8706,N_8471);
and U9290 (N_9290,N_8084,N_8286);
nand U9291 (N_9291,N_8263,N_8999);
and U9292 (N_9292,N_8929,N_8168);
and U9293 (N_9293,N_8637,N_8795);
xnor U9294 (N_9294,N_8989,N_8571);
or U9295 (N_9295,N_8805,N_8750);
nor U9296 (N_9296,N_8906,N_8169);
or U9297 (N_9297,N_8353,N_8843);
and U9298 (N_9298,N_8230,N_8133);
nor U9299 (N_9299,N_8431,N_8330);
and U9300 (N_9300,N_8755,N_8315);
nor U9301 (N_9301,N_8841,N_8803);
and U9302 (N_9302,N_8613,N_8175);
nor U9303 (N_9303,N_8146,N_8655);
or U9304 (N_9304,N_8959,N_8547);
nor U9305 (N_9305,N_8982,N_8451);
xnor U9306 (N_9306,N_8878,N_8413);
nand U9307 (N_9307,N_8153,N_8809);
nand U9308 (N_9308,N_8727,N_8564);
nand U9309 (N_9309,N_8749,N_8635);
nor U9310 (N_9310,N_8522,N_8662);
xor U9311 (N_9311,N_8823,N_8721);
xor U9312 (N_9312,N_8763,N_8627);
or U9313 (N_9313,N_8713,N_8254);
nor U9314 (N_9314,N_8494,N_8884);
or U9315 (N_9315,N_8556,N_8935);
xnor U9316 (N_9316,N_8406,N_8500);
xnor U9317 (N_9317,N_8908,N_8141);
nor U9318 (N_9318,N_8382,N_8882);
nand U9319 (N_9319,N_8577,N_8159);
or U9320 (N_9320,N_8534,N_8114);
xnor U9321 (N_9321,N_8893,N_8503);
nor U9322 (N_9322,N_8636,N_8005);
or U9323 (N_9323,N_8306,N_8840);
xnor U9324 (N_9324,N_8390,N_8080);
or U9325 (N_9325,N_8896,N_8796);
nor U9326 (N_9326,N_8752,N_8722);
and U9327 (N_9327,N_8282,N_8913);
or U9328 (N_9328,N_8446,N_8229);
xnor U9329 (N_9329,N_8665,N_8491);
and U9330 (N_9330,N_8404,N_8820);
and U9331 (N_9331,N_8456,N_8915);
nand U9332 (N_9332,N_8502,N_8191);
and U9333 (N_9333,N_8548,N_8715);
or U9334 (N_9334,N_8334,N_8029);
xor U9335 (N_9335,N_8623,N_8160);
xor U9336 (N_9336,N_8197,N_8072);
nor U9337 (N_9337,N_8606,N_8836);
xor U9338 (N_9338,N_8651,N_8113);
and U9339 (N_9339,N_8405,N_8041);
nand U9340 (N_9340,N_8003,N_8970);
and U9341 (N_9341,N_8815,N_8461);
xor U9342 (N_9342,N_8251,N_8681);
nor U9343 (N_9343,N_8324,N_8852);
nor U9344 (N_9344,N_8314,N_8206);
and U9345 (N_9345,N_8782,N_8161);
and U9346 (N_9346,N_8675,N_8768);
nand U9347 (N_9347,N_8115,N_8543);
and U9348 (N_9348,N_8121,N_8944);
xor U9349 (N_9349,N_8377,N_8237);
and U9350 (N_9350,N_8248,N_8625);
nand U9351 (N_9351,N_8995,N_8238);
xnor U9352 (N_9352,N_8744,N_8365);
nand U9353 (N_9353,N_8317,N_8650);
nor U9354 (N_9354,N_8198,N_8278);
nor U9355 (N_9355,N_8376,N_8174);
xnor U9356 (N_9356,N_8017,N_8952);
xnor U9357 (N_9357,N_8272,N_8081);
or U9358 (N_9358,N_8862,N_8210);
nor U9359 (N_9359,N_8881,N_8297);
nor U9360 (N_9360,N_8572,N_8053);
nor U9361 (N_9361,N_8667,N_8019);
nor U9362 (N_9362,N_8903,N_8265);
nand U9363 (N_9363,N_8747,N_8897);
and U9364 (N_9364,N_8774,N_8403);
nand U9365 (N_9365,N_8974,N_8464);
or U9366 (N_9366,N_8595,N_8791);
and U9367 (N_9367,N_8131,N_8889);
or U9368 (N_9368,N_8436,N_8562);
nor U9369 (N_9369,N_8614,N_8866);
nor U9370 (N_9370,N_8728,N_8661);
nor U9371 (N_9371,N_8301,N_8591);
or U9372 (N_9372,N_8515,N_8739);
nor U9373 (N_9373,N_8386,N_8452);
nand U9374 (N_9374,N_8099,N_8857);
nor U9375 (N_9375,N_8128,N_8162);
nor U9376 (N_9376,N_8459,N_8481);
nor U9377 (N_9377,N_8524,N_8111);
xnor U9378 (N_9378,N_8867,N_8666);
nand U9379 (N_9379,N_8870,N_8123);
or U9380 (N_9380,N_8762,N_8904);
nand U9381 (N_9381,N_8892,N_8444);
and U9382 (N_9382,N_8578,N_8876);
or U9383 (N_9383,N_8567,N_8554);
nand U9384 (N_9384,N_8842,N_8829);
or U9385 (N_9385,N_8589,N_8231);
xnor U9386 (N_9386,N_8599,N_8639);
xor U9387 (N_9387,N_8394,N_8388);
xnor U9388 (N_9388,N_8157,N_8078);
nor U9389 (N_9389,N_8259,N_8854);
nor U9390 (N_9390,N_8015,N_8262);
or U9391 (N_9391,N_8307,N_8056);
xor U9392 (N_9392,N_8646,N_8653);
nor U9393 (N_9393,N_8208,N_8907);
or U9394 (N_9394,N_8346,N_8563);
or U9395 (N_9395,N_8196,N_8801);
or U9396 (N_9396,N_8104,N_8241);
nor U9397 (N_9397,N_8853,N_8869);
nor U9398 (N_9398,N_8294,N_8071);
or U9399 (N_9399,N_8292,N_8190);
and U9400 (N_9400,N_8605,N_8998);
and U9401 (N_9401,N_8911,N_8427);
xor U9402 (N_9402,N_8022,N_8620);
nor U9403 (N_9403,N_8584,N_8073);
xnor U9404 (N_9404,N_8700,N_8879);
nor U9405 (N_9405,N_8976,N_8526);
xor U9406 (N_9406,N_8261,N_8192);
xor U9407 (N_9407,N_8939,N_8997);
xnor U9408 (N_9408,N_8531,N_8207);
or U9409 (N_9409,N_8226,N_8234);
xor U9410 (N_9410,N_8375,N_8676);
xor U9411 (N_9411,N_8741,N_8487);
or U9412 (N_9412,N_8373,N_8184);
nor U9413 (N_9413,N_8026,N_8000);
nand U9414 (N_9414,N_8410,N_8552);
or U9415 (N_9415,N_8771,N_8313);
or U9416 (N_9416,N_8445,N_8138);
xor U9417 (N_9417,N_8672,N_8568);
nor U9418 (N_9418,N_8112,N_8474);
nand U9419 (N_9419,N_8032,N_8002);
xor U9420 (N_9420,N_8692,N_8919);
or U9421 (N_9421,N_8082,N_8064);
xnor U9422 (N_9422,N_8256,N_8077);
xor U9423 (N_9423,N_8035,N_8220);
nor U9424 (N_9424,N_8385,N_8178);
nor U9425 (N_9425,N_8396,N_8921);
xnor U9426 (N_9426,N_8838,N_8579);
nor U9427 (N_9427,N_8544,N_8316);
and U9428 (N_9428,N_8090,N_8312);
nand U9429 (N_9429,N_8144,N_8609);
nand U9430 (N_9430,N_8575,N_8045);
nand U9431 (N_9431,N_8766,N_8289);
or U9432 (N_9432,N_8034,N_8305);
nor U9433 (N_9433,N_8630,N_8135);
nor U9434 (N_9434,N_8182,N_8189);
and U9435 (N_9435,N_8399,N_8828);
nand U9436 (N_9436,N_8601,N_8957);
xnor U9437 (N_9437,N_8785,N_8401);
nand U9438 (N_9438,N_8581,N_8290);
and U9439 (N_9439,N_8764,N_8284);
nor U9440 (N_9440,N_8040,N_8794);
or U9441 (N_9441,N_8668,N_8963);
nor U9442 (N_9442,N_8948,N_8697);
or U9443 (N_9443,N_8299,N_8106);
or U9444 (N_9444,N_8020,N_8943);
xnor U9445 (N_9445,N_8776,N_8699);
nor U9446 (N_9446,N_8338,N_8054);
or U9447 (N_9447,N_8734,N_8641);
nor U9448 (N_9448,N_8453,N_8789);
nor U9449 (N_9449,N_8057,N_8352);
and U9450 (N_9450,N_8310,N_8985);
nand U9451 (N_9451,N_8097,N_8967);
xnor U9452 (N_9452,N_8846,N_8743);
or U9453 (N_9453,N_8322,N_8185);
nor U9454 (N_9454,N_8532,N_8541);
and U9455 (N_9455,N_8521,N_8973);
nand U9456 (N_9456,N_8066,N_8654);
nor U9457 (N_9457,N_8356,N_8784);
nor U9458 (N_9458,N_8048,N_8209);
and U9459 (N_9459,N_8691,N_8440);
nand U9460 (N_9460,N_8204,N_8354);
or U9461 (N_9461,N_8250,N_8050);
xnor U9462 (N_9462,N_8193,N_8730);
nand U9463 (N_9463,N_8496,N_8922);
and U9464 (N_9464,N_8361,N_8302);
xor U9465 (N_9465,N_8108,N_8349);
nand U9466 (N_9466,N_8201,N_8972);
nor U9467 (N_9467,N_8143,N_8686);
and U9468 (N_9468,N_8802,N_8363);
nand U9469 (N_9469,N_8480,N_8411);
nand U9470 (N_9470,N_8102,N_8454);
nor U9471 (N_9471,N_8171,N_8395);
and U9472 (N_9472,N_8181,N_8649);
xor U9473 (N_9473,N_8754,N_8996);
nand U9474 (N_9474,N_8788,N_8746);
nor U9475 (N_9475,N_8092,N_8028);
nor U9476 (N_9476,N_8875,N_8083);
xnor U9477 (N_9477,N_8812,N_8219);
or U9478 (N_9478,N_8619,N_8304);
nand U9479 (N_9479,N_8332,N_8467);
nand U9480 (N_9480,N_8031,N_8530);
nand U9481 (N_9481,N_8618,N_8847);
and U9482 (N_9482,N_8428,N_8585);
or U9483 (N_9483,N_8300,N_8527);
or U9484 (N_9484,N_8049,N_8419);
xnor U9485 (N_9485,N_8617,N_8594);
and U9486 (N_9486,N_8400,N_8381);
nand U9487 (N_9487,N_8920,N_8993);
nor U9488 (N_9488,N_8696,N_8971);
and U9489 (N_9489,N_8116,N_8984);
or U9490 (N_9490,N_8888,N_8514);
nand U9491 (N_9491,N_8969,N_8006);
nand U9492 (N_9492,N_8709,N_8673);
nand U9493 (N_9493,N_8953,N_8014);
nor U9494 (N_9494,N_8243,N_8555);
or U9495 (N_9495,N_8910,N_8132);
nor U9496 (N_9496,N_8110,N_8227);
nor U9497 (N_9497,N_8808,N_8674);
nor U9498 (N_9498,N_8336,N_8366);
or U9499 (N_9499,N_8023,N_8435);
nand U9500 (N_9500,N_8568,N_8179);
nand U9501 (N_9501,N_8098,N_8787);
nand U9502 (N_9502,N_8365,N_8791);
or U9503 (N_9503,N_8632,N_8219);
nand U9504 (N_9504,N_8534,N_8916);
or U9505 (N_9505,N_8003,N_8889);
xor U9506 (N_9506,N_8642,N_8106);
nor U9507 (N_9507,N_8454,N_8857);
xnor U9508 (N_9508,N_8263,N_8753);
nor U9509 (N_9509,N_8027,N_8063);
xor U9510 (N_9510,N_8378,N_8733);
and U9511 (N_9511,N_8483,N_8657);
nor U9512 (N_9512,N_8532,N_8249);
xnor U9513 (N_9513,N_8652,N_8677);
and U9514 (N_9514,N_8672,N_8293);
and U9515 (N_9515,N_8128,N_8230);
nor U9516 (N_9516,N_8800,N_8671);
nor U9517 (N_9517,N_8455,N_8178);
and U9518 (N_9518,N_8855,N_8979);
and U9519 (N_9519,N_8590,N_8439);
or U9520 (N_9520,N_8968,N_8175);
xor U9521 (N_9521,N_8018,N_8094);
nand U9522 (N_9522,N_8806,N_8689);
xor U9523 (N_9523,N_8490,N_8263);
nor U9524 (N_9524,N_8458,N_8725);
nor U9525 (N_9525,N_8059,N_8609);
nand U9526 (N_9526,N_8329,N_8246);
nand U9527 (N_9527,N_8881,N_8506);
nor U9528 (N_9528,N_8877,N_8671);
or U9529 (N_9529,N_8258,N_8405);
nor U9530 (N_9530,N_8076,N_8129);
or U9531 (N_9531,N_8444,N_8205);
and U9532 (N_9532,N_8143,N_8526);
nor U9533 (N_9533,N_8676,N_8715);
or U9534 (N_9534,N_8208,N_8510);
or U9535 (N_9535,N_8301,N_8989);
and U9536 (N_9536,N_8584,N_8235);
or U9537 (N_9537,N_8531,N_8026);
nand U9538 (N_9538,N_8883,N_8474);
xor U9539 (N_9539,N_8896,N_8480);
nor U9540 (N_9540,N_8958,N_8354);
nand U9541 (N_9541,N_8160,N_8373);
or U9542 (N_9542,N_8204,N_8662);
nand U9543 (N_9543,N_8701,N_8968);
nand U9544 (N_9544,N_8800,N_8109);
xor U9545 (N_9545,N_8588,N_8797);
xnor U9546 (N_9546,N_8718,N_8242);
xnor U9547 (N_9547,N_8350,N_8943);
and U9548 (N_9548,N_8923,N_8096);
or U9549 (N_9549,N_8325,N_8525);
nor U9550 (N_9550,N_8045,N_8901);
nor U9551 (N_9551,N_8617,N_8297);
xor U9552 (N_9552,N_8596,N_8381);
and U9553 (N_9553,N_8076,N_8758);
nand U9554 (N_9554,N_8675,N_8873);
nor U9555 (N_9555,N_8150,N_8930);
xor U9556 (N_9556,N_8305,N_8568);
or U9557 (N_9557,N_8680,N_8486);
nor U9558 (N_9558,N_8584,N_8514);
xor U9559 (N_9559,N_8110,N_8621);
nand U9560 (N_9560,N_8946,N_8742);
or U9561 (N_9561,N_8064,N_8528);
or U9562 (N_9562,N_8872,N_8703);
xor U9563 (N_9563,N_8116,N_8437);
or U9564 (N_9564,N_8344,N_8228);
xor U9565 (N_9565,N_8731,N_8736);
nor U9566 (N_9566,N_8126,N_8686);
xnor U9567 (N_9567,N_8419,N_8191);
or U9568 (N_9568,N_8485,N_8070);
or U9569 (N_9569,N_8609,N_8071);
xor U9570 (N_9570,N_8231,N_8852);
and U9571 (N_9571,N_8541,N_8875);
or U9572 (N_9572,N_8734,N_8589);
nor U9573 (N_9573,N_8637,N_8310);
or U9574 (N_9574,N_8752,N_8515);
nand U9575 (N_9575,N_8278,N_8659);
nand U9576 (N_9576,N_8130,N_8763);
nand U9577 (N_9577,N_8476,N_8036);
and U9578 (N_9578,N_8392,N_8142);
and U9579 (N_9579,N_8510,N_8206);
nor U9580 (N_9580,N_8231,N_8673);
nor U9581 (N_9581,N_8386,N_8810);
nand U9582 (N_9582,N_8420,N_8215);
nor U9583 (N_9583,N_8605,N_8409);
nand U9584 (N_9584,N_8604,N_8734);
nor U9585 (N_9585,N_8768,N_8382);
and U9586 (N_9586,N_8141,N_8876);
and U9587 (N_9587,N_8286,N_8280);
nand U9588 (N_9588,N_8860,N_8253);
and U9589 (N_9589,N_8358,N_8140);
or U9590 (N_9590,N_8732,N_8415);
xnor U9591 (N_9591,N_8908,N_8396);
and U9592 (N_9592,N_8121,N_8070);
xor U9593 (N_9593,N_8793,N_8787);
nor U9594 (N_9594,N_8170,N_8526);
nor U9595 (N_9595,N_8999,N_8642);
and U9596 (N_9596,N_8554,N_8982);
nor U9597 (N_9597,N_8839,N_8747);
and U9598 (N_9598,N_8492,N_8524);
and U9599 (N_9599,N_8864,N_8836);
and U9600 (N_9600,N_8289,N_8448);
or U9601 (N_9601,N_8306,N_8686);
nand U9602 (N_9602,N_8177,N_8574);
or U9603 (N_9603,N_8514,N_8513);
or U9604 (N_9604,N_8060,N_8442);
xnor U9605 (N_9605,N_8492,N_8991);
nand U9606 (N_9606,N_8344,N_8714);
xor U9607 (N_9607,N_8690,N_8403);
xnor U9608 (N_9608,N_8870,N_8085);
xor U9609 (N_9609,N_8136,N_8616);
xnor U9610 (N_9610,N_8728,N_8990);
or U9611 (N_9611,N_8690,N_8500);
nor U9612 (N_9612,N_8490,N_8232);
nor U9613 (N_9613,N_8753,N_8150);
xnor U9614 (N_9614,N_8752,N_8391);
nor U9615 (N_9615,N_8562,N_8241);
and U9616 (N_9616,N_8833,N_8594);
and U9617 (N_9617,N_8365,N_8686);
xor U9618 (N_9618,N_8251,N_8249);
and U9619 (N_9619,N_8984,N_8030);
xor U9620 (N_9620,N_8754,N_8647);
or U9621 (N_9621,N_8739,N_8009);
or U9622 (N_9622,N_8073,N_8193);
xor U9623 (N_9623,N_8131,N_8108);
or U9624 (N_9624,N_8766,N_8442);
or U9625 (N_9625,N_8076,N_8260);
xor U9626 (N_9626,N_8406,N_8065);
nor U9627 (N_9627,N_8544,N_8409);
xor U9628 (N_9628,N_8778,N_8730);
nand U9629 (N_9629,N_8892,N_8841);
nor U9630 (N_9630,N_8741,N_8089);
nand U9631 (N_9631,N_8309,N_8200);
and U9632 (N_9632,N_8543,N_8291);
xor U9633 (N_9633,N_8687,N_8089);
nor U9634 (N_9634,N_8449,N_8901);
xnor U9635 (N_9635,N_8183,N_8985);
and U9636 (N_9636,N_8669,N_8995);
or U9637 (N_9637,N_8362,N_8123);
and U9638 (N_9638,N_8623,N_8085);
or U9639 (N_9639,N_8626,N_8054);
nor U9640 (N_9640,N_8645,N_8964);
xnor U9641 (N_9641,N_8848,N_8967);
nand U9642 (N_9642,N_8901,N_8626);
nor U9643 (N_9643,N_8250,N_8340);
or U9644 (N_9644,N_8904,N_8625);
xor U9645 (N_9645,N_8933,N_8593);
and U9646 (N_9646,N_8236,N_8361);
nand U9647 (N_9647,N_8047,N_8740);
nand U9648 (N_9648,N_8495,N_8378);
nand U9649 (N_9649,N_8833,N_8466);
nand U9650 (N_9650,N_8313,N_8208);
xor U9651 (N_9651,N_8117,N_8885);
nor U9652 (N_9652,N_8995,N_8422);
and U9653 (N_9653,N_8011,N_8933);
nor U9654 (N_9654,N_8913,N_8868);
xor U9655 (N_9655,N_8114,N_8495);
xor U9656 (N_9656,N_8630,N_8554);
and U9657 (N_9657,N_8745,N_8231);
and U9658 (N_9658,N_8085,N_8686);
xor U9659 (N_9659,N_8316,N_8221);
and U9660 (N_9660,N_8423,N_8247);
and U9661 (N_9661,N_8637,N_8261);
and U9662 (N_9662,N_8116,N_8431);
xnor U9663 (N_9663,N_8117,N_8352);
and U9664 (N_9664,N_8397,N_8377);
and U9665 (N_9665,N_8137,N_8911);
nand U9666 (N_9666,N_8260,N_8531);
or U9667 (N_9667,N_8318,N_8747);
and U9668 (N_9668,N_8379,N_8085);
and U9669 (N_9669,N_8686,N_8011);
xor U9670 (N_9670,N_8915,N_8384);
or U9671 (N_9671,N_8215,N_8075);
xor U9672 (N_9672,N_8110,N_8870);
nand U9673 (N_9673,N_8357,N_8719);
nand U9674 (N_9674,N_8906,N_8417);
xor U9675 (N_9675,N_8490,N_8304);
and U9676 (N_9676,N_8508,N_8251);
and U9677 (N_9677,N_8823,N_8555);
xnor U9678 (N_9678,N_8685,N_8090);
nor U9679 (N_9679,N_8497,N_8163);
xor U9680 (N_9680,N_8651,N_8983);
nor U9681 (N_9681,N_8984,N_8811);
or U9682 (N_9682,N_8628,N_8342);
and U9683 (N_9683,N_8680,N_8620);
nor U9684 (N_9684,N_8154,N_8021);
and U9685 (N_9685,N_8293,N_8939);
nor U9686 (N_9686,N_8933,N_8536);
and U9687 (N_9687,N_8508,N_8877);
xnor U9688 (N_9688,N_8171,N_8551);
nand U9689 (N_9689,N_8809,N_8262);
or U9690 (N_9690,N_8459,N_8222);
nor U9691 (N_9691,N_8590,N_8995);
and U9692 (N_9692,N_8678,N_8742);
nor U9693 (N_9693,N_8226,N_8673);
or U9694 (N_9694,N_8169,N_8354);
nor U9695 (N_9695,N_8426,N_8108);
or U9696 (N_9696,N_8380,N_8442);
nand U9697 (N_9697,N_8905,N_8108);
nand U9698 (N_9698,N_8267,N_8534);
nand U9699 (N_9699,N_8188,N_8004);
or U9700 (N_9700,N_8406,N_8165);
nand U9701 (N_9701,N_8922,N_8927);
nor U9702 (N_9702,N_8121,N_8208);
and U9703 (N_9703,N_8437,N_8199);
nor U9704 (N_9704,N_8778,N_8249);
and U9705 (N_9705,N_8230,N_8376);
and U9706 (N_9706,N_8114,N_8661);
xnor U9707 (N_9707,N_8841,N_8719);
and U9708 (N_9708,N_8695,N_8731);
or U9709 (N_9709,N_8090,N_8087);
nand U9710 (N_9710,N_8225,N_8918);
xnor U9711 (N_9711,N_8293,N_8812);
nand U9712 (N_9712,N_8114,N_8506);
nand U9713 (N_9713,N_8032,N_8188);
or U9714 (N_9714,N_8164,N_8803);
or U9715 (N_9715,N_8022,N_8356);
nor U9716 (N_9716,N_8519,N_8284);
nand U9717 (N_9717,N_8012,N_8114);
nand U9718 (N_9718,N_8357,N_8195);
xnor U9719 (N_9719,N_8370,N_8395);
xnor U9720 (N_9720,N_8806,N_8353);
or U9721 (N_9721,N_8249,N_8134);
nand U9722 (N_9722,N_8846,N_8212);
or U9723 (N_9723,N_8770,N_8823);
nor U9724 (N_9724,N_8661,N_8162);
xor U9725 (N_9725,N_8628,N_8868);
or U9726 (N_9726,N_8769,N_8525);
nand U9727 (N_9727,N_8760,N_8785);
or U9728 (N_9728,N_8523,N_8367);
or U9729 (N_9729,N_8898,N_8891);
nor U9730 (N_9730,N_8607,N_8068);
nor U9731 (N_9731,N_8077,N_8318);
and U9732 (N_9732,N_8680,N_8007);
nand U9733 (N_9733,N_8741,N_8509);
xor U9734 (N_9734,N_8777,N_8295);
xor U9735 (N_9735,N_8072,N_8297);
and U9736 (N_9736,N_8776,N_8524);
nor U9737 (N_9737,N_8983,N_8924);
or U9738 (N_9738,N_8294,N_8098);
nand U9739 (N_9739,N_8458,N_8163);
nand U9740 (N_9740,N_8620,N_8229);
nand U9741 (N_9741,N_8735,N_8333);
nor U9742 (N_9742,N_8662,N_8267);
nand U9743 (N_9743,N_8053,N_8305);
nor U9744 (N_9744,N_8879,N_8893);
xnor U9745 (N_9745,N_8895,N_8114);
and U9746 (N_9746,N_8844,N_8248);
or U9747 (N_9747,N_8991,N_8797);
or U9748 (N_9748,N_8725,N_8021);
and U9749 (N_9749,N_8636,N_8688);
xnor U9750 (N_9750,N_8994,N_8861);
xor U9751 (N_9751,N_8541,N_8523);
nand U9752 (N_9752,N_8232,N_8848);
nor U9753 (N_9753,N_8944,N_8712);
and U9754 (N_9754,N_8661,N_8307);
nor U9755 (N_9755,N_8168,N_8476);
xor U9756 (N_9756,N_8870,N_8569);
nand U9757 (N_9757,N_8216,N_8853);
xnor U9758 (N_9758,N_8871,N_8408);
or U9759 (N_9759,N_8146,N_8604);
xor U9760 (N_9760,N_8395,N_8180);
and U9761 (N_9761,N_8529,N_8780);
nor U9762 (N_9762,N_8639,N_8148);
and U9763 (N_9763,N_8010,N_8337);
or U9764 (N_9764,N_8286,N_8272);
and U9765 (N_9765,N_8638,N_8726);
and U9766 (N_9766,N_8595,N_8053);
xor U9767 (N_9767,N_8821,N_8847);
or U9768 (N_9768,N_8319,N_8781);
nor U9769 (N_9769,N_8460,N_8697);
nand U9770 (N_9770,N_8210,N_8263);
nand U9771 (N_9771,N_8216,N_8756);
nand U9772 (N_9772,N_8955,N_8377);
nand U9773 (N_9773,N_8585,N_8665);
nand U9774 (N_9774,N_8423,N_8049);
xnor U9775 (N_9775,N_8432,N_8225);
xnor U9776 (N_9776,N_8457,N_8936);
or U9777 (N_9777,N_8711,N_8449);
and U9778 (N_9778,N_8020,N_8796);
xnor U9779 (N_9779,N_8240,N_8658);
or U9780 (N_9780,N_8088,N_8590);
xor U9781 (N_9781,N_8857,N_8634);
nor U9782 (N_9782,N_8612,N_8641);
xnor U9783 (N_9783,N_8541,N_8610);
and U9784 (N_9784,N_8369,N_8269);
and U9785 (N_9785,N_8246,N_8288);
nand U9786 (N_9786,N_8961,N_8083);
nand U9787 (N_9787,N_8627,N_8745);
and U9788 (N_9788,N_8999,N_8384);
xnor U9789 (N_9789,N_8009,N_8229);
or U9790 (N_9790,N_8288,N_8154);
and U9791 (N_9791,N_8987,N_8786);
nand U9792 (N_9792,N_8549,N_8178);
nor U9793 (N_9793,N_8278,N_8544);
xnor U9794 (N_9794,N_8158,N_8843);
nor U9795 (N_9795,N_8455,N_8019);
nor U9796 (N_9796,N_8574,N_8524);
or U9797 (N_9797,N_8399,N_8687);
nand U9798 (N_9798,N_8232,N_8000);
nand U9799 (N_9799,N_8215,N_8877);
and U9800 (N_9800,N_8875,N_8519);
xor U9801 (N_9801,N_8053,N_8088);
nand U9802 (N_9802,N_8269,N_8994);
or U9803 (N_9803,N_8411,N_8999);
xnor U9804 (N_9804,N_8916,N_8354);
nor U9805 (N_9805,N_8538,N_8812);
or U9806 (N_9806,N_8210,N_8587);
nor U9807 (N_9807,N_8709,N_8513);
or U9808 (N_9808,N_8832,N_8132);
nand U9809 (N_9809,N_8483,N_8985);
or U9810 (N_9810,N_8166,N_8429);
and U9811 (N_9811,N_8241,N_8888);
nand U9812 (N_9812,N_8228,N_8282);
xnor U9813 (N_9813,N_8609,N_8912);
and U9814 (N_9814,N_8923,N_8282);
or U9815 (N_9815,N_8865,N_8951);
or U9816 (N_9816,N_8704,N_8621);
or U9817 (N_9817,N_8678,N_8090);
and U9818 (N_9818,N_8538,N_8084);
nor U9819 (N_9819,N_8390,N_8432);
and U9820 (N_9820,N_8002,N_8073);
or U9821 (N_9821,N_8078,N_8658);
and U9822 (N_9822,N_8734,N_8268);
and U9823 (N_9823,N_8254,N_8978);
nor U9824 (N_9824,N_8131,N_8444);
nor U9825 (N_9825,N_8453,N_8582);
and U9826 (N_9826,N_8420,N_8059);
and U9827 (N_9827,N_8432,N_8250);
nand U9828 (N_9828,N_8033,N_8979);
or U9829 (N_9829,N_8237,N_8697);
xnor U9830 (N_9830,N_8204,N_8024);
or U9831 (N_9831,N_8644,N_8326);
xnor U9832 (N_9832,N_8661,N_8901);
and U9833 (N_9833,N_8068,N_8091);
and U9834 (N_9834,N_8388,N_8641);
nor U9835 (N_9835,N_8831,N_8237);
nor U9836 (N_9836,N_8755,N_8325);
and U9837 (N_9837,N_8986,N_8652);
nor U9838 (N_9838,N_8088,N_8561);
or U9839 (N_9839,N_8788,N_8126);
nand U9840 (N_9840,N_8573,N_8655);
xor U9841 (N_9841,N_8399,N_8906);
xor U9842 (N_9842,N_8109,N_8613);
xnor U9843 (N_9843,N_8767,N_8071);
nand U9844 (N_9844,N_8535,N_8667);
nor U9845 (N_9845,N_8801,N_8103);
nor U9846 (N_9846,N_8591,N_8752);
nor U9847 (N_9847,N_8346,N_8041);
xor U9848 (N_9848,N_8064,N_8651);
nor U9849 (N_9849,N_8355,N_8027);
and U9850 (N_9850,N_8720,N_8609);
and U9851 (N_9851,N_8339,N_8892);
xnor U9852 (N_9852,N_8974,N_8053);
nand U9853 (N_9853,N_8185,N_8894);
xnor U9854 (N_9854,N_8689,N_8163);
nor U9855 (N_9855,N_8970,N_8183);
nand U9856 (N_9856,N_8010,N_8181);
nor U9857 (N_9857,N_8810,N_8186);
xnor U9858 (N_9858,N_8779,N_8294);
nor U9859 (N_9859,N_8785,N_8110);
or U9860 (N_9860,N_8274,N_8860);
or U9861 (N_9861,N_8611,N_8231);
and U9862 (N_9862,N_8674,N_8533);
xnor U9863 (N_9863,N_8237,N_8596);
or U9864 (N_9864,N_8986,N_8728);
or U9865 (N_9865,N_8253,N_8017);
and U9866 (N_9866,N_8879,N_8102);
or U9867 (N_9867,N_8638,N_8765);
xnor U9868 (N_9868,N_8587,N_8944);
or U9869 (N_9869,N_8503,N_8981);
xor U9870 (N_9870,N_8304,N_8263);
nor U9871 (N_9871,N_8376,N_8149);
and U9872 (N_9872,N_8991,N_8717);
xor U9873 (N_9873,N_8639,N_8401);
xnor U9874 (N_9874,N_8073,N_8334);
nand U9875 (N_9875,N_8915,N_8889);
and U9876 (N_9876,N_8787,N_8741);
xor U9877 (N_9877,N_8405,N_8839);
xnor U9878 (N_9878,N_8505,N_8976);
nor U9879 (N_9879,N_8645,N_8462);
nor U9880 (N_9880,N_8070,N_8642);
xor U9881 (N_9881,N_8228,N_8409);
nand U9882 (N_9882,N_8132,N_8883);
nor U9883 (N_9883,N_8800,N_8766);
or U9884 (N_9884,N_8057,N_8503);
xnor U9885 (N_9885,N_8340,N_8413);
nand U9886 (N_9886,N_8684,N_8795);
nor U9887 (N_9887,N_8855,N_8296);
xor U9888 (N_9888,N_8056,N_8063);
nand U9889 (N_9889,N_8716,N_8468);
nor U9890 (N_9890,N_8628,N_8321);
nand U9891 (N_9891,N_8551,N_8277);
nand U9892 (N_9892,N_8385,N_8135);
nand U9893 (N_9893,N_8293,N_8000);
or U9894 (N_9894,N_8566,N_8349);
or U9895 (N_9895,N_8978,N_8787);
and U9896 (N_9896,N_8132,N_8984);
nand U9897 (N_9897,N_8801,N_8150);
or U9898 (N_9898,N_8614,N_8772);
nand U9899 (N_9899,N_8248,N_8815);
nor U9900 (N_9900,N_8486,N_8600);
nand U9901 (N_9901,N_8744,N_8669);
xor U9902 (N_9902,N_8665,N_8608);
nand U9903 (N_9903,N_8862,N_8829);
xnor U9904 (N_9904,N_8003,N_8088);
or U9905 (N_9905,N_8519,N_8745);
or U9906 (N_9906,N_8187,N_8698);
and U9907 (N_9907,N_8615,N_8235);
nor U9908 (N_9908,N_8866,N_8921);
nor U9909 (N_9909,N_8145,N_8240);
nor U9910 (N_9910,N_8792,N_8563);
and U9911 (N_9911,N_8541,N_8554);
xor U9912 (N_9912,N_8680,N_8552);
or U9913 (N_9913,N_8073,N_8994);
nor U9914 (N_9914,N_8209,N_8986);
nand U9915 (N_9915,N_8584,N_8156);
xor U9916 (N_9916,N_8636,N_8514);
xor U9917 (N_9917,N_8346,N_8793);
nor U9918 (N_9918,N_8851,N_8543);
or U9919 (N_9919,N_8834,N_8644);
nor U9920 (N_9920,N_8488,N_8360);
or U9921 (N_9921,N_8389,N_8076);
or U9922 (N_9922,N_8875,N_8134);
xnor U9923 (N_9923,N_8490,N_8418);
and U9924 (N_9924,N_8694,N_8874);
or U9925 (N_9925,N_8576,N_8768);
and U9926 (N_9926,N_8968,N_8009);
or U9927 (N_9927,N_8169,N_8427);
or U9928 (N_9928,N_8863,N_8759);
nor U9929 (N_9929,N_8318,N_8651);
nand U9930 (N_9930,N_8209,N_8166);
or U9931 (N_9931,N_8381,N_8914);
nand U9932 (N_9932,N_8993,N_8543);
or U9933 (N_9933,N_8055,N_8203);
nor U9934 (N_9934,N_8697,N_8484);
nor U9935 (N_9935,N_8610,N_8459);
nor U9936 (N_9936,N_8654,N_8838);
nor U9937 (N_9937,N_8448,N_8577);
nor U9938 (N_9938,N_8391,N_8494);
nand U9939 (N_9939,N_8470,N_8774);
or U9940 (N_9940,N_8072,N_8995);
nor U9941 (N_9941,N_8311,N_8799);
nand U9942 (N_9942,N_8940,N_8284);
xor U9943 (N_9943,N_8530,N_8807);
and U9944 (N_9944,N_8040,N_8651);
or U9945 (N_9945,N_8015,N_8380);
and U9946 (N_9946,N_8047,N_8416);
nand U9947 (N_9947,N_8585,N_8618);
or U9948 (N_9948,N_8663,N_8418);
nand U9949 (N_9949,N_8623,N_8408);
or U9950 (N_9950,N_8613,N_8881);
xnor U9951 (N_9951,N_8514,N_8718);
or U9952 (N_9952,N_8683,N_8763);
nor U9953 (N_9953,N_8386,N_8827);
nand U9954 (N_9954,N_8515,N_8836);
nand U9955 (N_9955,N_8614,N_8694);
nand U9956 (N_9956,N_8350,N_8683);
and U9957 (N_9957,N_8458,N_8621);
or U9958 (N_9958,N_8600,N_8534);
nand U9959 (N_9959,N_8246,N_8556);
nand U9960 (N_9960,N_8266,N_8318);
nand U9961 (N_9961,N_8075,N_8336);
xor U9962 (N_9962,N_8524,N_8423);
or U9963 (N_9963,N_8912,N_8766);
or U9964 (N_9964,N_8076,N_8262);
nand U9965 (N_9965,N_8734,N_8444);
and U9966 (N_9966,N_8626,N_8919);
nor U9967 (N_9967,N_8018,N_8920);
and U9968 (N_9968,N_8177,N_8517);
nor U9969 (N_9969,N_8567,N_8328);
xor U9970 (N_9970,N_8435,N_8920);
nor U9971 (N_9971,N_8712,N_8186);
nor U9972 (N_9972,N_8849,N_8757);
or U9973 (N_9973,N_8533,N_8870);
or U9974 (N_9974,N_8966,N_8411);
nand U9975 (N_9975,N_8049,N_8524);
or U9976 (N_9976,N_8452,N_8026);
or U9977 (N_9977,N_8205,N_8650);
xor U9978 (N_9978,N_8965,N_8998);
and U9979 (N_9979,N_8125,N_8188);
xor U9980 (N_9980,N_8021,N_8887);
nor U9981 (N_9981,N_8348,N_8219);
xnor U9982 (N_9982,N_8467,N_8832);
or U9983 (N_9983,N_8217,N_8736);
nor U9984 (N_9984,N_8251,N_8687);
nand U9985 (N_9985,N_8836,N_8758);
or U9986 (N_9986,N_8140,N_8242);
nand U9987 (N_9987,N_8959,N_8534);
xor U9988 (N_9988,N_8250,N_8559);
xnor U9989 (N_9989,N_8407,N_8163);
nor U9990 (N_9990,N_8149,N_8632);
and U9991 (N_9991,N_8331,N_8143);
nor U9992 (N_9992,N_8411,N_8549);
and U9993 (N_9993,N_8469,N_8790);
and U9994 (N_9994,N_8174,N_8548);
or U9995 (N_9995,N_8287,N_8658);
and U9996 (N_9996,N_8489,N_8990);
nor U9997 (N_9997,N_8551,N_8318);
or U9998 (N_9998,N_8727,N_8645);
nor U9999 (N_9999,N_8254,N_8459);
nor U10000 (N_10000,N_9415,N_9026);
or U10001 (N_10001,N_9045,N_9465);
xor U10002 (N_10002,N_9241,N_9311);
xnor U10003 (N_10003,N_9214,N_9204);
nand U10004 (N_10004,N_9927,N_9551);
xnor U10005 (N_10005,N_9746,N_9928);
and U10006 (N_10006,N_9352,N_9323);
or U10007 (N_10007,N_9284,N_9560);
and U10008 (N_10008,N_9998,N_9036);
nand U10009 (N_10009,N_9754,N_9582);
or U10010 (N_10010,N_9179,N_9675);
and U10011 (N_10011,N_9930,N_9547);
nand U10012 (N_10012,N_9780,N_9375);
and U10013 (N_10013,N_9864,N_9115);
and U10014 (N_10014,N_9424,N_9795);
nand U10015 (N_10015,N_9227,N_9123);
and U10016 (N_10016,N_9859,N_9866);
and U10017 (N_10017,N_9345,N_9999);
nand U10018 (N_10018,N_9244,N_9163);
nor U10019 (N_10019,N_9049,N_9128);
nor U10020 (N_10020,N_9381,N_9138);
or U10021 (N_10021,N_9225,N_9702);
or U10022 (N_10022,N_9785,N_9704);
or U10023 (N_10023,N_9275,N_9805);
and U10024 (N_10024,N_9318,N_9578);
nand U10025 (N_10025,N_9621,N_9386);
or U10026 (N_10026,N_9694,N_9738);
or U10027 (N_10027,N_9836,N_9543);
or U10028 (N_10028,N_9639,N_9978);
xor U10029 (N_10029,N_9863,N_9800);
nand U10030 (N_10030,N_9692,N_9130);
nor U10031 (N_10031,N_9609,N_9382);
nand U10032 (N_10032,N_9467,N_9791);
or U10033 (N_10033,N_9807,N_9555);
or U10034 (N_10034,N_9257,N_9568);
nand U10035 (N_10035,N_9913,N_9797);
nor U10036 (N_10036,N_9983,N_9308);
and U10037 (N_10037,N_9945,N_9495);
xor U10038 (N_10038,N_9222,N_9814);
nor U10039 (N_10039,N_9679,N_9852);
and U10040 (N_10040,N_9843,N_9297);
and U10041 (N_10041,N_9909,N_9712);
xnor U10042 (N_10042,N_9078,N_9066);
xnor U10043 (N_10043,N_9321,N_9708);
and U10044 (N_10044,N_9444,N_9765);
nand U10045 (N_10045,N_9152,N_9292);
or U10046 (N_10046,N_9695,N_9678);
nor U10047 (N_10047,N_9970,N_9208);
nand U10048 (N_10048,N_9146,N_9087);
nand U10049 (N_10049,N_9725,N_9183);
nor U10050 (N_10050,N_9471,N_9728);
xor U10051 (N_10051,N_9887,N_9472);
or U10052 (N_10052,N_9389,N_9619);
nand U10053 (N_10053,N_9486,N_9340);
nand U10054 (N_10054,N_9083,N_9588);
nand U10055 (N_10055,N_9833,N_9359);
nor U10056 (N_10056,N_9688,N_9480);
nand U10057 (N_10057,N_9149,N_9764);
nand U10058 (N_10058,N_9406,N_9975);
xnor U10059 (N_10059,N_9203,N_9553);
nor U10060 (N_10060,N_9080,N_9372);
and U10061 (N_10061,N_9145,N_9507);
and U10062 (N_10062,N_9557,N_9035);
nor U10063 (N_10063,N_9865,N_9682);
nor U10064 (N_10064,N_9758,N_9501);
xor U10065 (N_10065,N_9918,N_9230);
xor U10066 (N_10066,N_9696,N_9339);
nand U10067 (N_10067,N_9460,N_9937);
or U10068 (N_10068,N_9388,N_9879);
nor U10069 (N_10069,N_9242,N_9656);
nor U10070 (N_10070,N_9925,N_9816);
nor U10071 (N_10071,N_9464,N_9629);
xor U10072 (N_10072,N_9569,N_9358);
or U10073 (N_10073,N_9623,N_9686);
and U10074 (N_10074,N_9029,N_9786);
and U10075 (N_10075,N_9170,N_9662);
xnor U10076 (N_10076,N_9707,N_9243);
nand U10077 (N_10077,N_9914,N_9544);
and U10078 (N_10078,N_9693,N_9260);
and U10079 (N_10079,N_9373,N_9427);
nor U10080 (N_10080,N_9458,N_9735);
nor U10081 (N_10081,N_9683,N_9261);
or U10082 (N_10082,N_9660,N_9484);
and U10083 (N_10083,N_9285,N_9191);
xor U10084 (N_10084,N_9393,N_9881);
nand U10085 (N_10085,N_9594,N_9302);
nand U10086 (N_10086,N_9575,N_9108);
and U10087 (N_10087,N_9605,N_9857);
or U10088 (N_10088,N_9690,N_9652);
nand U10089 (N_10089,N_9342,N_9479);
xnor U10090 (N_10090,N_9911,N_9270);
or U10091 (N_10091,N_9948,N_9752);
nor U10092 (N_10092,N_9198,N_9330);
xnor U10093 (N_10093,N_9538,N_9614);
and U10094 (N_10094,N_9360,N_9399);
nand U10095 (N_10095,N_9092,N_9396);
nand U10096 (N_10096,N_9132,N_9337);
nor U10097 (N_10097,N_9748,N_9942);
xnor U10098 (N_10098,N_9473,N_9417);
xnor U10099 (N_10099,N_9369,N_9400);
xor U10100 (N_10100,N_9653,N_9071);
nor U10101 (N_10101,N_9246,N_9030);
or U10102 (N_10102,N_9210,N_9371);
or U10103 (N_10103,N_9142,N_9434);
nand U10104 (N_10104,N_9809,N_9721);
nor U10105 (N_10105,N_9824,N_9563);
or U10106 (N_10106,N_9002,N_9182);
nand U10107 (N_10107,N_9118,N_9591);
or U10108 (N_10108,N_9338,N_9109);
or U10109 (N_10109,N_9901,N_9808);
or U10110 (N_10110,N_9353,N_9401);
nand U10111 (N_10111,N_9364,N_9583);
xnor U10112 (N_10112,N_9150,N_9095);
or U10113 (N_10113,N_9587,N_9554);
nand U10114 (N_10114,N_9559,N_9121);
xor U10115 (N_10115,N_9305,N_9412);
nand U10116 (N_10116,N_9477,N_9005);
xnor U10117 (N_10117,N_9516,N_9521);
nand U10118 (N_10118,N_9449,N_9732);
nor U10119 (N_10119,N_9453,N_9586);
or U10120 (N_10120,N_9295,N_9119);
nand U10121 (N_10121,N_9362,N_9985);
nor U10122 (N_10122,N_9485,N_9468);
nor U10123 (N_10123,N_9710,N_9154);
xor U10124 (N_10124,N_9319,N_9439);
nor U10125 (N_10125,N_9976,N_9221);
and U10126 (N_10126,N_9011,N_9552);
nor U10127 (N_10127,N_9205,N_9713);
and U10128 (N_10128,N_9954,N_9753);
and U10129 (N_10129,N_9193,N_9917);
nor U10130 (N_10130,N_9476,N_9056);
xor U10131 (N_10131,N_9403,N_9497);
or U10132 (N_10132,N_9428,N_9231);
nor U10133 (N_10133,N_9343,N_9736);
nand U10134 (N_10134,N_9291,N_9992);
nand U10135 (N_10135,N_9046,N_9788);
nand U10136 (N_10136,N_9531,N_9589);
or U10137 (N_10137,N_9896,N_9514);
or U10138 (N_10138,N_9000,N_9420);
xnor U10139 (N_10139,N_9768,N_9063);
or U10140 (N_10140,N_9633,N_9838);
nor U10141 (N_10141,N_9706,N_9831);
or U10142 (N_10142,N_9176,N_9745);
nand U10143 (N_10143,N_9466,N_9039);
and U10144 (N_10144,N_9689,N_9931);
xnor U10145 (N_10145,N_9934,N_9296);
nand U10146 (N_10146,N_9781,N_9116);
nand U10147 (N_10147,N_9067,N_9845);
and U10148 (N_10148,N_9168,N_9703);
nand U10149 (N_10149,N_9581,N_9050);
and U10150 (N_10150,N_9580,N_9136);
nand U10151 (N_10151,N_9237,N_9654);
or U10152 (N_10152,N_9778,N_9437);
nand U10153 (N_10153,N_9885,N_9442);
and U10154 (N_10154,N_9891,N_9405);
nor U10155 (N_10155,N_9895,N_9025);
nor U10156 (N_10156,N_9890,N_9929);
xor U10157 (N_10157,N_9487,N_9958);
xnor U10158 (N_10158,N_9209,N_9390);
nor U10159 (N_10159,N_9215,N_9515);
and U10160 (N_10160,N_9829,N_9332);
xnor U10161 (N_10161,N_9625,N_9532);
and U10162 (N_10162,N_9720,N_9189);
nor U10163 (N_10163,N_9613,N_9883);
nand U10164 (N_10164,N_9262,N_9317);
or U10165 (N_10165,N_9562,N_9445);
xor U10166 (N_10166,N_9938,N_9727);
nand U10167 (N_10167,N_9378,N_9894);
xnor U10168 (N_10168,N_9597,N_9610);
or U10169 (N_10169,N_9456,N_9787);
nand U10170 (N_10170,N_9631,N_9033);
or U10171 (N_10171,N_9777,N_9773);
xnor U10172 (N_10172,N_9411,N_9987);
nor U10173 (N_10173,N_9546,N_9640);
nor U10174 (N_10174,N_9069,N_9509);
nor U10175 (N_10175,N_9286,N_9091);
and U10176 (N_10176,N_9782,N_9641);
and U10177 (N_10177,N_9573,N_9212);
or U10178 (N_10178,N_9677,N_9137);
or U10179 (N_10179,N_9463,N_9734);
nor U10180 (N_10180,N_9001,N_9759);
xnor U10181 (N_10181,N_9065,N_9665);
and U10182 (N_10182,N_9774,N_9113);
or U10183 (N_10183,N_9974,N_9761);
nor U10184 (N_10184,N_9923,N_9847);
nor U10185 (N_10185,N_9264,N_9120);
and U10186 (N_10186,N_9726,N_9618);
xnor U10187 (N_10187,N_9632,N_9977);
or U10188 (N_10188,N_9825,N_9756);
nand U10189 (N_10189,N_9004,N_9889);
and U10190 (N_10190,N_9878,N_9117);
or U10191 (N_10191,N_9664,N_9964);
nand U10192 (N_10192,N_9714,N_9835);
nor U10193 (N_10193,N_9862,N_9548);
and U10194 (N_10194,N_9848,N_9638);
nor U10195 (N_10195,N_9572,N_9074);
or U10196 (N_10196,N_9705,N_9041);
and U10197 (N_10197,N_9169,N_9790);
and U10198 (N_10198,N_9634,N_9806);
and U10199 (N_10199,N_9523,N_9920);
and U10200 (N_10200,N_9147,N_9624);
nor U10201 (N_10201,N_9351,N_9248);
xor U10202 (N_10202,N_9022,N_9269);
xor U10203 (N_10203,N_9666,N_9658);
xor U10204 (N_10204,N_9851,N_9320);
or U10205 (N_10205,N_9616,N_9349);
nand U10206 (N_10206,N_9828,N_9853);
nor U10207 (N_10207,N_9892,N_9329);
and U10208 (N_10208,N_9126,N_9973);
xnor U10209 (N_10209,N_9195,N_9111);
xor U10210 (N_10210,N_9886,N_9558);
xor U10211 (N_10211,N_9024,N_9031);
nand U10212 (N_10212,N_9144,N_9194);
nand U10213 (N_10213,N_9966,N_9072);
nor U10214 (N_10214,N_9837,N_9379);
and U10215 (N_10215,N_9511,N_9939);
nor U10216 (N_10216,N_9850,N_9990);
nand U10217 (N_10217,N_9316,N_9483);
xnor U10218 (N_10218,N_9447,N_9893);
xnor U10219 (N_10219,N_9398,N_9579);
or U10220 (N_10220,N_9593,N_9419);
and U10221 (N_10221,N_9162,N_9627);
xor U10222 (N_10222,N_9187,N_9451);
xnor U10223 (N_10223,N_9238,N_9946);
and U10224 (N_10224,N_9141,N_9151);
xnor U10225 (N_10225,N_9902,N_9088);
nand U10226 (N_10226,N_9252,N_9414);
xor U10227 (N_10227,N_9549,N_9874);
nor U10228 (N_10228,N_9410,N_9153);
nand U10229 (N_10229,N_9073,N_9968);
xor U10230 (N_10230,N_9164,N_9489);
nand U10231 (N_10231,N_9438,N_9576);
xor U10232 (N_10232,N_9226,N_9470);
nand U10233 (N_10233,N_9770,N_9749);
or U10234 (N_10234,N_9611,N_9245);
xnor U10235 (N_10235,N_9094,N_9719);
nor U10236 (N_10236,N_9047,N_9076);
nand U10237 (N_10237,N_9960,N_9102);
or U10238 (N_10238,N_9490,N_9924);
xor U10239 (N_10239,N_9802,N_9839);
and U10240 (N_10240,N_9595,N_9969);
nand U10241 (N_10241,N_9919,N_9013);
nor U10242 (N_10242,N_9823,N_9249);
or U10243 (N_10243,N_9229,N_9667);
or U10244 (N_10244,N_9334,N_9742);
nand U10245 (N_10245,N_9328,N_9899);
xnor U10246 (N_10246,N_9635,N_9256);
xnor U10247 (N_10247,N_9645,N_9266);
and U10248 (N_10248,N_9180,N_9017);
or U10249 (N_10249,N_9644,N_9200);
or U10250 (N_10250,N_9160,N_9043);
or U10251 (N_10251,N_9124,N_9100);
or U10252 (N_10252,N_9028,N_9457);
and U10253 (N_10253,N_9980,N_9023);
or U10254 (N_10254,N_9085,N_9723);
and U10255 (N_10255,N_9963,N_9197);
nand U10256 (N_10256,N_9448,N_9407);
nand U10257 (N_10257,N_9769,N_9875);
and U10258 (N_10258,N_9139,N_9984);
xor U10259 (N_10259,N_9818,N_9167);
nor U10260 (N_10260,N_9674,N_9522);
xor U10261 (N_10261,N_9199,N_9661);
nand U10262 (N_10262,N_9630,N_9175);
and U10263 (N_10263,N_9293,N_9042);
nand U10264 (N_10264,N_9263,N_9481);
or U10265 (N_10265,N_9775,N_9133);
xnor U10266 (N_10266,N_9691,N_9190);
nand U10267 (N_10267,N_9812,N_9826);
nand U10268 (N_10268,N_9500,N_9733);
and U10269 (N_10269,N_9015,N_9622);
xnor U10270 (N_10270,N_9397,N_9161);
and U10271 (N_10271,N_9717,N_9815);
xor U10272 (N_10272,N_9997,N_9021);
and U10273 (N_10273,N_9620,N_9053);
and U10274 (N_10274,N_9129,N_9165);
nand U10275 (N_10275,N_9055,N_9273);
nor U10276 (N_10276,N_9647,N_9416);
xor U10277 (N_10277,N_9671,N_9213);
xnor U10278 (N_10278,N_9408,N_9265);
and U10279 (N_10279,N_9711,N_9143);
or U10280 (N_10280,N_9333,N_9981);
and U10281 (N_10281,N_9520,N_9492);
nand U10282 (N_10282,N_9910,N_9421);
xor U10283 (N_10283,N_9650,N_9166);
nand U10284 (N_10284,N_9821,N_9861);
xnor U10285 (N_10285,N_9432,N_9697);
and U10286 (N_10286,N_9668,N_9374);
or U10287 (N_10287,N_9680,N_9234);
and U10288 (N_10288,N_9377,N_9801);
or U10289 (N_10289,N_9536,N_9429);
nand U10290 (N_10290,N_9051,N_9599);
nand U10291 (N_10291,N_9057,N_9496);
or U10292 (N_10292,N_9217,N_9016);
or U10293 (N_10293,N_9955,N_9798);
and U10294 (N_10294,N_9426,N_9341);
and U10295 (N_10295,N_9643,N_9218);
and U10296 (N_10296,N_9882,N_9052);
or U10297 (N_10297,N_9959,N_9084);
nand U10298 (N_10298,N_9898,N_9953);
nor U10299 (N_10299,N_9988,N_9127);
nand U10300 (N_10300,N_9093,N_9433);
xor U10301 (N_10301,N_9903,N_9277);
or U10302 (N_10302,N_9729,N_9574);
and U10303 (N_10303,N_9505,N_9391);
nand U10304 (N_10304,N_9503,N_9979);
and U10305 (N_10305,N_9657,N_9409);
and U10306 (N_10306,N_9228,N_9075);
xor U10307 (N_10307,N_9799,N_9796);
nor U10308 (N_10308,N_9870,N_9300);
and U10309 (N_10309,N_9598,N_9646);
xnor U10310 (N_10310,N_9289,N_9418);
nor U10311 (N_10311,N_9268,N_9254);
nor U10312 (N_10312,N_9010,N_9037);
nor U10313 (N_10313,N_9335,N_9854);
nor U10314 (N_10314,N_9112,N_9856);
nor U10315 (N_10315,N_9125,N_9766);
xnor U10316 (N_10316,N_9982,N_9685);
nor U10317 (N_10317,N_9475,N_9659);
and U10318 (N_10318,N_9855,N_9820);
nor U10319 (N_10319,N_9994,N_9701);
xor U10320 (N_10320,N_9159,N_9207);
and U10321 (N_10321,N_9422,N_9699);
nand U10322 (N_10322,N_9304,N_9584);
or U10323 (N_10323,N_9669,N_9873);
nor U10324 (N_10324,N_9846,N_9684);
and U10325 (N_10325,N_9098,N_9904);
and U10326 (N_10326,N_9506,N_9608);
nand U10327 (N_10327,N_9965,N_9663);
nand U10328 (N_10328,N_9648,N_9709);
and U10329 (N_10329,N_9577,N_9601);
xor U10330 (N_10330,N_9283,N_9602);
nand U10331 (N_10331,N_9932,N_9615);
nand U10332 (N_10332,N_9216,N_9687);
xnor U10333 (N_10333,N_9792,N_9344);
or U10334 (N_10334,N_9279,N_9545);
nand U10335 (N_10335,N_9716,N_9804);
or U10336 (N_10336,N_9600,N_9681);
nor U10337 (N_10337,N_9003,N_9941);
and U10338 (N_10338,N_9274,N_9211);
or U10339 (N_10339,N_9431,N_9040);
nand U10340 (N_10340,N_9086,N_9949);
nand U10341 (N_10341,N_9097,N_9255);
and U10342 (N_10342,N_9915,N_9202);
or U10343 (N_10343,N_9858,N_9649);
or U10344 (N_10344,N_9077,N_9655);
xnor U10345 (N_10345,N_9430,N_9566);
or U10346 (N_10346,N_9474,N_9044);
and U10347 (N_10347,N_9530,N_9366);
and U10348 (N_10348,N_9177,N_9989);
and U10349 (N_10349,N_9060,N_9535);
nor U10350 (N_10350,N_9008,N_9884);
and U10351 (N_10351,N_9384,N_9306);
or U10352 (N_10352,N_9561,N_9957);
or U10353 (N_10353,N_9944,N_9355);
xnor U10354 (N_10354,N_9834,N_9900);
and U10355 (N_10355,N_9240,N_9223);
nor U10356 (N_10356,N_9592,N_9567);
and U10357 (N_10357,N_9533,N_9383);
xor U10358 (N_10358,N_9184,N_9868);
and U10359 (N_10359,N_9423,N_9518);
or U10360 (N_10360,N_9539,N_9730);
or U10361 (N_10361,N_9178,N_9722);
nor U10362 (N_10362,N_9744,N_9007);
nor U10363 (N_10363,N_9313,N_9922);
and U10364 (N_10364,N_9724,N_9096);
and U10365 (N_10365,N_9596,N_9443);
nor U10366 (N_10366,N_9247,N_9803);
and U10367 (N_10367,N_9534,N_9081);
xnor U10368 (N_10368,N_9068,N_9606);
nand U10369 (N_10369,N_9519,N_9188);
and U10370 (N_10370,N_9871,N_9811);
and U10371 (N_10371,N_9140,N_9012);
nor U10372 (N_10372,N_9440,N_9493);
nor U10373 (N_10373,N_9972,N_9488);
or U10374 (N_10374,N_9921,N_9258);
nor U10375 (N_10375,N_9089,N_9276);
and U10376 (N_10376,N_9491,N_9737);
nand U10377 (N_10377,N_9986,N_9196);
or U10378 (N_10378,N_9750,N_9387);
and U10379 (N_10379,N_9540,N_9590);
xnor U10380 (N_10380,N_9392,N_9844);
xor U10381 (N_10381,N_9110,N_9731);
or U10382 (N_10382,N_9478,N_9783);
nor U10383 (N_10383,N_9906,N_9916);
or U10384 (N_10384,N_9537,N_9206);
nor U10385 (N_10385,N_9469,N_9905);
and U10386 (N_10386,N_9779,N_9626);
xor U10387 (N_10387,N_9935,N_9019);
nor U10388 (N_10388,N_9933,N_9236);
nand U10389 (N_10389,N_9018,N_9054);
xor U10390 (N_10390,N_9526,N_9006);
nor U10391 (N_10391,N_9527,N_9103);
or U10392 (N_10392,N_9793,N_9715);
or U10393 (N_10393,N_9079,N_9517);
nor U10394 (N_10394,N_9395,N_9743);
or U10395 (N_10395,N_9385,N_9950);
and U10396 (N_10396,N_9114,N_9104);
nand U10397 (N_10397,N_9105,N_9185);
xnor U10398 (N_10398,N_9082,N_9700);
nor U10399 (N_10399,N_9336,N_9740);
or U10400 (N_10400,N_9441,N_9762);
and U10401 (N_10401,N_9872,N_9672);
and U10402 (N_10402,N_9842,N_9832);
xor U10403 (N_10403,N_9134,N_9027);
nor U10404 (N_10404,N_9288,N_9099);
and U10405 (N_10405,N_9789,N_9529);
and U10406 (N_10406,N_9331,N_9718);
or U10407 (N_10407,N_9757,N_9239);
nor U10408 (N_10408,N_9637,N_9897);
nand U10409 (N_10409,N_9524,N_9947);
xor U10410 (N_10410,N_9278,N_9310);
nand U10411 (N_10411,N_9281,N_9346);
and U10412 (N_10412,N_9219,N_9322);
xor U10413 (N_10413,N_9867,N_9309);
xnor U10414 (N_10414,N_9991,N_9435);
xor U10415 (N_10415,N_9698,N_9090);
nor U10416 (N_10416,N_9951,N_9172);
or U10417 (N_10417,N_9971,N_9763);
nor U10418 (N_10418,N_9357,N_9462);
or U10419 (N_10419,N_9993,N_9908);
and U10420 (N_10420,N_9327,N_9394);
or U10421 (N_10421,N_9186,N_9347);
nand U10422 (N_10422,N_9402,N_9528);
xor U10423 (N_10423,N_9038,N_9325);
or U10424 (N_10424,N_9361,N_9926);
and U10425 (N_10425,N_9158,N_9482);
or U10426 (N_10426,N_9751,N_9995);
or U10427 (N_10427,N_9363,N_9784);
nand U10428 (N_10428,N_9513,N_9413);
nand U10429 (N_10429,N_9106,N_9171);
or U10430 (N_10430,N_9822,N_9155);
and U10431 (N_10431,N_9425,N_9565);
nand U10432 (N_10432,N_9967,N_9354);
or U10433 (N_10433,N_9810,N_9282);
xor U10434 (N_10434,N_9512,N_9272);
nand U10435 (N_10435,N_9510,N_9251);
xnor U10436 (N_10436,N_9772,N_9499);
xnor U10437 (N_10437,N_9450,N_9636);
nand U10438 (N_10438,N_9131,N_9612);
and U10439 (N_10439,N_9446,N_9303);
nor U10440 (N_10440,N_9461,N_9014);
and U10441 (N_10441,N_9174,N_9869);
nor U10442 (N_10442,N_9301,N_9148);
nor U10443 (N_10443,N_9454,N_9290);
nor U10444 (N_10444,N_9267,N_9048);
nand U10445 (N_10445,N_9376,N_9767);
nand U10446 (N_10446,N_9287,N_9604);
nand U10447 (N_10447,N_9324,N_9760);
nor U10448 (N_10448,N_9181,N_9771);
nor U10449 (N_10449,N_9307,N_9494);
or U10450 (N_10450,N_9541,N_9061);
or U10451 (N_10451,N_9550,N_9617);
xor U10452 (N_10452,N_9508,N_9062);
nor U10453 (N_10453,N_9314,N_9259);
or U10454 (N_10454,N_9880,N_9628);
xor U10455 (N_10455,N_9996,N_9157);
and U10456 (N_10456,N_9830,N_9525);
nor U10457 (N_10457,N_9940,N_9294);
nor U10458 (N_10458,N_9235,N_9135);
and U10459 (N_10459,N_9356,N_9436);
xor U10460 (N_10460,N_9452,N_9961);
or U10461 (N_10461,N_9813,N_9849);
nand U10462 (N_10462,N_9502,N_9956);
nor U10463 (N_10463,N_9299,N_9840);
xnor U10464 (N_10464,N_9876,N_9192);
nor U10465 (N_10465,N_9542,N_9271);
and U10466 (N_10466,N_9952,N_9009);
or U10467 (N_10467,N_9201,N_9173);
xnor U10468 (N_10468,N_9348,N_9250);
xor U10469 (N_10469,N_9747,N_9404);
nand U10470 (N_10470,N_9156,N_9670);
nor U10471 (N_10471,N_9817,N_9370);
or U10472 (N_10472,N_9350,N_9962);
nand U10473 (N_10473,N_9367,N_9315);
nand U10474 (N_10474,N_9571,N_9607);
or U10475 (N_10475,N_9365,N_9101);
nor U10476 (N_10476,N_9741,N_9564);
xor U10477 (N_10477,N_9827,N_9651);
nor U10478 (N_10478,N_9912,N_9253);
nand U10479 (N_10479,N_9943,N_9860);
or U10480 (N_10480,N_9070,N_9642);
or U10481 (N_10481,N_9794,N_9380);
nand U10482 (N_10482,N_9224,N_9059);
nor U10483 (N_10483,N_9064,N_9556);
xor U10484 (N_10484,N_9232,N_9034);
or U10485 (N_10485,N_9755,N_9673);
or U10486 (N_10486,N_9819,N_9326);
nor U10487 (N_10487,N_9907,N_9498);
or U10488 (N_10488,N_9676,N_9058);
and U10489 (N_10489,N_9032,N_9220);
or U10490 (N_10490,N_9877,N_9312);
and U10491 (N_10491,N_9888,N_9776);
nand U10492 (N_10492,N_9122,N_9280);
nor U10493 (N_10493,N_9603,N_9936);
nor U10494 (N_10494,N_9841,N_9739);
nor U10495 (N_10495,N_9298,N_9570);
nor U10496 (N_10496,N_9459,N_9368);
xor U10497 (N_10497,N_9233,N_9455);
nor U10498 (N_10498,N_9107,N_9585);
nor U10499 (N_10499,N_9504,N_9020);
or U10500 (N_10500,N_9526,N_9229);
and U10501 (N_10501,N_9255,N_9182);
and U10502 (N_10502,N_9317,N_9912);
nand U10503 (N_10503,N_9582,N_9595);
and U10504 (N_10504,N_9399,N_9588);
nor U10505 (N_10505,N_9798,N_9559);
and U10506 (N_10506,N_9119,N_9622);
nand U10507 (N_10507,N_9895,N_9226);
xor U10508 (N_10508,N_9699,N_9030);
or U10509 (N_10509,N_9711,N_9506);
nand U10510 (N_10510,N_9712,N_9312);
nand U10511 (N_10511,N_9131,N_9309);
and U10512 (N_10512,N_9904,N_9227);
or U10513 (N_10513,N_9357,N_9448);
nor U10514 (N_10514,N_9247,N_9737);
nand U10515 (N_10515,N_9412,N_9350);
xnor U10516 (N_10516,N_9167,N_9737);
and U10517 (N_10517,N_9283,N_9114);
nand U10518 (N_10518,N_9873,N_9049);
nand U10519 (N_10519,N_9989,N_9916);
xor U10520 (N_10520,N_9708,N_9325);
or U10521 (N_10521,N_9211,N_9956);
and U10522 (N_10522,N_9193,N_9332);
nand U10523 (N_10523,N_9163,N_9737);
and U10524 (N_10524,N_9301,N_9257);
nor U10525 (N_10525,N_9016,N_9179);
nand U10526 (N_10526,N_9091,N_9298);
or U10527 (N_10527,N_9549,N_9135);
nand U10528 (N_10528,N_9689,N_9042);
and U10529 (N_10529,N_9522,N_9930);
and U10530 (N_10530,N_9811,N_9737);
and U10531 (N_10531,N_9298,N_9670);
and U10532 (N_10532,N_9860,N_9225);
nor U10533 (N_10533,N_9959,N_9265);
and U10534 (N_10534,N_9391,N_9273);
nand U10535 (N_10535,N_9462,N_9340);
nor U10536 (N_10536,N_9196,N_9594);
or U10537 (N_10537,N_9970,N_9946);
or U10538 (N_10538,N_9877,N_9392);
xor U10539 (N_10539,N_9625,N_9035);
or U10540 (N_10540,N_9680,N_9045);
and U10541 (N_10541,N_9346,N_9111);
or U10542 (N_10542,N_9433,N_9189);
nor U10543 (N_10543,N_9735,N_9470);
xnor U10544 (N_10544,N_9717,N_9566);
nor U10545 (N_10545,N_9748,N_9014);
nand U10546 (N_10546,N_9024,N_9404);
or U10547 (N_10547,N_9505,N_9905);
nand U10548 (N_10548,N_9249,N_9216);
nand U10549 (N_10549,N_9125,N_9445);
nand U10550 (N_10550,N_9147,N_9126);
xnor U10551 (N_10551,N_9622,N_9139);
nand U10552 (N_10552,N_9956,N_9210);
and U10553 (N_10553,N_9868,N_9347);
nand U10554 (N_10554,N_9670,N_9116);
and U10555 (N_10555,N_9013,N_9019);
nand U10556 (N_10556,N_9406,N_9735);
nand U10557 (N_10557,N_9126,N_9941);
and U10558 (N_10558,N_9493,N_9903);
xnor U10559 (N_10559,N_9963,N_9327);
nand U10560 (N_10560,N_9043,N_9787);
xor U10561 (N_10561,N_9586,N_9594);
and U10562 (N_10562,N_9034,N_9706);
nor U10563 (N_10563,N_9304,N_9533);
or U10564 (N_10564,N_9112,N_9382);
xnor U10565 (N_10565,N_9690,N_9501);
nand U10566 (N_10566,N_9694,N_9740);
nand U10567 (N_10567,N_9514,N_9690);
nor U10568 (N_10568,N_9390,N_9938);
or U10569 (N_10569,N_9000,N_9073);
nand U10570 (N_10570,N_9031,N_9380);
or U10571 (N_10571,N_9289,N_9530);
and U10572 (N_10572,N_9484,N_9661);
nand U10573 (N_10573,N_9205,N_9655);
nand U10574 (N_10574,N_9274,N_9406);
nor U10575 (N_10575,N_9696,N_9624);
nor U10576 (N_10576,N_9273,N_9657);
xor U10577 (N_10577,N_9361,N_9872);
nand U10578 (N_10578,N_9069,N_9978);
nor U10579 (N_10579,N_9368,N_9413);
or U10580 (N_10580,N_9571,N_9919);
xnor U10581 (N_10581,N_9828,N_9226);
xnor U10582 (N_10582,N_9882,N_9378);
xor U10583 (N_10583,N_9623,N_9769);
xnor U10584 (N_10584,N_9622,N_9668);
nand U10585 (N_10585,N_9999,N_9957);
and U10586 (N_10586,N_9354,N_9344);
xor U10587 (N_10587,N_9806,N_9592);
nand U10588 (N_10588,N_9240,N_9608);
and U10589 (N_10589,N_9480,N_9391);
nor U10590 (N_10590,N_9742,N_9743);
nand U10591 (N_10591,N_9394,N_9796);
nand U10592 (N_10592,N_9569,N_9979);
nand U10593 (N_10593,N_9334,N_9024);
nor U10594 (N_10594,N_9950,N_9141);
and U10595 (N_10595,N_9118,N_9039);
and U10596 (N_10596,N_9190,N_9857);
nor U10597 (N_10597,N_9608,N_9904);
and U10598 (N_10598,N_9548,N_9303);
nand U10599 (N_10599,N_9054,N_9914);
nor U10600 (N_10600,N_9042,N_9113);
nand U10601 (N_10601,N_9169,N_9150);
and U10602 (N_10602,N_9092,N_9173);
and U10603 (N_10603,N_9664,N_9436);
or U10604 (N_10604,N_9117,N_9400);
xor U10605 (N_10605,N_9068,N_9945);
nand U10606 (N_10606,N_9418,N_9754);
nand U10607 (N_10607,N_9377,N_9943);
nand U10608 (N_10608,N_9947,N_9877);
nand U10609 (N_10609,N_9261,N_9543);
and U10610 (N_10610,N_9617,N_9149);
nor U10611 (N_10611,N_9101,N_9654);
nand U10612 (N_10612,N_9355,N_9291);
nand U10613 (N_10613,N_9224,N_9230);
or U10614 (N_10614,N_9350,N_9897);
nor U10615 (N_10615,N_9354,N_9840);
nor U10616 (N_10616,N_9707,N_9937);
or U10617 (N_10617,N_9593,N_9423);
nand U10618 (N_10618,N_9971,N_9800);
and U10619 (N_10619,N_9685,N_9862);
nor U10620 (N_10620,N_9494,N_9976);
xor U10621 (N_10621,N_9358,N_9388);
or U10622 (N_10622,N_9174,N_9316);
and U10623 (N_10623,N_9627,N_9346);
and U10624 (N_10624,N_9415,N_9268);
or U10625 (N_10625,N_9923,N_9139);
nor U10626 (N_10626,N_9923,N_9685);
or U10627 (N_10627,N_9479,N_9347);
xor U10628 (N_10628,N_9464,N_9463);
xor U10629 (N_10629,N_9327,N_9488);
nor U10630 (N_10630,N_9825,N_9607);
and U10631 (N_10631,N_9891,N_9952);
and U10632 (N_10632,N_9982,N_9860);
xnor U10633 (N_10633,N_9065,N_9581);
nand U10634 (N_10634,N_9087,N_9187);
nand U10635 (N_10635,N_9471,N_9501);
and U10636 (N_10636,N_9114,N_9910);
or U10637 (N_10637,N_9824,N_9513);
xor U10638 (N_10638,N_9611,N_9388);
nor U10639 (N_10639,N_9385,N_9367);
xor U10640 (N_10640,N_9871,N_9608);
and U10641 (N_10641,N_9316,N_9144);
or U10642 (N_10642,N_9444,N_9809);
and U10643 (N_10643,N_9911,N_9802);
or U10644 (N_10644,N_9829,N_9306);
nand U10645 (N_10645,N_9877,N_9584);
and U10646 (N_10646,N_9254,N_9765);
and U10647 (N_10647,N_9869,N_9365);
nor U10648 (N_10648,N_9007,N_9768);
nand U10649 (N_10649,N_9515,N_9296);
xor U10650 (N_10650,N_9778,N_9238);
nand U10651 (N_10651,N_9369,N_9302);
and U10652 (N_10652,N_9833,N_9918);
xnor U10653 (N_10653,N_9076,N_9083);
nor U10654 (N_10654,N_9104,N_9791);
xor U10655 (N_10655,N_9987,N_9273);
xor U10656 (N_10656,N_9599,N_9061);
or U10657 (N_10657,N_9901,N_9449);
or U10658 (N_10658,N_9467,N_9559);
xnor U10659 (N_10659,N_9565,N_9078);
or U10660 (N_10660,N_9627,N_9182);
or U10661 (N_10661,N_9782,N_9562);
or U10662 (N_10662,N_9119,N_9704);
nor U10663 (N_10663,N_9620,N_9918);
xnor U10664 (N_10664,N_9764,N_9681);
nor U10665 (N_10665,N_9968,N_9003);
xor U10666 (N_10666,N_9933,N_9006);
or U10667 (N_10667,N_9480,N_9628);
and U10668 (N_10668,N_9361,N_9934);
nor U10669 (N_10669,N_9435,N_9641);
nor U10670 (N_10670,N_9245,N_9174);
and U10671 (N_10671,N_9972,N_9647);
and U10672 (N_10672,N_9148,N_9143);
and U10673 (N_10673,N_9323,N_9784);
nand U10674 (N_10674,N_9271,N_9961);
and U10675 (N_10675,N_9412,N_9000);
nor U10676 (N_10676,N_9149,N_9294);
or U10677 (N_10677,N_9594,N_9961);
xor U10678 (N_10678,N_9338,N_9143);
or U10679 (N_10679,N_9725,N_9513);
or U10680 (N_10680,N_9160,N_9652);
or U10681 (N_10681,N_9152,N_9739);
and U10682 (N_10682,N_9975,N_9609);
xor U10683 (N_10683,N_9383,N_9090);
or U10684 (N_10684,N_9436,N_9944);
or U10685 (N_10685,N_9620,N_9080);
or U10686 (N_10686,N_9246,N_9943);
nor U10687 (N_10687,N_9283,N_9585);
nor U10688 (N_10688,N_9889,N_9952);
and U10689 (N_10689,N_9886,N_9094);
or U10690 (N_10690,N_9466,N_9181);
and U10691 (N_10691,N_9653,N_9443);
xor U10692 (N_10692,N_9670,N_9739);
xor U10693 (N_10693,N_9760,N_9277);
xor U10694 (N_10694,N_9124,N_9905);
nand U10695 (N_10695,N_9702,N_9943);
nand U10696 (N_10696,N_9839,N_9375);
or U10697 (N_10697,N_9972,N_9759);
xor U10698 (N_10698,N_9036,N_9594);
nand U10699 (N_10699,N_9346,N_9272);
nor U10700 (N_10700,N_9837,N_9558);
or U10701 (N_10701,N_9484,N_9643);
xor U10702 (N_10702,N_9093,N_9577);
nand U10703 (N_10703,N_9199,N_9445);
xnor U10704 (N_10704,N_9456,N_9179);
xor U10705 (N_10705,N_9340,N_9042);
and U10706 (N_10706,N_9427,N_9597);
or U10707 (N_10707,N_9932,N_9705);
and U10708 (N_10708,N_9969,N_9000);
or U10709 (N_10709,N_9579,N_9254);
nand U10710 (N_10710,N_9314,N_9380);
and U10711 (N_10711,N_9827,N_9979);
xnor U10712 (N_10712,N_9650,N_9091);
xor U10713 (N_10713,N_9949,N_9396);
or U10714 (N_10714,N_9547,N_9013);
nor U10715 (N_10715,N_9893,N_9409);
nor U10716 (N_10716,N_9858,N_9358);
or U10717 (N_10717,N_9426,N_9540);
xnor U10718 (N_10718,N_9637,N_9941);
nor U10719 (N_10719,N_9115,N_9186);
or U10720 (N_10720,N_9441,N_9993);
or U10721 (N_10721,N_9739,N_9740);
and U10722 (N_10722,N_9691,N_9656);
nand U10723 (N_10723,N_9525,N_9271);
or U10724 (N_10724,N_9438,N_9513);
nand U10725 (N_10725,N_9737,N_9646);
xor U10726 (N_10726,N_9627,N_9484);
xor U10727 (N_10727,N_9429,N_9882);
nor U10728 (N_10728,N_9756,N_9266);
nand U10729 (N_10729,N_9524,N_9570);
and U10730 (N_10730,N_9324,N_9637);
or U10731 (N_10731,N_9134,N_9800);
nand U10732 (N_10732,N_9518,N_9729);
nor U10733 (N_10733,N_9032,N_9700);
or U10734 (N_10734,N_9377,N_9952);
or U10735 (N_10735,N_9963,N_9549);
xnor U10736 (N_10736,N_9712,N_9526);
or U10737 (N_10737,N_9836,N_9225);
nand U10738 (N_10738,N_9964,N_9234);
and U10739 (N_10739,N_9766,N_9045);
or U10740 (N_10740,N_9636,N_9600);
and U10741 (N_10741,N_9328,N_9272);
or U10742 (N_10742,N_9935,N_9379);
xnor U10743 (N_10743,N_9035,N_9229);
or U10744 (N_10744,N_9381,N_9353);
nand U10745 (N_10745,N_9214,N_9824);
and U10746 (N_10746,N_9581,N_9446);
xor U10747 (N_10747,N_9479,N_9858);
and U10748 (N_10748,N_9035,N_9111);
xor U10749 (N_10749,N_9410,N_9875);
or U10750 (N_10750,N_9500,N_9171);
nand U10751 (N_10751,N_9434,N_9016);
xnor U10752 (N_10752,N_9235,N_9499);
and U10753 (N_10753,N_9819,N_9396);
nor U10754 (N_10754,N_9788,N_9985);
nand U10755 (N_10755,N_9963,N_9477);
or U10756 (N_10756,N_9346,N_9443);
or U10757 (N_10757,N_9023,N_9128);
nor U10758 (N_10758,N_9839,N_9317);
nand U10759 (N_10759,N_9750,N_9214);
nor U10760 (N_10760,N_9084,N_9367);
nor U10761 (N_10761,N_9542,N_9622);
and U10762 (N_10762,N_9769,N_9562);
nand U10763 (N_10763,N_9747,N_9832);
and U10764 (N_10764,N_9718,N_9768);
nand U10765 (N_10765,N_9068,N_9693);
nand U10766 (N_10766,N_9248,N_9204);
nand U10767 (N_10767,N_9174,N_9153);
and U10768 (N_10768,N_9655,N_9446);
and U10769 (N_10769,N_9536,N_9983);
nor U10770 (N_10770,N_9453,N_9237);
or U10771 (N_10771,N_9831,N_9236);
and U10772 (N_10772,N_9688,N_9105);
nand U10773 (N_10773,N_9329,N_9894);
or U10774 (N_10774,N_9280,N_9638);
and U10775 (N_10775,N_9035,N_9859);
nor U10776 (N_10776,N_9071,N_9244);
nor U10777 (N_10777,N_9519,N_9090);
xnor U10778 (N_10778,N_9806,N_9699);
nand U10779 (N_10779,N_9900,N_9973);
nand U10780 (N_10780,N_9146,N_9566);
or U10781 (N_10781,N_9733,N_9838);
and U10782 (N_10782,N_9657,N_9607);
xor U10783 (N_10783,N_9591,N_9692);
and U10784 (N_10784,N_9316,N_9988);
xor U10785 (N_10785,N_9169,N_9468);
nand U10786 (N_10786,N_9824,N_9674);
nor U10787 (N_10787,N_9198,N_9238);
or U10788 (N_10788,N_9895,N_9229);
xor U10789 (N_10789,N_9469,N_9045);
nand U10790 (N_10790,N_9908,N_9371);
or U10791 (N_10791,N_9089,N_9334);
nor U10792 (N_10792,N_9169,N_9728);
xnor U10793 (N_10793,N_9073,N_9251);
and U10794 (N_10794,N_9531,N_9486);
xnor U10795 (N_10795,N_9017,N_9585);
and U10796 (N_10796,N_9677,N_9540);
or U10797 (N_10797,N_9580,N_9093);
nand U10798 (N_10798,N_9009,N_9770);
nor U10799 (N_10799,N_9412,N_9858);
nor U10800 (N_10800,N_9749,N_9122);
nor U10801 (N_10801,N_9249,N_9778);
xnor U10802 (N_10802,N_9242,N_9725);
xnor U10803 (N_10803,N_9149,N_9028);
and U10804 (N_10804,N_9370,N_9077);
nand U10805 (N_10805,N_9703,N_9655);
or U10806 (N_10806,N_9891,N_9308);
xor U10807 (N_10807,N_9366,N_9464);
or U10808 (N_10808,N_9296,N_9353);
xor U10809 (N_10809,N_9308,N_9464);
nor U10810 (N_10810,N_9619,N_9834);
or U10811 (N_10811,N_9282,N_9362);
and U10812 (N_10812,N_9859,N_9007);
or U10813 (N_10813,N_9291,N_9272);
nor U10814 (N_10814,N_9264,N_9437);
nor U10815 (N_10815,N_9967,N_9618);
and U10816 (N_10816,N_9220,N_9632);
or U10817 (N_10817,N_9742,N_9376);
and U10818 (N_10818,N_9397,N_9349);
nor U10819 (N_10819,N_9513,N_9206);
xor U10820 (N_10820,N_9415,N_9759);
or U10821 (N_10821,N_9673,N_9613);
and U10822 (N_10822,N_9955,N_9920);
nand U10823 (N_10823,N_9416,N_9559);
or U10824 (N_10824,N_9629,N_9354);
or U10825 (N_10825,N_9974,N_9890);
xnor U10826 (N_10826,N_9025,N_9172);
xnor U10827 (N_10827,N_9136,N_9946);
xor U10828 (N_10828,N_9112,N_9805);
and U10829 (N_10829,N_9844,N_9753);
nand U10830 (N_10830,N_9060,N_9943);
or U10831 (N_10831,N_9817,N_9130);
or U10832 (N_10832,N_9652,N_9618);
nor U10833 (N_10833,N_9350,N_9549);
nand U10834 (N_10834,N_9164,N_9317);
nor U10835 (N_10835,N_9388,N_9998);
nor U10836 (N_10836,N_9144,N_9318);
or U10837 (N_10837,N_9910,N_9832);
xor U10838 (N_10838,N_9831,N_9657);
nor U10839 (N_10839,N_9544,N_9354);
nand U10840 (N_10840,N_9286,N_9114);
nand U10841 (N_10841,N_9284,N_9147);
or U10842 (N_10842,N_9886,N_9060);
and U10843 (N_10843,N_9218,N_9327);
nor U10844 (N_10844,N_9014,N_9255);
or U10845 (N_10845,N_9389,N_9054);
nor U10846 (N_10846,N_9163,N_9384);
or U10847 (N_10847,N_9120,N_9560);
nand U10848 (N_10848,N_9494,N_9280);
nor U10849 (N_10849,N_9555,N_9502);
nor U10850 (N_10850,N_9350,N_9093);
nor U10851 (N_10851,N_9891,N_9151);
xor U10852 (N_10852,N_9932,N_9147);
nand U10853 (N_10853,N_9259,N_9558);
xnor U10854 (N_10854,N_9050,N_9693);
nor U10855 (N_10855,N_9395,N_9768);
and U10856 (N_10856,N_9461,N_9371);
nor U10857 (N_10857,N_9127,N_9564);
and U10858 (N_10858,N_9375,N_9209);
nor U10859 (N_10859,N_9900,N_9299);
nor U10860 (N_10860,N_9015,N_9749);
nand U10861 (N_10861,N_9182,N_9522);
nor U10862 (N_10862,N_9457,N_9958);
and U10863 (N_10863,N_9734,N_9488);
xnor U10864 (N_10864,N_9893,N_9397);
or U10865 (N_10865,N_9323,N_9891);
xor U10866 (N_10866,N_9663,N_9439);
or U10867 (N_10867,N_9601,N_9033);
or U10868 (N_10868,N_9808,N_9159);
xor U10869 (N_10869,N_9126,N_9981);
nand U10870 (N_10870,N_9869,N_9231);
nor U10871 (N_10871,N_9671,N_9633);
or U10872 (N_10872,N_9623,N_9377);
xor U10873 (N_10873,N_9284,N_9723);
nand U10874 (N_10874,N_9702,N_9133);
nor U10875 (N_10875,N_9291,N_9514);
and U10876 (N_10876,N_9739,N_9242);
or U10877 (N_10877,N_9038,N_9136);
xor U10878 (N_10878,N_9453,N_9960);
nor U10879 (N_10879,N_9647,N_9575);
nor U10880 (N_10880,N_9300,N_9213);
and U10881 (N_10881,N_9248,N_9274);
or U10882 (N_10882,N_9464,N_9138);
and U10883 (N_10883,N_9549,N_9757);
and U10884 (N_10884,N_9605,N_9973);
xnor U10885 (N_10885,N_9068,N_9801);
or U10886 (N_10886,N_9354,N_9057);
or U10887 (N_10887,N_9929,N_9354);
and U10888 (N_10888,N_9438,N_9313);
nand U10889 (N_10889,N_9686,N_9524);
or U10890 (N_10890,N_9043,N_9898);
and U10891 (N_10891,N_9036,N_9681);
nand U10892 (N_10892,N_9275,N_9910);
nand U10893 (N_10893,N_9406,N_9106);
nand U10894 (N_10894,N_9063,N_9980);
nor U10895 (N_10895,N_9989,N_9134);
or U10896 (N_10896,N_9132,N_9322);
nor U10897 (N_10897,N_9386,N_9326);
nand U10898 (N_10898,N_9482,N_9111);
nand U10899 (N_10899,N_9796,N_9719);
xnor U10900 (N_10900,N_9508,N_9142);
and U10901 (N_10901,N_9368,N_9367);
or U10902 (N_10902,N_9959,N_9810);
nand U10903 (N_10903,N_9480,N_9828);
or U10904 (N_10904,N_9305,N_9107);
xor U10905 (N_10905,N_9735,N_9308);
nor U10906 (N_10906,N_9645,N_9872);
or U10907 (N_10907,N_9856,N_9129);
xnor U10908 (N_10908,N_9534,N_9849);
and U10909 (N_10909,N_9207,N_9000);
and U10910 (N_10910,N_9231,N_9366);
xnor U10911 (N_10911,N_9383,N_9106);
and U10912 (N_10912,N_9766,N_9755);
and U10913 (N_10913,N_9870,N_9798);
nor U10914 (N_10914,N_9631,N_9981);
nor U10915 (N_10915,N_9133,N_9780);
nor U10916 (N_10916,N_9688,N_9596);
xor U10917 (N_10917,N_9438,N_9377);
or U10918 (N_10918,N_9132,N_9900);
or U10919 (N_10919,N_9453,N_9519);
nand U10920 (N_10920,N_9731,N_9811);
or U10921 (N_10921,N_9352,N_9134);
nor U10922 (N_10922,N_9032,N_9355);
nand U10923 (N_10923,N_9321,N_9873);
xnor U10924 (N_10924,N_9466,N_9689);
nand U10925 (N_10925,N_9176,N_9598);
or U10926 (N_10926,N_9393,N_9940);
nand U10927 (N_10927,N_9819,N_9478);
nand U10928 (N_10928,N_9264,N_9299);
and U10929 (N_10929,N_9309,N_9333);
nand U10930 (N_10930,N_9538,N_9001);
or U10931 (N_10931,N_9110,N_9298);
or U10932 (N_10932,N_9268,N_9286);
nand U10933 (N_10933,N_9002,N_9109);
and U10934 (N_10934,N_9000,N_9885);
nor U10935 (N_10935,N_9241,N_9295);
and U10936 (N_10936,N_9756,N_9411);
and U10937 (N_10937,N_9606,N_9795);
nor U10938 (N_10938,N_9514,N_9946);
and U10939 (N_10939,N_9497,N_9688);
or U10940 (N_10940,N_9916,N_9249);
or U10941 (N_10941,N_9870,N_9632);
and U10942 (N_10942,N_9009,N_9804);
or U10943 (N_10943,N_9608,N_9759);
and U10944 (N_10944,N_9781,N_9099);
xnor U10945 (N_10945,N_9244,N_9867);
nor U10946 (N_10946,N_9677,N_9824);
xnor U10947 (N_10947,N_9842,N_9037);
nor U10948 (N_10948,N_9022,N_9700);
and U10949 (N_10949,N_9334,N_9540);
or U10950 (N_10950,N_9891,N_9628);
nand U10951 (N_10951,N_9266,N_9441);
nor U10952 (N_10952,N_9755,N_9887);
nand U10953 (N_10953,N_9162,N_9513);
xor U10954 (N_10954,N_9824,N_9719);
nand U10955 (N_10955,N_9201,N_9387);
nor U10956 (N_10956,N_9021,N_9100);
xnor U10957 (N_10957,N_9511,N_9737);
xor U10958 (N_10958,N_9392,N_9724);
nor U10959 (N_10959,N_9135,N_9913);
xor U10960 (N_10960,N_9548,N_9503);
nand U10961 (N_10961,N_9370,N_9010);
xor U10962 (N_10962,N_9150,N_9766);
and U10963 (N_10963,N_9953,N_9210);
nor U10964 (N_10964,N_9441,N_9934);
nor U10965 (N_10965,N_9706,N_9891);
nand U10966 (N_10966,N_9559,N_9655);
or U10967 (N_10967,N_9704,N_9280);
nand U10968 (N_10968,N_9070,N_9875);
nand U10969 (N_10969,N_9614,N_9309);
or U10970 (N_10970,N_9377,N_9794);
nor U10971 (N_10971,N_9007,N_9910);
and U10972 (N_10972,N_9251,N_9339);
and U10973 (N_10973,N_9106,N_9860);
nand U10974 (N_10974,N_9495,N_9915);
nor U10975 (N_10975,N_9022,N_9751);
nor U10976 (N_10976,N_9139,N_9280);
nor U10977 (N_10977,N_9711,N_9827);
or U10978 (N_10978,N_9359,N_9240);
nand U10979 (N_10979,N_9461,N_9293);
and U10980 (N_10980,N_9396,N_9109);
and U10981 (N_10981,N_9917,N_9716);
or U10982 (N_10982,N_9288,N_9490);
nor U10983 (N_10983,N_9659,N_9355);
xor U10984 (N_10984,N_9355,N_9881);
and U10985 (N_10985,N_9257,N_9395);
xnor U10986 (N_10986,N_9367,N_9853);
or U10987 (N_10987,N_9625,N_9475);
nor U10988 (N_10988,N_9078,N_9316);
and U10989 (N_10989,N_9021,N_9300);
or U10990 (N_10990,N_9633,N_9854);
xnor U10991 (N_10991,N_9248,N_9653);
or U10992 (N_10992,N_9458,N_9371);
nand U10993 (N_10993,N_9475,N_9177);
nor U10994 (N_10994,N_9907,N_9707);
xnor U10995 (N_10995,N_9552,N_9216);
and U10996 (N_10996,N_9623,N_9596);
nand U10997 (N_10997,N_9739,N_9752);
nand U10998 (N_10998,N_9327,N_9586);
and U10999 (N_10999,N_9601,N_9055);
nand U11000 (N_11000,N_10840,N_10711);
or U11001 (N_11001,N_10142,N_10956);
nand U11002 (N_11002,N_10568,N_10601);
and U11003 (N_11003,N_10229,N_10726);
xnor U11004 (N_11004,N_10903,N_10429);
or U11005 (N_11005,N_10853,N_10282);
nor U11006 (N_11006,N_10397,N_10108);
xor U11007 (N_11007,N_10343,N_10374);
nand U11008 (N_11008,N_10713,N_10953);
or U11009 (N_11009,N_10471,N_10611);
or U11010 (N_11010,N_10731,N_10881);
or U11011 (N_11011,N_10905,N_10749);
and U11012 (N_11012,N_10136,N_10984);
or U11013 (N_11013,N_10486,N_10402);
or U11014 (N_11014,N_10944,N_10216);
xor U11015 (N_11015,N_10697,N_10365);
nand U11016 (N_11016,N_10173,N_10442);
and U11017 (N_11017,N_10570,N_10519);
or U11018 (N_11018,N_10597,N_10513);
nor U11019 (N_11019,N_10144,N_10764);
nor U11020 (N_11020,N_10464,N_10633);
and U11021 (N_11021,N_10854,N_10192);
nand U11022 (N_11022,N_10813,N_10991);
and U11023 (N_11023,N_10129,N_10950);
or U11024 (N_11024,N_10819,N_10494);
nand U11025 (N_11025,N_10544,N_10244);
nor U11026 (N_11026,N_10561,N_10013);
and U11027 (N_11027,N_10790,N_10123);
or U11028 (N_11028,N_10795,N_10566);
and U11029 (N_11029,N_10565,N_10349);
xnor U11030 (N_11030,N_10933,N_10985);
and U11031 (N_11031,N_10255,N_10051);
or U11032 (N_11032,N_10098,N_10980);
or U11033 (N_11033,N_10341,N_10109);
nand U11034 (N_11034,N_10317,N_10434);
nand U11035 (N_11035,N_10882,N_10850);
and U11036 (N_11036,N_10484,N_10163);
and U11037 (N_11037,N_10578,N_10902);
and U11038 (N_11038,N_10678,N_10584);
and U11039 (N_11039,N_10065,N_10973);
nor U11040 (N_11040,N_10497,N_10211);
nor U11041 (N_11041,N_10396,N_10480);
and U11042 (N_11042,N_10030,N_10663);
and U11043 (N_11043,N_10910,N_10859);
xor U11044 (N_11044,N_10828,N_10280);
or U11045 (N_11045,N_10212,N_10080);
nor U11046 (N_11046,N_10485,N_10914);
and U11047 (N_11047,N_10862,N_10846);
nand U11048 (N_11048,N_10745,N_10313);
or U11049 (N_11049,N_10206,N_10072);
and U11050 (N_11050,N_10208,N_10572);
or U11051 (N_11051,N_10182,N_10391);
nand U11052 (N_11052,N_10703,N_10405);
nor U11053 (N_11053,N_10028,N_10390);
nor U11054 (N_11054,N_10997,N_10553);
nand U11055 (N_11055,N_10929,N_10281);
xor U11056 (N_11056,N_10094,N_10372);
or U11057 (N_11057,N_10151,N_10474);
nor U11058 (N_11058,N_10976,N_10571);
and U11059 (N_11059,N_10930,N_10367);
xor U11060 (N_11060,N_10079,N_10863);
nand U11061 (N_11061,N_10945,N_10665);
nor U11062 (N_11062,N_10575,N_10753);
and U11063 (N_11063,N_10202,N_10406);
nand U11064 (N_11064,N_10761,N_10931);
nor U11065 (N_11065,N_10201,N_10783);
nand U11066 (N_11066,N_10059,N_10185);
xnor U11067 (N_11067,N_10638,N_10856);
or U11068 (N_11068,N_10619,N_10320);
and U11069 (N_11069,N_10132,N_10298);
nand U11070 (N_11070,N_10603,N_10730);
and U11071 (N_11071,N_10803,N_10545);
or U11072 (N_11072,N_10149,N_10009);
or U11073 (N_11073,N_10082,N_10137);
nand U11074 (N_11074,N_10838,N_10453);
or U11075 (N_11075,N_10467,N_10912);
xor U11076 (N_11076,N_10135,N_10509);
nand U11077 (N_11077,N_10071,N_10878);
nand U11078 (N_11078,N_10772,N_10528);
nor U11079 (N_11079,N_10841,N_10807);
xnor U11080 (N_11080,N_10554,N_10284);
or U11081 (N_11081,N_10380,N_10252);
nand U11082 (N_11082,N_10555,N_10928);
or U11083 (N_11083,N_10225,N_10200);
xnor U11084 (N_11084,N_10830,N_10010);
nor U11085 (N_11085,N_10037,N_10334);
nand U11086 (N_11086,N_10412,N_10337);
nor U11087 (N_11087,N_10630,N_10256);
xnor U11088 (N_11088,N_10270,N_10112);
and U11089 (N_11089,N_10117,N_10737);
xor U11090 (N_11090,N_10787,N_10768);
or U11091 (N_11091,N_10250,N_10696);
and U11092 (N_11092,N_10971,N_10034);
nor U11093 (N_11093,N_10851,N_10982);
nand U11094 (N_11094,N_10981,N_10829);
nand U11095 (N_11095,N_10750,N_10328);
xnor U11096 (N_11096,N_10056,N_10567);
or U11097 (N_11097,N_10877,N_10809);
and U11098 (N_11098,N_10530,N_10475);
and U11099 (N_11099,N_10789,N_10101);
and U11100 (N_11100,N_10860,N_10331);
and U11101 (N_11101,N_10427,N_10277);
nor U11102 (N_11102,N_10029,N_10265);
and U11103 (N_11103,N_10375,N_10677);
nor U11104 (N_11104,N_10360,N_10869);
and U11105 (N_11105,N_10573,N_10539);
nor U11106 (N_11106,N_10383,N_10230);
xor U11107 (N_11107,N_10004,N_10574);
and U11108 (N_11108,N_10063,N_10636);
xnor U11109 (N_11109,N_10249,N_10125);
and U11110 (N_11110,N_10319,N_10156);
and U11111 (N_11111,N_10818,N_10607);
or U11112 (N_11112,N_10322,N_10826);
and U11113 (N_11113,N_10552,N_10569);
and U11114 (N_11114,N_10248,N_10140);
xnor U11115 (N_11115,N_10801,N_10055);
xor U11116 (N_11116,N_10704,N_10295);
nor U11117 (N_11117,N_10189,N_10222);
xnor U11118 (N_11118,N_10089,N_10077);
nor U11119 (N_11119,N_10147,N_10235);
and U11120 (N_11120,N_10096,N_10060);
or U11121 (N_11121,N_10264,N_10806);
nand U11122 (N_11122,N_10747,N_10844);
or U11123 (N_11123,N_10420,N_10490);
or U11124 (N_11124,N_10836,N_10642);
xnor U11125 (N_11125,N_10213,N_10348);
nor U11126 (N_11126,N_10674,N_10487);
and U11127 (N_11127,N_10363,N_10968);
nand U11128 (N_11128,N_10289,N_10918);
nor U11129 (N_11129,N_10947,N_10445);
nor U11130 (N_11130,N_10033,N_10018);
nand U11131 (N_11131,N_10935,N_10825);
xnor U11132 (N_11132,N_10027,N_10651);
and U11133 (N_11133,N_10304,N_10162);
or U11134 (N_11134,N_10241,N_10259);
and U11135 (N_11135,N_10771,N_10128);
and U11136 (N_11136,N_10989,N_10158);
or U11137 (N_11137,N_10915,N_10439);
or U11138 (N_11138,N_10253,N_10754);
xnor U11139 (N_11139,N_10515,N_10612);
xor U11140 (N_11140,N_10352,N_10632);
xor U11141 (N_11141,N_10791,N_10917);
xnor U11142 (N_11142,N_10261,N_10164);
nor U11143 (N_11143,N_10451,N_10624);
xor U11144 (N_11144,N_10269,N_10350);
xnor U11145 (N_11145,N_10675,N_10450);
nand U11146 (N_11146,N_10623,N_10873);
or U11147 (N_11147,N_10078,N_10880);
nor U11148 (N_11148,N_10816,N_10001);
and U11149 (N_11149,N_10934,N_10291);
or U11150 (N_11150,N_10410,N_10488);
nor U11151 (N_11151,N_10088,N_10026);
nor U11152 (N_11152,N_10035,N_10534);
xor U11153 (N_11153,N_10314,N_10837);
and U11154 (N_11154,N_10141,N_10047);
xor U11155 (N_11155,N_10338,N_10738);
nand U11156 (N_11156,N_10344,N_10522);
xnor U11157 (N_11157,N_10583,N_10591);
nor U11158 (N_11158,N_10900,N_10994);
nor U11159 (N_11159,N_10462,N_10921);
and U11160 (N_11160,N_10146,N_10833);
or U11161 (N_11161,N_10786,N_10458);
nand U11162 (N_11162,N_10822,N_10045);
or U11163 (N_11163,N_10942,N_10274);
xor U11164 (N_11164,N_10385,N_10735);
xor U11165 (N_11165,N_10395,N_10233);
and U11166 (N_11166,N_10303,N_10710);
or U11167 (N_11167,N_10774,N_10231);
or U11168 (N_11168,N_10058,N_10776);
and U11169 (N_11169,N_10657,N_10872);
nor U11170 (N_11170,N_10742,N_10118);
nor U11171 (N_11171,N_10955,N_10207);
xor U11172 (N_11172,N_10381,N_10316);
nor U11173 (N_11173,N_10884,N_10170);
xnor U11174 (N_11174,N_10242,N_10852);
nor U11175 (N_11175,N_10700,N_10422);
nor U11176 (N_11176,N_10014,N_10021);
nor U11177 (N_11177,N_10105,N_10031);
xor U11178 (N_11178,N_10111,N_10389);
nand U11179 (N_11179,N_10861,N_10650);
and U11180 (N_11180,N_10048,N_10911);
nor U11181 (N_11181,N_10551,N_10378);
nor U11182 (N_11182,N_10020,N_10898);
nor U11183 (N_11183,N_10007,N_10218);
xor U11184 (N_11184,N_10237,N_10647);
or U11185 (N_11185,N_10689,N_10533);
xnor U11186 (N_11186,N_10549,N_10062);
xor U11187 (N_11187,N_10679,N_10699);
nand U11188 (N_11188,N_10901,N_10336);
xnor U11189 (N_11189,N_10329,N_10963);
or U11190 (N_11190,N_10325,N_10986);
and U11191 (N_11191,N_10682,N_10763);
or U11192 (N_11192,N_10040,N_10845);
nor U11193 (N_11193,N_10318,N_10784);
nand U11194 (N_11194,N_10649,N_10932);
or U11195 (N_11195,N_10906,N_10215);
nor U11196 (N_11196,N_10472,N_10746);
and U11197 (N_11197,N_10416,N_10017);
nor U11198 (N_11198,N_10413,N_10300);
or U11199 (N_11199,N_10924,N_10376);
nor U11200 (N_11200,N_10187,N_10660);
or U11201 (N_11201,N_10672,N_10262);
nor U11202 (N_11202,N_10195,N_10073);
nand U11203 (N_11203,N_10401,N_10110);
nand U11204 (N_11204,N_10645,N_10996);
nand U11205 (N_11205,N_10245,N_10181);
nand U11206 (N_11206,N_10210,N_10805);
xnor U11207 (N_11207,N_10547,N_10686);
and U11208 (N_11208,N_10688,N_10639);
or U11209 (N_11209,N_10617,N_10448);
xnor U11210 (N_11210,N_10523,N_10941);
xnor U11211 (N_11211,N_10143,N_10558);
nor U11212 (N_11212,N_10708,N_10150);
xor U11213 (N_11213,N_10719,N_10512);
nor U11214 (N_11214,N_10342,N_10099);
xor U11215 (N_11215,N_10011,N_10122);
xnor U11216 (N_11216,N_10526,N_10812);
nor U11217 (N_11217,N_10449,N_10600);
nor U11218 (N_11218,N_10925,N_10097);
or U11219 (N_11219,N_10590,N_10693);
xnor U11220 (N_11220,N_10899,N_10946);
xnor U11221 (N_11221,N_10543,N_10839);
xnor U11222 (N_11222,N_10793,N_10171);
or U11223 (N_11223,N_10762,N_10960);
xor U11224 (N_11224,N_10564,N_10827);
or U11225 (N_11225,N_10423,N_10891);
and U11226 (N_11226,N_10246,N_10532);
or U11227 (N_11227,N_10114,N_10279);
and U11228 (N_11228,N_10066,N_10894);
and U11229 (N_11229,N_10585,N_10967);
or U11230 (N_11230,N_10267,N_10174);
nand U11231 (N_11231,N_10823,N_10508);
nor U11232 (N_11232,N_10667,N_10668);
nand U11233 (N_11233,N_10384,N_10404);
and U11234 (N_11234,N_10373,N_10323);
xor U11235 (N_11235,N_10428,N_10436);
xnor U11236 (N_11236,N_10788,N_10635);
and U11237 (N_11237,N_10294,N_10000);
nand U11238 (N_11238,N_10580,N_10596);
nor U11239 (N_11239,N_10039,N_10223);
nand U11240 (N_11240,N_10609,N_10054);
xor U11241 (N_11241,N_10759,N_10479);
or U11242 (N_11242,N_10907,N_10936);
and U11243 (N_11243,N_10362,N_10036);
or U11244 (N_11244,N_10496,N_10714);
nor U11245 (N_11245,N_10897,N_10507);
and U11246 (N_11246,N_10705,N_10770);
xnor U11247 (N_11247,N_10736,N_10315);
nand U11248 (N_11248,N_10403,N_10979);
nand U11249 (N_11249,N_10115,N_10271);
xnor U11250 (N_11250,N_10081,N_10832);
nand U11251 (N_11251,N_10593,N_10411);
nor U11252 (N_11252,N_10874,N_10346);
and U11253 (N_11253,N_10452,N_10721);
nand U11254 (N_11254,N_10870,N_10516);
or U11255 (N_11255,N_10104,N_10556);
nand U11256 (N_11256,N_10415,N_10893);
or U11257 (N_11257,N_10425,N_10370);
or U11258 (N_11258,N_10327,N_10919);
xnor U11259 (N_11259,N_10306,N_10292);
xnor U11260 (N_11260,N_10501,N_10003);
nor U11261 (N_11261,N_10998,N_10684);
xnor U11262 (N_11262,N_10157,N_10371);
nor U11263 (N_11263,N_10975,N_10399);
and U11264 (N_11264,N_10866,N_10042);
xor U11265 (N_11265,N_10871,N_10278);
and U11266 (N_11266,N_10247,N_10356);
nand U11267 (N_11267,N_10527,N_10550);
xnor U11268 (N_11268,N_10625,N_10068);
or U11269 (N_11269,N_10160,N_10161);
nand U11270 (N_11270,N_10477,N_10126);
or U11271 (N_11271,N_10469,N_10444);
nand U11272 (N_11272,N_10312,N_10419);
and U11273 (N_11273,N_10086,N_10627);
and U11274 (N_11274,N_10426,N_10116);
nand U11275 (N_11275,N_10727,N_10299);
nor U11276 (N_11276,N_10521,N_10433);
nor U11277 (N_11277,N_10070,N_10199);
xnor U11278 (N_11278,N_10992,N_10514);
and U11279 (N_11279,N_10308,N_10085);
or U11280 (N_11280,N_10706,N_10400);
nor U11281 (N_11281,N_10032,N_10722);
and U11282 (N_11282,N_10307,N_10510);
nand U11283 (N_11283,N_10364,N_10780);
and U11284 (N_11284,N_10493,N_10226);
or U11285 (N_11285,N_10186,N_10131);
and U11286 (N_11286,N_10432,N_10922);
nand U11287 (N_11287,N_10709,N_10361);
or U11288 (N_11288,N_10120,N_10666);
and U11289 (N_11289,N_10015,N_10948);
nand U11290 (N_11290,N_10172,N_10379);
or U11291 (N_11291,N_10301,N_10579);
or U11292 (N_11292,N_10755,N_10858);
or U11293 (N_11293,N_10610,N_10197);
nand U11294 (N_11294,N_10440,N_10606);
nor U11295 (N_11295,N_10531,N_10814);
or U11296 (N_11296,N_10848,N_10061);
and U11297 (N_11297,N_10330,N_10938);
and U11298 (N_11298,N_10408,N_10655);
xnor U11299 (N_11299,N_10798,N_10430);
nor U11300 (N_11300,N_10498,N_10683);
or U11301 (N_11301,N_10712,N_10103);
or U11302 (N_11302,N_10481,N_10069);
nand U11303 (N_11303,N_10810,N_10634);
and U11304 (N_11304,N_10100,N_10889);
or U11305 (N_11305,N_10263,N_10053);
or U11306 (N_11306,N_10254,N_10599);
xnor U11307 (N_11307,N_10723,N_10811);
xnor U11308 (N_11308,N_10366,N_10733);
nor U11309 (N_11309,N_10022,N_10865);
nand U11310 (N_11310,N_10221,N_10691);
xnor U11311 (N_11311,N_10431,N_10618);
xnor U11312 (N_11312,N_10064,N_10559);
or U11313 (N_11313,N_10951,N_10890);
and U11314 (N_11314,N_10418,N_10987);
nand U11315 (N_11315,N_10969,N_10417);
and U11316 (N_11316,N_10359,N_10382);
nand U11317 (N_11317,N_10744,N_10626);
or U11318 (N_11318,N_10855,N_10305);
nor U11319 (N_11319,N_10659,N_10339);
nor U11320 (N_11320,N_10926,N_10023);
or U11321 (N_11321,N_10817,N_10978);
nor U11322 (N_11322,N_10756,N_10847);
nand U11323 (N_11323,N_10463,N_10052);
and U11324 (N_11324,N_10455,N_10748);
nand U11325 (N_11325,N_10074,N_10243);
and U11326 (N_11326,N_10228,N_10183);
nor U11327 (N_11327,N_10155,N_10133);
and U11328 (N_11328,N_10868,N_10091);
and U11329 (N_11329,N_10615,N_10658);
nand U11330 (N_11330,N_10130,N_10760);
nand U11331 (N_11331,N_10190,N_10286);
and U11332 (N_11332,N_10113,N_10562);
and U11333 (N_11333,N_10751,N_10005);
and U11334 (N_11334,N_10652,N_10165);
nor U11335 (N_11335,N_10729,N_10808);
nand U11336 (N_11336,N_10757,N_10489);
or U11337 (N_11337,N_10191,N_10275);
nor U11338 (N_11338,N_10717,N_10664);
xor U11339 (N_11339,N_10090,N_10916);
nand U11340 (N_11340,N_10205,N_10044);
nand U11341 (N_11341,N_10293,N_10589);
nand U11342 (N_11342,N_10196,N_10608);
and U11343 (N_11343,N_10258,N_10369);
xnor U11344 (N_11344,N_10224,N_10598);
and U11345 (N_11345,N_10209,N_10257);
nor U11346 (N_11346,N_10613,N_10188);
nand U11347 (N_11347,N_10025,N_10824);
nand U11348 (N_11348,N_10669,N_10506);
or U11349 (N_11349,N_10456,N_10057);
xor U11350 (N_11350,N_10707,N_10139);
nor U11351 (N_11351,N_10990,N_10127);
nand U11352 (N_11352,N_10377,N_10092);
and U11353 (N_11353,N_10725,N_10896);
nor U11354 (N_11354,N_10831,N_10518);
nand U11355 (N_11355,N_10876,N_10957);
nor U11356 (N_11356,N_10690,N_10888);
xnor U11357 (N_11357,N_10266,N_10084);
and U11358 (N_11358,N_10016,N_10121);
nor U11359 (N_11359,N_10517,N_10387);
nand U11360 (N_11360,N_10954,N_10715);
and U11361 (N_11361,N_10076,N_10198);
and U11362 (N_11362,N_10287,N_10093);
nor U11363 (N_11363,N_10581,N_10106);
or U11364 (N_11364,N_10240,N_10662);
xnor U11365 (N_11365,N_10961,N_10538);
and U11366 (N_11366,N_10283,N_10184);
nor U11367 (N_11367,N_10177,N_10168);
and U11368 (N_11368,N_10692,N_10680);
nand U11369 (N_11369,N_10435,N_10214);
nor U11370 (N_11370,N_10145,N_10049);
nor U11371 (N_11371,N_10779,N_10794);
or U11372 (N_11372,N_10504,N_10796);
or U11373 (N_11373,N_10491,N_10309);
nor U11374 (N_11374,N_10966,N_10778);
and U11375 (N_11375,N_10804,N_10075);
nand U11376 (N_11376,N_10993,N_10716);
nand U11377 (N_11377,N_10019,N_10698);
nor U11378 (N_11378,N_10179,N_10333);
and U11379 (N_11379,N_10886,N_10785);
xnor U11380 (N_11380,N_10476,N_10604);
nand U11381 (N_11381,N_10766,N_10276);
or U11382 (N_11382,N_10576,N_10459);
nor U11383 (N_11383,N_10637,N_10653);
nand U11384 (N_11384,N_10398,N_10648);
xor U11385 (N_11385,N_10102,N_10909);
nand U11386 (N_11386,N_10701,N_10927);
nor U11387 (N_11387,N_10499,N_10193);
nor U11388 (N_11388,N_10622,N_10482);
xor U11389 (N_11389,N_10483,N_10478);
nand U11390 (N_11390,N_10694,N_10765);
nor U11391 (N_11391,N_10937,N_10273);
nand U11392 (N_11392,N_10446,N_10238);
xor U11393 (N_11393,N_10466,N_10166);
nand U11394 (N_11394,N_10169,N_10834);
nor U11395 (N_11395,N_10268,N_10867);
nor U11396 (N_11396,N_10180,N_10536);
nand U11397 (N_11397,N_10849,N_10964);
nor U11398 (N_11398,N_10388,N_10671);
and U11399 (N_11399,N_10883,N_10904);
nor U11400 (N_11400,N_10232,N_10525);
nor U11401 (N_11401,N_10353,N_10656);
nor U11402 (N_11402,N_10792,N_10176);
nand U11403 (N_11403,N_10702,N_10724);
xnor U11404 (N_11404,N_10815,N_10773);
or U11405 (N_11405,N_10326,N_10620);
or U11406 (N_11406,N_10718,N_10394);
or U11407 (N_11407,N_10586,N_10821);
or U11408 (N_11408,N_10332,N_10043);
nand U11409 (N_11409,N_10802,N_10970);
nand U11410 (N_11410,N_10438,N_10740);
or U11411 (N_11411,N_10782,N_10468);
and U11412 (N_11412,N_10473,N_10687);
nor U11413 (N_11413,N_10194,N_10594);
nor U11414 (N_11414,N_10743,N_10050);
nor U11415 (N_11415,N_10628,N_10441);
nand U11416 (N_11416,N_10119,N_10977);
nand U11417 (N_11417,N_10217,N_10087);
nor U11418 (N_11418,N_10843,N_10386);
or U11419 (N_11419,N_10560,N_10272);
nor U11420 (N_11420,N_10465,N_10260);
xnor U11421 (N_11421,N_10347,N_10939);
nor U11422 (N_11422,N_10175,N_10949);
xor U11423 (N_11423,N_10321,N_10546);
xor U11424 (N_11424,N_10952,N_10414);
nor U11425 (N_11425,N_10443,N_10879);
nand U11426 (N_11426,N_10392,N_10124);
nand U11427 (N_11427,N_10038,N_10741);
nor U11428 (N_11428,N_10354,N_10605);
nand U11429 (N_11429,N_10767,N_10524);
xnor U11430 (N_11430,N_10542,N_10797);
and U11431 (N_11431,N_10520,N_10288);
or U11432 (N_11432,N_10958,N_10582);
or U11433 (N_11433,N_10540,N_10368);
xor U11434 (N_11434,N_10592,N_10324);
and U11435 (N_11435,N_10357,N_10204);
and U11436 (N_11436,N_10999,N_10335);
xor U11437 (N_11437,N_10457,N_10138);
and U11438 (N_11438,N_10437,N_10227);
and U11439 (N_11439,N_10351,N_10885);
or U11440 (N_11440,N_10752,N_10407);
nor U11441 (N_11441,N_10974,N_10908);
xor U11442 (N_11442,N_10548,N_10892);
nor U11443 (N_11443,N_10393,N_10159);
nor U11444 (N_11444,N_10732,N_10920);
or U11445 (N_11445,N_10621,N_10563);
xnor U11446 (N_11446,N_10895,N_10681);
nand U11447 (N_11447,N_10775,N_10421);
xnor U11448 (N_11448,N_10923,N_10988);
nand U11449 (N_11449,N_10024,N_10875);
xnor U11450 (N_11450,N_10345,N_10219);
nor U11451 (N_11451,N_10629,N_10153);
nor U11452 (N_11452,N_10500,N_10447);
nor U11453 (N_11453,N_10643,N_10577);
and U11454 (N_11454,N_10537,N_10857);
and U11455 (N_11455,N_10148,N_10234);
and U11456 (N_11456,N_10820,N_10959);
xnor U11457 (N_11457,N_10535,N_10640);
nor U11458 (N_11458,N_10424,N_10887);
nor U11459 (N_11459,N_10769,N_10503);
and U11460 (N_11460,N_10670,N_10492);
xnor U11461 (N_11461,N_10154,N_10178);
nand U11462 (N_11462,N_10734,N_10239);
and U11463 (N_11463,N_10541,N_10460);
nor U11464 (N_11464,N_10470,N_10654);
nand U11465 (N_11465,N_10728,N_10220);
or U11466 (N_11466,N_10006,N_10461);
xor U11467 (N_11467,N_10134,N_10777);
nor U11468 (N_11468,N_10983,N_10673);
xor U11469 (N_11469,N_10913,N_10962);
and U11470 (N_11470,N_10614,N_10781);
nand U11471 (N_11471,N_10940,N_10758);
nand U11472 (N_11472,N_10012,N_10587);
nor U11473 (N_11473,N_10236,N_10529);
nand U11474 (N_11474,N_10557,N_10641);
or U11475 (N_11475,N_10631,N_10505);
or U11476 (N_11476,N_10409,N_10454);
or U11477 (N_11477,N_10285,N_10835);
xnor U11478 (N_11478,N_10588,N_10297);
or U11479 (N_11479,N_10965,N_10661);
xor U11480 (N_11480,N_10646,N_10083);
and U11481 (N_11481,N_10203,N_10676);
nand U11482 (N_11482,N_10695,N_10616);
nand U11483 (N_11483,N_10495,N_10067);
or U11484 (N_11484,N_10800,N_10167);
xor U11485 (N_11485,N_10340,N_10972);
and U11486 (N_11486,N_10644,N_10355);
and U11487 (N_11487,N_10152,N_10502);
and U11488 (N_11488,N_10842,N_10511);
nand U11489 (N_11489,N_10302,N_10311);
nand U11490 (N_11490,N_10095,N_10995);
nor U11491 (N_11491,N_10046,N_10943);
or U11492 (N_11492,N_10602,N_10685);
xor U11493 (N_11493,N_10799,N_10002);
and U11494 (N_11494,N_10008,N_10041);
or U11495 (N_11495,N_10739,N_10720);
or U11496 (N_11496,N_10107,N_10358);
and U11497 (N_11497,N_10290,N_10864);
nor U11498 (N_11498,N_10310,N_10595);
xnor U11499 (N_11499,N_10251,N_10296);
nand U11500 (N_11500,N_10231,N_10901);
nor U11501 (N_11501,N_10078,N_10383);
nand U11502 (N_11502,N_10372,N_10958);
xor U11503 (N_11503,N_10151,N_10305);
or U11504 (N_11504,N_10000,N_10987);
and U11505 (N_11505,N_10915,N_10049);
xor U11506 (N_11506,N_10887,N_10686);
or U11507 (N_11507,N_10024,N_10877);
or U11508 (N_11508,N_10356,N_10677);
or U11509 (N_11509,N_10813,N_10379);
or U11510 (N_11510,N_10105,N_10120);
and U11511 (N_11511,N_10288,N_10028);
and U11512 (N_11512,N_10818,N_10470);
and U11513 (N_11513,N_10184,N_10985);
or U11514 (N_11514,N_10434,N_10903);
nand U11515 (N_11515,N_10101,N_10133);
and U11516 (N_11516,N_10255,N_10260);
nand U11517 (N_11517,N_10569,N_10184);
and U11518 (N_11518,N_10861,N_10220);
and U11519 (N_11519,N_10357,N_10330);
nor U11520 (N_11520,N_10250,N_10494);
nor U11521 (N_11521,N_10577,N_10805);
and U11522 (N_11522,N_10310,N_10623);
or U11523 (N_11523,N_10073,N_10637);
nand U11524 (N_11524,N_10146,N_10736);
and U11525 (N_11525,N_10843,N_10871);
xnor U11526 (N_11526,N_10483,N_10538);
xor U11527 (N_11527,N_10877,N_10335);
xnor U11528 (N_11528,N_10602,N_10663);
nand U11529 (N_11529,N_10298,N_10945);
and U11530 (N_11530,N_10355,N_10660);
or U11531 (N_11531,N_10348,N_10316);
nor U11532 (N_11532,N_10367,N_10839);
and U11533 (N_11533,N_10570,N_10883);
nand U11534 (N_11534,N_10507,N_10583);
xnor U11535 (N_11535,N_10606,N_10698);
or U11536 (N_11536,N_10951,N_10865);
and U11537 (N_11537,N_10897,N_10481);
and U11538 (N_11538,N_10528,N_10891);
or U11539 (N_11539,N_10012,N_10496);
xor U11540 (N_11540,N_10426,N_10527);
nand U11541 (N_11541,N_10121,N_10448);
nor U11542 (N_11542,N_10353,N_10102);
nor U11543 (N_11543,N_10885,N_10207);
or U11544 (N_11544,N_10224,N_10689);
or U11545 (N_11545,N_10505,N_10138);
nand U11546 (N_11546,N_10952,N_10873);
and U11547 (N_11547,N_10651,N_10421);
and U11548 (N_11548,N_10739,N_10741);
nand U11549 (N_11549,N_10664,N_10628);
xnor U11550 (N_11550,N_10291,N_10820);
xor U11551 (N_11551,N_10804,N_10422);
xor U11552 (N_11552,N_10796,N_10486);
or U11553 (N_11553,N_10589,N_10156);
nor U11554 (N_11554,N_10629,N_10749);
or U11555 (N_11555,N_10025,N_10390);
nor U11556 (N_11556,N_10044,N_10308);
or U11557 (N_11557,N_10826,N_10125);
and U11558 (N_11558,N_10726,N_10986);
or U11559 (N_11559,N_10237,N_10732);
nand U11560 (N_11560,N_10001,N_10145);
and U11561 (N_11561,N_10159,N_10126);
nand U11562 (N_11562,N_10429,N_10057);
xor U11563 (N_11563,N_10912,N_10418);
or U11564 (N_11564,N_10648,N_10796);
nand U11565 (N_11565,N_10995,N_10880);
nor U11566 (N_11566,N_10247,N_10843);
nand U11567 (N_11567,N_10489,N_10792);
xnor U11568 (N_11568,N_10860,N_10088);
or U11569 (N_11569,N_10516,N_10981);
or U11570 (N_11570,N_10552,N_10085);
and U11571 (N_11571,N_10519,N_10503);
or U11572 (N_11572,N_10410,N_10137);
or U11573 (N_11573,N_10170,N_10134);
xor U11574 (N_11574,N_10903,N_10304);
and U11575 (N_11575,N_10768,N_10030);
nand U11576 (N_11576,N_10168,N_10682);
nand U11577 (N_11577,N_10852,N_10874);
xnor U11578 (N_11578,N_10237,N_10004);
or U11579 (N_11579,N_10277,N_10223);
nand U11580 (N_11580,N_10078,N_10455);
and U11581 (N_11581,N_10823,N_10425);
and U11582 (N_11582,N_10844,N_10153);
and U11583 (N_11583,N_10432,N_10695);
xnor U11584 (N_11584,N_10585,N_10878);
nand U11585 (N_11585,N_10745,N_10605);
or U11586 (N_11586,N_10303,N_10475);
and U11587 (N_11587,N_10135,N_10455);
xor U11588 (N_11588,N_10246,N_10355);
nor U11589 (N_11589,N_10433,N_10001);
nand U11590 (N_11590,N_10020,N_10418);
xnor U11591 (N_11591,N_10239,N_10423);
or U11592 (N_11592,N_10576,N_10334);
and U11593 (N_11593,N_10479,N_10561);
nand U11594 (N_11594,N_10722,N_10639);
and U11595 (N_11595,N_10426,N_10576);
xor U11596 (N_11596,N_10885,N_10972);
and U11597 (N_11597,N_10994,N_10422);
nor U11598 (N_11598,N_10591,N_10502);
and U11599 (N_11599,N_10730,N_10274);
or U11600 (N_11600,N_10496,N_10727);
nor U11601 (N_11601,N_10610,N_10618);
or U11602 (N_11602,N_10881,N_10796);
and U11603 (N_11603,N_10117,N_10177);
and U11604 (N_11604,N_10321,N_10621);
xnor U11605 (N_11605,N_10833,N_10932);
xnor U11606 (N_11606,N_10712,N_10054);
and U11607 (N_11607,N_10306,N_10231);
nand U11608 (N_11608,N_10819,N_10331);
or U11609 (N_11609,N_10154,N_10456);
or U11610 (N_11610,N_10837,N_10158);
nor U11611 (N_11611,N_10761,N_10602);
or U11612 (N_11612,N_10157,N_10687);
nor U11613 (N_11613,N_10026,N_10601);
or U11614 (N_11614,N_10117,N_10300);
nand U11615 (N_11615,N_10704,N_10687);
or U11616 (N_11616,N_10201,N_10800);
or U11617 (N_11617,N_10005,N_10368);
xnor U11618 (N_11618,N_10922,N_10464);
nand U11619 (N_11619,N_10410,N_10339);
xor U11620 (N_11620,N_10564,N_10573);
nand U11621 (N_11621,N_10204,N_10460);
xor U11622 (N_11622,N_10039,N_10893);
and U11623 (N_11623,N_10835,N_10034);
and U11624 (N_11624,N_10801,N_10001);
xor U11625 (N_11625,N_10193,N_10070);
and U11626 (N_11626,N_10962,N_10929);
and U11627 (N_11627,N_10198,N_10417);
or U11628 (N_11628,N_10577,N_10972);
or U11629 (N_11629,N_10468,N_10274);
nor U11630 (N_11630,N_10300,N_10689);
or U11631 (N_11631,N_10694,N_10163);
and U11632 (N_11632,N_10401,N_10763);
and U11633 (N_11633,N_10323,N_10281);
nand U11634 (N_11634,N_10674,N_10390);
and U11635 (N_11635,N_10705,N_10563);
xor U11636 (N_11636,N_10513,N_10425);
or U11637 (N_11637,N_10768,N_10595);
and U11638 (N_11638,N_10844,N_10042);
nor U11639 (N_11639,N_10152,N_10614);
or U11640 (N_11640,N_10453,N_10006);
xor U11641 (N_11641,N_10168,N_10992);
nand U11642 (N_11642,N_10627,N_10263);
nor U11643 (N_11643,N_10678,N_10114);
nand U11644 (N_11644,N_10512,N_10300);
and U11645 (N_11645,N_10237,N_10637);
or U11646 (N_11646,N_10522,N_10406);
and U11647 (N_11647,N_10463,N_10083);
nand U11648 (N_11648,N_10123,N_10647);
and U11649 (N_11649,N_10326,N_10145);
nor U11650 (N_11650,N_10597,N_10769);
nand U11651 (N_11651,N_10489,N_10373);
nor U11652 (N_11652,N_10526,N_10981);
and U11653 (N_11653,N_10546,N_10956);
nor U11654 (N_11654,N_10230,N_10534);
nor U11655 (N_11655,N_10841,N_10936);
or U11656 (N_11656,N_10603,N_10516);
xor U11657 (N_11657,N_10828,N_10396);
or U11658 (N_11658,N_10651,N_10386);
nor U11659 (N_11659,N_10150,N_10588);
and U11660 (N_11660,N_10875,N_10122);
or U11661 (N_11661,N_10569,N_10331);
nor U11662 (N_11662,N_10594,N_10026);
nand U11663 (N_11663,N_10234,N_10380);
and U11664 (N_11664,N_10772,N_10204);
nand U11665 (N_11665,N_10088,N_10069);
nor U11666 (N_11666,N_10756,N_10589);
and U11667 (N_11667,N_10136,N_10341);
nand U11668 (N_11668,N_10361,N_10956);
and U11669 (N_11669,N_10929,N_10222);
and U11670 (N_11670,N_10328,N_10697);
or U11671 (N_11671,N_10642,N_10688);
xnor U11672 (N_11672,N_10505,N_10230);
xor U11673 (N_11673,N_10204,N_10312);
or U11674 (N_11674,N_10768,N_10445);
and U11675 (N_11675,N_10917,N_10579);
xnor U11676 (N_11676,N_10046,N_10689);
xnor U11677 (N_11677,N_10247,N_10204);
xor U11678 (N_11678,N_10009,N_10131);
xnor U11679 (N_11679,N_10285,N_10139);
nor U11680 (N_11680,N_10335,N_10449);
and U11681 (N_11681,N_10308,N_10347);
xor U11682 (N_11682,N_10991,N_10992);
or U11683 (N_11683,N_10963,N_10007);
nor U11684 (N_11684,N_10463,N_10819);
and U11685 (N_11685,N_10601,N_10226);
or U11686 (N_11686,N_10187,N_10550);
nand U11687 (N_11687,N_10410,N_10032);
xor U11688 (N_11688,N_10447,N_10806);
or U11689 (N_11689,N_10721,N_10120);
nor U11690 (N_11690,N_10079,N_10988);
and U11691 (N_11691,N_10629,N_10782);
and U11692 (N_11692,N_10067,N_10513);
nand U11693 (N_11693,N_10722,N_10204);
or U11694 (N_11694,N_10761,N_10433);
nand U11695 (N_11695,N_10293,N_10544);
or U11696 (N_11696,N_10272,N_10216);
or U11697 (N_11697,N_10143,N_10698);
nor U11698 (N_11698,N_10527,N_10729);
and U11699 (N_11699,N_10407,N_10184);
nor U11700 (N_11700,N_10588,N_10343);
xnor U11701 (N_11701,N_10719,N_10343);
or U11702 (N_11702,N_10575,N_10150);
nand U11703 (N_11703,N_10981,N_10260);
xor U11704 (N_11704,N_10663,N_10703);
and U11705 (N_11705,N_10768,N_10183);
and U11706 (N_11706,N_10793,N_10986);
nor U11707 (N_11707,N_10473,N_10326);
nor U11708 (N_11708,N_10188,N_10909);
nor U11709 (N_11709,N_10559,N_10346);
and U11710 (N_11710,N_10430,N_10859);
and U11711 (N_11711,N_10164,N_10330);
xor U11712 (N_11712,N_10951,N_10472);
and U11713 (N_11713,N_10671,N_10658);
xor U11714 (N_11714,N_10143,N_10681);
and U11715 (N_11715,N_10136,N_10849);
or U11716 (N_11716,N_10091,N_10096);
or U11717 (N_11717,N_10772,N_10343);
xor U11718 (N_11718,N_10144,N_10195);
nor U11719 (N_11719,N_10777,N_10318);
and U11720 (N_11720,N_10007,N_10923);
and U11721 (N_11721,N_10699,N_10191);
xor U11722 (N_11722,N_10684,N_10744);
nand U11723 (N_11723,N_10419,N_10562);
or U11724 (N_11724,N_10492,N_10299);
xor U11725 (N_11725,N_10916,N_10010);
nor U11726 (N_11726,N_10067,N_10928);
and U11727 (N_11727,N_10100,N_10163);
xor U11728 (N_11728,N_10080,N_10921);
or U11729 (N_11729,N_10945,N_10606);
nor U11730 (N_11730,N_10256,N_10835);
xnor U11731 (N_11731,N_10615,N_10796);
or U11732 (N_11732,N_10650,N_10616);
and U11733 (N_11733,N_10836,N_10499);
or U11734 (N_11734,N_10862,N_10051);
xnor U11735 (N_11735,N_10288,N_10223);
xnor U11736 (N_11736,N_10966,N_10265);
xnor U11737 (N_11737,N_10571,N_10557);
nand U11738 (N_11738,N_10819,N_10686);
nor U11739 (N_11739,N_10981,N_10655);
xnor U11740 (N_11740,N_10381,N_10895);
and U11741 (N_11741,N_10226,N_10127);
xor U11742 (N_11742,N_10221,N_10184);
or U11743 (N_11743,N_10913,N_10021);
nor U11744 (N_11744,N_10762,N_10879);
nand U11745 (N_11745,N_10286,N_10775);
and U11746 (N_11746,N_10540,N_10476);
and U11747 (N_11747,N_10475,N_10876);
nand U11748 (N_11748,N_10264,N_10392);
and U11749 (N_11749,N_10410,N_10634);
and U11750 (N_11750,N_10052,N_10898);
nor U11751 (N_11751,N_10549,N_10944);
and U11752 (N_11752,N_10149,N_10224);
nand U11753 (N_11753,N_10262,N_10243);
or U11754 (N_11754,N_10396,N_10195);
xnor U11755 (N_11755,N_10588,N_10793);
and U11756 (N_11756,N_10000,N_10586);
or U11757 (N_11757,N_10130,N_10488);
nand U11758 (N_11758,N_10394,N_10601);
and U11759 (N_11759,N_10630,N_10573);
nand U11760 (N_11760,N_10964,N_10599);
and U11761 (N_11761,N_10947,N_10418);
or U11762 (N_11762,N_10512,N_10142);
xor U11763 (N_11763,N_10066,N_10598);
nand U11764 (N_11764,N_10275,N_10881);
or U11765 (N_11765,N_10609,N_10801);
xor U11766 (N_11766,N_10401,N_10892);
or U11767 (N_11767,N_10986,N_10758);
or U11768 (N_11768,N_10736,N_10024);
xnor U11769 (N_11769,N_10318,N_10914);
and U11770 (N_11770,N_10470,N_10708);
nand U11771 (N_11771,N_10609,N_10780);
and U11772 (N_11772,N_10442,N_10688);
nor U11773 (N_11773,N_10913,N_10093);
nand U11774 (N_11774,N_10265,N_10377);
nor U11775 (N_11775,N_10754,N_10152);
or U11776 (N_11776,N_10568,N_10406);
nor U11777 (N_11777,N_10972,N_10411);
nand U11778 (N_11778,N_10180,N_10669);
and U11779 (N_11779,N_10914,N_10404);
or U11780 (N_11780,N_10268,N_10227);
nor U11781 (N_11781,N_10950,N_10741);
and U11782 (N_11782,N_10124,N_10532);
nor U11783 (N_11783,N_10842,N_10009);
and U11784 (N_11784,N_10310,N_10492);
nor U11785 (N_11785,N_10304,N_10413);
nor U11786 (N_11786,N_10013,N_10343);
nand U11787 (N_11787,N_10508,N_10810);
nor U11788 (N_11788,N_10291,N_10899);
xnor U11789 (N_11789,N_10998,N_10704);
or U11790 (N_11790,N_10056,N_10458);
nand U11791 (N_11791,N_10328,N_10620);
xor U11792 (N_11792,N_10620,N_10356);
nor U11793 (N_11793,N_10867,N_10810);
nor U11794 (N_11794,N_10745,N_10624);
nor U11795 (N_11795,N_10982,N_10479);
nand U11796 (N_11796,N_10530,N_10545);
and U11797 (N_11797,N_10984,N_10286);
xor U11798 (N_11798,N_10920,N_10844);
nor U11799 (N_11799,N_10602,N_10815);
xor U11800 (N_11800,N_10960,N_10259);
xor U11801 (N_11801,N_10854,N_10568);
xor U11802 (N_11802,N_10823,N_10291);
nand U11803 (N_11803,N_10938,N_10353);
and U11804 (N_11804,N_10818,N_10815);
and U11805 (N_11805,N_10673,N_10145);
xnor U11806 (N_11806,N_10841,N_10703);
and U11807 (N_11807,N_10539,N_10327);
xnor U11808 (N_11808,N_10329,N_10177);
or U11809 (N_11809,N_10753,N_10443);
nor U11810 (N_11810,N_10045,N_10487);
or U11811 (N_11811,N_10063,N_10340);
or U11812 (N_11812,N_10436,N_10225);
nand U11813 (N_11813,N_10992,N_10211);
and U11814 (N_11814,N_10331,N_10241);
or U11815 (N_11815,N_10550,N_10460);
nand U11816 (N_11816,N_10395,N_10007);
or U11817 (N_11817,N_10086,N_10991);
nor U11818 (N_11818,N_10637,N_10823);
nand U11819 (N_11819,N_10321,N_10168);
nor U11820 (N_11820,N_10149,N_10330);
xnor U11821 (N_11821,N_10651,N_10970);
nor U11822 (N_11822,N_10457,N_10008);
and U11823 (N_11823,N_10750,N_10222);
xor U11824 (N_11824,N_10222,N_10709);
nand U11825 (N_11825,N_10035,N_10791);
nand U11826 (N_11826,N_10016,N_10070);
or U11827 (N_11827,N_10611,N_10610);
xnor U11828 (N_11828,N_10023,N_10378);
or U11829 (N_11829,N_10348,N_10446);
and U11830 (N_11830,N_10252,N_10814);
and U11831 (N_11831,N_10375,N_10119);
nand U11832 (N_11832,N_10445,N_10384);
and U11833 (N_11833,N_10000,N_10258);
nor U11834 (N_11834,N_10506,N_10931);
xor U11835 (N_11835,N_10488,N_10709);
and U11836 (N_11836,N_10351,N_10255);
nand U11837 (N_11837,N_10592,N_10090);
and U11838 (N_11838,N_10927,N_10844);
and U11839 (N_11839,N_10334,N_10836);
nand U11840 (N_11840,N_10518,N_10514);
nand U11841 (N_11841,N_10675,N_10089);
and U11842 (N_11842,N_10201,N_10266);
and U11843 (N_11843,N_10503,N_10890);
or U11844 (N_11844,N_10709,N_10859);
xnor U11845 (N_11845,N_10598,N_10712);
nand U11846 (N_11846,N_10305,N_10689);
nor U11847 (N_11847,N_10185,N_10274);
nand U11848 (N_11848,N_10582,N_10118);
nor U11849 (N_11849,N_10378,N_10416);
or U11850 (N_11850,N_10694,N_10872);
or U11851 (N_11851,N_10157,N_10021);
nor U11852 (N_11852,N_10501,N_10978);
nand U11853 (N_11853,N_10254,N_10047);
and U11854 (N_11854,N_10946,N_10905);
and U11855 (N_11855,N_10859,N_10846);
or U11856 (N_11856,N_10497,N_10631);
or U11857 (N_11857,N_10523,N_10852);
xnor U11858 (N_11858,N_10887,N_10347);
xor U11859 (N_11859,N_10155,N_10204);
nor U11860 (N_11860,N_10781,N_10523);
nor U11861 (N_11861,N_10589,N_10056);
or U11862 (N_11862,N_10814,N_10545);
xnor U11863 (N_11863,N_10519,N_10406);
or U11864 (N_11864,N_10023,N_10826);
nand U11865 (N_11865,N_10104,N_10021);
and U11866 (N_11866,N_10758,N_10176);
and U11867 (N_11867,N_10003,N_10115);
nand U11868 (N_11868,N_10291,N_10011);
nor U11869 (N_11869,N_10542,N_10817);
and U11870 (N_11870,N_10960,N_10802);
or U11871 (N_11871,N_10146,N_10579);
and U11872 (N_11872,N_10153,N_10299);
and U11873 (N_11873,N_10295,N_10557);
or U11874 (N_11874,N_10569,N_10522);
xnor U11875 (N_11875,N_10944,N_10686);
nand U11876 (N_11876,N_10471,N_10407);
nor U11877 (N_11877,N_10292,N_10778);
and U11878 (N_11878,N_10567,N_10219);
xnor U11879 (N_11879,N_10633,N_10593);
or U11880 (N_11880,N_10007,N_10379);
nand U11881 (N_11881,N_10749,N_10030);
nor U11882 (N_11882,N_10163,N_10143);
nand U11883 (N_11883,N_10945,N_10610);
nand U11884 (N_11884,N_10033,N_10364);
nor U11885 (N_11885,N_10922,N_10598);
and U11886 (N_11886,N_10253,N_10417);
and U11887 (N_11887,N_10006,N_10280);
nand U11888 (N_11888,N_10395,N_10796);
or U11889 (N_11889,N_10385,N_10170);
nor U11890 (N_11890,N_10281,N_10993);
xor U11891 (N_11891,N_10626,N_10443);
or U11892 (N_11892,N_10078,N_10158);
or U11893 (N_11893,N_10183,N_10885);
nor U11894 (N_11894,N_10564,N_10642);
and U11895 (N_11895,N_10903,N_10220);
nand U11896 (N_11896,N_10993,N_10685);
nand U11897 (N_11897,N_10954,N_10953);
nand U11898 (N_11898,N_10054,N_10434);
nor U11899 (N_11899,N_10814,N_10377);
and U11900 (N_11900,N_10028,N_10493);
xnor U11901 (N_11901,N_10068,N_10619);
nor U11902 (N_11902,N_10856,N_10316);
and U11903 (N_11903,N_10280,N_10252);
and U11904 (N_11904,N_10223,N_10768);
and U11905 (N_11905,N_10094,N_10319);
or U11906 (N_11906,N_10219,N_10690);
nand U11907 (N_11907,N_10690,N_10064);
nand U11908 (N_11908,N_10319,N_10179);
nand U11909 (N_11909,N_10229,N_10088);
or U11910 (N_11910,N_10726,N_10072);
nand U11911 (N_11911,N_10243,N_10943);
xnor U11912 (N_11912,N_10445,N_10264);
and U11913 (N_11913,N_10240,N_10533);
nor U11914 (N_11914,N_10400,N_10141);
and U11915 (N_11915,N_10252,N_10384);
nor U11916 (N_11916,N_10118,N_10431);
and U11917 (N_11917,N_10802,N_10888);
xor U11918 (N_11918,N_10235,N_10464);
nor U11919 (N_11919,N_10263,N_10758);
xor U11920 (N_11920,N_10841,N_10635);
or U11921 (N_11921,N_10160,N_10152);
xnor U11922 (N_11922,N_10627,N_10316);
and U11923 (N_11923,N_10800,N_10814);
or U11924 (N_11924,N_10220,N_10471);
and U11925 (N_11925,N_10680,N_10315);
and U11926 (N_11926,N_10713,N_10968);
nor U11927 (N_11927,N_10338,N_10781);
and U11928 (N_11928,N_10549,N_10138);
nand U11929 (N_11929,N_10274,N_10227);
or U11930 (N_11930,N_10943,N_10830);
xor U11931 (N_11931,N_10839,N_10605);
xor U11932 (N_11932,N_10556,N_10337);
nor U11933 (N_11933,N_10613,N_10130);
nand U11934 (N_11934,N_10966,N_10026);
nor U11935 (N_11935,N_10809,N_10790);
nor U11936 (N_11936,N_10516,N_10841);
nor U11937 (N_11937,N_10625,N_10735);
nand U11938 (N_11938,N_10414,N_10089);
nand U11939 (N_11939,N_10619,N_10213);
nor U11940 (N_11940,N_10307,N_10501);
nand U11941 (N_11941,N_10522,N_10769);
and U11942 (N_11942,N_10076,N_10624);
or U11943 (N_11943,N_10543,N_10100);
and U11944 (N_11944,N_10323,N_10933);
xnor U11945 (N_11945,N_10691,N_10589);
xor U11946 (N_11946,N_10430,N_10505);
xnor U11947 (N_11947,N_10548,N_10037);
nand U11948 (N_11948,N_10065,N_10631);
xor U11949 (N_11949,N_10338,N_10897);
or U11950 (N_11950,N_10621,N_10122);
nor U11951 (N_11951,N_10266,N_10687);
nand U11952 (N_11952,N_10514,N_10714);
and U11953 (N_11953,N_10289,N_10567);
or U11954 (N_11954,N_10232,N_10777);
xnor U11955 (N_11955,N_10870,N_10700);
or U11956 (N_11956,N_10664,N_10888);
xor U11957 (N_11957,N_10181,N_10264);
xnor U11958 (N_11958,N_10592,N_10392);
nor U11959 (N_11959,N_10939,N_10780);
and U11960 (N_11960,N_10804,N_10458);
and U11961 (N_11961,N_10080,N_10176);
nor U11962 (N_11962,N_10895,N_10240);
xnor U11963 (N_11963,N_10639,N_10144);
or U11964 (N_11964,N_10966,N_10551);
or U11965 (N_11965,N_10363,N_10150);
or U11966 (N_11966,N_10618,N_10860);
nor U11967 (N_11967,N_10421,N_10926);
or U11968 (N_11968,N_10063,N_10047);
xor U11969 (N_11969,N_10173,N_10860);
nand U11970 (N_11970,N_10311,N_10035);
and U11971 (N_11971,N_10213,N_10488);
or U11972 (N_11972,N_10483,N_10200);
or U11973 (N_11973,N_10492,N_10458);
or U11974 (N_11974,N_10237,N_10714);
and U11975 (N_11975,N_10781,N_10991);
or U11976 (N_11976,N_10310,N_10477);
nand U11977 (N_11977,N_10962,N_10887);
nor U11978 (N_11978,N_10757,N_10238);
nand U11979 (N_11979,N_10088,N_10842);
xnor U11980 (N_11980,N_10066,N_10481);
nand U11981 (N_11981,N_10258,N_10930);
nand U11982 (N_11982,N_10602,N_10333);
xnor U11983 (N_11983,N_10537,N_10538);
nor U11984 (N_11984,N_10263,N_10655);
and U11985 (N_11985,N_10974,N_10929);
nand U11986 (N_11986,N_10682,N_10133);
nand U11987 (N_11987,N_10618,N_10273);
nand U11988 (N_11988,N_10625,N_10342);
xor U11989 (N_11989,N_10176,N_10608);
xor U11990 (N_11990,N_10898,N_10292);
xor U11991 (N_11991,N_10424,N_10674);
xnor U11992 (N_11992,N_10987,N_10110);
xor U11993 (N_11993,N_10765,N_10818);
or U11994 (N_11994,N_10613,N_10679);
nor U11995 (N_11995,N_10957,N_10046);
nand U11996 (N_11996,N_10969,N_10184);
nor U11997 (N_11997,N_10052,N_10621);
or U11998 (N_11998,N_10934,N_10509);
or U11999 (N_11999,N_10823,N_10619);
nand U12000 (N_12000,N_11956,N_11831);
xor U12001 (N_12001,N_11420,N_11302);
nand U12002 (N_12002,N_11224,N_11691);
or U12003 (N_12003,N_11776,N_11978);
nor U12004 (N_12004,N_11267,N_11493);
or U12005 (N_12005,N_11836,N_11027);
and U12006 (N_12006,N_11929,N_11479);
and U12007 (N_12007,N_11094,N_11835);
nor U12008 (N_12008,N_11780,N_11883);
and U12009 (N_12009,N_11706,N_11939);
and U12010 (N_12010,N_11797,N_11312);
nand U12011 (N_12011,N_11904,N_11033);
nand U12012 (N_12012,N_11752,N_11503);
nand U12013 (N_12013,N_11018,N_11363);
nor U12014 (N_12014,N_11130,N_11171);
nand U12015 (N_12015,N_11671,N_11062);
and U12016 (N_12016,N_11680,N_11807);
nand U12017 (N_12017,N_11458,N_11051);
nand U12018 (N_12018,N_11150,N_11377);
or U12019 (N_12019,N_11481,N_11976);
nand U12020 (N_12020,N_11996,N_11136);
or U12021 (N_12021,N_11915,N_11186);
nor U12022 (N_12022,N_11057,N_11974);
nor U12023 (N_12023,N_11355,N_11176);
or U12024 (N_12024,N_11554,N_11701);
and U12025 (N_12025,N_11007,N_11813);
and U12026 (N_12026,N_11060,N_11622);
xor U12027 (N_12027,N_11669,N_11046);
nand U12028 (N_12028,N_11574,N_11991);
and U12029 (N_12029,N_11360,N_11695);
or U12030 (N_12030,N_11812,N_11958);
xor U12031 (N_12031,N_11521,N_11153);
nor U12032 (N_12032,N_11539,N_11488);
xnor U12033 (N_12033,N_11876,N_11860);
and U12034 (N_12034,N_11029,N_11205);
nor U12035 (N_12035,N_11855,N_11803);
or U12036 (N_12036,N_11347,N_11160);
xnor U12037 (N_12037,N_11453,N_11167);
xor U12038 (N_12038,N_11228,N_11432);
nand U12039 (N_12039,N_11074,N_11700);
nor U12040 (N_12040,N_11418,N_11945);
or U12041 (N_12041,N_11576,N_11044);
or U12042 (N_12042,N_11537,N_11102);
nand U12043 (N_12043,N_11424,N_11278);
nand U12044 (N_12044,N_11392,N_11485);
and U12045 (N_12045,N_11291,N_11705);
xnor U12046 (N_12046,N_11200,N_11838);
and U12047 (N_12047,N_11848,N_11529);
nor U12048 (N_12048,N_11384,N_11082);
xnor U12049 (N_12049,N_11623,N_11567);
nand U12050 (N_12050,N_11434,N_11282);
xnor U12051 (N_12051,N_11548,N_11744);
xnor U12052 (N_12052,N_11353,N_11947);
nand U12053 (N_12053,N_11735,N_11506);
nand U12054 (N_12054,N_11526,N_11229);
nor U12055 (N_12055,N_11533,N_11842);
or U12056 (N_12056,N_11024,N_11422);
nand U12057 (N_12057,N_11988,N_11818);
and U12058 (N_12058,N_11568,N_11254);
or U12059 (N_12059,N_11294,N_11239);
xor U12060 (N_12060,N_11374,N_11937);
and U12061 (N_12061,N_11115,N_11206);
xnor U12062 (N_12062,N_11452,N_11738);
and U12063 (N_12063,N_11647,N_11689);
nor U12064 (N_12064,N_11138,N_11483);
nand U12065 (N_12065,N_11620,N_11091);
or U12066 (N_12066,N_11764,N_11183);
xnor U12067 (N_12067,N_11522,N_11199);
and U12068 (N_12068,N_11238,N_11581);
and U12069 (N_12069,N_11314,N_11050);
and U12070 (N_12070,N_11072,N_11354);
and U12071 (N_12071,N_11447,N_11646);
or U12072 (N_12072,N_11069,N_11362);
xnor U12073 (N_12073,N_11014,N_11677);
and U12074 (N_12074,N_11968,N_11605);
or U12075 (N_12075,N_11149,N_11310);
and U12076 (N_12076,N_11070,N_11356);
or U12077 (N_12077,N_11435,N_11955);
or U12078 (N_12078,N_11441,N_11092);
nor U12079 (N_12079,N_11553,N_11110);
nand U12080 (N_12080,N_11970,N_11196);
nand U12081 (N_12081,N_11467,N_11711);
nor U12082 (N_12082,N_11963,N_11967);
and U12083 (N_12083,N_11656,N_11035);
nand U12084 (N_12084,N_11165,N_11340);
nand U12085 (N_12085,N_11657,N_11575);
or U12086 (N_12086,N_11473,N_11728);
nor U12087 (N_12087,N_11437,N_11376);
nand U12088 (N_12088,N_11566,N_11882);
or U12089 (N_12089,N_11515,N_11607);
or U12090 (N_12090,N_11837,N_11075);
nand U12091 (N_12091,N_11665,N_11564);
xnor U12092 (N_12092,N_11109,N_11008);
nand U12093 (N_12093,N_11962,N_11013);
and U12094 (N_12094,N_11081,N_11920);
nand U12095 (N_12095,N_11852,N_11667);
and U12096 (N_12096,N_11468,N_11182);
nand U12097 (N_12097,N_11120,N_11864);
xor U12098 (N_12098,N_11459,N_11442);
or U12099 (N_12099,N_11819,N_11048);
nor U12100 (N_12100,N_11993,N_11439);
and U12101 (N_12101,N_11732,N_11663);
and U12102 (N_12102,N_11843,N_11536);
xor U12103 (N_12103,N_11193,N_11785);
nand U12104 (N_12104,N_11794,N_11839);
nand U12105 (N_12105,N_11147,N_11272);
nor U12106 (N_12106,N_11042,N_11664);
nor U12107 (N_12107,N_11219,N_11233);
or U12108 (N_12108,N_11543,N_11604);
nor U12109 (N_12109,N_11719,N_11713);
xnor U12110 (N_12110,N_11260,N_11203);
and U12111 (N_12111,N_11132,N_11119);
or U12112 (N_12112,N_11561,N_11723);
or U12113 (N_12113,N_11884,N_11757);
nor U12114 (N_12114,N_11270,N_11565);
nor U12115 (N_12115,N_11402,N_11651);
xor U12116 (N_12116,N_11192,N_11103);
xor U12117 (N_12117,N_11379,N_11817);
or U12118 (N_12118,N_11005,N_11635);
nand U12119 (N_12119,N_11530,N_11710);
or U12120 (N_12120,N_11873,N_11313);
nand U12121 (N_12121,N_11389,N_11342);
or U12122 (N_12122,N_11734,N_11375);
or U12123 (N_12123,N_11403,N_11068);
nand U12124 (N_12124,N_11600,N_11134);
nor U12125 (N_12125,N_11430,N_11358);
xnor U12126 (N_12126,N_11912,N_11867);
nor U12127 (N_12127,N_11261,N_11888);
or U12128 (N_12128,N_11778,N_11639);
or U12129 (N_12129,N_11509,N_11391);
and U12130 (N_12130,N_11930,N_11318);
nand U12131 (N_12131,N_11045,N_11933);
and U12132 (N_12132,N_11792,N_11682);
xnor U12133 (N_12133,N_11084,N_11385);
and U12134 (N_12134,N_11077,N_11015);
nor U12135 (N_12135,N_11862,N_11804);
nor U12136 (N_12136,N_11230,N_11612);
or U12137 (N_12137,N_11498,N_11053);
or U12138 (N_12138,N_11531,N_11316);
or U12139 (N_12139,N_11184,N_11357);
xor U12140 (N_12140,N_11501,N_11104);
or U12141 (N_12141,N_11919,N_11984);
nand U12142 (N_12142,N_11025,N_11683);
nor U12143 (N_12143,N_11268,N_11129);
xor U12144 (N_12144,N_11809,N_11673);
and U12145 (N_12145,N_11088,N_11383);
or U12146 (N_12146,N_11999,N_11801);
nor U12147 (N_12147,N_11777,N_11252);
nor U12148 (N_12148,N_11298,N_11514);
and U12149 (N_12149,N_11692,N_11582);
and U12150 (N_12150,N_11246,N_11512);
nor U12151 (N_12151,N_11517,N_11440);
xor U12152 (N_12152,N_11629,N_11262);
or U12153 (N_12153,N_11480,N_11257);
and U12154 (N_12154,N_11649,N_11159);
or U12155 (N_12155,N_11162,N_11688);
or U12156 (N_12156,N_11779,N_11758);
nand U12157 (N_12157,N_11551,N_11197);
or U12158 (N_12158,N_11627,N_11825);
xnor U12159 (N_12159,N_11903,N_11908);
or U12160 (N_12160,N_11398,N_11000);
and U12161 (N_12161,N_11405,N_11766);
nand U12162 (N_12162,N_11305,N_11118);
or U12163 (N_12163,N_11917,N_11660);
and U12164 (N_12164,N_11731,N_11293);
or U12165 (N_12165,N_11321,N_11423);
xor U12166 (N_12166,N_11059,N_11227);
xor U12167 (N_12167,N_11065,N_11387);
nand U12168 (N_12168,N_11887,N_11889);
nor U12169 (N_12169,N_11063,N_11407);
or U12170 (N_12170,N_11408,N_11460);
xor U12171 (N_12171,N_11528,N_11943);
nand U12172 (N_12172,N_11796,N_11388);
nor U12173 (N_12173,N_11614,N_11854);
and U12174 (N_12174,N_11087,N_11940);
nand U12175 (N_12175,N_11726,N_11634);
xor U12176 (N_12176,N_11821,N_11122);
and U12177 (N_12177,N_11212,N_11832);
and U12178 (N_12178,N_11306,N_11499);
xnor U12179 (N_12179,N_11210,N_11031);
and U12180 (N_12180,N_11093,N_11608);
and U12181 (N_12181,N_11644,N_11214);
nor U12182 (N_12182,N_11168,N_11849);
or U12183 (N_12183,N_11469,N_11433);
xor U12184 (N_12184,N_11096,N_11964);
or U12185 (N_12185,N_11489,N_11411);
nor U12186 (N_12186,N_11679,N_11995);
and U12187 (N_12187,N_11948,N_11790);
nor U12188 (N_12188,N_11444,N_11263);
nor U12189 (N_12189,N_11906,N_11463);
nand U12190 (N_12190,N_11966,N_11187);
or U12191 (N_12191,N_11343,N_11108);
and U12192 (N_12192,N_11983,N_11365);
nand U12193 (N_12193,N_11676,N_11942);
nor U12194 (N_12194,N_11275,N_11658);
nand U12195 (N_12195,N_11350,N_11470);
xnor U12196 (N_12196,N_11894,N_11341);
and U12197 (N_12197,N_11339,N_11421);
nand U12198 (N_12198,N_11451,N_11002);
nand U12199 (N_12199,N_11519,N_11870);
or U12200 (N_12200,N_11768,N_11715);
nand U12201 (N_12201,N_11220,N_11934);
nor U12202 (N_12202,N_11351,N_11751);
or U12203 (N_12203,N_11532,N_11559);
nor U12204 (N_12204,N_11325,N_11895);
and U12205 (N_12205,N_11822,N_11164);
xnor U12206 (N_12206,N_11253,N_11204);
and U12207 (N_12207,N_11626,N_11924);
and U12208 (N_12208,N_11897,N_11127);
and U12209 (N_12209,N_11979,N_11753);
xnor U12210 (N_12210,N_11021,N_11240);
xor U12211 (N_12211,N_11793,N_11017);
nor U12212 (N_12212,N_11425,N_11041);
and U12213 (N_12213,N_11880,N_11178);
and U12214 (N_12214,N_11678,N_11638);
nand U12215 (N_12215,N_11874,N_11218);
or U12216 (N_12216,N_11180,N_11875);
nand U12217 (N_12217,N_11834,N_11382);
xnor U12218 (N_12218,N_11580,N_11959);
xnor U12219 (N_12219,N_11949,N_11207);
xnor U12220 (N_12220,N_11798,N_11429);
xor U12221 (N_12221,N_11586,N_11390);
nor U12222 (N_12222,N_11098,N_11139);
nor U12223 (N_12223,N_11012,N_11058);
xor U12224 (N_12224,N_11598,N_11630);
xnor U12225 (N_12225,N_11300,N_11513);
or U12226 (N_12226,N_11456,N_11789);
nor U12227 (N_12227,N_11386,N_11724);
and U12228 (N_12228,N_11795,N_11685);
and U12229 (N_12229,N_11280,N_11370);
nor U12230 (N_12230,N_11173,N_11327);
nor U12231 (N_12231,N_11893,N_11292);
nand U12232 (N_12232,N_11938,N_11787);
xor U12233 (N_12233,N_11289,N_11116);
xor U12234 (N_12234,N_11188,N_11428);
xor U12235 (N_12235,N_11556,N_11808);
xnor U12236 (N_12236,N_11538,N_11410);
nor U12237 (N_12237,N_11284,N_11746);
nand U12238 (N_12238,N_11918,N_11805);
or U12239 (N_12239,N_11953,N_11201);
xnor U12240 (N_12240,N_11992,N_11563);
or U12241 (N_12241,N_11117,N_11043);
xor U12242 (N_12242,N_11694,N_11571);
and U12243 (N_12243,N_11121,N_11475);
or U12244 (N_12244,N_11064,N_11181);
and U12245 (N_12245,N_11047,N_11668);
nor U12246 (N_12246,N_11511,N_11040);
nor U12247 (N_12247,N_11814,N_11401);
nor U12248 (N_12248,N_11765,N_11237);
and U12249 (N_12249,N_11800,N_11923);
nor U12250 (N_12250,N_11890,N_11523);
nand U12251 (N_12251,N_11247,N_11223);
and U12252 (N_12252,N_11037,N_11461);
and U12253 (N_12253,N_11902,N_11345);
xor U12254 (N_12254,N_11759,N_11823);
or U12255 (N_12255,N_11857,N_11816);
nor U12256 (N_12256,N_11319,N_11592);
and U12257 (N_12257,N_11935,N_11535);
xor U12258 (N_12258,N_11965,N_11546);
nand U12259 (N_12259,N_11969,N_11226);
or U12260 (N_12260,N_11085,N_11232);
nand U12261 (N_12261,N_11415,N_11806);
xnor U12262 (N_12262,N_11359,N_11335);
xor U12263 (N_12263,N_11741,N_11844);
or U12264 (N_12264,N_11898,N_11648);
or U12265 (N_12265,N_11020,N_11455);
nor U12266 (N_12266,N_11621,N_11258);
nor U12267 (N_12267,N_11245,N_11578);
xor U12268 (N_12268,N_11961,N_11328);
and U12269 (N_12269,N_11006,N_11799);
xor U12270 (N_12270,N_11975,N_11443);
nand U12271 (N_12271,N_11869,N_11144);
nor U12272 (N_12272,N_11113,N_11954);
or U12273 (N_12273,N_11073,N_11562);
nand U12274 (N_12274,N_11960,N_11169);
or U12275 (N_12275,N_11552,N_11703);
or U12276 (N_12276,N_11846,N_11775);
nor U12277 (N_12277,N_11739,N_11885);
nor U12278 (N_12278,N_11445,N_11010);
or U12279 (N_12279,N_11255,N_11427);
nor U12280 (N_12280,N_11004,N_11476);
and U12281 (N_12281,N_11631,N_11277);
nand U12282 (N_12282,N_11769,N_11772);
nor U12283 (N_12283,N_11802,N_11722);
or U12284 (N_12284,N_11097,N_11507);
nand U12285 (N_12285,N_11315,N_11185);
nand U12286 (N_12286,N_11672,N_11235);
xor U12287 (N_12287,N_11426,N_11454);
or U12288 (N_12288,N_11859,N_11055);
xnor U12289 (N_12289,N_11079,N_11881);
nor U12290 (N_12290,N_11770,N_11003);
nand U12291 (N_12291,N_11404,N_11827);
nor U12292 (N_12292,N_11718,N_11613);
xor U12293 (N_12293,N_11783,N_11071);
nand U12294 (N_12294,N_11866,N_11727);
xor U12295 (N_12295,N_11448,N_11901);
nor U12296 (N_12296,N_11242,N_11332);
and U12297 (N_12297,N_11001,N_11610);
nand U12298 (N_12298,N_11952,N_11251);
nor U12299 (N_12299,N_11140,N_11449);
and U12300 (N_12300,N_11491,N_11594);
and U12301 (N_12301,N_11926,N_11364);
nor U12302 (N_12302,N_11891,N_11419);
nor U12303 (N_12303,N_11583,N_11083);
xor U12304 (N_12304,N_11865,N_11555);
nand U12305 (N_12305,N_11299,N_11290);
and U12306 (N_12306,N_11348,N_11244);
xnor U12307 (N_12307,N_11393,N_11763);
or U12308 (N_12308,N_11011,N_11640);
and U12309 (N_12309,N_11811,N_11740);
and U12310 (N_12310,N_11266,N_11283);
nor U12311 (N_12311,N_11527,N_11215);
nand U12312 (N_12312,N_11494,N_11907);
xor U12313 (N_12313,N_11928,N_11100);
and U12314 (N_12314,N_11861,N_11756);
nand U12315 (N_12315,N_11076,N_11438);
or U12316 (N_12316,N_11484,N_11380);
or U12317 (N_12317,N_11932,N_11191);
nor U12318 (N_12318,N_11322,N_11981);
or U12319 (N_12319,N_11023,N_11372);
or U12320 (N_12320,N_11308,N_11324);
or U12321 (N_12321,N_11708,N_11274);
and U12322 (N_12322,N_11736,N_11972);
or U12323 (N_12323,N_11516,N_11154);
or U12324 (N_12324,N_11899,N_11684);
nor U12325 (N_12325,N_11107,N_11659);
or U12326 (N_12326,N_11208,N_11369);
xor U12327 (N_12327,N_11141,N_11161);
and U12328 (N_12328,N_11826,N_11256);
or U12329 (N_12329,N_11090,N_11986);
xor U12330 (N_12330,N_11782,N_11311);
and U12331 (N_12331,N_11510,N_11784);
xnor U12332 (N_12332,N_11137,N_11397);
nand U12333 (N_12333,N_11155,N_11520);
and U12334 (N_12334,N_11337,N_11286);
or U12335 (N_12335,N_11720,N_11755);
nand U12336 (N_12336,N_11569,N_11276);
or U12337 (N_12337,N_11269,N_11466);
and U12338 (N_12338,N_11450,N_11927);
or U12339 (N_12339,N_11095,N_11541);
nand U12340 (N_12340,N_11518,N_11591);
nor U12341 (N_12341,N_11525,N_11288);
xor U12342 (N_12342,N_11222,N_11016);
and U12343 (N_12343,N_11086,N_11845);
and U12344 (N_12344,N_11707,N_11641);
nand U12345 (N_12345,N_11396,N_11307);
or U12346 (N_12346,N_11971,N_11587);
and U12347 (N_12347,N_11317,N_11414);
and U12348 (N_12348,N_11590,N_11271);
xnor U12349 (N_12349,N_11371,N_11601);
or U12350 (N_12350,N_11497,N_11209);
and U12351 (N_12351,N_11241,N_11714);
or U12352 (N_12352,N_11504,N_11540);
nand U12353 (N_12353,N_11747,N_11599);
and U12354 (N_12354,N_11824,N_11297);
or U12355 (N_12355,N_11815,N_11544);
nand U12356 (N_12356,N_11654,N_11616);
or U12357 (N_12357,N_11304,N_11381);
xor U12358 (N_12358,N_11990,N_11287);
nand U12359 (N_12359,N_11330,N_11052);
and U12360 (N_12360,N_11754,N_11645);
and U12361 (N_12361,N_11774,N_11886);
nand U12362 (N_12362,N_11417,N_11236);
nor U12363 (N_12363,N_11211,N_11124);
nor U12364 (N_12364,N_11436,N_11056);
xor U12365 (N_12365,N_11039,N_11061);
or U12366 (N_12366,N_11344,N_11112);
xor U12367 (N_12367,N_11609,N_11911);
nand U12368 (N_12368,N_11702,N_11295);
xnor U12369 (N_12369,N_11950,N_11858);
or U12370 (N_12370,N_11550,N_11851);
xnor U12371 (N_12371,N_11265,N_11101);
xnor U12372 (N_12372,N_11279,N_11570);
nor U12373 (N_12373,N_11748,N_11737);
xor U12374 (N_12374,N_11745,N_11603);
nand U12375 (N_12375,N_11573,N_11549);
or U12376 (N_12376,N_11189,N_11847);
and U12377 (N_12377,N_11145,N_11878);
xnor U12378 (N_12378,N_11259,N_11547);
and U12379 (N_12379,N_11951,N_11394);
xnor U12380 (N_12380,N_11416,N_11030);
nor U12381 (N_12381,N_11464,N_11472);
or U12382 (N_12382,N_11152,N_11326);
or U12383 (N_12383,N_11067,N_11632);
or U12384 (N_12384,N_11980,N_11697);
and U12385 (N_12385,N_11166,N_11944);
and U12386 (N_12386,N_11361,N_11490);
or U12387 (N_12387,N_11213,N_11833);
nand U12388 (N_12388,N_11704,N_11243);
nor U12389 (N_12389,N_11914,N_11596);
xnor U12390 (N_12390,N_11123,N_11977);
nand U12391 (N_12391,N_11301,N_11593);
or U12392 (N_12392,N_11099,N_11773);
and U12393 (N_12393,N_11666,N_11588);
nand U12394 (N_12394,N_11111,N_11309);
and U12395 (N_12395,N_11760,N_11133);
xnor U12396 (N_12396,N_11431,N_11721);
nand U12397 (N_12397,N_11221,N_11333);
and U12398 (N_12398,N_11749,N_11693);
nor U12399 (N_12399,N_11346,N_11655);
nor U12400 (N_12400,N_11628,N_11670);
nor U12401 (N_12401,N_11791,N_11032);
nor U12402 (N_12402,N_11500,N_11633);
and U12403 (N_12403,N_11892,N_11661);
nand U12404 (N_12404,N_11643,N_11399);
xnor U12405 (N_12405,N_11249,N_11368);
or U12406 (N_12406,N_11653,N_11636);
or U12407 (N_12407,N_11615,N_11496);
or U12408 (N_12408,N_11172,N_11717);
and U12409 (N_12409,N_11413,N_11577);
nand U12410 (N_12410,N_11925,N_11997);
xor U12411 (N_12411,N_11611,N_11687);
nand U12412 (N_12412,N_11323,N_11373);
or U12413 (N_12413,N_11409,N_11151);
nand U12414 (N_12414,N_11681,N_11148);
and U12415 (N_12415,N_11457,N_11202);
xnor U12416 (N_12416,N_11146,N_11482);
nor U12417 (N_12417,N_11872,N_11126);
xnor U12418 (N_12418,N_11877,N_11524);
nand U12419 (N_12419,N_11725,N_11036);
xor U12420 (N_12420,N_11198,N_11114);
nor U12421 (N_12421,N_11019,N_11856);
xnor U12422 (N_12422,N_11595,N_11941);
xnor U12423 (N_12423,N_11998,N_11026);
or U12424 (N_12424,N_11840,N_11495);
xor U12425 (N_12425,N_11973,N_11248);
or U12426 (N_12426,N_11982,N_11828);
and U12427 (N_12427,N_11131,N_11618);
xnor U12428 (N_12428,N_11989,N_11675);
and U12429 (N_12429,N_11909,N_11853);
xor U12430 (N_12430,N_11125,N_11698);
xnor U12431 (N_12431,N_11089,N_11128);
and U12432 (N_12432,N_11462,N_11028);
and U12433 (N_12433,N_11195,N_11788);
nor U12434 (N_12434,N_11771,N_11743);
or U12435 (N_12435,N_11395,N_11686);
xor U12436 (N_12436,N_11352,N_11579);
or U12437 (N_12437,N_11810,N_11009);
or U12438 (N_12438,N_11066,N_11850);
and U12439 (N_12439,N_11054,N_11225);
and U12440 (N_12440,N_11730,N_11508);
and U12441 (N_12441,N_11637,N_11366);
or U12442 (N_12442,N_11994,N_11762);
xnor U12443 (N_12443,N_11285,N_11879);
xnor U12444 (N_12444,N_11320,N_11820);
and U12445 (N_12445,N_11156,N_11916);
or U12446 (N_12446,N_11690,N_11331);
xor U12447 (N_12447,N_11135,N_11830);
nand U12448 (N_12448,N_11696,N_11896);
or U12449 (N_12449,N_11742,N_11250);
or U12450 (N_12450,N_11662,N_11617);
or U12451 (N_12451,N_11194,N_11190);
and U12452 (N_12452,N_11913,N_11841);
and U12453 (N_12453,N_11158,N_11534);
nor U12454 (N_12454,N_11143,N_11625);
nand U12455 (N_12455,N_11558,N_11105);
xor U12456 (N_12456,N_11985,N_11175);
or U12457 (N_12457,N_11652,N_11400);
xor U12458 (N_12458,N_11922,N_11905);
or U12459 (N_12459,N_11987,N_11446);
nand U12460 (N_12460,N_11336,N_11022);
or U12461 (N_12461,N_11157,N_11412);
or U12462 (N_12462,N_11231,N_11699);
or U12463 (N_12463,N_11281,N_11786);
and U12464 (N_12464,N_11750,N_11624);
nand U12465 (N_12465,N_11584,N_11589);
nand U12466 (N_12466,N_11273,N_11367);
or U12467 (N_12467,N_11871,N_11163);
xnor U12468 (N_12468,N_11557,N_11303);
xnor U12469 (N_12469,N_11709,N_11329);
nand U12470 (N_12470,N_11761,N_11034);
nor U12471 (N_12471,N_11900,N_11406);
nand U12472 (N_12472,N_11602,N_11910);
xor U12473 (N_12473,N_11936,N_11619);
nand U12474 (N_12474,N_11572,N_11585);
nor U12475 (N_12475,N_11349,N_11921);
and U12476 (N_12476,N_11868,N_11216);
xor U12477 (N_12477,N_11142,N_11650);
nor U12478 (N_12478,N_11486,N_11174);
or U12479 (N_12479,N_11767,N_11674);
nor U12480 (N_12480,N_11560,N_11234);
nor U12481 (N_12481,N_11106,N_11946);
and U12482 (N_12482,N_11492,N_11378);
and U12483 (N_12483,N_11487,N_11957);
and U12484 (N_12484,N_11642,N_11217);
nand U12485 (N_12485,N_11863,N_11477);
and U12486 (N_12486,N_11177,N_11829);
or U12487 (N_12487,N_11545,N_11505);
or U12488 (N_12488,N_11729,N_11542);
nor U12489 (N_12489,N_11465,N_11179);
xor U12490 (N_12490,N_11502,N_11597);
or U12491 (N_12491,N_11038,N_11080);
nand U12492 (N_12492,N_11078,N_11471);
nor U12493 (N_12493,N_11049,N_11712);
and U12494 (N_12494,N_11478,N_11733);
nor U12495 (N_12495,N_11606,N_11474);
xnor U12496 (N_12496,N_11716,N_11264);
nor U12497 (N_12497,N_11170,N_11781);
nand U12498 (N_12498,N_11338,N_11296);
nor U12499 (N_12499,N_11334,N_11931);
and U12500 (N_12500,N_11225,N_11299);
and U12501 (N_12501,N_11316,N_11878);
or U12502 (N_12502,N_11856,N_11451);
xor U12503 (N_12503,N_11576,N_11789);
xor U12504 (N_12504,N_11210,N_11770);
xnor U12505 (N_12505,N_11318,N_11372);
and U12506 (N_12506,N_11332,N_11627);
or U12507 (N_12507,N_11613,N_11735);
nand U12508 (N_12508,N_11711,N_11397);
xor U12509 (N_12509,N_11554,N_11887);
nand U12510 (N_12510,N_11791,N_11839);
nand U12511 (N_12511,N_11373,N_11079);
or U12512 (N_12512,N_11824,N_11594);
or U12513 (N_12513,N_11237,N_11755);
or U12514 (N_12514,N_11329,N_11679);
xor U12515 (N_12515,N_11398,N_11324);
nand U12516 (N_12516,N_11494,N_11790);
nor U12517 (N_12517,N_11561,N_11936);
nor U12518 (N_12518,N_11957,N_11712);
nand U12519 (N_12519,N_11460,N_11900);
xnor U12520 (N_12520,N_11614,N_11645);
nor U12521 (N_12521,N_11791,N_11842);
or U12522 (N_12522,N_11718,N_11156);
or U12523 (N_12523,N_11942,N_11080);
nand U12524 (N_12524,N_11201,N_11317);
nand U12525 (N_12525,N_11599,N_11904);
or U12526 (N_12526,N_11599,N_11134);
nor U12527 (N_12527,N_11066,N_11860);
or U12528 (N_12528,N_11908,N_11227);
and U12529 (N_12529,N_11969,N_11669);
xnor U12530 (N_12530,N_11349,N_11380);
xnor U12531 (N_12531,N_11986,N_11012);
and U12532 (N_12532,N_11876,N_11047);
or U12533 (N_12533,N_11033,N_11286);
nand U12534 (N_12534,N_11144,N_11841);
xor U12535 (N_12535,N_11174,N_11619);
or U12536 (N_12536,N_11349,N_11785);
nand U12537 (N_12537,N_11618,N_11916);
xor U12538 (N_12538,N_11564,N_11861);
or U12539 (N_12539,N_11298,N_11262);
nor U12540 (N_12540,N_11371,N_11925);
and U12541 (N_12541,N_11397,N_11550);
or U12542 (N_12542,N_11146,N_11827);
or U12543 (N_12543,N_11440,N_11388);
or U12544 (N_12544,N_11428,N_11443);
nor U12545 (N_12545,N_11239,N_11486);
or U12546 (N_12546,N_11915,N_11732);
xor U12547 (N_12547,N_11543,N_11157);
nand U12548 (N_12548,N_11789,N_11203);
and U12549 (N_12549,N_11422,N_11229);
and U12550 (N_12550,N_11435,N_11379);
and U12551 (N_12551,N_11876,N_11605);
xor U12552 (N_12552,N_11881,N_11544);
or U12553 (N_12553,N_11121,N_11542);
nor U12554 (N_12554,N_11740,N_11502);
nand U12555 (N_12555,N_11347,N_11995);
xnor U12556 (N_12556,N_11099,N_11012);
nor U12557 (N_12557,N_11573,N_11991);
nor U12558 (N_12558,N_11682,N_11170);
and U12559 (N_12559,N_11267,N_11620);
or U12560 (N_12560,N_11047,N_11242);
nor U12561 (N_12561,N_11951,N_11644);
or U12562 (N_12562,N_11919,N_11834);
xor U12563 (N_12563,N_11025,N_11978);
or U12564 (N_12564,N_11064,N_11818);
and U12565 (N_12565,N_11893,N_11641);
or U12566 (N_12566,N_11567,N_11366);
nand U12567 (N_12567,N_11657,N_11209);
xnor U12568 (N_12568,N_11870,N_11020);
nand U12569 (N_12569,N_11717,N_11493);
xnor U12570 (N_12570,N_11273,N_11666);
and U12571 (N_12571,N_11339,N_11490);
and U12572 (N_12572,N_11355,N_11071);
nor U12573 (N_12573,N_11279,N_11692);
and U12574 (N_12574,N_11970,N_11264);
nand U12575 (N_12575,N_11007,N_11632);
nand U12576 (N_12576,N_11282,N_11544);
nand U12577 (N_12577,N_11479,N_11395);
or U12578 (N_12578,N_11010,N_11634);
xnor U12579 (N_12579,N_11673,N_11791);
and U12580 (N_12580,N_11507,N_11878);
xor U12581 (N_12581,N_11421,N_11017);
xor U12582 (N_12582,N_11834,N_11650);
nor U12583 (N_12583,N_11934,N_11289);
and U12584 (N_12584,N_11817,N_11540);
xnor U12585 (N_12585,N_11690,N_11111);
nand U12586 (N_12586,N_11181,N_11711);
nand U12587 (N_12587,N_11307,N_11854);
xor U12588 (N_12588,N_11382,N_11072);
or U12589 (N_12589,N_11340,N_11401);
or U12590 (N_12590,N_11490,N_11461);
or U12591 (N_12591,N_11483,N_11160);
nor U12592 (N_12592,N_11556,N_11043);
or U12593 (N_12593,N_11278,N_11415);
and U12594 (N_12594,N_11360,N_11935);
or U12595 (N_12595,N_11063,N_11315);
or U12596 (N_12596,N_11233,N_11781);
or U12597 (N_12597,N_11518,N_11617);
xor U12598 (N_12598,N_11816,N_11404);
or U12599 (N_12599,N_11926,N_11307);
or U12600 (N_12600,N_11902,N_11523);
nand U12601 (N_12601,N_11558,N_11170);
nand U12602 (N_12602,N_11382,N_11792);
nor U12603 (N_12603,N_11188,N_11950);
and U12604 (N_12604,N_11037,N_11976);
or U12605 (N_12605,N_11408,N_11702);
nor U12606 (N_12606,N_11041,N_11889);
nor U12607 (N_12607,N_11060,N_11369);
and U12608 (N_12608,N_11235,N_11540);
nor U12609 (N_12609,N_11945,N_11295);
and U12610 (N_12610,N_11965,N_11405);
or U12611 (N_12611,N_11271,N_11959);
xor U12612 (N_12612,N_11983,N_11308);
or U12613 (N_12613,N_11276,N_11986);
nand U12614 (N_12614,N_11160,N_11647);
nand U12615 (N_12615,N_11580,N_11573);
xnor U12616 (N_12616,N_11832,N_11284);
and U12617 (N_12617,N_11248,N_11303);
or U12618 (N_12618,N_11959,N_11485);
and U12619 (N_12619,N_11675,N_11425);
nor U12620 (N_12620,N_11415,N_11121);
xor U12621 (N_12621,N_11493,N_11687);
nor U12622 (N_12622,N_11367,N_11445);
xor U12623 (N_12623,N_11457,N_11034);
and U12624 (N_12624,N_11205,N_11964);
xnor U12625 (N_12625,N_11177,N_11037);
or U12626 (N_12626,N_11132,N_11959);
nor U12627 (N_12627,N_11695,N_11084);
and U12628 (N_12628,N_11856,N_11414);
or U12629 (N_12629,N_11858,N_11937);
and U12630 (N_12630,N_11278,N_11343);
nor U12631 (N_12631,N_11303,N_11541);
nor U12632 (N_12632,N_11719,N_11004);
and U12633 (N_12633,N_11964,N_11659);
nand U12634 (N_12634,N_11183,N_11051);
xnor U12635 (N_12635,N_11414,N_11688);
nand U12636 (N_12636,N_11467,N_11071);
nand U12637 (N_12637,N_11631,N_11357);
nand U12638 (N_12638,N_11180,N_11339);
and U12639 (N_12639,N_11500,N_11048);
and U12640 (N_12640,N_11166,N_11782);
and U12641 (N_12641,N_11476,N_11371);
and U12642 (N_12642,N_11441,N_11410);
or U12643 (N_12643,N_11112,N_11852);
nor U12644 (N_12644,N_11617,N_11542);
xor U12645 (N_12645,N_11197,N_11392);
xnor U12646 (N_12646,N_11844,N_11808);
nand U12647 (N_12647,N_11990,N_11555);
and U12648 (N_12648,N_11874,N_11684);
and U12649 (N_12649,N_11707,N_11683);
xor U12650 (N_12650,N_11013,N_11448);
or U12651 (N_12651,N_11783,N_11806);
and U12652 (N_12652,N_11877,N_11779);
xnor U12653 (N_12653,N_11279,N_11632);
and U12654 (N_12654,N_11512,N_11152);
xnor U12655 (N_12655,N_11067,N_11964);
xor U12656 (N_12656,N_11765,N_11083);
or U12657 (N_12657,N_11456,N_11734);
nand U12658 (N_12658,N_11263,N_11971);
or U12659 (N_12659,N_11884,N_11877);
nand U12660 (N_12660,N_11784,N_11464);
or U12661 (N_12661,N_11607,N_11680);
nor U12662 (N_12662,N_11937,N_11318);
xor U12663 (N_12663,N_11669,N_11409);
nand U12664 (N_12664,N_11525,N_11217);
nor U12665 (N_12665,N_11671,N_11474);
or U12666 (N_12666,N_11278,N_11962);
nor U12667 (N_12667,N_11529,N_11514);
nor U12668 (N_12668,N_11914,N_11699);
nor U12669 (N_12669,N_11514,N_11453);
nand U12670 (N_12670,N_11123,N_11196);
xor U12671 (N_12671,N_11531,N_11318);
and U12672 (N_12672,N_11183,N_11874);
nand U12673 (N_12673,N_11257,N_11886);
nor U12674 (N_12674,N_11356,N_11629);
xor U12675 (N_12675,N_11803,N_11044);
and U12676 (N_12676,N_11070,N_11863);
nand U12677 (N_12677,N_11884,N_11576);
nor U12678 (N_12678,N_11882,N_11775);
and U12679 (N_12679,N_11423,N_11052);
xnor U12680 (N_12680,N_11627,N_11454);
or U12681 (N_12681,N_11640,N_11580);
nor U12682 (N_12682,N_11757,N_11674);
and U12683 (N_12683,N_11475,N_11626);
nor U12684 (N_12684,N_11486,N_11702);
and U12685 (N_12685,N_11977,N_11568);
xor U12686 (N_12686,N_11408,N_11741);
nand U12687 (N_12687,N_11894,N_11513);
or U12688 (N_12688,N_11000,N_11809);
nand U12689 (N_12689,N_11532,N_11979);
or U12690 (N_12690,N_11146,N_11483);
xnor U12691 (N_12691,N_11242,N_11384);
xor U12692 (N_12692,N_11024,N_11407);
xnor U12693 (N_12693,N_11281,N_11873);
nor U12694 (N_12694,N_11013,N_11922);
nand U12695 (N_12695,N_11646,N_11093);
and U12696 (N_12696,N_11136,N_11517);
nand U12697 (N_12697,N_11526,N_11075);
or U12698 (N_12698,N_11511,N_11508);
nor U12699 (N_12699,N_11904,N_11298);
nor U12700 (N_12700,N_11035,N_11659);
and U12701 (N_12701,N_11589,N_11172);
nand U12702 (N_12702,N_11026,N_11482);
nor U12703 (N_12703,N_11256,N_11773);
and U12704 (N_12704,N_11916,N_11370);
and U12705 (N_12705,N_11995,N_11463);
xor U12706 (N_12706,N_11381,N_11376);
or U12707 (N_12707,N_11941,N_11303);
nand U12708 (N_12708,N_11526,N_11783);
nand U12709 (N_12709,N_11291,N_11780);
nand U12710 (N_12710,N_11952,N_11993);
and U12711 (N_12711,N_11483,N_11637);
xor U12712 (N_12712,N_11453,N_11794);
nand U12713 (N_12713,N_11432,N_11868);
nor U12714 (N_12714,N_11703,N_11586);
nand U12715 (N_12715,N_11091,N_11496);
or U12716 (N_12716,N_11149,N_11973);
and U12717 (N_12717,N_11142,N_11740);
nor U12718 (N_12718,N_11648,N_11480);
nand U12719 (N_12719,N_11832,N_11778);
nor U12720 (N_12720,N_11255,N_11494);
xnor U12721 (N_12721,N_11162,N_11505);
xnor U12722 (N_12722,N_11461,N_11992);
nand U12723 (N_12723,N_11710,N_11897);
nor U12724 (N_12724,N_11348,N_11453);
or U12725 (N_12725,N_11125,N_11427);
nor U12726 (N_12726,N_11092,N_11889);
or U12727 (N_12727,N_11406,N_11462);
nand U12728 (N_12728,N_11353,N_11827);
xor U12729 (N_12729,N_11175,N_11840);
nand U12730 (N_12730,N_11794,N_11856);
xor U12731 (N_12731,N_11406,N_11452);
nor U12732 (N_12732,N_11507,N_11094);
nand U12733 (N_12733,N_11022,N_11289);
and U12734 (N_12734,N_11935,N_11323);
nor U12735 (N_12735,N_11595,N_11112);
xor U12736 (N_12736,N_11619,N_11829);
nand U12737 (N_12737,N_11552,N_11204);
nor U12738 (N_12738,N_11560,N_11714);
nand U12739 (N_12739,N_11019,N_11490);
nand U12740 (N_12740,N_11636,N_11735);
nor U12741 (N_12741,N_11544,N_11089);
nor U12742 (N_12742,N_11785,N_11825);
and U12743 (N_12743,N_11745,N_11242);
nor U12744 (N_12744,N_11397,N_11147);
xor U12745 (N_12745,N_11938,N_11198);
xor U12746 (N_12746,N_11355,N_11131);
nand U12747 (N_12747,N_11160,N_11947);
xor U12748 (N_12748,N_11719,N_11876);
or U12749 (N_12749,N_11810,N_11360);
or U12750 (N_12750,N_11459,N_11193);
nor U12751 (N_12751,N_11636,N_11674);
xor U12752 (N_12752,N_11532,N_11701);
nand U12753 (N_12753,N_11499,N_11256);
nor U12754 (N_12754,N_11361,N_11286);
and U12755 (N_12755,N_11574,N_11945);
nand U12756 (N_12756,N_11764,N_11775);
nand U12757 (N_12757,N_11124,N_11950);
nand U12758 (N_12758,N_11734,N_11276);
nand U12759 (N_12759,N_11567,N_11909);
nand U12760 (N_12760,N_11081,N_11163);
xor U12761 (N_12761,N_11861,N_11316);
or U12762 (N_12762,N_11709,N_11102);
or U12763 (N_12763,N_11928,N_11596);
or U12764 (N_12764,N_11018,N_11433);
or U12765 (N_12765,N_11015,N_11293);
nand U12766 (N_12766,N_11192,N_11273);
and U12767 (N_12767,N_11773,N_11619);
nand U12768 (N_12768,N_11194,N_11892);
or U12769 (N_12769,N_11245,N_11353);
and U12770 (N_12770,N_11554,N_11009);
or U12771 (N_12771,N_11956,N_11162);
and U12772 (N_12772,N_11243,N_11188);
and U12773 (N_12773,N_11661,N_11440);
nand U12774 (N_12774,N_11958,N_11780);
and U12775 (N_12775,N_11693,N_11759);
nand U12776 (N_12776,N_11641,N_11768);
nand U12777 (N_12777,N_11436,N_11420);
xor U12778 (N_12778,N_11500,N_11497);
xor U12779 (N_12779,N_11068,N_11776);
xor U12780 (N_12780,N_11274,N_11452);
and U12781 (N_12781,N_11909,N_11049);
nor U12782 (N_12782,N_11171,N_11828);
xor U12783 (N_12783,N_11165,N_11666);
and U12784 (N_12784,N_11451,N_11602);
xor U12785 (N_12785,N_11429,N_11591);
nor U12786 (N_12786,N_11643,N_11937);
and U12787 (N_12787,N_11683,N_11211);
or U12788 (N_12788,N_11452,N_11034);
nand U12789 (N_12789,N_11001,N_11475);
nor U12790 (N_12790,N_11563,N_11684);
xnor U12791 (N_12791,N_11655,N_11372);
xor U12792 (N_12792,N_11843,N_11997);
and U12793 (N_12793,N_11025,N_11024);
or U12794 (N_12794,N_11009,N_11311);
nand U12795 (N_12795,N_11782,N_11145);
nor U12796 (N_12796,N_11583,N_11299);
and U12797 (N_12797,N_11970,N_11347);
nand U12798 (N_12798,N_11570,N_11021);
nor U12799 (N_12799,N_11931,N_11488);
nand U12800 (N_12800,N_11010,N_11829);
or U12801 (N_12801,N_11254,N_11028);
nor U12802 (N_12802,N_11961,N_11957);
and U12803 (N_12803,N_11927,N_11127);
xor U12804 (N_12804,N_11120,N_11809);
xor U12805 (N_12805,N_11035,N_11498);
xnor U12806 (N_12806,N_11367,N_11682);
or U12807 (N_12807,N_11102,N_11184);
nor U12808 (N_12808,N_11745,N_11991);
or U12809 (N_12809,N_11503,N_11447);
or U12810 (N_12810,N_11617,N_11013);
and U12811 (N_12811,N_11261,N_11153);
and U12812 (N_12812,N_11832,N_11251);
nand U12813 (N_12813,N_11136,N_11409);
or U12814 (N_12814,N_11168,N_11654);
or U12815 (N_12815,N_11347,N_11826);
nor U12816 (N_12816,N_11104,N_11283);
and U12817 (N_12817,N_11523,N_11055);
and U12818 (N_12818,N_11389,N_11504);
and U12819 (N_12819,N_11272,N_11028);
or U12820 (N_12820,N_11137,N_11754);
nand U12821 (N_12821,N_11487,N_11543);
nor U12822 (N_12822,N_11736,N_11502);
nand U12823 (N_12823,N_11070,N_11969);
nor U12824 (N_12824,N_11580,N_11577);
or U12825 (N_12825,N_11957,N_11371);
xor U12826 (N_12826,N_11084,N_11703);
xor U12827 (N_12827,N_11061,N_11955);
nand U12828 (N_12828,N_11096,N_11329);
xnor U12829 (N_12829,N_11452,N_11626);
nor U12830 (N_12830,N_11780,N_11971);
xor U12831 (N_12831,N_11624,N_11274);
nor U12832 (N_12832,N_11196,N_11392);
or U12833 (N_12833,N_11017,N_11132);
xor U12834 (N_12834,N_11449,N_11874);
or U12835 (N_12835,N_11389,N_11889);
nand U12836 (N_12836,N_11371,N_11197);
nor U12837 (N_12837,N_11395,N_11361);
nand U12838 (N_12838,N_11279,N_11731);
or U12839 (N_12839,N_11261,N_11838);
xnor U12840 (N_12840,N_11312,N_11502);
nand U12841 (N_12841,N_11452,N_11615);
and U12842 (N_12842,N_11028,N_11269);
xnor U12843 (N_12843,N_11623,N_11164);
nand U12844 (N_12844,N_11130,N_11111);
and U12845 (N_12845,N_11848,N_11812);
and U12846 (N_12846,N_11814,N_11943);
and U12847 (N_12847,N_11058,N_11796);
nand U12848 (N_12848,N_11724,N_11960);
or U12849 (N_12849,N_11678,N_11701);
nand U12850 (N_12850,N_11863,N_11199);
nor U12851 (N_12851,N_11979,N_11529);
nand U12852 (N_12852,N_11681,N_11868);
xnor U12853 (N_12853,N_11386,N_11030);
xnor U12854 (N_12854,N_11457,N_11912);
nor U12855 (N_12855,N_11260,N_11966);
nand U12856 (N_12856,N_11254,N_11718);
nor U12857 (N_12857,N_11645,N_11652);
or U12858 (N_12858,N_11725,N_11069);
xor U12859 (N_12859,N_11961,N_11691);
or U12860 (N_12860,N_11485,N_11081);
nand U12861 (N_12861,N_11656,N_11451);
nand U12862 (N_12862,N_11787,N_11306);
or U12863 (N_12863,N_11323,N_11857);
nor U12864 (N_12864,N_11001,N_11878);
nand U12865 (N_12865,N_11627,N_11235);
nor U12866 (N_12866,N_11175,N_11749);
nand U12867 (N_12867,N_11535,N_11427);
xor U12868 (N_12868,N_11306,N_11657);
and U12869 (N_12869,N_11397,N_11476);
nand U12870 (N_12870,N_11931,N_11695);
xor U12871 (N_12871,N_11222,N_11499);
and U12872 (N_12872,N_11856,N_11611);
nand U12873 (N_12873,N_11336,N_11240);
and U12874 (N_12874,N_11869,N_11274);
nor U12875 (N_12875,N_11490,N_11392);
and U12876 (N_12876,N_11612,N_11725);
or U12877 (N_12877,N_11123,N_11221);
nor U12878 (N_12878,N_11993,N_11346);
xnor U12879 (N_12879,N_11468,N_11434);
nand U12880 (N_12880,N_11372,N_11219);
and U12881 (N_12881,N_11916,N_11476);
nand U12882 (N_12882,N_11272,N_11165);
and U12883 (N_12883,N_11111,N_11497);
and U12884 (N_12884,N_11365,N_11635);
and U12885 (N_12885,N_11158,N_11223);
and U12886 (N_12886,N_11063,N_11314);
nand U12887 (N_12887,N_11717,N_11610);
nand U12888 (N_12888,N_11022,N_11080);
xnor U12889 (N_12889,N_11259,N_11898);
and U12890 (N_12890,N_11641,N_11200);
nor U12891 (N_12891,N_11536,N_11271);
or U12892 (N_12892,N_11423,N_11883);
or U12893 (N_12893,N_11108,N_11716);
and U12894 (N_12894,N_11887,N_11219);
nand U12895 (N_12895,N_11878,N_11045);
nand U12896 (N_12896,N_11101,N_11880);
xor U12897 (N_12897,N_11947,N_11810);
and U12898 (N_12898,N_11170,N_11510);
nor U12899 (N_12899,N_11575,N_11151);
xor U12900 (N_12900,N_11411,N_11483);
and U12901 (N_12901,N_11566,N_11890);
or U12902 (N_12902,N_11521,N_11709);
xnor U12903 (N_12903,N_11151,N_11884);
and U12904 (N_12904,N_11427,N_11598);
xor U12905 (N_12905,N_11780,N_11220);
or U12906 (N_12906,N_11010,N_11574);
nand U12907 (N_12907,N_11445,N_11562);
and U12908 (N_12908,N_11748,N_11272);
and U12909 (N_12909,N_11392,N_11122);
and U12910 (N_12910,N_11975,N_11070);
xor U12911 (N_12911,N_11855,N_11209);
xor U12912 (N_12912,N_11962,N_11829);
nand U12913 (N_12913,N_11882,N_11273);
nand U12914 (N_12914,N_11187,N_11168);
and U12915 (N_12915,N_11561,N_11624);
and U12916 (N_12916,N_11408,N_11961);
nand U12917 (N_12917,N_11744,N_11313);
and U12918 (N_12918,N_11935,N_11491);
nor U12919 (N_12919,N_11881,N_11386);
nand U12920 (N_12920,N_11087,N_11002);
nor U12921 (N_12921,N_11752,N_11722);
nand U12922 (N_12922,N_11528,N_11979);
nand U12923 (N_12923,N_11374,N_11056);
nor U12924 (N_12924,N_11494,N_11101);
nor U12925 (N_12925,N_11469,N_11397);
nand U12926 (N_12926,N_11314,N_11392);
nor U12927 (N_12927,N_11312,N_11616);
or U12928 (N_12928,N_11802,N_11520);
xnor U12929 (N_12929,N_11635,N_11326);
nand U12930 (N_12930,N_11385,N_11874);
and U12931 (N_12931,N_11989,N_11521);
or U12932 (N_12932,N_11492,N_11386);
and U12933 (N_12933,N_11519,N_11308);
or U12934 (N_12934,N_11576,N_11235);
and U12935 (N_12935,N_11265,N_11293);
nand U12936 (N_12936,N_11026,N_11332);
nand U12937 (N_12937,N_11596,N_11397);
nand U12938 (N_12938,N_11121,N_11336);
nand U12939 (N_12939,N_11511,N_11284);
and U12940 (N_12940,N_11073,N_11257);
nor U12941 (N_12941,N_11721,N_11711);
or U12942 (N_12942,N_11888,N_11402);
xor U12943 (N_12943,N_11576,N_11269);
or U12944 (N_12944,N_11346,N_11986);
or U12945 (N_12945,N_11391,N_11082);
nand U12946 (N_12946,N_11326,N_11485);
xor U12947 (N_12947,N_11385,N_11575);
and U12948 (N_12948,N_11850,N_11103);
nor U12949 (N_12949,N_11256,N_11093);
nand U12950 (N_12950,N_11768,N_11400);
xor U12951 (N_12951,N_11050,N_11853);
nor U12952 (N_12952,N_11474,N_11732);
nor U12953 (N_12953,N_11560,N_11067);
or U12954 (N_12954,N_11105,N_11217);
and U12955 (N_12955,N_11762,N_11342);
and U12956 (N_12956,N_11420,N_11341);
nand U12957 (N_12957,N_11628,N_11814);
xnor U12958 (N_12958,N_11400,N_11018);
xnor U12959 (N_12959,N_11463,N_11886);
or U12960 (N_12960,N_11720,N_11901);
nor U12961 (N_12961,N_11193,N_11701);
nand U12962 (N_12962,N_11785,N_11750);
xnor U12963 (N_12963,N_11532,N_11356);
and U12964 (N_12964,N_11987,N_11125);
xor U12965 (N_12965,N_11974,N_11417);
nor U12966 (N_12966,N_11934,N_11277);
xnor U12967 (N_12967,N_11174,N_11686);
xor U12968 (N_12968,N_11678,N_11104);
xor U12969 (N_12969,N_11716,N_11926);
or U12970 (N_12970,N_11826,N_11841);
and U12971 (N_12971,N_11609,N_11233);
or U12972 (N_12972,N_11588,N_11824);
and U12973 (N_12973,N_11813,N_11553);
and U12974 (N_12974,N_11848,N_11788);
xnor U12975 (N_12975,N_11254,N_11085);
nor U12976 (N_12976,N_11957,N_11697);
nand U12977 (N_12977,N_11813,N_11550);
nor U12978 (N_12978,N_11742,N_11613);
and U12979 (N_12979,N_11496,N_11257);
nor U12980 (N_12980,N_11827,N_11389);
and U12981 (N_12981,N_11727,N_11966);
nor U12982 (N_12982,N_11995,N_11606);
nand U12983 (N_12983,N_11377,N_11049);
or U12984 (N_12984,N_11571,N_11163);
nor U12985 (N_12985,N_11941,N_11590);
or U12986 (N_12986,N_11514,N_11124);
xnor U12987 (N_12987,N_11820,N_11805);
nand U12988 (N_12988,N_11463,N_11324);
nand U12989 (N_12989,N_11007,N_11119);
nand U12990 (N_12990,N_11572,N_11794);
nand U12991 (N_12991,N_11968,N_11104);
xnor U12992 (N_12992,N_11199,N_11347);
nand U12993 (N_12993,N_11879,N_11544);
and U12994 (N_12994,N_11851,N_11890);
nand U12995 (N_12995,N_11113,N_11999);
or U12996 (N_12996,N_11707,N_11467);
and U12997 (N_12997,N_11282,N_11149);
xnor U12998 (N_12998,N_11326,N_11610);
xnor U12999 (N_12999,N_11469,N_11773);
and U13000 (N_13000,N_12700,N_12372);
or U13001 (N_13001,N_12616,N_12104);
nand U13002 (N_13002,N_12362,N_12980);
nand U13003 (N_13003,N_12872,N_12525);
or U13004 (N_13004,N_12510,N_12472);
nor U13005 (N_13005,N_12086,N_12975);
and U13006 (N_13006,N_12971,N_12060);
or U13007 (N_13007,N_12192,N_12860);
and U13008 (N_13008,N_12325,N_12940);
xnor U13009 (N_13009,N_12549,N_12809);
and U13010 (N_13010,N_12215,N_12571);
or U13011 (N_13011,N_12850,N_12076);
and U13012 (N_13012,N_12339,N_12529);
and U13013 (N_13013,N_12686,N_12461);
and U13014 (N_13014,N_12012,N_12394);
or U13015 (N_13015,N_12098,N_12369);
and U13016 (N_13016,N_12122,N_12693);
and U13017 (N_13017,N_12828,N_12918);
nand U13018 (N_13018,N_12143,N_12785);
and U13019 (N_13019,N_12226,N_12958);
xor U13020 (N_13020,N_12757,N_12795);
and U13021 (N_13021,N_12044,N_12799);
nand U13022 (N_13022,N_12987,N_12405);
or U13023 (N_13023,N_12560,N_12422);
and U13024 (N_13024,N_12488,N_12313);
or U13025 (N_13025,N_12552,N_12855);
nor U13026 (N_13026,N_12434,N_12807);
xnor U13027 (N_13027,N_12195,N_12985);
and U13028 (N_13028,N_12661,N_12917);
nor U13029 (N_13029,N_12846,N_12223);
or U13030 (N_13030,N_12285,N_12703);
nor U13031 (N_13031,N_12894,N_12006);
xnor U13032 (N_13032,N_12252,N_12901);
nor U13033 (N_13033,N_12508,N_12874);
or U13034 (N_13034,N_12484,N_12026);
nand U13035 (N_13035,N_12966,N_12648);
nand U13036 (N_13036,N_12146,N_12833);
or U13037 (N_13037,N_12897,N_12256);
and U13038 (N_13038,N_12296,N_12355);
nand U13039 (N_13039,N_12704,N_12916);
and U13040 (N_13040,N_12443,N_12038);
nor U13041 (N_13041,N_12915,N_12269);
nor U13042 (N_13042,N_12534,N_12125);
or U13043 (N_13043,N_12806,N_12589);
and U13044 (N_13044,N_12793,N_12290);
and U13045 (N_13045,N_12007,N_12132);
nor U13046 (N_13046,N_12638,N_12567);
nor U13047 (N_13047,N_12227,N_12191);
xor U13048 (N_13048,N_12249,N_12332);
nand U13049 (N_13049,N_12818,N_12194);
xor U13050 (N_13050,N_12716,N_12726);
nand U13051 (N_13051,N_12999,N_12278);
or U13052 (N_13052,N_12625,N_12156);
xor U13053 (N_13053,N_12555,N_12084);
nor U13054 (N_13054,N_12517,N_12691);
nor U13055 (N_13055,N_12336,N_12615);
nor U13056 (N_13056,N_12509,N_12870);
nor U13057 (N_13057,N_12713,N_12882);
nand U13058 (N_13058,N_12939,N_12664);
nand U13059 (N_13059,N_12646,N_12028);
nor U13060 (N_13060,N_12974,N_12457);
and U13061 (N_13061,N_12129,N_12174);
xnor U13062 (N_13062,N_12873,N_12655);
nand U13063 (N_13063,N_12139,N_12030);
nand U13064 (N_13064,N_12024,N_12896);
and U13065 (N_13065,N_12979,N_12930);
or U13066 (N_13066,N_12074,N_12016);
nand U13067 (N_13067,N_12432,N_12933);
and U13068 (N_13068,N_12193,N_12468);
or U13069 (N_13069,N_12852,N_12690);
nand U13070 (N_13070,N_12724,N_12891);
nor U13071 (N_13071,N_12264,N_12388);
or U13072 (N_13072,N_12692,N_12527);
nor U13073 (N_13073,N_12665,N_12328);
nand U13074 (N_13074,N_12546,N_12063);
xor U13075 (N_13075,N_12454,N_12922);
nor U13076 (N_13076,N_12165,N_12617);
xnor U13077 (N_13077,N_12747,N_12566);
nand U13078 (N_13078,N_12340,N_12229);
or U13079 (N_13079,N_12298,N_12014);
xnor U13080 (N_13080,N_12358,N_12554);
nor U13081 (N_13081,N_12613,N_12556);
xnor U13082 (N_13082,N_12118,N_12823);
or U13083 (N_13083,N_12059,N_12236);
and U13084 (N_13084,N_12277,N_12420);
nor U13085 (N_13085,N_12113,N_12418);
nor U13086 (N_13086,N_12456,N_12723);
nand U13087 (N_13087,N_12889,N_12380);
and U13088 (N_13088,N_12473,N_12900);
xnor U13089 (N_13089,N_12768,N_12387);
or U13090 (N_13090,N_12498,N_12600);
and U13091 (N_13091,N_12198,N_12159);
nor U13092 (N_13092,N_12920,N_12748);
nor U13093 (N_13093,N_12588,N_12424);
xor U13094 (N_13094,N_12389,N_12611);
nand U13095 (N_13095,N_12984,N_12295);
nand U13096 (N_13096,N_12449,N_12003);
or U13097 (N_13097,N_12265,N_12234);
nor U13098 (N_13098,N_12992,N_12591);
and U13099 (N_13099,N_12138,N_12145);
nand U13100 (N_13100,N_12276,N_12144);
and U13101 (N_13101,N_12097,N_12272);
or U13102 (N_13102,N_12733,N_12013);
xnor U13103 (N_13103,N_12208,N_12307);
nand U13104 (N_13104,N_12801,N_12157);
nand U13105 (N_13105,N_12969,N_12950);
or U13106 (N_13106,N_12819,N_12354);
nor U13107 (N_13107,N_12303,N_12242);
and U13108 (N_13108,N_12004,N_12490);
or U13109 (N_13109,N_12385,N_12993);
nand U13110 (N_13110,N_12957,N_12426);
and U13111 (N_13111,N_12210,N_12034);
nand U13112 (N_13112,N_12240,N_12927);
nand U13113 (N_13113,N_12904,N_12634);
xnor U13114 (N_13114,N_12452,N_12049);
or U13115 (N_13115,N_12671,N_12645);
nand U13116 (N_13116,N_12268,N_12730);
and U13117 (N_13117,N_12347,N_12124);
or U13118 (N_13118,N_12140,N_12323);
xor U13119 (N_13119,N_12649,N_12180);
nand U13120 (N_13120,N_12366,N_12926);
nor U13121 (N_13121,N_12414,N_12261);
nand U13122 (N_13122,N_12696,N_12953);
or U13123 (N_13123,N_12792,N_12941);
and U13124 (N_13124,N_12319,N_12618);
or U13125 (N_13125,N_12479,N_12031);
nor U13126 (N_13126,N_12598,N_12599);
or U13127 (N_13127,N_12438,N_12831);
nor U13128 (N_13128,N_12105,N_12722);
nand U13129 (N_13129,N_12844,N_12341);
or U13130 (N_13130,N_12856,N_12458);
and U13131 (N_13131,N_12575,N_12382);
and U13132 (N_13132,N_12899,N_12910);
nand U13133 (N_13133,N_12353,N_12288);
nand U13134 (N_13134,N_12944,N_12908);
nand U13135 (N_13135,N_12160,N_12550);
nand U13136 (N_13136,N_12885,N_12417);
nor U13137 (N_13137,N_12482,N_12005);
nand U13138 (N_13138,N_12250,N_12330);
nor U13139 (N_13139,N_12907,N_12116);
xor U13140 (N_13140,N_12780,N_12286);
nor U13141 (N_13141,N_12131,N_12172);
or U13142 (N_13142,N_12441,N_12150);
nor U13143 (N_13143,N_12720,N_12346);
nand U13144 (N_13144,N_12676,N_12994);
and U13145 (N_13145,N_12043,N_12214);
nor U13146 (N_13146,N_12167,N_12022);
or U13147 (N_13147,N_12535,N_12090);
xnor U13148 (N_13148,N_12688,N_12868);
or U13149 (N_13149,N_12756,N_12919);
or U13150 (N_13150,N_12786,N_12155);
nand U13151 (N_13151,N_12083,N_12370);
nand U13152 (N_13152,N_12364,N_12861);
nor U13153 (N_13153,N_12365,N_12800);
and U13154 (N_13154,N_12112,N_12875);
and U13155 (N_13155,N_12141,N_12854);
or U13156 (N_13156,N_12762,N_12179);
xor U13157 (N_13157,N_12647,N_12789);
nor U13158 (N_13158,N_12310,N_12238);
or U13159 (N_13159,N_12080,N_12462);
and U13160 (N_13160,N_12357,N_12830);
or U13161 (N_13161,N_12841,N_12936);
and U13162 (N_13162,N_12672,N_12128);
xnor U13163 (N_13163,N_12121,N_12469);
xnor U13164 (N_13164,N_12185,N_12400);
xor U13165 (N_13165,N_12674,N_12981);
and U13166 (N_13166,N_12796,N_12053);
nand U13167 (N_13167,N_12858,N_12173);
xor U13168 (N_13168,N_12072,N_12437);
or U13169 (N_13169,N_12623,N_12453);
xor U13170 (N_13170,N_12597,N_12565);
xnor U13171 (N_13171,N_12843,N_12130);
or U13172 (N_13172,N_12204,N_12867);
nor U13173 (N_13173,N_12622,N_12101);
nor U13174 (N_13174,N_12551,N_12512);
xnor U13175 (N_13175,N_12660,N_12052);
and U13176 (N_13176,N_12518,N_12317);
or U13177 (N_13177,N_12408,N_12188);
and U13178 (N_13178,N_12849,N_12879);
nand U13179 (N_13179,N_12574,N_12989);
xnor U13180 (N_13180,N_12224,N_12048);
nor U13181 (N_13181,N_12959,N_12189);
xnor U13182 (N_13182,N_12563,N_12318);
and U13183 (N_13183,N_12784,N_12183);
xor U13184 (N_13184,N_12531,N_12501);
nand U13185 (N_13185,N_12521,N_12862);
or U13186 (N_13186,N_12390,N_12311);
nand U13187 (N_13187,N_12371,N_12302);
or U13188 (N_13188,N_12562,N_12375);
nand U13189 (N_13189,N_12892,N_12668);
or U13190 (N_13190,N_12478,N_12399);
or U13191 (N_13191,N_12816,N_12621);
nor U13192 (N_13192,N_12094,N_12911);
and U13193 (N_13193,N_12769,N_12175);
nor U13194 (N_13194,N_12883,N_12241);
nand U13195 (N_13195,N_12106,N_12763);
nor U13196 (N_13196,N_12754,N_12292);
nor U13197 (N_13197,N_12678,N_12243);
or U13198 (N_13198,N_12091,N_12759);
and U13199 (N_13199,N_12036,N_12503);
xnor U13200 (N_13200,N_12176,N_12836);
and U13201 (N_13201,N_12281,N_12778);
xnor U13202 (N_13202,N_12471,N_12761);
or U13203 (N_13203,N_12320,N_12440);
nand U13204 (N_13204,N_12134,N_12973);
and U13205 (N_13205,N_12628,N_12804);
or U13206 (N_13206,N_12201,N_12069);
nand U13207 (N_13207,N_12218,N_12886);
and U13208 (N_13208,N_12502,N_12564);
nand U13209 (N_13209,N_12573,N_12702);
or U13210 (N_13210,N_12271,N_12865);
or U13211 (N_13211,N_12071,N_12935);
or U13212 (N_13212,N_12835,N_12612);
and U13213 (N_13213,N_12120,N_12041);
nor U13214 (N_13214,N_12480,N_12802);
and U13215 (N_13215,N_12656,N_12058);
nor U13216 (N_13216,N_12913,N_12871);
nand U13217 (N_13217,N_12220,N_12682);
nor U13218 (N_13218,N_12051,N_12496);
and U13219 (N_13219,N_12148,N_12499);
or U13220 (N_13220,N_12329,N_12744);
xnor U13221 (N_13221,N_12297,N_12368);
nor U13222 (N_13222,N_12609,N_12620);
or U13223 (N_13223,N_12078,N_12570);
or U13224 (N_13224,N_12951,N_12988);
nor U13225 (N_13225,N_12548,N_12301);
nand U13226 (N_13226,N_12881,N_12832);
or U13227 (N_13227,N_12783,N_12603);
or U13228 (N_13228,N_12685,N_12137);
or U13229 (N_13229,N_12349,N_12779);
and U13230 (N_13230,N_12075,N_12280);
xor U13231 (N_13231,N_12864,N_12406);
or U13232 (N_13232,N_12244,N_12639);
xor U13233 (N_13233,N_12251,N_12359);
xnor U13234 (N_13234,N_12465,N_12746);
or U13235 (N_13235,N_12827,N_12593);
nor U13236 (N_13236,N_12629,N_12483);
nand U13237 (N_13237,N_12197,N_12532);
xor U13238 (N_13238,N_12898,N_12035);
or U13239 (N_13239,N_12445,N_12111);
nand U13240 (N_13240,N_12990,N_12367);
xor U13241 (N_13241,N_12247,N_12729);
xnor U13242 (N_13242,N_12151,N_12263);
nand U13243 (N_13243,N_12632,N_12558);
nor U13244 (N_13244,N_12513,N_12798);
and U13245 (N_13245,N_12859,N_12230);
xor U13246 (N_13246,N_12333,N_12519);
xnor U13247 (N_13247,N_12109,N_12579);
and U13248 (N_13248,N_12299,N_12636);
or U13249 (N_13249,N_12163,N_12960);
xor U13250 (N_13250,N_12978,N_12409);
or U13251 (N_13251,N_12228,N_12415);
or U13252 (N_13252,N_12103,N_12115);
nor U13253 (N_13253,N_12196,N_12212);
and U13254 (N_13254,N_12863,N_12381);
xnor U13255 (N_13255,N_12705,N_12395);
xnor U13256 (N_13256,N_12110,N_12001);
or U13257 (N_13257,N_12717,N_12711);
nor U13258 (N_13258,N_12351,N_12963);
and U13259 (N_13259,N_12644,N_12543);
and U13260 (N_13260,N_12102,N_12050);
or U13261 (N_13261,N_12100,N_12853);
nand U13262 (N_13262,N_12507,N_12650);
nor U13263 (N_13263,N_12460,N_12039);
xnor U13264 (N_13264,N_12493,N_12516);
xor U13265 (N_13265,N_12123,N_12184);
nand U13266 (N_13266,N_12787,N_12710);
nor U13267 (N_13267,N_12133,N_12736);
and U13268 (N_13268,N_12169,N_12257);
nor U13269 (N_13269,N_12652,N_12360);
and U13270 (N_13270,N_12475,N_12530);
xor U13271 (N_13271,N_12755,N_12350);
nand U13272 (N_13272,N_12986,N_12938);
and U13273 (N_13273,N_12055,N_12291);
or U13274 (N_13274,N_12547,N_12222);
or U13275 (N_13275,N_12680,N_12178);
and U13276 (N_13276,N_12338,N_12061);
nor U13277 (N_13277,N_12029,N_12595);
or U13278 (N_13278,N_12221,N_12187);
and U13279 (N_13279,N_12011,N_12834);
xor U13280 (N_13280,N_12970,N_12170);
and U13281 (N_13281,N_12315,N_12497);
nand U13282 (N_13282,N_12738,N_12316);
xor U13283 (N_13283,N_12135,N_12166);
or U13284 (N_13284,N_12663,N_12539);
nand U13285 (N_13285,N_12177,N_12033);
or U13286 (N_13286,N_12162,N_12514);
nor U13287 (N_13287,N_12734,N_12342);
xnor U13288 (N_13288,N_12758,N_12237);
nor U13289 (N_13289,N_12253,N_12965);
or U13290 (N_13290,N_12377,N_12925);
xor U13291 (N_13291,N_12020,N_12056);
xnor U13292 (N_13292,N_12293,N_12119);
xor U13293 (N_13293,N_12439,N_12594);
and U13294 (N_13294,N_12995,N_12066);
xor U13295 (N_13295,N_12096,N_12450);
and U13296 (N_13296,N_12997,N_12699);
and U13297 (N_13297,N_12707,N_12486);
xnor U13298 (N_13298,N_12423,N_12088);
and U13299 (N_13299,N_12814,N_12383);
nand U13300 (N_13300,N_12413,N_12147);
and U13301 (N_13301,N_12949,N_12255);
nor U13302 (N_13302,N_12335,N_12605);
nand U13303 (N_13303,N_12721,N_12666);
nor U13304 (N_13304,N_12374,N_12495);
nor U13305 (N_13305,N_12630,N_12283);
and U13306 (N_13306,N_12444,N_12675);
nand U13307 (N_13307,N_12967,N_12829);
or U13308 (N_13308,N_12258,N_12402);
xnor U13309 (N_13309,N_12087,N_12662);
nor U13310 (N_13310,N_12081,N_12270);
and U13311 (N_13311,N_12403,N_12765);
and U13312 (N_13312,N_12714,N_12541);
and U13313 (N_13313,N_12817,N_12659);
and U13314 (N_13314,N_12407,N_12373);
and U13315 (N_13315,N_12474,N_12749);
xor U13316 (N_13316,N_12766,N_12770);
or U13317 (N_13317,N_12544,N_12481);
or U13318 (N_13318,N_12037,N_12945);
nand U13319 (N_13319,N_12337,N_12876);
xnor U13320 (N_13320,N_12500,N_12788);
or U13321 (N_13321,N_12154,N_12248);
nand U13322 (N_13322,N_12794,N_12308);
xnor U13323 (N_13323,N_12489,N_12209);
or U13324 (N_13324,N_12455,N_12851);
and U13325 (N_13325,N_12824,N_12379);
nand U13326 (N_13326,N_12322,N_12306);
or U13327 (N_13327,N_12740,N_12586);
and U13328 (N_13328,N_12932,N_12673);
nand U13329 (N_13329,N_12528,N_12895);
or U13330 (N_13330,N_12089,N_12062);
or U13331 (N_13331,N_12866,N_12576);
xor U13332 (N_13332,N_12181,N_12421);
xnor U13333 (N_13333,N_12186,N_12903);
nand U13334 (N_13334,N_12772,N_12040);
or U13335 (N_13335,N_12274,N_12905);
nor U13336 (N_13336,N_12822,N_12679);
nand U13337 (N_13337,N_12750,N_12976);
xnor U13338 (N_13338,N_12182,N_12411);
xor U13339 (N_13339,N_12961,N_12161);
or U13340 (N_13340,N_12206,N_12401);
nor U13341 (N_13341,N_12027,N_12677);
xnor U13342 (N_13342,N_12654,N_12614);
or U13343 (N_13343,N_12893,N_12641);
or U13344 (N_13344,N_12568,N_12924);
and U13345 (N_13345,N_12448,N_12604);
or U13346 (N_13346,N_12619,N_12718);
nor U13347 (N_13347,N_12538,N_12376);
or U13348 (N_13348,N_12929,N_12643);
and U13349 (N_13349,N_12937,N_12515);
or U13350 (N_13350,N_12781,N_12466);
nor U13351 (N_13351,N_12309,N_12777);
xnor U13352 (N_13352,N_12398,N_12735);
nand U13353 (N_13353,N_12108,N_12343);
xnor U13354 (N_13354,N_12153,N_12085);
and U13355 (N_13355,N_12239,N_12869);
or U13356 (N_13356,N_12931,N_12719);
xnor U13357 (N_13357,N_12631,N_12695);
nor U13358 (N_13358,N_12943,N_12300);
and U13359 (N_13359,N_12542,N_12136);
and U13360 (N_13360,N_12741,N_12259);
nor U13361 (N_13361,N_12942,N_12447);
nor U13362 (N_13362,N_12627,N_12972);
or U13363 (N_13363,N_12267,N_12235);
and U13364 (N_13364,N_12021,N_12392);
or U13365 (N_13365,N_12934,N_12569);
and U13366 (N_13366,N_12845,N_12289);
xor U13367 (N_13367,N_12689,N_12838);
nor U13368 (N_13368,N_12045,N_12331);
xor U13369 (N_13369,N_12523,N_12312);
and U13370 (N_13370,N_12429,N_12419);
nand U13371 (N_13371,N_12275,N_12470);
or U13372 (N_13372,N_12171,N_12524);
nor U13373 (N_13373,N_12393,N_12266);
nand U13374 (N_13374,N_12065,N_12077);
or U13375 (N_13375,N_12168,N_12811);
nand U13376 (N_13376,N_12808,N_12397);
nor U13377 (N_13377,N_12912,N_12533);
and U13378 (N_13378,N_12706,N_12287);
xor U13379 (N_13379,N_12522,N_12092);
nand U13380 (N_13380,N_12219,N_12459);
xor U13381 (N_13381,N_12887,N_12428);
nor U13382 (N_13382,N_12812,N_12624);
nor U13383 (N_13383,N_12391,N_12260);
and U13384 (N_13384,N_12626,N_12923);
nor U13385 (N_13385,N_12070,N_12216);
and U13386 (N_13386,N_12504,N_12494);
nor U13387 (N_13387,N_12982,N_12590);
and U13388 (N_13388,N_12584,N_12142);
nand U13389 (N_13389,N_12540,N_12964);
and U13390 (N_13390,N_12431,N_12667);
nand U13391 (N_13391,N_12737,N_12651);
nor U13392 (N_13392,N_12361,N_12760);
or U13393 (N_13393,N_12890,N_12412);
nand U13394 (N_13394,N_12637,N_12902);
xor U13395 (N_13395,N_12436,N_12334);
nor U13396 (N_13396,N_12996,N_12246);
nor U13397 (N_13397,N_12505,N_12775);
xnor U13398 (N_13398,N_12245,N_12492);
or U13399 (N_13399,N_12577,N_12203);
and U13400 (N_13400,N_12683,N_12487);
and U13401 (N_13401,N_12463,N_12345);
nor U13402 (N_13402,N_12363,N_12233);
and U13403 (N_13403,N_12709,N_12327);
and U13404 (N_13404,N_12653,N_12553);
nand U13405 (N_13405,N_12506,N_12752);
xnor U13406 (N_13406,N_12199,N_12149);
and U13407 (N_13407,N_12213,N_12114);
or U13408 (N_13408,N_12324,N_12821);
xnor U13409 (N_13409,N_12745,N_12742);
and U13410 (N_13410,N_12545,N_12888);
or U13411 (N_13411,N_12921,N_12476);
and U13412 (N_13412,N_12670,N_12410);
nand U13413 (N_13413,N_12581,N_12602);
nand U13414 (N_13414,N_12764,N_12294);
or U13415 (N_13415,N_12557,N_12232);
nor U13416 (N_13416,N_12073,N_12607);
or U13417 (N_13417,N_12946,N_12608);
xor U13418 (N_13418,N_12694,N_12606);
nor U13419 (N_13419,N_12158,N_12042);
or U13420 (N_13420,N_12202,N_12190);
xor U13421 (N_13421,N_12751,N_12725);
xor U13422 (N_13422,N_12842,N_12848);
xnor U13423 (N_13423,N_12803,N_12928);
or U13424 (N_13424,N_12047,N_12767);
nor U13425 (N_13425,N_12825,N_12321);
nor U13426 (N_13426,N_12010,N_12712);
and U13427 (N_13427,N_12715,N_12314);
or U13428 (N_13428,N_12023,N_12352);
or U13429 (N_13429,N_12435,N_12082);
nor U13430 (N_13430,N_12464,N_12017);
and U13431 (N_13431,N_12107,N_12776);
nor U13432 (N_13432,N_12231,N_12633);
nor U13433 (N_13433,N_12991,N_12743);
nor U13434 (N_13434,N_12728,N_12000);
xor U13435 (N_13435,N_12791,N_12384);
and U13436 (N_13436,N_12977,N_12537);
or U13437 (N_13437,N_12520,N_12305);
nor U13438 (N_13438,N_12284,N_12810);
nand U13439 (N_13439,N_12727,N_12610);
or U13440 (N_13440,N_12947,N_12536);
or U13441 (N_13441,N_12687,N_12559);
and U13442 (N_13442,N_12378,N_12304);
and U13443 (N_13443,N_12009,N_12561);
nor U13444 (N_13444,N_12442,N_12592);
nor U13445 (N_13445,N_12127,N_12254);
xor U13446 (N_13446,N_12279,N_12878);
and U13447 (N_13447,N_12356,N_12032);
nand U13448 (N_13448,N_12467,N_12093);
or U13449 (N_13449,N_12477,N_12914);
or U13450 (N_13450,N_12732,N_12774);
nor U13451 (N_13451,N_12580,N_12095);
nand U13452 (N_13452,N_12805,N_12948);
nor U13453 (N_13453,N_12344,N_12698);
nor U13454 (N_13454,N_12046,N_12954);
xnor U13455 (N_13455,N_12425,N_12684);
xnor U13456 (N_13456,N_12526,N_12446);
and U13457 (N_13457,N_12731,N_12273);
nand U13458 (N_13458,N_12152,N_12955);
nor U13459 (N_13459,N_12164,N_12857);
xor U13460 (N_13460,N_12815,N_12416);
nand U13461 (N_13461,N_12642,N_12396);
xnor U13462 (N_13462,N_12217,N_12681);
and U13463 (N_13463,N_12054,N_12739);
nor U13464 (N_13464,N_12433,N_12906);
nor U13465 (N_13465,N_12983,N_12404);
nand U13466 (N_13466,N_12826,N_12596);
nand U13467 (N_13467,N_12386,N_12200);
nor U13468 (N_13468,N_12813,N_12582);
nor U13469 (N_13469,N_12635,N_12773);
and U13470 (N_13470,N_12601,N_12585);
nor U13471 (N_13471,N_12968,N_12225);
nor U13472 (N_13472,N_12820,N_12326);
or U13473 (N_13473,N_12282,N_12877);
and U13474 (N_13474,N_12797,N_12657);
nor U13475 (N_13475,N_12956,N_12511);
or U13476 (N_13476,N_12430,N_12099);
xnor U13477 (N_13477,N_12067,N_12952);
or U13478 (N_13478,N_12782,N_12998);
nand U13479 (N_13479,N_12701,N_12205);
and U13480 (N_13480,N_12583,N_12207);
nand U13481 (N_13481,N_12771,N_12572);
and U13482 (N_13482,N_12491,N_12790);
xnor U13483 (N_13483,N_12909,N_12880);
xnor U13484 (N_13484,N_12708,N_12587);
nand U13485 (N_13485,N_12126,N_12840);
or U13486 (N_13486,N_12117,N_12079);
or U13487 (N_13487,N_12019,N_12847);
and U13488 (N_13488,N_12485,N_12018);
xnor U13489 (N_13489,N_12427,N_12578);
or U13490 (N_13490,N_12211,N_12837);
nor U13491 (N_13491,N_12669,N_12002);
nor U13492 (N_13492,N_12008,N_12962);
nor U13493 (N_13493,N_12015,N_12640);
nor U13494 (N_13494,N_12839,N_12068);
xnor U13495 (N_13495,N_12753,N_12658);
or U13496 (N_13496,N_12025,N_12697);
and U13497 (N_13497,N_12451,N_12262);
or U13498 (N_13498,N_12348,N_12884);
or U13499 (N_13499,N_12064,N_12057);
or U13500 (N_13500,N_12071,N_12994);
nor U13501 (N_13501,N_12501,N_12210);
xor U13502 (N_13502,N_12886,N_12363);
or U13503 (N_13503,N_12656,N_12974);
nand U13504 (N_13504,N_12915,N_12107);
xnor U13505 (N_13505,N_12090,N_12922);
nor U13506 (N_13506,N_12515,N_12098);
nand U13507 (N_13507,N_12782,N_12308);
or U13508 (N_13508,N_12498,N_12594);
nand U13509 (N_13509,N_12629,N_12913);
xor U13510 (N_13510,N_12440,N_12529);
nand U13511 (N_13511,N_12771,N_12177);
or U13512 (N_13512,N_12544,N_12780);
xnor U13513 (N_13513,N_12321,N_12012);
or U13514 (N_13514,N_12121,N_12324);
xor U13515 (N_13515,N_12472,N_12156);
and U13516 (N_13516,N_12695,N_12952);
and U13517 (N_13517,N_12765,N_12465);
or U13518 (N_13518,N_12869,N_12469);
nor U13519 (N_13519,N_12845,N_12473);
or U13520 (N_13520,N_12515,N_12492);
and U13521 (N_13521,N_12721,N_12708);
nand U13522 (N_13522,N_12618,N_12742);
nand U13523 (N_13523,N_12495,N_12886);
nor U13524 (N_13524,N_12568,N_12853);
or U13525 (N_13525,N_12195,N_12659);
or U13526 (N_13526,N_12667,N_12606);
or U13527 (N_13527,N_12391,N_12548);
or U13528 (N_13528,N_12389,N_12235);
nor U13529 (N_13529,N_12246,N_12393);
or U13530 (N_13530,N_12348,N_12483);
or U13531 (N_13531,N_12404,N_12227);
nor U13532 (N_13532,N_12692,N_12046);
and U13533 (N_13533,N_12523,N_12423);
xor U13534 (N_13534,N_12394,N_12926);
and U13535 (N_13535,N_12152,N_12735);
and U13536 (N_13536,N_12186,N_12551);
nand U13537 (N_13537,N_12410,N_12931);
nand U13538 (N_13538,N_12669,N_12133);
nor U13539 (N_13539,N_12486,N_12119);
xnor U13540 (N_13540,N_12206,N_12375);
nand U13541 (N_13541,N_12963,N_12677);
xor U13542 (N_13542,N_12446,N_12256);
nor U13543 (N_13543,N_12495,N_12341);
xnor U13544 (N_13544,N_12356,N_12776);
nor U13545 (N_13545,N_12305,N_12416);
xnor U13546 (N_13546,N_12738,N_12856);
or U13547 (N_13547,N_12719,N_12070);
nand U13548 (N_13548,N_12536,N_12007);
nor U13549 (N_13549,N_12997,N_12993);
nand U13550 (N_13550,N_12133,N_12027);
nand U13551 (N_13551,N_12296,N_12683);
nand U13552 (N_13552,N_12689,N_12251);
nand U13553 (N_13553,N_12105,N_12107);
nor U13554 (N_13554,N_12067,N_12220);
xnor U13555 (N_13555,N_12405,N_12247);
and U13556 (N_13556,N_12262,N_12032);
or U13557 (N_13557,N_12522,N_12140);
and U13558 (N_13558,N_12093,N_12821);
or U13559 (N_13559,N_12067,N_12443);
nor U13560 (N_13560,N_12543,N_12544);
and U13561 (N_13561,N_12337,N_12150);
or U13562 (N_13562,N_12701,N_12585);
and U13563 (N_13563,N_12778,N_12838);
xnor U13564 (N_13564,N_12033,N_12063);
nor U13565 (N_13565,N_12606,N_12281);
nand U13566 (N_13566,N_12845,N_12910);
and U13567 (N_13567,N_12087,N_12214);
nor U13568 (N_13568,N_12717,N_12231);
xor U13569 (N_13569,N_12759,N_12825);
or U13570 (N_13570,N_12608,N_12794);
or U13571 (N_13571,N_12836,N_12004);
nor U13572 (N_13572,N_12931,N_12025);
nor U13573 (N_13573,N_12118,N_12167);
and U13574 (N_13574,N_12021,N_12442);
xnor U13575 (N_13575,N_12661,N_12035);
nand U13576 (N_13576,N_12596,N_12279);
or U13577 (N_13577,N_12405,N_12983);
xnor U13578 (N_13578,N_12940,N_12316);
or U13579 (N_13579,N_12891,N_12930);
nand U13580 (N_13580,N_12531,N_12951);
xnor U13581 (N_13581,N_12232,N_12655);
xor U13582 (N_13582,N_12228,N_12138);
nand U13583 (N_13583,N_12961,N_12948);
or U13584 (N_13584,N_12827,N_12698);
or U13585 (N_13585,N_12087,N_12955);
xor U13586 (N_13586,N_12430,N_12580);
and U13587 (N_13587,N_12595,N_12813);
or U13588 (N_13588,N_12971,N_12050);
xnor U13589 (N_13589,N_12102,N_12340);
and U13590 (N_13590,N_12201,N_12542);
nor U13591 (N_13591,N_12693,N_12403);
xor U13592 (N_13592,N_12060,N_12253);
nand U13593 (N_13593,N_12083,N_12298);
xnor U13594 (N_13594,N_12172,N_12302);
or U13595 (N_13595,N_12767,N_12065);
nand U13596 (N_13596,N_12984,N_12103);
or U13597 (N_13597,N_12184,N_12513);
xor U13598 (N_13598,N_12320,N_12076);
and U13599 (N_13599,N_12828,N_12070);
nor U13600 (N_13600,N_12756,N_12807);
or U13601 (N_13601,N_12551,N_12584);
nor U13602 (N_13602,N_12980,N_12161);
nor U13603 (N_13603,N_12284,N_12015);
or U13604 (N_13604,N_12998,N_12734);
xor U13605 (N_13605,N_12018,N_12763);
xnor U13606 (N_13606,N_12575,N_12041);
xor U13607 (N_13607,N_12577,N_12092);
or U13608 (N_13608,N_12309,N_12452);
xor U13609 (N_13609,N_12170,N_12486);
nand U13610 (N_13610,N_12706,N_12666);
nor U13611 (N_13611,N_12293,N_12507);
nor U13612 (N_13612,N_12418,N_12465);
nand U13613 (N_13613,N_12786,N_12729);
nor U13614 (N_13614,N_12165,N_12177);
nor U13615 (N_13615,N_12279,N_12669);
or U13616 (N_13616,N_12450,N_12489);
and U13617 (N_13617,N_12516,N_12111);
and U13618 (N_13618,N_12545,N_12818);
nor U13619 (N_13619,N_12509,N_12723);
xor U13620 (N_13620,N_12072,N_12091);
and U13621 (N_13621,N_12578,N_12104);
xnor U13622 (N_13622,N_12365,N_12899);
xnor U13623 (N_13623,N_12881,N_12821);
nand U13624 (N_13624,N_12592,N_12782);
and U13625 (N_13625,N_12591,N_12534);
nor U13626 (N_13626,N_12031,N_12485);
and U13627 (N_13627,N_12074,N_12145);
and U13628 (N_13628,N_12379,N_12883);
xor U13629 (N_13629,N_12396,N_12702);
xnor U13630 (N_13630,N_12695,N_12762);
nor U13631 (N_13631,N_12252,N_12590);
nor U13632 (N_13632,N_12212,N_12250);
nand U13633 (N_13633,N_12866,N_12371);
nand U13634 (N_13634,N_12997,N_12640);
and U13635 (N_13635,N_12325,N_12065);
and U13636 (N_13636,N_12800,N_12663);
xnor U13637 (N_13637,N_12858,N_12680);
or U13638 (N_13638,N_12323,N_12334);
nand U13639 (N_13639,N_12136,N_12574);
or U13640 (N_13640,N_12705,N_12980);
and U13641 (N_13641,N_12526,N_12733);
and U13642 (N_13642,N_12209,N_12602);
or U13643 (N_13643,N_12548,N_12353);
nand U13644 (N_13644,N_12323,N_12317);
nand U13645 (N_13645,N_12143,N_12818);
or U13646 (N_13646,N_12409,N_12754);
and U13647 (N_13647,N_12837,N_12424);
nand U13648 (N_13648,N_12707,N_12463);
or U13649 (N_13649,N_12905,N_12606);
and U13650 (N_13650,N_12636,N_12389);
xor U13651 (N_13651,N_12298,N_12045);
nor U13652 (N_13652,N_12893,N_12053);
nor U13653 (N_13653,N_12351,N_12493);
nor U13654 (N_13654,N_12553,N_12489);
and U13655 (N_13655,N_12619,N_12429);
nor U13656 (N_13656,N_12195,N_12840);
or U13657 (N_13657,N_12944,N_12084);
nand U13658 (N_13658,N_12417,N_12675);
and U13659 (N_13659,N_12269,N_12822);
and U13660 (N_13660,N_12469,N_12452);
and U13661 (N_13661,N_12053,N_12300);
nand U13662 (N_13662,N_12645,N_12600);
nand U13663 (N_13663,N_12169,N_12967);
or U13664 (N_13664,N_12488,N_12557);
or U13665 (N_13665,N_12842,N_12803);
nand U13666 (N_13666,N_12034,N_12732);
nor U13667 (N_13667,N_12013,N_12961);
nor U13668 (N_13668,N_12279,N_12323);
xor U13669 (N_13669,N_12604,N_12808);
nand U13670 (N_13670,N_12968,N_12194);
xor U13671 (N_13671,N_12037,N_12091);
or U13672 (N_13672,N_12495,N_12358);
xor U13673 (N_13673,N_12556,N_12292);
or U13674 (N_13674,N_12217,N_12476);
nor U13675 (N_13675,N_12889,N_12811);
and U13676 (N_13676,N_12753,N_12870);
nor U13677 (N_13677,N_12084,N_12429);
or U13678 (N_13678,N_12073,N_12553);
nor U13679 (N_13679,N_12176,N_12369);
nand U13680 (N_13680,N_12214,N_12318);
and U13681 (N_13681,N_12832,N_12616);
and U13682 (N_13682,N_12962,N_12511);
nand U13683 (N_13683,N_12906,N_12796);
nor U13684 (N_13684,N_12555,N_12733);
and U13685 (N_13685,N_12697,N_12600);
and U13686 (N_13686,N_12799,N_12868);
nand U13687 (N_13687,N_12148,N_12941);
and U13688 (N_13688,N_12057,N_12199);
nor U13689 (N_13689,N_12081,N_12795);
or U13690 (N_13690,N_12592,N_12112);
nand U13691 (N_13691,N_12856,N_12373);
or U13692 (N_13692,N_12126,N_12758);
or U13693 (N_13693,N_12590,N_12995);
or U13694 (N_13694,N_12113,N_12866);
xnor U13695 (N_13695,N_12601,N_12943);
nor U13696 (N_13696,N_12581,N_12789);
xnor U13697 (N_13697,N_12738,N_12676);
nand U13698 (N_13698,N_12241,N_12285);
or U13699 (N_13699,N_12309,N_12493);
nand U13700 (N_13700,N_12927,N_12050);
and U13701 (N_13701,N_12736,N_12760);
and U13702 (N_13702,N_12239,N_12073);
nor U13703 (N_13703,N_12424,N_12379);
or U13704 (N_13704,N_12192,N_12105);
or U13705 (N_13705,N_12693,N_12212);
and U13706 (N_13706,N_12873,N_12215);
xor U13707 (N_13707,N_12376,N_12191);
xor U13708 (N_13708,N_12344,N_12457);
and U13709 (N_13709,N_12809,N_12250);
nor U13710 (N_13710,N_12403,N_12599);
nand U13711 (N_13711,N_12082,N_12981);
nand U13712 (N_13712,N_12223,N_12076);
or U13713 (N_13713,N_12997,N_12162);
and U13714 (N_13714,N_12614,N_12930);
xor U13715 (N_13715,N_12557,N_12192);
and U13716 (N_13716,N_12111,N_12106);
or U13717 (N_13717,N_12398,N_12139);
nor U13718 (N_13718,N_12839,N_12816);
xor U13719 (N_13719,N_12225,N_12910);
nand U13720 (N_13720,N_12463,N_12186);
and U13721 (N_13721,N_12307,N_12662);
nor U13722 (N_13722,N_12725,N_12028);
nand U13723 (N_13723,N_12080,N_12786);
xor U13724 (N_13724,N_12352,N_12231);
and U13725 (N_13725,N_12727,N_12293);
nor U13726 (N_13726,N_12516,N_12204);
nor U13727 (N_13727,N_12073,N_12716);
nand U13728 (N_13728,N_12063,N_12287);
nand U13729 (N_13729,N_12830,N_12689);
nor U13730 (N_13730,N_12166,N_12411);
nand U13731 (N_13731,N_12841,N_12454);
nand U13732 (N_13732,N_12111,N_12808);
nor U13733 (N_13733,N_12127,N_12140);
xnor U13734 (N_13734,N_12206,N_12291);
xor U13735 (N_13735,N_12732,N_12483);
nand U13736 (N_13736,N_12093,N_12204);
nor U13737 (N_13737,N_12832,N_12110);
nand U13738 (N_13738,N_12621,N_12407);
xnor U13739 (N_13739,N_12583,N_12972);
or U13740 (N_13740,N_12181,N_12888);
nor U13741 (N_13741,N_12473,N_12718);
nor U13742 (N_13742,N_12251,N_12169);
nor U13743 (N_13743,N_12181,N_12455);
nor U13744 (N_13744,N_12015,N_12394);
nand U13745 (N_13745,N_12073,N_12752);
or U13746 (N_13746,N_12637,N_12504);
nor U13747 (N_13747,N_12489,N_12146);
and U13748 (N_13748,N_12860,N_12388);
and U13749 (N_13749,N_12862,N_12436);
nor U13750 (N_13750,N_12216,N_12257);
xor U13751 (N_13751,N_12421,N_12846);
nor U13752 (N_13752,N_12658,N_12354);
nor U13753 (N_13753,N_12920,N_12709);
nor U13754 (N_13754,N_12376,N_12315);
xor U13755 (N_13755,N_12488,N_12563);
nor U13756 (N_13756,N_12792,N_12311);
or U13757 (N_13757,N_12695,N_12170);
nand U13758 (N_13758,N_12736,N_12374);
or U13759 (N_13759,N_12098,N_12251);
xor U13760 (N_13760,N_12882,N_12781);
nand U13761 (N_13761,N_12562,N_12629);
or U13762 (N_13762,N_12424,N_12957);
or U13763 (N_13763,N_12833,N_12441);
nor U13764 (N_13764,N_12961,N_12343);
nor U13765 (N_13765,N_12991,N_12334);
and U13766 (N_13766,N_12469,N_12622);
or U13767 (N_13767,N_12504,N_12174);
nor U13768 (N_13768,N_12288,N_12489);
or U13769 (N_13769,N_12591,N_12876);
or U13770 (N_13770,N_12536,N_12531);
or U13771 (N_13771,N_12735,N_12902);
and U13772 (N_13772,N_12830,N_12471);
and U13773 (N_13773,N_12425,N_12640);
xnor U13774 (N_13774,N_12655,N_12716);
nand U13775 (N_13775,N_12622,N_12094);
nor U13776 (N_13776,N_12383,N_12550);
xnor U13777 (N_13777,N_12704,N_12131);
or U13778 (N_13778,N_12069,N_12641);
nand U13779 (N_13779,N_12620,N_12378);
or U13780 (N_13780,N_12149,N_12205);
nand U13781 (N_13781,N_12301,N_12251);
xor U13782 (N_13782,N_12657,N_12350);
or U13783 (N_13783,N_12162,N_12047);
xor U13784 (N_13784,N_12644,N_12042);
or U13785 (N_13785,N_12522,N_12899);
nand U13786 (N_13786,N_12535,N_12579);
nor U13787 (N_13787,N_12939,N_12068);
and U13788 (N_13788,N_12848,N_12514);
or U13789 (N_13789,N_12955,N_12268);
and U13790 (N_13790,N_12586,N_12401);
and U13791 (N_13791,N_12388,N_12022);
xnor U13792 (N_13792,N_12435,N_12255);
and U13793 (N_13793,N_12245,N_12902);
xor U13794 (N_13794,N_12119,N_12015);
nand U13795 (N_13795,N_12859,N_12511);
nand U13796 (N_13796,N_12757,N_12907);
nor U13797 (N_13797,N_12946,N_12376);
nand U13798 (N_13798,N_12139,N_12218);
nor U13799 (N_13799,N_12957,N_12384);
xnor U13800 (N_13800,N_12910,N_12750);
nand U13801 (N_13801,N_12396,N_12300);
nand U13802 (N_13802,N_12078,N_12229);
nor U13803 (N_13803,N_12020,N_12954);
and U13804 (N_13804,N_12242,N_12218);
and U13805 (N_13805,N_12042,N_12230);
nand U13806 (N_13806,N_12950,N_12992);
nor U13807 (N_13807,N_12346,N_12447);
xor U13808 (N_13808,N_12735,N_12453);
nor U13809 (N_13809,N_12421,N_12016);
xnor U13810 (N_13810,N_12952,N_12494);
nand U13811 (N_13811,N_12642,N_12143);
nor U13812 (N_13812,N_12955,N_12751);
nor U13813 (N_13813,N_12226,N_12660);
nor U13814 (N_13814,N_12792,N_12080);
and U13815 (N_13815,N_12221,N_12179);
xnor U13816 (N_13816,N_12628,N_12149);
and U13817 (N_13817,N_12776,N_12191);
nand U13818 (N_13818,N_12455,N_12726);
xor U13819 (N_13819,N_12941,N_12720);
and U13820 (N_13820,N_12206,N_12459);
nor U13821 (N_13821,N_12323,N_12151);
nor U13822 (N_13822,N_12034,N_12066);
or U13823 (N_13823,N_12495,N_12530);
and U13824 (N_13824,N_12316,N_12905);
xnor U13825 (N_13825,N_12872,N_12935);
nand U13826 (N_13826,N_12042,N_12656);
or U13827 (N_13827,N_12834,N_12377);
nand U13828 (N_13828,N_12409,N_12985);
and U13829 (N_13829,N_12069,N_12252);
nand U13830 (N_13830,N_12862,N_12285);
xor U13831 (N_13831,N_12102,N_12851);
nand U13832 (N_13832,N_12968,N_12832);
nor U13833 (N_13833,N_12998,N_12664);
nand U13834 (N_13834,N_12040,N_12474);
and U13835 (N_13835,N_12186,N_12134);
nor U13836 (N_13836,N_12300,N_12409);
and U13837 (N_13837,N_12665,N_12083);
nand U13838 (N_13838,N_12963,N_12295);
xor U13839 (N_13839,N_12369,N_12030);
nand U13840 (N_13840,N_12900,N_12323);
nor U13841 (N_13841,N_12634,N_12554);
and U13842 (N_13842,N_12542,N_12649);
and U13843 (N_13843,N_12411,N_12902);
and U13844 (N_13844,N_12246,N_12634);
xor U13845 (N_13845,N_12898,N_12332);
nand U13846 (N_13846,N_12592,N_12626);
xor U13847 (N_13847,N_12042,N_12552);
nand U13848 (N_13848,N_12831,N_12943);
or U13849 (N_13849,N_12445,N_12501);
xor U13850 (N_13850,N_12433,N_12873);
nor U13851 (N_13851,N_12295,N_12524);
or U13852 (N_13852,N_12499,N_12294);
nor U13853 (N_13853,N_12592,N_12107);
nand U13854 (N_13854,N_12918,N_12433);
nand U13855 (N_13855,N_12296,N_12773);
xnor U13856 (N_13856,N_12843,N_12000);
or U13857 (N_13857,N_12510,N_12893);
xor U13858 (N_13858,N_12855,N_12624);
xnor U13859 (N_13859,N_12706,N_12879);
nand U13860 (N_13860,N_12718,N_12727);
or U13861 (N_13861,N_12289,N_12854);
and U13862 (N_13862,N_12316,N_12260);
xor U13863 (N_13863,N_12644,N_12461);
xnor U13864 (N_13864,N_12246,N_12791);
nor U13865 (N_13865,N_12148,N_12112);
or U13866 (N_13866,N_12691,N_12485);
nor U13867 (N_13867,N_12714,N_12732);
nand U13868 (N_13868,N_12157,N_12026);
xor U13869 (N_13869,N_12140,N_12004);
or U13870 (N_13870,N_12190,N_12591);
xnor U13871 (N_13871,N_12786,N_12090);
nor U13872 (N_13872,N_12163,N_12303);
or U13873 (N_13873,N_12228,N_12265);
xor U13874 (N_13874,N_12432,N_12398);
nand U13875 (N_13875,N_12470,N_12956);
nand U13876 (N_13876,N_12287,N_12737);
and U13877 (N_13877,N_12021,N_12223);
or U13878 (N_13878,N_12032,N_12185);
xor U13879 (N_13879,N_12319,N_12981);
nand U13880 (N_13880,N_12930,N_12625);
or U13881 (N_13881,N_12227,N_12238);
or U13882 (N_13882,N_12711,N_12693);
nand U13883 (N_13883,N_12009,N_12551);
and U13884 (N_13884,N_12733,N_12990);
and U13885 (N_13885,N_12729,N_12083);
xnor U13886 (N_13886,N_12821,N_12867);
nand U13887 (N_13887,N_12558,N_12758);
or U13888 (N_13888,N_12583,N_12514);
nand U13889 (N_13889,N_12661,N_12140);
nand U13890 (N_13890,N_12991,N_12489);
xnor U13891 (N_13891,N_12113,N_12871);
nand U13892 (N_13892,N_12361,N_12848);
or U13893 (N_13893,N_12276,N_12263);
and U13894 (N_13894,N_12322,N_12058);
xor U13895 (N_13895,N_12226,N_12978);
and U13896 (N_13896,N_12071,N_12327);
and U13897 (N_13897,N_12541,N_12131);
nor U13898 (N_13898,N_12183,N_12059);
and U13899 (N_13899,N_12406,N_12915);
nand U13900 (N_13900,N_12450,N_12454);
xnor U13901 (N_13901,N_12474,N_12537);
nor U13902 (N_13902,N_12093,N_12723);
and U13903 (N_13903,N_12375,N_12816);
or U13904 (N_13904,N_12494,N_12396);
nand U13905 (N_13905,N_12073,N_12811);
xor U13906 (N_13906,N_12084,N_12926);
or U13907 (N_13907,N_12818,N_12778);
xor U13908 (N_13908,N_12433,N_12553);
nand U13909 (N_13909,N_12223,N_12346);
nor U13910 (N_13910,N_12338,N_12799);
nand U13911 (N_13911,N_12492,N_12039);
xnor U13912 (N_13912,N_12708,N_12673);
xnor U13913 (N_13913,N_12097,N_12975);
xnor U13914 (N_13914,N_12044,N_12596);
and U13915 (N_13915,N_12854,N_12416);
and U13916 (N_13916,N_12982,N_12510);
or U13917 (N_13917,N_12313,N_12090);
nor U13918 (N_13918,N_12436,N_12631);
or U13919 (N_13919,N_12575,N_12747);
and U13920 (N_13920,N_12632,N_12404);
or U13921 (N_13921,N_12048,N_12974);
nor U13922 (N_13922,N_12383,N_12712);
nor U13923 (N_13923,N_12810,N_12635);
or U13924 (N_13924,N_12900,N_12015);
nand U13925 (N_13925,N_12843,N_12413);
nor U13926 (N_13926,N_12333,N_12582);
and U13927 (N_13927,N_12850,N_12067);
nand U13928 (N_13928,N_12106,N_12941);
nand U13929 (N_13929,N_12228,N_12010);
nand U13930 (N_13930,N_12090,N_12202);
nor U13931 (N_13931,N_12770,N_12971);
nand U13932 (N_13932,N_12960,N_12703);
xnor U13933 (N_13933,N_12613,N_12044);
or U13934 (N_13934,N_12816,N_12485);
nor U13935 (N_13935,N_12351,N_12469);
and U13936 (N_13936,N_12548,N_12248);
nor U13937 (N_13937,N_12540,N_12347);
nor U13938 (N_13938,N_12603,N_12697);
xor U13939 (N_13939,N_12531,N_12039);
or U13940 (N_13940,N_12785,N_12343);
xnor U13941 (N_13941,N_12402,N_12660);
and U13942 (N_13942,N_12210,N_12945);
or U13943 (N_13943,N_12322,N_12908);
xnor U13944 (N_13944,N_12187,N_12039);
nand U13945 (N_13945,N_12472,N_12876);
and U13946 (N_13946,N_12893,N_12205);
nand U13947 (N_13947,N_12376,N_12540);
or U13948 (N_13948,N_12860,N_12455);
nand U13949 (N_13949,N_12639,N_12587);
xor U13950 (N_13950,N_12271,N_12784);
nand U13951 (N_13951,N_12644,N_12428);
and U13952 (N_13952,N_12589,N_12366);
nor U13953 (N_13953,N_12576,N_12971);
nor U13954 (N_13954,N_12550,N_12522);
and U13955 (N_13955,N_12584,N_12878);
and U13956 (N_13956,N_12163,N_12478);
nand U13957 (N_13957,N_12548,N_12427);
or U13958 (N_13958,N_12055,N_12056);
or U13959 (N_13959,N_12019,N_12225);
and U13960 (N_13960,N_12798,N_12246);
and U13961 (N_13961,N_12155,N_12428);
nand U13962 (N_13962,N_12839,N_12079);
and U13963 (N_13963,N_12175,N_12679);
nor U13964 (N_13964,N_12830,N_12677);
nor U13965 (N_13965,N_12171,N_12363);
xor U13966 (N_13966,N_12082,N_12342);
and U13967 (N_13967,N_12477,N_12997);
or U13968 (N_13968,N_12279,N_12063);
nand U13969 (N_13969,N_12077,N_12470);
nor U13970 (N_13970,N_12431,N_12699);
xor U13971 (N_13971,N_12104,N_12774);
nand U13972 (N_13972,N_12882,N_12012);
xor U13973 (N_13973,N_12867,N_12111);
nor U13974 (N_13974,N_12545,N_12058);
and U13975 (N_13975,N_12118,N_12769);
and U13976 (N_13976,N_12943,N_12669);
xor U13977 (N_13977,N_12976,N_12195);
and U13978 (N_13978,N_12910,N_12081);
nand U13979 (N_13979,N_12222,N_12943);
xor U13980 (N_13980,N_12866,N_12809);
or U13981 (N_13981,N_12467,N_12018);
nor U13982 (N_13982,N_12888,N_12463);
nor U13983 (N_13983,N_12104,N_12670);
xnor U13984 (N_13984,N_12121,N_12899);
and U13985 (N_13985,N_12974,N_12722);
xnor U13986 (N_13986,N_12017,N_12031);
nand U13987 (N_13987,N_12936,N_12238);
xnor U13988 (N_13988,N_12504,N_12778);
or U13989 (N_13989,N_12685,N_12539);
or U13990 (N_13990,N_12705,N_12284);
xor U13991 (N_13991,N_12749,N_12895);
and U13992 (N_13992,N_12379,N_12634);
or U13993 (N_13993,N_12077,N_12746);
xor U13994 (N_13994,N_12280,N_12599);
xnor U13995 (N_13995,N_12519,N_12688);
nand U13996 (N_13996,N_12649,N_12877);
and U13997 (N_13997,N_12104,N_12756);
or U13998 (N_13998,N_12353,N_12951);
or U13999 (N_13999,N_12731,N_12663);
and U14000 (N_14000,N_13343,N_13102);
or U14001 (N_14001,N_13719,N_13607);
and U14002 (N_14002,N_13562,N_13693);
or U14003 (N_14003,N_13299,N_13634);
or U14004 (N_14004,N_13797,N_13799);
nand U14005 (N_14005,N_13967,N_13982);
xor U14006 (N_14006,N_13162,N_13254);
or U14007 (N_14007,N_13042,N_13457);
nor U14008 (N_14008,N_13603,N_13574);
or U14009 (N_14009,N_13216,N_13208);
or U14010 (N_14010,N_13902,N_13110);
or U14011 (N_14011,N_13297,N_13853);
nand U14012 (N_14012,N_13304,N_13375);
nand U14013 (N_14013,N_13534,N_13941);
or U14014 (N_14014,N_13316,N_13252);
nor U14015 (N_14015,N_13218,N_13688);
nor U14016 (N_14016,N_13761,N_13883);
or U14017 (N_14017,N_13073,N_13080);
and U14018 (N_14018,N_13178,N_13636);
nor U14019 (N_14019,N_13029,N_13579);
xor U14020 (N_14020,N_13917,N_13262);
nand U14021 (N_14021,N_13597,N_13054);
xor U14022 (N_14022,N_13478,N_13240);
nand U14023 (N_14023,N_13847,N_13135);
xnor U14024 (N_14024,N_13676,N_13094);
xor U14025 (N_14025,N_13253,N_13849);
or U14026 (N_14026,N_13349,N_13625);
or U14027 (N_14027,N_13663,N_13837);
nand U14028 (N_14028,N_13128,N_13602);
or U14029 (N_14029,N_13116,N_13325);
nor U14030 (N_14030,N_13929,N_13228);
or U14031 (N_14031,N_13845,N_13322);
nand U14032 (N_14032,N_13736,N_13449);
or U14033 (N_14033,N_13113,N_13842);
and U14034 (N_14034,N_13956,N_13266);
or U14035 (N_14035,N_13996,N_13337);
nand U14036 (N_14036,N_13541,N_13631);
xnor U14037 (N_14037,N_13239,N_13923);
nand U14038 (N_14038,N_13918,N_13209);
nand U14039 (N_14039,N_13458,N_13238);
nor U14040 (N_14040,N_13168,N_13021);
or U14041 (N_14041,N_13617,N_13695);
nand U14042 (N_14042,N_13418,N_13740);
or U14043 (N_14043,N_13700,N_13900);
nor U14044 (N_14044,N_13437,N_13646);
or U14045 (N_14045,N_13757,N_13839);
or U14046 (N_14046,N_13058,N_13207);
xnor U14047 (N_14047,N_13188,N_13427);
nor U14048 (N_14048,N_13417,N_13392);
nand U14049 (N_14049,N_13801,N_13777);
xor U14050 (N_14050,N_13914,N_13721);
and U14051 (N_14051,N_13764,N_13624);
xnor U14052 (N_14052,N_13743,N_13015);
and U14053 (N_14053,N_13598,N_13893);
or U14054 (N_14054,N_13729,N_13287);
or U14055 (N_14055,N_13599,N_13187);
nor U14056 (N_14056,N_13660,N_13683);
nor U14057 (N_14057,N_13480,N_13482);
xor U14058 (N_14058,N_13023,N_13694);
xnor U14059 (N_14059,N_13069,N_13426);
nor U14060 (N_14060,N_13925,N_13994);
xor U14061 (N_14061,N_13014,N_13547);
and U14062 (N_14062,N_13711,N_13750);
nor U14063 (N_14063,N_13226,N_13463);
xnor U14064 (N_14064,N_13867,N_13552);
nand U14065 (N_14065,N_13792,N_13862);
or U14066 (N_14066,N_13855,N_13546);
nor U14067 (N_14067,N_13749,N_13785);
or U14068 (N_14068,N_13136,N_13537);
nor U14069 (N_14069,N_13024,N_13788);
xnor U14070 (N_14070,N_13555,N_13440);
nor U14071 (N_14071,N_13870,N_13583);
nor U14072 (N_14072,N_13858,N_13059);
and U14073 (N_14073,N_13513,N_13500);
and U14074 (N_14074,N_13576,N_13886);
or U14075 (N_14075,N_13214,N_13143);
or U14076 (N_14076,N_13985,N_13072);
nand U14077 (N_14077,N_13442,N_13255);
or U14078 (N_14078,N_13303,N_13123);
or U14079 (N_14079,N_13045,N_13079);
nand U14080 (N_14080,N_13860,N_13780);
nor U14081 (N_14081,N_13909,N_13974);
and U14082 (N_14082,N_13488,N_13869);
and U14083 (N_14083,N_13654,N_13250);
and U14084 (N_14084,N_13114,N_13578);
xnor U14085 (N_14085,N_13259,N_13521);
xnor U14086 (N_14086,N_13532,N_13321);
or U14087 (N_14087,N_13436,N_13413);
and U14088 (N_14088,N_13318,N_13822);
nand U14089 (N_14089,N_13610,N_13717);
and U14090 (N_14090,N_13510,N_13682);
nor U14091 (N_14091,N_13789,N_13157);
and U14092 (N_14092,N_13553,N_13728);
xor U14093 (N_14093,N_13542,N_13924);
or U14094 (N_14094,N_13489,N_13336);
nand U14095 (N_14095,N_13211,N_13629);
nor U14096 (N_14096,N_13366,N_13600);
nand U14097 (N_14097,N_13469,N_13456);
nand U14098 (N_14098,N_13410,N_13137);
nand U14099 (N_14099,N_13601,N_13774);
xnor U14100 (N_14100,N_13109,N_13233);
or U14101 (N_14101,N_13008,N_13000);
or U14102 (N_14102,N_13466,N_13222);
nor U14103 (N_14103,N_13907,N_13248);
xnor U14104 (N_14104,N_13174,N_13212);
and U14105 (N_14105,N_13086,N_13151);
xnor U14106 (N_14106,N_13702,N_13868);
or U14107 (N_14107,N_13698,N_13888);
nand U14108 (N_14108,N_13594,N_13235);
nor U14109 (N_14109,N_13081,N_13258);
and U14110 (N_14110,N_13887,N_13519);
nor U14111 (N_14111,N_13754,N_13840);
nor U14112 (N_14112,N_13285,N_13219);
or U14113 (N_14113,N_13751,N_13828);
and U14114 (N_14114,N_13882,N_13389);
xnor U14115 (N_14115,N_13429,N_13354);
or U14116 (N_14116,N_13346,N_13147);
nand U14117 (N_14117,N_13639,N_13311);
xor U14118 (N_14118,N_13390,N_13661);
nor U14119 (N_14119,N_13190,N_13380);
xnor U14120 (N_14120,N_13739,N_13644);
nand U14121 (N_14121,N_13411,N_13089);
xnor U14122 (N_14122,N_13768,N_13529);
or U14123 (N_14123,N_13567,N_13747);
and U14124 (N_14124,N_13955,N_13166);
nand U14125 (N_14125,N_13388,N_13498);
or U14126 (N_14126,N_13485,N_13913);
or U14127 (N_14127,N_13328,N_13612);
nor U14128 (N_14128,N_13505,N_13834);
nand U14129 (N_14129,N_13460,N_13405);
xor U14130 (N_14130,N_13097,N_13635);
xnor U14131 (N_14131,N_13971,N_13439);
and U14132 (N_14132,N_13675,N_13424);
or U14133 (N_14133,N_13824,N_13581);
and U14134 (N_14134,N_13001,N_13384);
or U14135 (N_14135,N_13916,N_13278);
or U14136 (N_14136,N_13904,N_13118);
xor U14137 (N_14137,N_13658,N_13310);
and U14138 (N_14138,N_13100,N_13261);
nor U14139 (N_14139,N_13181,N_13999);
nand U14140 (N_14140,N_13367,N_13078);
xnor U14141 (N_14141,N_13815,N_13674);
and U14142 (N_14142,N_13920,N_13350);
xnor U14143 (N_14143,N_13712,N_13025);
xnor U14144 (N_14144,N_13650,N_13645);
or U14145 (N_14145,N_13225,N_13351);
xor U14146 (N_14146,N_13707,N_13129);
nor U14147 (N_14147,N_13221,N_13517);
or U14148 (N_14148,N_13103,N_13813);
and U14149 (N_14149,N_13127,N_13085);
and U14150 (N_14150,N_13386,N_13782);
and U14151 (N_14151,N_13926,N_13535);
and U14152 (N_14152,N_13179,N_13525);
xnor U14153 (N_14153,N_13627,N_13334);
nor U14154 (N_14154,N_13672,N_13203);
nor U14155 (N_14155,N_13313,N_13461);
and U14156 (N_14156,N_13007,N_13575);
xor U14157 (N_14157,N_13082,N_13708);
nor U14158 (N_14158,N_13165,N_13016);
and U14159 (N_14159,N_13606,N_13308);
and U14160 (N_14160,N_13752,N_13279);
nand U14161 (N_14161,N_13964,N_13898);
nand U14162 (N_14162,N_13372,N_13856);
nor U14163 (N_14163,N_13809,N_13910);
xnor U14164 (N_14164,N_13479,N_13807);
xor U14165 (N_14165,N_13859,N_13486);
nand U14166 (N_14166,N_13538,N_13141);
xnor U14167 (N_14167,N_13951,N_13516);
and U14168 (N_14168,N_13531,N_13957);
or U14169 (N_14169,N_13395,N_13364);
nor U14170 (N_14170,N_13473,N_13229);
nor U14171 (N_14171,N_13382,N_13998);
xor U14172 (N_14172,N_13767,N_13043);
nor U14173 (N_14173,N_13560,N_13563);
and U14174 (N_14174,N_13342,N_13966);
nor U14175 (N_14175,N_13686,N_13671);
and U14176 (N_14176,N_13468,N_13787);
xor U14177 (N_14177,N_13591,N_13997);
nor U14178 (N_14178,N_13746,N_13159);
nand U14179 (N_14179,N_13154,N_13783);
nor U14180 (N_14180,N_13470,N_13573);
or U14181 (N_14181,N_13864,N_13111);
nor U14182 (N_14182,N_13087,N_13192);
or U14183 (N_14183,N_13194,N_13432);
or U14184 (N_14184,N_13160,N_13755);
nand U14185 (N_14185,N_13105,N_13611);
xnor U14186 (N_14186,N_13309,N_13851);
and U14187 (N_14187,N_13185,N_13186);
xor U14188 (N_14188,N_13294,N_13528);
and U14189 (N_14189,N_13040,N_13383);
or U14190 (N_14190,N_13202,N_13451);
xor U14191 (N_14191,N_13501,N_13170);
and U14192 (N_14192,N_13613,N_13009);
and U14193 (N_14193,N_13444,N_13067);
nand U14194 (N_14194,N_13090,N_13398);
xnor U14195 (N_14195,N_13199,N_13359);
and U14196 (N_14196,N_13450,N_13302);
and U14197 (N_14197,N_13829,N_13275);
nand U14198 (N_14198,N_13298,N_13465);
nand U14199 (N_14199,N_13282,N_13992);
nor U14200 (N_14200,N_13032,N_13565);
and U14201 (N_14201,N_13177,N_13246);
or U14202 (N_14202,N_13475,N_13935);
xor U14203 (N_14203,N_13561,N_13140);
or U14204 (N_14204,N_13134,N_13051);
and U14205 (N_14205,N_13846,N_13585);
nor U14206 (N_14206,N_13795,N_13234);
nor U14207 (N_14207,N_13317,N_13257);
nor U14208 (N_14208,N_13877,N_13520);
nor U14209 (N_14209,N_13741,N_13422);
nand U14210 (N_14210,N_13976,N_13580);
nand U14211 (N_14211,N_13987,N_13121);
xnor U14212 (N_14212,N_13980,N_13836);
or U14213 (N_14213,N_13706,N_13092);
xor U14214 (N_14214,N_13655,N_13830);
xnor U14215 (N_14215,N_13182,N_13524);
nand U14216 (N_14216,N_13270,N_13854);
nor U14217 (N_14217,N_13609,N_13290);
xor U14218 (N_14218,N_13930,N_13037);
or U14219 (N_14219,N_13831,N_13329);
or U14220 (N_14220,N_13604,N_13699);
xnor U14221 (N_14221,N_13263,N_13048);
and U14222 (N_14222,N_13738,N_13512);
xnor U14223 (N_14223,N_13802,N_13582);
or U14224 (N_14224,N_13377,N_13758);
or U14225 (N_14225,N_13133,N_13280);
xnor U14226 (N_14226,N_13175,N_13107);
nand U14227 (N_14227,N_13476,N_13430);
or U14228 (N_14228,N_13545,N_13816);
or U14229 (N_14229,N_13731,N_13713);
nor U14230 (N_14230,N_13622,N_13112);
and U14231 (N_14231,N_13288,N_13876);
nor U14232 (N_14232,N_13577,N_13215);
nand U14233 (N_14233,N_13903,N_13818);
or U14234 (N_14234,N_13863,N_13835);
and U14235 (N_14235,N_13471,N_13668);
or U14236 (N_14236,N_13419,N_13276);
nand U14237 (N_14237,N_13905,N_13673);
nand U14238 (N_14238,N_13339,N_13927);
nor U14239 (N_14239,N_13734,N_13514);
xnor U14240 (N_14240,N_13268,N_13791);
nand U14241 (N_14241,N_13393,N_13044);
nand U14242 (N_14242,N_13088,N_13231);
and U14243 (N_14243,N_13651,N_13352);
xnor U14244 (N_14244,N_13908,N_13568);
or U14245 (N_14245,N_13989,N_13369);
or U14246 (N_14246,N_13407,N_13446);
nand U14247 (N_14247,N_13333,N_13832);
nand U14248 (N_14248,N_13453,N_13838);
xor U14249 (N_14249,N_13742,N_13459);
and U14250 (N_14250,N_13643,N_13119);
nor U14251 (N_14251,N_13821,N_13195);
and U14252 (N_14252,N_13335,N_13251);
or U14253 (N_14253,N_13915,N_13361);
nor U14254 (N_14254,N_13931,N_13124);
or U14255 (N_14255,N_13628,N_13933);
and U14256 (N_14256,N_13669,N_13649);
xnor U14257 (N_14257,N_13176,N_13748);
and U14258 (N_14258,N_13245,N_13028);
and U14259 (N_14259,N_13036,N_13763);
nor U14260 (N_14260,N_13244,N_13362);
nand U14261 (N_14261,N_13569,N_13084);
xnor U14262 (N_14262,N_13979,N_13833);
or U14263 (N_14263,N_13656,N_13949);
nand U14264 (N_14264,N_13327,N_13723);
nand U14265 (N_14265,N_13968,N_13973);
nor U14266 (N_14266,N_13132,N_13047);
nand U14267 (N_14267,N_13269,N_13850);
nand U14268 (N_14268,N_13083,N_13551);
nor U14269 (N_14269,N_13070,N_13496);
xnor U14270 (N_14270,N_13066,N_13623);
xor U14271 (N_14271,N_13106,N_13183);
or U14272 (N_14272,N_13232,N_13452);
or U14273 (N_14273,N_13184,N_13098);
nand U14274 (N_14274,N_13356,N_13892);
xor U14275 (N_14275,N_13950,N_13156);
or U14276 (N_14276,N_13247,N_13928);
xor U14277 (N_14277,N_13527,N_13122);
nand U14278 (N_14278,N_13161,N_13705);
and U14279 (N_14279,N_13031,N_13472);
nor U14280 (N_14280,N_13690,N_13368);
xor U14281 (N_14281,N_13919,N_13626);
nand U14282 (N_14282,N_13875,N_13533);
or U14283 (N_14283,N_13891,N_13415);
nand U14284 (N_14284,N_13305,N_13387);
or U14285 (N_14285,N_13873,N_13138);
xnor U14286 (N_14286,N_13198,N_13434);
and U14287 (N_14287,N_13020,N_13117);
nand U14288 (N_14288,N_13588,N_13096);
and U14289 (N_14289,N_13293,N_13507);
or U14290 (N_14290,N_13556,N_13786);
nor U14291 (N_14291,N_13984,N_13074);
nor U14292 (N_14292,N_13895,N_13204);
or U14293 (N_14293,N_13213,N_13306);
nand U14294 (N_14294,N_13130,N_13068);
nand U14295 (N_14295,N_13848,N_13495);
or U14296 (N_14296,N_13331,N_13811);
nand U14297 (N_14297,N_13732,N_13227);
nor U14298 (N_14298,N_13491,N_13952);
nand U14299 (N_14299,N_13332,N_13314);
xnor U14300 (N_14300,N_13421,N_13614);
or U14301 (N_14301,N_13374,N_13618);
nor U14302 (N_14302,N_13959,N_13277);
nand U14303 (N_14303,N_13590,N_13237);
xnor U14304 (N_14304,N_13131,N_13091);
and U14305 (N_14305,N_13806,N_13400);
or U14306 (N_14306,N_13053,N_13722);
nor U14307 (N_14307,N_13477,N_13243);
nor U14308 (N_14308,N_13689,N_13771);
nor U14309 (N_14309,N_13353,N_13911);
xor U14310 (N_14310,N_13046,N_13381);
nor U14311 (N_14311,N_13800,N_13071);
nand U14312 (N_14312,N_13616,N_13544);
and U14313 (N_14313,N_13664,N_13633);
nor U14314 (N_14314,N_13050,N_13206);
or U14315 (N_14315,N_13249,N_13358);
and U14316 (N_14316,N_13104,N_13724);
or U14317 (N_14317,N_13572,N_13936);
or U14318 (N_14318,N_13338,N_13522);
nand U14319 (N_14319,N_13173,N_13049);
nand U14320 (N_14320,N_13587,N_13385);
nand U14321 (N_14321,N_13200,N_13093);
nand U14322 (N_14322,N_13993,N_13820);
or U14323 (N_14323,N_13283,N_13790);
xnor U14324 (N_14324,N_13265,N_13760);
nor U14325 (N_14325,N_13146,N_13005);
xnor U14326 (N_14326,N_13433,N_13497);
and U14327 (N_14327,N_13586,N_13158);
nor U14328 (N_14328,N_13281,N_13943);
nand U14329 (N_14329,N_13125,N_13896);
nand U14330 (N_14330,N_13013,N_13615);
or U14331 (N_14331,N_13798,N_13172);
xnor U14332 (N_14332,N_13564,N_13355);
xnor U14333 (N_14333,N_13536,N_13220);
and U14334 (N_14334,N_13487,N_13592);
nor U14335 (N_14335,N_13378,N_13938);
nand U14336 (N_14336,N_13484,N_13953);
xnor U14337 (N_14337,N_13144,N_13197);
and U14338 (N_14338,N_13523,N_13063);
nor U14339 (N_14339,N_13230,N_13735);
or U14340 (N_14340,N_13733,N_13778);
and U14341 (N_14341,N_13812,N_13167);
nor U14342 (N_14342,N_13554,N_13145);
and U14343 (N_14343,N_13946,N_13504);
xnor U14344 (N_14344,N_13697,N_13120);
nor U14345 (N_14345,N_13435,N_13503);
xnor U14346 (N_14346,N_13637,N_13150);
nand U14347 (N_14347,N_13765,N_13295);
xor U14348 (N_14348,N_13970,N_13944);
or U14349 (N_14349,N_13394,N_13670);
xor U14350 (N_14350,N_13320,N_13360);
nor U14351 (N_14351,N_13819,N_13019);
nor U14352 (N_14352,N_13937,N_13940);
or U14353 (N_14353,N_13978,N_13737);
or U14354 (N_14354,N_13155,N_13657);
nand U14355 (N_14355,N_13906,N_13681);
nor U14356 (N_14356,N_13678,N_13912);
or U14357 (N_14357,N_13954,N_13776);
nand U14358 (N_14358,N_13217,N_13704);
or U14359 (N_14359,N_13017,N_13990);
or U14360 (N_14360,N_13710,N_13559);
and U14361 (N_14361,N_13201,N_13960);
nand U14362 (N_14362,N_13866,N_13324);
and U14363 (N_14363,N_13301,N_13718);
nand U14364 (N_14364,N_13267,N_13163);
or U14365 (N_14365,N_13589,N_13630);
nor U14366 (N_14366,N_13271,N_13416);
nor U14367 (N_14367,N_13865,N_13810);
and U14368 (N_14368,N_13223,N_13030);
xor U14369 (N_14369,N_13494,N_13077);
or U14370 (N_14370,N_13880,N_13399);
or U14371 (N_14371,N_13148,N_13558);
xnor U14372 (N_14372,N_13961,N_13852);
nand U14373 (N_14373,N_13402,N_13945);
xor U14374 (N_14374,N_13779,N_13391);
xor U14375 (N_14375,N_13431,N_13289);
and U14376 (N_14376,N_13539,N_13344);
and U14377 (N_14377,N_13345,N_13784);
nand U14378 (N_14378,N_13052,N_13481);
nor U14379 (N_14379,N_13341,N_13942);
xnor U14380 (N_14380,N_13502,N_13483);
or U14381 (N_14381,N_13376,N_13679);
nor U14382 (N_14382,N_13115,N_13841);
and U14383 (N_14383,N_13680,N_13224);
or U14384 (N_14384,N_13793,N_13315);
and U14385 (N_14385,N_13152,N_13493);
nor U14386 (N_14386,N_13803,N_13035);
or U14387 (N_14387,N_13593,N_13241);
and U14388 (N_14388,N_13404,N_13894);
nand U14389 (N_14389,N_13753,N_13844);
or U14390 (N_14390,N_13595,N_13142);
or U14391 (N_14391,N_13447,N_13348);
and U14392 (N_14392,N_13814,N_13843);
nor U14393 (N_14393,N_13995,N_13284);
nor U14394 (N_14394,N_13164,N_13191);
nand U14395 (N_14395,N_13823,N_13180);
nor U14396 (N_14396,N_13897,N_13423);
or U14397 (N_14397,N_13991,N_13621);
or U14398 (N_14398,N_13871,N_13884);
nor U14399 (N_14399,N_13526,N_13441);
nor U14400 (N_14400,N_13730,N_13947);
xor U14401 (N_14401,N_13981,N_13330);
and U14402 (N_14402,N_13062,N_13126);
nand U14403 (N_14403,N_13584,N_13566);
and U14404 (N_14404,N_13323,N_13770);
nor U14405 (N_14405,N_13057,N_13260);
and U14406 (N_14406,N_13861,N_13027);
xnor U14407 (N_14407,N_13041,N_13881);
or U14408 (N_14408,N_13638,N_13756);
xnor U14409 (N_14409,N_13291,N_13781);
nor U14410 (N_14410,N_13703,N_13292);
xor U14411 (N_14411,N_13605,N_13641);
nor U14412 (N_14412,N_13509,N_13804);
nor U14413 (N_14413,N_13726,N_13038);
xor U14414 (N_14414,N_13548,N_13455);
and U14415 (N_14415,N_13508,N_13922);
and U14416 (N_14416,N_13939,N_13363);
xor U14417 (N_14417,N_13518,N_13026);
nor U14418 (N_14418,N_13766,N_13659);
or U14419 (N_14419,N_13033,N_13205);
or U14420 (N_14420,N_13099,N_13196);
nand U14421 (N_14421,N_13901,N_13759);
nor U14422 (N_14422,N_13492,N_13632);
and U14423 (N_14423,N_13108,N_13006);
or U14424 (N_14424,N_13357,N_13011);
nor U14425 (N_14425,N_13715,N_13653);
or U14426 (N_14426,N_13499,N_13454);
nor U14427 (N_14427,N_13879,N_13061);
xnor U14428 (N_14428,N_13236,N_13640);
xnor U14429 (N_14429,N_13462,N_13808);
nand U14430 (N_14430,N_13506,N_13921);
xor U14431 (N_14431,N_13720,N_13319);
or U14432 (N_14432,N_13665,N_13003);
nand U14433 (N_14433,N_13307,N_13401);
nand U14434 (N_14434,N_13448,N_13725);
and U14435 (N_14435,N_13296,N_13264);
nor U14436 (N_14436,N_13958,N_13169);
nand U14437 (N_14437,N_13932,N_13666);
xnor U14438 (N_14438,N_13714,N_13825);
nor U14439 (N_14439,N_13744,N_13242);
nor U14440 (N_14440,N_13691,N_13648);
or U14441 (N_14441,N_13340,N_13256);
nand U14442 (N_14442,N_13969,N_13425);
or U14443 (N_14443,N_13312,N_13065);
and U14444 (N_14444,N_13370,N_13010);
xnor U14445 (N_14445,N_13857,N_13769);
xor U14446 (N_14446,N_13550,N_13826);
or U14447 (N_14447,N_13445,N_13139);
nand U14448 (N_14448,N_13975,N_13530);
nand U14449 (N_14449,N_13193,N_13012);
nand U14450 (N_14450,N_13608,N_13620);
and U14451 (N_14451,N_13983,N_13474);
or U14452 (N_14452,N_13397,N_13667);
or U14453 (N_14453,N_13412,N_13075);
xnor U14454 (N_14454,N_13889,N_13874);
or U14455 (N_14455,N_13543,N_13414);
or U14456 (N_14456,N_13428,N_13326);
or U14457 (N_14457,N_13076,N_13002);
or U14458 (N_14458,N_13677,N_13004);
nor U14459 (N_14459,N_13962,N_13687);
nand U14460 (N_14460,N_13701,N_13948);
or U14461 (N_14461,N_13977,N_13064);
nor U14462 (N_14462,N_13596,N_13467);
nor U14463 (N_14463,N_13696,N_13056);
and U14464 (N_14464,N_13406,N_13986);
nor U14465 (N_14465,N_13273,N_13642);
xnor U14466 (N_14466,N_13773,N_13272);
and U14467 (N_14467,N_13210,N_13647);
xor U14468 (N_14468,N_13373,N_13055);
nor U14469 (N_14469,N_13570,N_13403);
nand U14470 (N_14470,N_13420,N_13652);
or U14471 (N_14471,N_13443,N_13018);
and U14472 (N_14472,N_13727,N_13101);
nor U14473 (N_14473,N_13662,N_13365);
nor U14474 (N_14474,N_13885,N_13396);
and U14475 (N_14475,N_13963,N_13409);
nor U14476 (N_14476,N_13692,N_13464);
xnor U14477 (N_14477,N_13685,N_13511);
xnor U14478 (N_14478,N_13772,N_13300);
or U14479 (N_14479,N_13149,N_13762);
xnor U14480 (N_14480,N_13034,N_13805);
nand U14481 (N_14481,N_13796,N_13371);
or U14482 (N_14482,N_13171,N_13557);
or U14483 (N_14483,N_13189,N_13988);
nand U14484 (N_14484,N_13684,N_13934);
nor U14485 (N_14485,N_13095,N_13540);
nand U14486 (N_14486,N_13745,N_13153);
xnor U14487 (N_14487,N_13716,N_13775);
xnor U14488 (N_14488,N_13965,N_13274);
xnor U14489 (N_14489,N_13794,N_13872);
or U14490 (N_14490,N_13817,N_13878);
or U14491 (N_14491,N_13379,N_13899);
or U14492 (N_14492,N_13619,N_13022);
or U14493 (N_14493,N_13827,N_13347);
xnor U14494 (N_14494,N_13286,N_13972);
xor U14495 (N_14495,N_13438,N_13039);
xnor U14496 (N_14496,N_13490,N_13060);
or U14497 (N_14497,N_13890,N_13549);
or U14498 (N_14498,N_13709,N_13571);
and U14499 (N_14499,N_13408,N_13515);
or U14500 (N_14500,N_13902,N_13569);
or U14501 (N_14501,N_13806,N_13906);
and U14502 (N_14502,N_13928,N_13730);
and U14503 (N_14503,N_13968,N_13945);
nand U14504 (N_14504,N_13206,N_13949);
xnor U14505 (N_14505,N_13854,N_13885);
or U14506 (N_14506,N_13069,N_13460);
or U14507 (N_14507,N_13052,N_13255);
nor U14508 (N_14508,N_13666,N_13220);
xnor U14509 (N_14509,N_13241,N_13239);
or U14510 (N_14510,N_13420,N_13882);
and U14511 (N_14511,N_13407,N_13543);
nand U14512 (N_14512,N_13102,N_13922);
and U14513 (N_14513,N_13466,N_13978);
or U14514 (N_14514,N_13321,N_13196);
and U14515 (N_14515,N_13287,N_13371);
nor U14516 (N_14516,N_13495,N_13983);
and U14517 (N_14517,N_13433,N_13795);
and U14518 (N_14518,N_13799,N_13478);
and U14519 (N_14519,N_13189,N_13207);
and U14520 (N_14520,N_13533,N_13878);
xor U14521 (N_14521,N_13885,N_13912);
and U14522 (N_14522,N_13587,N_13592);
and U14523 (N_14523,N_13640,N_13149);
nand U14524 (N_14524,N_13172,N_13882);
nand U14525 (N_14525,N_13685,N_13617);
nand U14526 (N_14526,N_13056,N_13690);
or U14527 (N_14527,N_13677,N_13389);
nand U14528 (N_14528,N_13873,N_13455);
nor U14529 (N_14529,N_13354,N_13211);
nand U14530 (N_14530,N_13226,N_13693);
nand U14531 (N_14531,N_13410,N_13918);
nor U14532 (N_14532,N_13157,N_13277);
nor U14533 (N_14533,N_13312,N_13986);
or U14534 (N_14534,N_13648,N_13892);
nand U14535 (N_14535,N_13040,N_13878);
nor U14536 (N_14536,N_13823,N_13558);
xor U14537 (N_14537,N_13813,N_13965);
nor U14538 (N_14538,N_13438,N_13312);
nand U14539 (N_14539,N_13175,N_13237);
or U14540 (N_14540,N_13147,N_13587);
nand U14541 (N_14541,N_13444,N_13310);
xnor U14542 (N_14542,N_13743,N_13585);
or U14543 (N_14543,N_13265,N_13387);
xor U14544 (N_14544,N_13160,N_13279);
nand U14545 (N_14545,N_13528,N_13725);
or U14546 (N_14546,N_13274,N_13972);
and U14547 (N_14547,N_13544,N_13881);
or U14548 (N_14548,N_13972,N_13835);
or U14549 (N_14549,N_13754,N_13869);
or U14550 (N_14550,N_13142,N_13466);
xnor U14551 (N_14551,N_13378,N_13088);
or U14552 (N_14552,N_13245,N_13552);
xor U14553 (N_14553,N_13435,N_13810);
xnor U14554 (N_14554,N_13266,N_13092);
nor U14555 (N_14555,N_13508,N_13883);
xnor U14556 (N_14556,N_13162,N_13295);
xnor U14557 (N_14557,N_13252,N_13006);
or U14558 (N_14558,N_13595,N_13818);
and U14559 (N_14559,N_13168,N_13851);
xor U14560 (N_14560,N_13906,N_13757);
or U14561 (N_14561,N_13240,N_13196);
and U14562 (N_14562,N_13042,N_13375);
nor U14563 (N_14563,N_13786,N_13995);
nor U14564 (N_14564,N_13848,N_13941);
or U14565 (N_14565,N_13373,N_13534);
xnor U14566 (N_14566,N_13842,N_13964);
xnor U14567 (N_14567,N_13470,N_13495);
or U14568 (N_14568,N_13706,N_13360);
or U14569 (N_14569,N_13707,N_13325);
and U14570 (N_14570,N_13154,N_13241);
or U14571 (N_14571,N_13932,N_13966);
nand U14572 (N_14572,N_13116,N_13108);
or U14573 (N_14573,N_13989,N_13585);
nand U14574 (N_14574,N_13354,N_13303);
or U14575 (N_14575,N_13657,N_13652);
nand U14576 (N_14576,N_13904,N_13535);
and U14577 (N_14577,N_13228,N_13850);
or U14578 (N_14578,N_13436,N_13555);
nor U14579 (N_14579,N_13732,N_13005);
xor U14580 (N_14580,N_13871,N_13966);
nor U14581 (N_14581,N_13626,N_13937);
nor U14582 (N_14582,N_13053,N_13403);
nor U14583 (N_14583,N_13355,N_13474);
xor U14584 (N_14584,N_13844,N_13929);
and U14585 (N_14585,N_13995,N_13864);
or U14586 (N_14586,N_13509,N_13727);
nand U14587 (N_14587,N_13262,N_13000);
and U14588 (N_14588,N_13428,N_13144);
and U14589 (N_14589,N_13501,N_13939);
and U14590 (N_14590,N_13726,N_13418);
nand U14591 (N_14591,N_13109,N_13102);
or U14592 (N_14592,N_13481,N_13496);
and U14593 (N_14593,N_13739,N_13183);
and U14594 (N_14594,N_13773,N_13173);
xor U14595 (N_14595,N_13960,N_13647);
nand U14596 (N_14596,N_13945,N_13536);
or U14597 (N_14597,N_13121,N_13569);
and U14598 (N_14598,N_13332,N_13771);
nand U14599 (N_14599,N_13149,N_13903);
or U14600 (N_14600,N_13397,N_13815);
xor U14601 (N_14601,N_13573,N_13652);
nor U14602 (N_14602,N_13573,N_13581);
xor U14603 (N_14603,N_13778,N_13672);
xnor U14604 (N_14604,N_13093,N_13216);
nor U14605 (N_14605,N_13323,N_13786);
nand U14606 (N_14606,N_13074,N_13847);
or U14607 (N_14607,N_13900,N_13447);
and U14608 (N_14608,N_13369,N_13077);
xnor U14609 (N_14609,N_13202,N_13483);
and U14610 (N_14610,N_13170,N_13915);
xor U14611 (N_14611,N_13404,N_13403);
nand U14612 (N_14612,N_13179,N_13560);
xnor U14613 (N_14613,N_13982,N_13949);
and U14614 (N_14614,N_13775,N_13729);
nor U14615 (N_14615,N_13547,N_13487);
and U14616 (N_14616,N_13674,N_13170);
xor U14617 (N_14617,N_13775,N_13064);
nor U14618 (N_14618,N_13672,N_13639);
nand U14619 (N_14619,N_13329,N_13814);
nand U14620 (N_14620,N_13960,N_13641);
nand U14621 (N_14621,N_13297,N_13041);
nor U14622 (N_14622,N_13796,N_13573);
or U14623 (N_14623,N_13999,N_13173);
or U14624 (N_14624,N_13928,N_13002);
and U14625 (N_14625,N_13295,N_13890);
nand U14626 (N_14626,N_13364,N_13600);
nand U14627 (N_14627,N_13660,N_13166);
and U14628 (N_14628,N_13802,N_13247);
nor U14629 (N_14629,N_13720,N_13042);
nand U14630 (N_14630,N_13626,N_13270);
xnor U14631 (N_14631,N_13126,N_13579);
xor U14632 (N_14632,N_13715,N_13012);
and U14633 (N_14633,N_13693,N_13240);
xor U14634 (N_14634,N_13444,N_13565);
nand U14635 (N_14635,N_13322,N_13790);
or U14636 (N_14636,N_13165,N_13265);
or U14637 (N_14637,N_13161,N_13236);
and U14638 (N_14638,N_13009,N_13403);
or U14639 (N_14639,N_13698,N_13145);
or U14640 (N_14640,N_13279,N_13583);
xor U14641 (N_14641,N_13795,N_13382);
and U14642 (N_14642,N_13820,N_13990);
or U14643 (N_14643,N_13696,N_13686);
nor U14644 (N_14644,N_13768,N_13482);
and U14645 (N_14645,N_13756,N_13612);
nand U14646 (N_14646,N_13852,N_13111);
xor U14647 (N_14647,N_13009,N_13600);
xnor U14648 (N_14648,N_13293,N_13411);
and U14649 (N_14649,N_13830,N_13715);
xnor U14650 (N_14650,N_13984,N_13663);
or U14651 (N_14651,N_13032,N_13253);
nand U14652 (N_14652,N_13600,N_13427);
xor U14653 (N_14653,N_13194,N_13378);
and U14654 (N_14654,N_13393,N_13740);
nand U14655 (N_14655,N_13223,N_13638);
nor U14656 (N_14656,N_13649,N_13292);
nor U14657 (N_14657,N_13485,N_13342);
xnor U14658 (N_14658,N_13702,N_13663);
nor U14659 (N_14659,N_13263,N_13447);
or U14660 (N_14660,N_13276,N_13848);
nand U14661 (N_14661,N_13518,N_13070);
nand U14662 (N_14662,N_13075,N_13081);
nor U14663 (N_14663,N_13941,N_13589);
and U14664 (N_14664,N_13301,N_13878);
and U14665 (N_14665,N_13067,N_13511);
xnor U14666 (N_14666,N_13359,N_13879);
nor U14667 (N_14667,N_13687,N_13286);
xnor U14668 (N_14668,N_13426,N_13421);
xnor U14669 (N_14669,N_13767,N_13592);
xor U14670 (N_14670,N_13208,N_13164);
nor U14671 (N_14671,N_13627,N_13271);
or U14672 (N_14672,N_13397,N_13553);
nor U14673 (N_14673,N_13932,N_13885);
nor U14674 (N_14674,N_13240,N_13995);
and U14675 (N_14675,N_13643,N_13371);
xor U14676 (N_14676,N_13017,N_13773);
nand U14677 (N_14677,N_13701,N_13305);
or U14678 (N_14678,N_13284,N_13318);
and U14679 (N_14679,N_13472,N_13961);
nand U14680 (N_14680,N_13576,N_13819);
nor U14681 (N_14681,N_13376,N_13464);
nor U14682 (N_14682,N_13766,N_13141);
nor U14683 (N_14683,N_13870,N_13880);
xor U14684 (N_14684,N_13039,N_13499);
xor U14685 (N_14685,N_13079,N_13595);
nor U14686 (N_14686,N_13346,N_13688);
and U14687 (N_14687,N_13924,N_13300);
xor U14688 (N_14688,N_13972,N_13903);
nand U14689 (N_14689,N_13969,N_13740);
nor U14690 (N_14690,N_13875,N_13225);
xor U14691 (N_14691,N_13417,N_13247);
nor U14692 (N_14692,N_13482,N_13244);
nor U14693 (N_14693,N_13999,N_13790);
nand U14694 (N_14694,N_13803,N_13057);
nor U14695 (N_14695,N_13545,N_13747);
nand U14696 (N_14696,N_13334,N_13863);
and U14697 (N_14697,N_13082,N_13844);
nor U14698 (N_14698,N_13716,N_13486);
nor U14699 (N_14699,N_13403,N_13659);
and U14700 (N_14700,N_13872,N_13422);
and U14701 (N_14701,N_13452,N_13029);
or U14702 (N_14702,N_13989,N_13401);
and U14703 (N_14703,N_13846,N_13047);
or U14704 (N_14704,N_13364,N_13991);
nor U14705 (N_14705,N_13242,N_13606);
and U14706 (N_14706,N_13819,N_13785);
nand U14707 (N_14707,N_13148,N_13207);
nand U14708 (N_14708,N_13546,N_13553);
and U14709 (N_14709,N_13784,N_13775);
or U14710 (N_14710,N_13574,N_13353);
and U14711 (N_14711,N_13521,N_13118);
xnor U14712 (N_14712,N_13754,N_13573);
xnor U14713 (N_14713,N_13123,N_13600);
and U14714 (N_14714,N_13059,N_13958);
or U14715 (N_14715,N_13811,N_13474);
or U14716 (N_14716,N_13991,N_13920);
and U14717 (N_14717,N_13273,N_13900);
nand U14718 (N_14718,N_13049,N_13275);
or U14719 (N_14719,N_13263,N_13053);
or U14720 (N_14720,N_13597,N_13437);
and U14721 (N_14721,N_13713,N_13248);
xor U14722 (N_14722,N_13128,N_13748);
nand U14723 (N_14723,N_13478,N_13643);
and U14724 (N_14724,N_13055,N_13202);
and U14725 (N_14725,N_13191,N_13657);
nor U14726 (N_14726,N_13764,N_13714);
or U14727 (N_14727,N_13271,N_13551);
xnor U14728 (N_14728,N_13508,N_13724);
and U14729 (N_14729,N_13701,N_13821);
nand U14730 (N_14730,N_13993,N_13909);
or U14731 (N_14731,N_13282,N_13563);
nand U14732 (N_14732,N_13821,N_13091);
xnor U14733 (N_14733,N_13748,N_13204);
nor U14734 (N_14734,N_13659,N_13931);
nor U14735 (N_14735,N_13416,N_13034);
xor U14736 (N_14736,N_13812,N_13608);
xor U14737 (N_14737,N_13661,N_13816);
nand U14738 (N_14738,N_13907,N_13780);
or U14739 (N_14739,N_13316,N_13201);
xor U14740 (N_14740,N_13217,N_13799);
and U14741 (N_14741,N_13482,N_13765);
nor U14742 (N_14742,N_13559,N_13057);
nand U14743 (N_14743,N_13786,N_13284);
nand U14744 (N_14744,N_13231,N_13814);
xnor U14745 (N_14745,N_13025,N_13766);
xnor U14746 (N_14746,N_13387,N_13552);
and U14747 (N_14747,N_13247,N_13286);
nand U14748 (N_14748,N_13876,N_13106);
nor U14749 (N_14749,N_13852,N_13607);
or U14750 (N_14750,N_13799,N_13641);
nand U14751 (N_14751,N_13214,N_13595);
xnor U14752 (N_14752,N_13680,N_13306);
and U14753 (N_14753,N_13412,N_13974);
xnor U14754 (N_14754,N_13320,N_13977);
and U14755 (N_14755,N_13831,N_13962);
and U14756 (N_14756,N_13501,N_13575);
or U14757 (N_14757,N_13329,N_13680);
and U14758 (N_14758,N_13369,N_13056);
xnor U14759 (N_14759,N_13073,N_13077);
or U14760 (N_14760,N_13009,N_13646);
and U14761 (N_14761,N_13217,N_13555);
nor U14762 (N_14762,N_13533,N_13064);
and U14763 (N_14763,N_13784,N_13135);
and U14764 (N_14764,N_13331,N_13513);
nand U14765 (N_14765,N_13427,N_13562);
xor U14766 (N_14766,N_13967,N_13133);
nor U14767 (N_14767,N_13612,N_13752);
xor U14768 (N_14768,N_13418,N_13777);
or U14769 (N_14769,N_13812,N_13133);
and U14770 (N_14770,N_13748,N_13658);
nor U14771 (N_14771,N_13653,N_13251);
nor U14772 (N_14772,N_13123,N_13698);
and U14773 (N_14773,N_13772,N_13507);
and U14774 (N_14774,N_13843,N_13011);
and U14775 (N_14775,N_13773,N_13776);
and U14776 (N_14776,N_13360,N_13685);
nor U14777 (N_14777,N_13443,N_13577);
or U14778 (N_14778,N_13170,N_13035);
xnor U14779 (N_14779,N_13867,N_13639);
nor U14780 (N_14780,N_13282,N_13152);
nand U14781 (N_14781,N_13278,N_13047);
xnor U14782 (N_14782,N_13582,N_13958);
or U14783 (N_14783,N_13932,N_13802);
and U14784 (N_14784,N_13158,N_13468);
nand U14785 (N_14785,N_13040,N_13882);
nor U14786 (N_14786,N_13681,N_13195);
or U14787 (N_14787,N_13953,N_13403);
nand U14788 (N_14788,N_13472,N_13906);
nand U14789 (N_14789,N_13420,N_13702);
and U14790 (N_14790,N_13044,N_13845);
nor U14791 (N_14791,N_13884,N_13621);
xnor U14792 (N_14792,N_13189,N_13060);
and U14793 (N_14793,N_13978,N_13017);
nand U14794 (N_14794,N_13004,N_13174);
nand U14795 (N_14795,N_13556,N_13638);
nand U14796 (N_14796,N_13624,N_13010);
xnor U14797 (N_14797,N_13317,N_13343);
or U14798 (N_14798,N_13862,N_13916);
nand U14799 (N_14799,N_13041,N_13034);
or U14800 (N_14800,N_13965,N_13716);
xor U14801 (N_14801,N_13780,N_13369);
xor U14802 (N_14802,N_13086,N_13903);
xor U14803 (N_14803,N_13731,N_13966);
nor U14804 (N_14804,N_13046,N_13687);
and U14805 (N_14805,N_13989,N_13901);
or U14806 (N_14806,N_13285,N_13794);
nor U14807 (N_14807,N_13262,N_13153);
and U14808 (N_14808,N_13030,N_13137);
nor U14809 (N_14809,N_13709,N_13796);
or U14810 (N_14810,N_13120,N_13602);
nor U14811 (N_14811,N_13559,N_13690);
xor U14812 (N_14812,N_13384,N_13033);
xnor U14813 (N_14813,N_13919,N_13999);
xnor U14814 (N_14814,N_13147,N_13648);
or U14815 (N_14815,N_13649,N_13393);
nor U14816 (N_14816,N_13149,N_13185);
xor U14817 (N_14817,N_13046,N_13026);
or U14818 (N_14818,N_13022,N_13506);
nand U14819 (N_14819,N_13661,N_13437);
xor U14820 (N_14820,N_13257,N_13565);
and U14821 (N_14821,N_13447,N_13149);
or U14822 (N_14822,N_13559,N_13818);
nor U14823 (N_14823,N_13569,N_13600);
or U14824 (N_14824,N_13794,N_13351);
and U14825 (N_14825,N_13130,N_13695);
xnor U14826 (N_14826,N_13287,N_13579);
or U14827 (N_14827,N_13877,N_13024);
nand U14828 (N_14828,N_13491,N_13291);
and U14829 (N_14829,N_13751,N_13561);
nor U14830 (N_14830,N_13383,N_13340);
nor U14831 (N_14831,N_13557,N_13475);
or U14832 (N_14832,N_13501,N_13956);
xor U14833 (N_14833,N_13802,N_13450);
nand U14834 (N_14834,N_13574,N_13516);
nor U14835 (N_14835,N_13166,N_13729);
nand U14836 (N_14836,N_13006,N_13999);
xnor U14837 (N_14837,N_13343,N_13348);
xnor U14838 (N_14838,N_13790,N_13206);
and U14839 (N_14839,N_13810,N_13679);
nor U14840 (N_14840,N_13431,N_13752);
and U14841 (N_14841,N_13052,N_13576);
nand U14842 (N_14842,N_13715,N_13738);
nand U14843 (N_14843,N_13090,N_13221);
nor U14844 (N_14844,N_13482,N_13350);
or U14845 (N_14845,N_13031,N_13881);
nor U14846 (N_14846,N_13897,N_13065);
nand U14847 (N_14847,N_13078,N_13832);
nor U14848 (N_14848,N_13786,N_13228);
and U14849 (N_14849,N_13673,N_13109);
and U14850 (N_14850,N_13594,N_13530);
or U14851 (N_14851,N_13520,N_13945);
nand U14852 (N_14852,N_13424,N_13248);
and U14853 (N_14853,N_13696,N_13346);
or U14854 (N_14854,N_13936,N_13003);
or U14855 (N_14855,N_13514,N_13036);
or U14856 (N_14856,N_13598,N_13995);
xnor U14857 (N_14857,N_13216,N_13877);
or U14858 (N_14858,N_13614,N_13095);
or U14859 (N_14859,N_13404,N_13180);
and U14860 (N_14860,N_13521,N_13052);
nand U14861 (N_14861,N_13456,N_13844);
nor U14862 (N_14862,N_13071,N_13283);
nor U14863 (N_14863,N_13061,N_13389);
and U14864 (N_14864,N_13664,N_13580);
and U14865 (N_14865,N_13394,N_13510);
nor U14866 (N_14866,N_13603,N_13980);
or U14867 (N_14867,N_13263,N_13399);
nor U14868 (N_14868,N_13842,N_13201);
or U14869 (N_14869,N_13773,N_13802);
xnor U14870 (N_14870,N_13476,N_13334);
xnor U14871 (N_14871,N_13246,N_13850);
or U14872 (N_14872,N_13318,N_13826);
nor U14873 (N_14873,N_13564,N_13234);
and U14874 (N_14874,N_13026,N_13588);
nor U14875 (N_14875,N_13852,N_13000);
and U14876 (N_14876,N_13086,N_13861);
and U14877 (N_14877,N_13315,N_13294);
or U14878 (N_14878,N_13294,N_13093);
nor U14879 (N_14879,N_13210,N_13202);
or U14880 (N_14880,N_13151,N_13165);
nor U14881 (N_14881,N_13801,N_13619);
or U14882 (N_14882,N_13182,N_13419);
or U14883 (N_14883,N_13797,N_13107);
or U14884 (N_14884,N_13335,N_13984);
nand U14885 (N_14885,N_13000,N_13476);
or U14886 (N_14886,N_13692,N_13560);
and U14887 (N_14887,N_13265,N_13095);
nand U14888 (N_14888,N_13761,N_13342);
and U14889 (N_14889,N_13174,N_13068);
nand U14890 (N_14890,N_13147,N_13369);
xnor U14891 (N_14891,N_13990,N_13375);
or U14892 (N_14892,N_13878,N_13677);
nor U14893 (N_14893,N_13106,N_13036);
or U14894 (N_14894,N_13720,N_13674);
and U14895 (N_14895,N_13969,N_13530);
xor U14896 (N_14896,N_13902,N_13657);
and U14897 (N_14897,N_13992,N_13152);
nor U14898 (N_14898,N_13478,N_13559);
nor U14899 (N_14899,N_13683,N_13261);
and U14900 (N_14900,N_13316,N_13662);
or U14901 (N_14901,N_13276,N_13475);
nor U14902 (N_14902,N_13755,N_13248);
or U14903 (N_14903,N_13548,N_13073);
xnor U14904 (N_14904,N_13436,N_13767);
or U14905 (N_14905,N_13812,N_13298);
nor U14906 (N_14906,N_13171,N_13572);
xor U14907 (N_14907,N_13239,N_13152);
nand U14908 (N_14908,N_13116,N_13704);
nand U14909 (N_14909,N_13568,N_13087);
nor U14910 (N_14910,N_13855,N_13153);
and U14911 (N_14911,N_13250,N_13191);
nand U14912 (N_14912,N_13806,N_13797);
or U14913 (N_14913,N_13200,N_13567);
nand U14914 (N_14914,N_13885,N_13809);
nor U14915 (N_14915,N_13832,N_13982);
nand U14916 (N_14916,N_13567,N_13706);
nor U14917 (N_14917,N_13755,N_13536);
or U14918 (N_14918,N_13290,N_13349);
nor U14919 (N_14919,N_13924,N_13404);
or U14920 (N_14920,N_13014,N_13466);
and U14921 (N_14921,N_13497,N_13152);
and U14922 (N_14922,N_13029,N_13423);
or U14923 (N_14923,N_13344,N_13334);
nor U14924 (N_14924,N_13982,N_13109);
nand U14925 (N_14925,N_13432,N_13029);
nor U14926 (N_14926,N_13980,N_13843);
xor U14927 (N_14927,N_13583,N_13837);
or U14928 (N_14928,N_13180,N_13552);
xnor U14929 (N_14929,N_13730,N_13006);
or U14930 (N_14930,N_13509,N_13726);
and U14931 (N_14931,N_13645,N_13814);
nand U14932 (N_14932,N_13133,N_13403);
and U14933 (N_14933,N_13467,N_13201);
nor U14934 (N_14934,N_13842,N_13828);
nand U14935 (N_14935,N_13999,N_13857);
nand U14936 (N_14936,N_13118,N_13566);
nor U14937 (N_14937,N_13303,N_13232);
nand U14938 (N_14938,N_13477,N_13442);
and U14939 (N_14939,N_13604,N_13166);
nor U14940 (N_14940,N_13222,N_13339);
xor U14941 (N_14941,N_13288,N_13551);
nor U14942 (N_14942,N_13316,N_13135);
nand U14943 (N_14943,N_13951,N_13561);
nor U14944 (N_14944,N_13595,N_13111);
and U14945 (N_14945,N_13453,N_13821);
and U14946 (N_14946,N_13662,N_13359);
nor U14947 (N_14947,N_13454,N_13796);
nor U14948 (N_14948,N_13648,N_13142);
or U14949 (N_14949,N_13236,N_13187);
or U14950 (N_14950,N_13458,N_13696);
nor U14951 (N_14951,N_13170,N_13469);
nor U14952 (N_14952,N_13532,N_13037);
or U14953 (N_14953,N_13372,N_13667);
nor U14954 (N_14954,N_13718,N_13114);
and U14955 (N_14955,N_13023,N_13233);
xnor U14956 (N_14956,N_13124,N_13173);
nor U14957 (N_14957,N_13209,N_13542);
xnor U14958 (N_14958,N_13820,N_13605);
xor U14959 (N_14959,N_13773,N_13246);
nor U14960 (N_14960,N_13207,N_13619);
or U14961 (N_14961,N_13567,N_13039);
nand U14962 (N_14962,N_13581,N_13480);
or U14963 (N_14963,N_13154,N_13681);
nand U14964 (N_14964,N_13181,N_13786);
nor U14965 (N_14965,N_13809,N_13460);
xor U14966 (N_14966,N_13009,N_13846);
nor U14967 (N_14967,N_13719,N_13350);
xor U14968 (N_14968,N_13032,N_13210);
and U14969 (N_14969,N_13046,N_13129);
xor U14970 (N_14970,N_13140,N_13496);
nor U14971 (N_14971,N_13621,N_13241);
and U14972 (N_14972,N_13490,N_13007);
xor U14973 (N_14973,N_13325,N_13035);
xor U14974 (N_14974,N_13005,N_13331);
or U14975 (N_14975,N_13480,N_13010);
or U14976 (N_14976,N_13830,N_13270);
xor U14977 (N_14977,N_13938,N_13824);
and U14978 (N_14978,N_13929,N_13750);
nor U14979 (N_14979,N_13681,N_13645);
nor U14980 (N_14980,N_13033,N_13178);
nand U14981 (N_14981,N_13056,N_13019);
and U14982 (N_14982,N_13413,N_13428);
nor U14983 (N_14983,N_13109,N_13008);
or U14984 (N_14984,N_13260,N_13049);
nand U14985 (N_14985,N_13037,N_13042);
or U14986 (N_14986,N_13999,N_13527);
nand U14987 (N_14987,N_13355,N_13284);
xor U14988 (N_14988,N_13732,N_13773);
or U14989 (N_14989,N_13832,N_13267);
and U14990 (N_14990,N_13537,N_13382);
or U14991 (N_14991,N_13605,N_13240);
nor U14992 (N_14992,N_13665,N_13685);
and U14993 (N_14993,N_13475,N_13713);
nand U14994 (N_14994,N_13152,N_13333);
xor U14995 (N_14995,N_13310,N_13879);
xnor U14996 (N_14996,N_13148,N_13468);
and U14997 (N_14997,N_13473,N_13135);
or U14998 (N_14998,N_13264,N_13809);
and U14999 (N_14999,N_13407,N_13142);
xnor U15000 (N_15000,N_14890,N_14395);
and U15001 (N_15001,N_14753,N_14829);
and U15002 (N_15002,N_14081,N_14728);
xnor U15003 (N_15003,N_14387,N_14489);
xor U15004 (N_15004,N_14096,N_14652);
or U15005 (N_15005,N_14146,N_14915);
nand U15006 (N_15006,N_14271,N_14595);
xor U15007 (N_15007,N_14956,N_14476);
xnor U15008 (N_15008,N_14340,N_14721);
or U15009 (N_15009,N_14708,N_14206);
nor U15010 (N_15010,N_14083,N_14738);
or U15011 (N_15011,N_14825,N_14002);
nand U15012 (N_15012,N_14255,N_14840);
xor U15013 (N_15013,N_14628,N_14657);
and U15014 (N_15014,N_14541,N_14132);
xnor U15015 (N_15015,N_14943,N_14016);
xnor U15016 (N_15016,N_14671,N_14803);
nor U15017 (N_15017,N_14209,N_14061);
xnor U15018 (N_15018,N_14348,N_14591);
xor U15019 (N_15019,N_14008,N_14996);
and U15020 (N_15020,N_14375,N_14337);
nor U15021 (N_15021,N_14195,N_14951);
nor U15022 (N_15022,N_14226,N_14100);
or U15023 (N_15023,N_14553,N_14438);
and U15024 (N_15024,N_14424,N_14783);
or U15025 (N_15025,N_14586,N_14357);
or U15026 (N_15026,N_14344,N_14169);
xor U15027 (N_15027,N_14958,N_14185);
xor U15028 (N_15028,N_14309,N_14510);
nand U15029 (N_15029,N_14318,N_14412);
nor U15030 (N_15030,N_14150,N_14297);
xor U15031 (N_15031,N_14334,N_14775);
xor U15032 (N_15032,N_14361,N_14937);
xor U15033 (N_15033,N_14291,N_14048);
xor U15034 (N_15034,N_14114,N_14874);
nand U15035 (N_15035,N_14976,N_14192);
nand U15036 (N_15036,N_14715,N_14091);
nand U15037 (N_15037,N_14716,N_14784);
nor U15038 (N_15038,N_14522,N_14046);
xor U15039 (N_15039,N_14953,N_14243);
xor U15040 (N_15040,N_14161,N_14518);
nor U15041 (N_15041,N_14741,N_14842);
xnor U15042 (N_15042,N_14734,N_14866);
and U15043 (N_15043,N_14449,N_14149);
xnor U15044 (N_15044,N_14520,N_14062);
nand U15045 (N_15045,N_14286,N_14848);
nor U15046 (N_15046,N_14440,N_14969);
or U15047 (N_15047,N_14214,N_14270);
nand U15048 (N_15048,N_14408,N_14078);
or U15049 (N_15049,N_14121,N_14622);
nand U15050 (N_15050,N_14273,N_14979);
or U15051 (N_15051,N_14780,N_14362);
or U15052 (N_15052,N_14802,N_14679);
xor U15053 (N_15053,N_14576,N_14148);
or U15054 (N_15054,N_14278,N_14488);
nor U15055 (N_15055,N_14985,N_14939);
nand U15056 (N_15056,N_14798,N_14913);
nor U15057 (N_15057,N_14792,N_14170);
nor U15058 (N_15058,N_14551,N_14727);
nand U15059 (N_15059,N_14515,N_14112);
and U15060 (N_15060,N_14963,N_14656);
nand U15061 (N_15061,N_14367,N_14154);
nor U15062 (N_15062,N_14805,N_14025);
or U15063 (N_15063,N_14856,N_14460);
nor U15064 (N_15064,N_14314,N_14852);
nor U15065 (N_15065,N_14131,N_14099);
nor U15066 (N_15066,N_14266,N_14364);
nor U15067 (N_15067,N_14631,N_14350);
xor U15068 (N_15068,N_14673,N_14228);
nor U15069 (N_15069,N_14880,N_14421);
xnor U15070 (N_15070,N_14946,N_14392);
xor U15071 (N_15071,N_14027,N_14499);
nand U15072 (N_15072,N_14846,N_14279);
and U15073 (N_15073,N_14503,N_14588);
nor U15074 (N_15074,N_14332,N_14974);
nand U15075 (N_15075,N_14101,N_14767);
nand U15076 (N_15076,N_14066,N_14247);
and U15077 (N_15077,N_14481,N_14687);
or U15078 (N_15078,N_14794,N_14638);
or U15079 (N_15079,N_14152,N_14335);
or U15080 (N_15080,N_14820,N_14675);
nor U15081 (N_15081,N_14873,N_14417);
nor U15082 (N_15082,N_14057,N_14198);
xnor U15083 (N_15083,N_14033,N_14843);
or U15084 (N_15084,N_14265,N_14063);
xnor U15085 (N_15085,N_14117,N_14982);
nand U15086 (N_15086,N_14865,N_14039);
nor U15087 (N_15087,N_14213,N_14160);
and U15088 (N_15088,N_14282,N_14024);
nand U15089 (N_15089,N_14621,N_14744);
xnor U15090 (N_15090,N_14137,N_14556);
and U15091 (N_15091,N_14277,N_14135);
nor U15092 (N_15092,N_14486,N_14513);
and U15093 (N_15093,N_14042,N_14186);
or U15094 (N_15094,N_14754,N_14818);
or U15095 (N_15095,N_14087,N_14686);
and U15096 (N_15096,N_14017,N_14069);
xor U15097 (N_15097,N_14891,N_14190);
and U15098 (N_15098,N_14237,N_14911);
and U15099 (N_15099,N_14324,N_14952);
or U15100 (N_15100,N_14623,N_14593);
or U15101 (N_15101,N_14352,N_14179);
or U15102 (N_15102,N_14723,N_14140);
xnor U15103 (N_15103,N_14126,N_14264);
nand U15104 (N_15104,N_14700,N_14872);
and U15105 (N_15105,N_14244,N_14181);
or U15106 (N_15106,N_14549,N_14750);
and U15107 (N_15107,N_14363,N_14110);
and U15108 (N_15108,N_14685,N_14225);
nand U15109 (N_15109,N_14756,N_14821);
or U15110 (N_15110,N_14430,N_14163);
nor U15111 (N_15111,N_14933,N_14581);
and U15112 (N_15112,N_14074,N_14054);
nor U15113 (N_15113,N_14116,N_14702);
xor U15114 (N_15114,N_14938,N_14568);
or U15115 (N_15115,N_14125,N_14659);
xor U15116 (N_15116,N_14105,N_14844);
and U15117 (N_15117,N_14498,N_14076);
nor U15118 (N_15118,N_14524,N_14761);
or U15119 (N_15119,N_14040,N_14322);
nand U15120 (N_15120,N_14766,N_14118);
nor U15121 (N_15121,N_14431,N_14372);
nor U15122 (N_15122,N_14875,N_14560);
nor U15123 (N_15123,N_14808,N_14639);
xor U15124 (N_15124,N_14910,N_14134);
xor U15125 (N_15125,N_14067,N_14323);
xor U15126 (N_15126,N_14159,N_14480);
xnor U15127 (N_15127,N_14407,N_14123);
nand U15128 (N_15128,N_14292,N_14053);
or U15129 (N_15129,N_14647,N_14834);
nand U15130 (N_15130,N_14954,N_14883);
nor U15131 (N_15131,N_14582,N_14535);
or U15132 (N_15132,N_14590,N_14109);
xnor U15133 (N_15133,N_14572,N_14287);
and U15134 (N_15134,N_14471,N_14947);
nor U15135 (N_15135,N_14534,N_14696);
or U15136 (N_15136,N_14165,N_14060);
nor U15137 (N_15137,N_14651,N_14763);
or U15138 (N_15138,N_14172,N_14859);
and U15139 (N_15139,N_14177,N_14986);
and U15140 (N_15140,N_14598,N_14563);
nor U15141 (N_15141,N_14980,N_14272);
and U15142 (N_15142,N_14092,N_14626);
and U15143 (N_15143,N_14878,N_14661);
and U15144 (N_15144,N_14786,N_14701);
xnor U15145 (N_15145,N_14837,N_14569);
nand U15146 (N_15146,N_14962,N_14385);
nand U15147 (N_15147,N_14887,N_14399);
nor U15148 (N_15148,N_14406,N_14683);
and U15149 (N_15149,N_14059,N_14311);
nor U15150 (N_15150,N_14839,N_14832);
nand U15151 (N_15151,N_14220,N_14461);
or U15152 (N_15152,N_14615,N_14609);
nor U15153 (N_15153,N_14787,N_14075);
xor U15154 (N_15154,N_14235,N_14779);
and U15155 (N_15155,N_14474,N_14381);
nand U15156 (N_15156,N_14012,N_14454);
and U15157 (N_15157,N_14436,N_14023);
xnor U15158 (N_15158,N_14442,N_14175);
nand U15159 (N_15159,N_14772,N_14119);
and U15160 (N_15160,N_14014,N_14452);
or U15161 (N_15161,N_14536,N_14793);
or U15162 (N_15162,N_14538,N_14371);
nand U15163 (N_15163,N_14690,N_14253);
or U15164 (N_15164,N_14819,N_14000);
nor U15165 (N_15165,N_14594,N_14705);
xor U15166 (N_15166,N_14936,N_14869);
nor U15167 (N_15167,N_14104,N_14166);
and U15168 (N_15168,N_14932,N_14703);
nand U15169 (N_15169,N_14566,N_14722);
nor U15170 (N_15170,N_14799,N_14633);
xnor U15171 (N_15171,N_14306,N_14851);
and U15172 (N_15172,N_14571,N_14712);
nor U15173 (N_15173,N_14575,N_14774);
nand U15174 (N_15174,N_14508,N_14815);
nand U15175 (N_15175,N_14307,N_14393);
and U15176 (N_15176,N_14885,N_14022);
or U15177 (N_15177,N_14677,N_14707);
and U15178 (N_15178,N_14713,N_14250);
and U15179 (N_15179,N_14216,N_14469);
and U15180 (N_15180,N_14330,N_14732);
nor U15181 (N_15181,N_14525,N_14240);
nor U15182 (N_15182,N_14669,N_14428);
xnor U15183 (N_15183,N_14580,N_14426);
and U15184 (N_15184,N_14302,N_14504);
nor U15185 (N_15185,N_14655,N_14317);
nor U15186 (N_15186,N_14989,N_14296);
xnor U15187 (N_15187,N_14196,N_14044);
or U15188 (N_15188,N_14251,N_14736);
xor U15189 (N_15189,N_14695,N_14212);
nand U15190 (N_15190,N_14710,N_14577);
xnor U15191 (N_15191,N_14811,N_14781);
nand U15192 (N_15192,N_14411,N_14258);
or U15193 (N_15193,N_14434,N_14725);
or U15194 (N_15194,N_14379,N_14382);
xor U15195 (N_15195,N_14992,N_14031);
nand U15196 (N_15196,N_14433,N_14618);
nand U15197 (N_15197,N_14831,N_14923);
nand U15198 (N_15198,N_14472,N_14111);
nor U15199 (N_15199,N_14429,N_14011);
nand U15200 (N_15200,N_14740,N_14927);
xor U15201 (N_15201,N_14005,N_14562);
xnor U15202 (N_15202,N_14051,N_14280);
and U15203 (N_15203,N_14122,N_14574);
and U15204 (N_15204,N_14338,N_14550);
and U15205 (N_15205,N_14868,N_14174);
xor U15206 (N_15206,N_14315,N_14545);
nand U15207 (N_15207,N_14863,N_14441);
xor U15208 (N_15208,N_14288,N_14689);
nor U15209 (N_15209,N_14648,N_14584);
nor U15210 (N_15210,N_14353,N_14448);
or U15211 (N_15211,N_14635,N_14403);
and U15212 (N_15212,N_14446,N_14966);
nand U15213 (N_15213,N_14641,N_14463);
and U15214 (N_15214,N_14726,N_14573);
or U15215 (N_15215,N_14972,N_14400);
or U15216 (N_15216,N_14490,N_14398);
nand U15217 (N_15217,N_14373,N_14804);
nand U15218 (N_15218,N_14080,N_14435);
and U15219 (N_15219,N_14529,N_14711);
and U15220 (N_15220,N_14293,N_14893);
or U15221 (N_15221,N_14778,N_14339);
and U15222 (N_15222,N_14917,N_14298);
or U15223 (N_15223,N_14743,N_14924);
nand U15224 (N_15224,N_14931,N_14506);
or U15225 (N_15225,N_14475,N_14329);
nor U15226 (N_15226,N_14877,N_14079);
and U15227 (N_15227,N_14791,N_14482);
or U15228 (N_15228,N_14055,N_14351);
nor U15229 (N_15229,N_14833,N_14785);
xor U15230 (N_15230,N_14564,N_14139);
nor U15231 (N_15231,N_14864,N_14967);
or U15232 (N_15232,N_14672,N_14610);
nor U15233 (N_15233,N_14261,N_14369);
and U15234 (N_15234,N_14456,N_14926);
xnor U15235 (N_15235,N_14483,N_14903);
xnor U15236 (N_15236,N_14465,N_14285);
nor U15237 (N_15237,N_14233,N_14236);
nor U15238 (N_15238,N_14902,N_14128);
nand U15239 (N_15239,N_14921,N_14642);
nand U15240 (N_15240,N_14627,N_14814);
xor U15241 (N_15241,N_14035,N_14645);
nand U15242 (N_15242,N_14603,N_14180);
or U15243 (N_15243,N_14771,N_14664);
nand U15244 (N_15244,N_14867,N_14276);
xnor U15245 (N_15245,N_14444,N_14912);
xor U15246 (N_15246,N_14420,N_14245);
xor U15247 (N_15247,N_14602,N_14445);
or U15248 (N_15248,N_14559,N_14082);
nand U15249 (N_15249,N_14994,N_14222);
nand U15250 (N_15250,N_14491,N_14879);
nor U15251 (N_15251,N_14171,N_14800);
nand U15252 (N_15252,N_14283,N_14770);
or U15253 (N_15253,N_14983,N_14227);
xor U15254 (N_15254,N_14733,N_14527);
nand U15255 (N_15255,N_14145,N_14300);
nor U15256 (N_15256,N_14409,N_14987);
nand U15257 (N_15257,N_14384,N_14796);
nor U15258 (N_15258,N_14028,N_14208);
nand U15259 (N_15259,N_14305,N_14684);
and U15260 (N_15260,N_14319,N_14935);
nand U15261 (N_15261,N_14467,N_14606);
or U15262 (N_15262,N_14530,N_14533);
nand U15263 (N_15263,N_14904,N_14760);
xor U15264 (N_15264,N_14698,N_14676);
or U15265 (N_15265,N_14519,N_14681);
or U15266 (N_15266,N_14678,N_14528);
and U15267 (N_15267,N_14432,N_14151);
xnor U15268 (N_15268,N_14516,N_14094);
and U15269 (N_15269,N_14202,N_14630);
and U15270 (N_15270,N_14167,N_14548);
and U15271 (N_15271,N_14929,N_14249);
nor U15272 (N_15272,N_14049,N_14719);
and U15273 (N_15273,N_14437,N_14223);
or U15274 (N_15274,N_14036,N_14341);
xor U15275 (N_15275,N_14680,N_14977);
nor U15276 (N_15276,N_14397,N_14999);
and U15277 (N_15277,N_14493,N_14130);
and U15278 (N_15278,N_14136,N_14898);
xnor U15279 (N_15279,N_14897,N_14200);
and U15280 (N_15280,N_14817,N_14579);
and U15281 (N_15281,N_14295,N_14459);
or U15282 (N_15282,N_14876,N_14824);
nand U15283 (N_15283,N_14532,N_14260);
or U15284 (N_15284,N_14047,N_14084);
xnor U15285 (N_15285,N_14103,N_14546);
nor U15286 (N_15286,N_14201,N_14289);
xnor U15287 (N_15287,N_14758,N_14089);
or U15288 (N_15288,N_14592,N_14355);
and U15289 (N_15289,N_14555,N_14252);
nand U15290 (N_15290,N_14512,N_14178);
nand U15291 (N_15291,N_14841,N_14451);
and U15292 (N_15292,N_14823,N_14826);
nor U15293 (N_15293,N_14138,N_14997);
or U15294 (N_15294,N_14404,N_14410);
xor U15295 (N_15295,N_14995,N_14973);
xor U15296 (N_15296,N_14349,N_14511);
and U15297 (N_15297,N_14124,N_14102);
and U15298 (N_15298,N_14718,N_14658);
or U15299 (N_15299,N_14182,N_14144);
nand U15300 (N_15300,N_14269,N_14360);
or U15301 (N_15301,N_14120,N_14850);
nand U15302 (N_15302,N_14540,N_14347);
xnor U15303 (N_15303,N_14210,N_14735);
xnor U15304 (N_15304,N_14849,N_14782);
xnor U15305 (N_15305,N_14906,N_14514);
nor U15306 (N_15306,N_14523,N_14968);
or U15307 (N_15307,N_14961,N_14881);
nor U15308 (N_15308,N_14773,N_14356);
and U15309 (N_15309,N_14199,N_14855);
nor U15310 (N_15310,N_14238,N_14313);
nand U15311 (N_15311,N_14162,N_14729);
or U15312 (N_15312,N_14345,N_14617);
and U15313 (N_15313,N_14714,N_14401);
and U15314 (N_15314,N_14242,N_14884);
nand U15315 (N_15315,N_14164,N_14071);
nand U15316 (N_15316,N_14359,N_14693);
xor U15317 (N_15317,N_14405,N_14965);
or U15318 (N_15318,N_14427,N_14263);
xnor U15319 (N_15319,N_14558,N_14919);
or U15320 (N_15320,N_14697,N_14991);
or U15321 (N_15321,N_14653,N_14959);
xor U15322 (N_15322,N_14466,N_14207);
or U15323 (N_15323,N_14045,N_14640);
nor U15324 (N_15324,N_14717,N_14422);
or U15325 (N_15325,N_14343,N_14517);
and U15326 (N_15326,N_14674,N_14981);
or U15327 (N_15327,N_14443,N_14239);
nand U15328 (N_15328,N_14215,N_14205);
nor U15329 (N_15329,N_14248,N_14497);
or U15330 (N_15330,N_14757,N_14822);
or U15331 (N_15331,N_14870,N_14189);
nand U15332 (N_15332,N_14905,N_14739);
or U15333 (N_15333,N_14468,N_14604);
or U15334 (N_15334,N_14464,N_14414);
xor U15335 (N_15335,N_14462,N_14458);
or U15336 (N_15336,N_14203,N_14896);
nand U15337 (N_15337,N_14147,N_14453);
or U15338 (N_15338,N_14388,N_14900);
xnor U15339 (N_15339,N_14599,N_14095);
nand U15340 (N_15340,N_14644,N_14886);
xnor U15341 (N_15341,N_14478,N_14742);
nand U15342 (N_15342,N_14004,N_14806);
or U15343 (N_15343,N_14663,N_14037);
and U15344 (N_15344,N_14988,N_14133);
and U15345 (N_15345,N_14336,N_14041);
xnor U15346 (N_15346,N_14015,N_14984);
nand U15347 (N_15347,N_14835,N_14378);
xnor U15348 (N_15348,N_14221,N_14231);
nor U15349 (N_15349,N_14386,N_14026);
or U15350 (N_15350,N_14376,N_14762);
or U15351 (N_15351,N_14749,N_14812);
nor U15352 (N_15352,N_14667,N_14457);
nor U15353 (N_15353,N_14747,N_14502);
xor U15354 (N_15354,N_14485,N_14888);
and U15355 (N_15355,N_14328,N_14807);
nor U15356 (N_15356,N_14050,N_14585);
and U15357 (N_15357,N_14234,N_14380);
or U15358 (N_15358,N_14646,N_14847);
xor U15359 (N_15359,N_14521,N_14899);
xor U15360 (N_15360,N_14043,N_14542);
or U15361 (N_15361,N_14613,N_14854);
nor U15362 (N_15362,N_14290,N_14871);
nand U15363 (N_15363,N_14157,N_14281);
nand U15364 (N_15364,N_14254,N_14724);
nand U15365 (N_15365,N_14601,N_14745);
nand U15366 (N_15366,N_14990,N_14187);
and U15367 (N_15367,N_14326,N_14916);
and U15368 (N_15368,N_14731,N_14629);
and U15369 (N_15369,N_14415,N_14570);
or U15370 (N_15370,N_14383,N_14097);
nand U15371 (N_15371,N_14267,N_14666);
nand U15372 (N_15372,N_14193,N_14746);
or U15373 (N_15373,N_14670,N_14940);
or U15374 (N_15374,N_14583,N_14034);
and U15375 (N_15375,N_14224,N_14509);
and U15376 (N_15376,N_14001,N_14975);
or U15377 (N_15377,N_14567,N_14776);
and U15378 (N_15378,N_14788,N_14816);
xnor U15379 (N_15379,N_14544,N_14003);
nand U15380 (N_15380,N_14423,N_14882);
nor U15381 (N_15381,N_14636,N_14925);
xor U15382 (N_15382,N_14068,N_14611);
nor U15383 (N_15383,N_14030,N_14010);
or U15384 (N_15384,N_14777,N_14668);
and U15385 (N_15385,N_14908,N_14557);
and U15386 (N_15386,N_14346,N_14769);
nor U15387 (N_15387,N_14971,N_14143);
nor U15388 (N_15388,N_14928,N_14909);
or U15389 (N_15389,N_14184,N_14256);
xnor U15390 (N_15390,N_14934,N_14688);
and U15391 (N_15391,N_14013,N_14539);
xnor U15392 (N_15392,N_14470,N_14643);
or U15393 (N_15393,N_14194,N_14065);
nand U15394 (N_15394,N_14077,N_14625);
nor U15395 (N_15395,N_14587,N_14993);
nand U15396 (N_15396,N_14416,N_14914);
xor U15397 (N_15397,N_14704,N_14894);
nand U15398 (N_15398,N_14790,N_14321);
xor U15399 (N_15399,N_14402,N_14107);
nor U15400 (N_15400,N_14183,N_14419);
xnor U15401 (N_15401,N_14191,N_14494);
xor U15402 (N_15402,N_14608,N_14246);
xor U15403 (N_15403,N_14391,N_14316);
and U15404 (N_15404,N_14358,N_14920);
nand U15405 (N_15405,N_14021,N_14970);
nand U15406 (N_15406,N_14861,N_14365);
xor U15407 (N_15407,N_14945,N_14377);
and U15408 (N_15408,N_14978,N_14605);
nand U15409 (N_15409,N_14058,N_14230);
nor U15410 (N_15410,N_14662,N_14860);
xor U15411 (N_15411,N_14578,N_14115);
or U15412 (N_15412,N_14699,N_14998);
and U15413 (N_15413,N_14895,N_14614);
and U15414 (N_15414,N_14838,N_14052);
nand U15415 (N_15415,N_14554,N_14070);
nand U15416 (N_15416,N_14537,N_14211);
xor U15417 (N_15417,N_14168,N_14907);
nand U15418 (N_15418,N_14032,N_14730);
or U15419 (N_15419,N_14129,N_14156);
or U15420 (N_15420,N_14142,N_14692);
or U15421 (N_15421,N_14531,N_14217);
and U15422 (N_15422,N_14176,N_14301);
nor U15423 (N_15423,N_14304,N_14492);
xor U15424 (N_15424,N_14901,N_14589);
or U15425 (N_15425,N_14764,N_14331);
nor U15426 (N_15426,N_14197,N_14543);
nor U15427 (N_15427,N_14596,N_14862);
xor U15428 (N_15428,N_14942,N_14188);
nor U15429 (N_15429,N_14484,N_14706);
and U15430 (N_15430,N_14098,N_14085);
nand U15431 (N_15431,N_14072,N_14394);
xor U15432 (N_15432,N_14845,N_14858);
xnor U15433 (N_15433,N_14552,N_14964);
and U15434 (N_15434,N_14836,N_14370);
nand U15435 (N_15435,N_14694,N_14634);
xor U15436 (N_15436,N_14827,N_14607);
nand U15437 (N_15437,N_14038,N_14654);
nand U15438 (N_15438,N_14957,N_14294);
xnor U15439 (N_15439,N_14018,N_14029);
xnor U15440 (N_15440,N_14616,N_14450);
nor U15441 (N_15441,N_14413,N_14158);
nor U15442 (N_15442,N_14073,N_14765);
or U15443 (N_15443,N_14828,N_14241);
or U15444 (N_15444,N_14056,N_14310);
or U15445 (N_15445,N_14299,N_14950);
and U15446 (N_15446,N_14561,N_14853);
and U15447 (N_15447,N_14141,N_14325);
nand U15448 (N_15448,N_14086,N_14219);
nor U15449 (N_15449,N_14624,N_14650);
nor U15450 (N_15450,N_14487,N_14789);
xnor U15451 (N_15451,N_14389,N_14333);
and U15452 (N_15452,N_14153,N_14455);
nand U15453 (N_15453,N_14709,N_14303);
xor U15454 (N_15454,N_14009,N_14108);
and U15455 (N_15455,N_14955,N_14374);
xor U15456 (N_15456,N_14795,N_14944);
xor U15457 (N_15457,N_14390,N_14797);
or U15458 (N_15458,N_14660,N_14007);
xnor U15459 (N_15459,N_14597,N_14006);
or U15460 (N_15460,N_14889,N_14752);
and U15461 (N_15461,N_14755,N_14892);
nor U15462 (N_15462,N_14366,N_14759);
nand U15463 (N_15463,N_14275,N_14801);
or U15464 (N_15464,N_14809,N_14020);
and U15465 (N_15465,N_14477,N_14501);
nand U15466 (N_15466,N_14632,N_14064);
and U15467 (N_15467,N_14751,N_14682);
and U15468 (N_15468,N_14768,N_14857);
nor U15469 (N_15469,N_14259,N_14665);
nor U15470 (N_15470,N_14418,N_14620);
or U15471 (N_15471,N_14930,N_14257);
xor U15472 (N_15472,N_14619,N_14218);
xor U15473 (N_15473,N_14500,N_14425);
nor U15474 (N_15474,N_14127,N_14830);
nand U15475 (N_15475,N_14810,N_14691);
and U15476 (N_15476,N_14439,N_14565);
nand U15477 (N_15477,N_14106,N_14396);
or U15478 (N_15478,N_14342,N_14948);
and U15479 (N_15479,N_14547,N_14268);
xnor U15480 (N_15480,N_14720,N_14612);
nand U15481 (N_15481,N_14507,N_14949);
nor U15482 (N_15482,N_14496,N_14173);
and U15483 (N_15483,N_14232,N_14368);
or U15484 (N_15484,N_14113,N_14922);
nand U15485 (N_15485,N_14505,N_14473);
or U15486 (N_15486,N_14090,N_14155);
nand U15487 (N_15487,N_14941,N_14479);
xnor U15488 (N_15488,N_14019,N_14320);
nand U15489 (N_15489,N_14737,N_14447);
nand U15490 (N_15490,N_14649,N_14229);
or U15491 (N_15491,N_14918,N_14748);
and U15492 (N_15492,N_14093,N_14600);
or U15493 (N_15493,N_14308,N_14960);
xnor U15494 (N_15494,N_14312,N_14813);
nor U15495 (N_15495,N_14262,N_14204);
xor U15496 (N_15496,N_14327,N_14495);
or U15497 (N_15497,N_14274,N_14088);
nand U15498 (N_15498,N_14284,N_14526);
nand U15499 (N_15499,N_14354,N_14637);
xnor U15500 (N_15500,N_14644,N_14854);
xor U15501 (N_15501,N_14705,N_14554);
and U15502 (N_15502,N_14953,N_14458);
and U15503 (N_15503,N_14375,N_14364);
or U15504 (N_15504,N_14927,N_14426);
nand U15505 (N_15505,N_14997,N_14235);
nor U15506 (N_15506,N_14259,N_14595);
and U15507 (N_15507,N_14982,N_14166);
xnor U15508 (N_15508,N_14693,N_14835);
nand U15509 (N_15509,N_14558,N_14719);
and U15510 (N_15510,N_14937,N_14054);
xnor U15511 (N_15511,N_14178,N_14391);
nand U15512 (N_15512,N_14683,N_14630);
xnor U15513 (N_15513,N_14860,N_14595);
or U15514 (N_15514,N_14413,N_14007);
and U15515 (N_15515,N_14358,N_14977);
nor U15516 (N_15516,N_14844,N_14679);
xor U15517 (N_15517,N_14447,N_14632);
or U15518 (N_15518,N_14355,N_14533);
and U15519 (N_15519,N_14865,N_14425);
xor U15520 (N_15520,N_14634,N_14000);
xnor U15521 (N_15521,N_14660,N_14270);
nand U15522 (N_15522,N_14279,N_14490);
xnor U15523 (N_15523,N_14783,N_14298);
or U15524 (N_15524,N_14115,N_14588);
xnor U15525 (N_15525,N_14356,N_14646);
nor U15526 (N_15526,N_14204,N_14071);
and U15527 (N_15527,N_14529,N_14795);
and U15528 (N_15528,N_14366,N_14031);
nor U15529 (N_15529,N_14379,N_14515);
and U15530 (N_15530,N_14527,N_14392);
or U15531 (N_15531,N_14730,N_14599);
or U15532 (N_15532,N_14818,N_14000);
or U15533 (N_15533,N_14760,N_14624);
xnor U15534 (N_15534,N_14068,N_14465);
nor U15535 (N_15535,N_14307,N_14566);
xor U15536 (N_15536,N_14614,N_14266);
xnor U15537 (N_15537,N_14656,N_14477);
and U15538 (N_15538,N_14716,N_14391);
nor U15539 (N_15539,N_14391,N_14435);
or U15540 (N_15540,N_14209,N_14560);
and U15541 (N_15541,N_14717,N_14558);
nand U15542 (N_15542,N_14447,N_14228);
nor U15543 (N_15543,N_14700,N_14530);
nor U15544 (N_15544,N_14804,N_14873);
nand U15545 (N_15545,N_14189,N_14623);
and U15546 (N_15546,N_14407,N_14792);
nand U15547 (N_15547,N_14428,N_14389);
or U15548 (N_15548,N_14129,N_14248);
or U15549 (N_15549,N_14308,N_14111);
nand U15550 (N_15550,N_14801,N_14956);
or U15551 (N_15551,N_14713,N_14149);
xnor U15552 (N_15552,N_14577,N_14119);
nor U15553 (N_15553,N_14426,N_14216);
or U15554 (N_15554,N_14042,N_14657);
xor U15555 (N_15555,N_14887,N_14392);
or U15556 (N_15556,N_14085,N_14158);
or U15557 (N_15557,N_14687,N_14079);
nor U15558 (N_15558,N_14433,N_14688);
xnor U15559 (N_15559,N_14705,N_14886);
and U15560 (N_15560,N_14033,N_14516);
or U15561 (N_15561,N_14940,N_14792);
or U15562 (N_15562,N_14851,N_14675);
and U15563 (N_15563,N_14566,N_14447);
nor U15564 (N_15564,N_14798,N_14627);
nand U15565 (N_15565,N_14410,N_14423);
or U15566 (N_15566,N_14803,N_14810);
nor U15567 (N_15567,N_14522,N_14211);
or U15568 (N_15568,N_14904,N_14003);
or U15569 (N_15569,N_14877,N_14343);
nand U15570 (N_15570,N_14288,N_14404);
or U15571 (N_15571,N_14423,N_14548);
nand U15572 (N_15572,N_14875,N_14558);
nand U15573 (N_15573,N_14487,N_14398);
xnor U15574 (N_15574,N_14924,N_14574);
nand U15575 (N_15575,N_14297,N_14139);
nand U15576 (N_15576,N_14368,N_14481);
and U15577 (N_15577,N_14117,N_14647);
and U15578 (N_15578,N_14042,N_14350);
nor U15579 (N_15579,N_14476,N_14415);
and U15580 (N_15580,N_14347,N_14092);
xnor U15581 (N_15581,N_14746,N_14719);
nor U15582 (N_15582,N_14206,N_14361);
nor U15583 (N_15583,N_14948,N_14136);
xnor U15584 (N_15584,N_14674,N_14110);
and U15585 (N_15585,N_14717,N_14294);
and U15586 (N_15586,N_14660,N_14658);
or U15587 (N_15587,N_14683,N_14455);
nor U15588 (N_15588,N_14239,N_14116);
nand U15589 (N_15589,N_14026,N_14182);
or U15590 (N_15590,N_14584,N_14216);
or U15591 (N_15591,N_14959,N_14314);
or U15592 (N_15592,N_14696,N_14717);
or U15593 (N_15593,N_14076,N_14242);
nor U15594 (N_15594,N_14808,N_14656);
nor U15595 (N_15595,N_14553,N_14295);
nand U15596 (N_15596,N_14862,N_14799);
or U15597 (N_15597,N_14386,N_14549);
or U15598 (N_15598,N_14419,N_14648);
nor U15599 (N_15599,N_14629,N_14557);
nand U15600 (N_15600,N_14405,N_14003);
nand U15601 (N_15601,N_14954,N_14670);
xor U15602 (N_15602,N_14488,N_14601);
xnor U15603 (N_15603,N_14192,N_14338);
xnor U15604 (N_15604,N_14861,N_14515);
xor U15605 (N_15605,N_14774,N_14579);
nor U15606 (N_15606,N_14531,N_14743);
xor U15607 (N_15607,N_14038,N_14487);
or U15608 (N_15608,N_14594,N_14787);
nor U15609 (N_15609,N_14261,N_14266);
and U15610 (N_15610,N_14863,N_14374);
or U15611 (N_15611,N_14808,N_14024);
or U15612 (N_15612,N_14092,N_14849);
xor U15613 (N_15613,N_14096,N_14957);
xor U15614 (N_15614,N_14350,N_14257);
and U15615 (N_15615,N_14116,N_14692);
nor U15616 (N_15616,N_14604,N_14685);
nand U15617 (N_15617,N_14392,N_14461);
or U15618 (N_15618,N_14633,N_14230);
or U15619 (N_15619,N_14352,N_14499);
nand U15620 (N_15620,N_14281,N_14820);
xor U15621 (N_15621,N_14567,N_14973);
or U15622 (N_15622,N_14248,N_14684);
nand U15623 (N_15623,N_14204,N_14271);
xor U15624 (N_15624,N_14014,N_14017);
nand U15625 (N_15625,N_14332,N_14648);
or U15626 (N_15626,N_14924,N_14271);
and U15627 (N_15627,N_14099,N_14496);
and U15628 (N_15628,N_14540,N_14199);
or U15629 (N_15629,N_14523,N_14143);
xnor U15630 (N_15630,N_14619,N_14581);
and U15631 (N_15631,N_14707,N_14697);
nor U15632 (N_15632,N_14093,N_14070);
and U15633 (N_15633,N_14952,N_14988);
and U15634 (N_15634,N_14930,N_14534);
nor U15635 (N_15635,N_14762,N_14283);
or U15636 (N_15636,N_14133,N_14395);
xor U15637 (N_15637,N_14630,N_14478);
xnor U15638 (N_15638,N_14841,N_14457);
and U15639 (N_15639,N_14029,N_14709);
xor U15640 (N_15640,N_14993,N_14913);
or U15641 (N_15641,N_14253,N_14332);
and U15642 (N_15642,N_14343,N_14684);
or U15643 (N_15643,N_14779,N_14214);
nor U15644 (N_15644,N_14045,N_14176);
nand U15645 (N_15645,N_14470,N_14707);
xnor U15646 (N_15646,N_14174,N_14352);
nand U15647 (N_15647,N_14544,N_14245);
xor U15648 (N_15648,N_14590,N_14215);
xor U15649 (N_15649,N_14833,N_14989);
and U15650 (N_15650,N_14555,N_14340);
nand U15651 (N_15651,N_14743,N_14303);
nor U15652 (N_15652,N_14456,N_14289);
or U15653 (N_15653,N_14325,N_14066);
xnor U15654 (N_15654,N_14914,N_14167);
and U15655 (N_15655,N_14567,N_14286);
and U15656 (N_15656,N_14367,N_14052);
nor U15657 (N_15657,N_14602,N_14079);
nor U15658 (N_15658,N_14689,N_14554);
or U15659 (N_15659,N_14141,N_14005);
nor U15660 (N_15660,N_14956,N_14260);
and U15661 (N_15661,N_14304,N_14178);
nand U15662 (N_15662,N_14582,N_14148);
nor U15663 (N_15663,N_14050,N_14511);
or U15664 (N_15664,N_14677,N_14236);
xnor U15665 (N_15665,N_14166,N_14713);
or U15666 (N_15666,N_14077,N_14830);
nand U15667 (N_15667,N_14831,N_14694);
nand U15668 (N_15668,N_14105,N_14470);
xor U15669 (N_15669,N_14576,N_14868);
or U15670 (N_15670,N_14086,N_14963);
nand U15671 (N_15671,N_14140,N_14687);
nor U15672 (N_15672,N_14278,N_14491);
and U15673 (N_15673,N_14120,N_14138);
nand U15674 (N_15674,N_14878,N_14142);
or U15675 (N_15675,N_14412,N_14544);
nor U15676 (N_15676,N_14182,N_14007);
nor U15677 (N_15677,N_14508,N_14433);
xnor U15678 (N_15678,N_14604,N_14757);
nand U15679 (N_15679,N_14313,N_14784);
xor U15680 (N_15680,N_14991,N_14484);
xor U15681 (N_15681,N_14182,N_14524);
nand U15682 (N_15682,N_14682,N_14542);
nand U15683 (N_15683,N_14703,N_14677);
nand U15684 (N_15684,N_14233,N_14103);
and U15685 (N_15685,N_14533,N_14399);
xor U15686 (N_15686,N_14311,N_14102);
nor U15687 (N_15687,N_14729,N_14210);
and U15688 (N_15688,N_14942,N_14400);
nand U15689 (N_15689,N_14452,N_14618);
or U15690 (N_15690,N_14030,N_14936);
or U15691 (N_15691,N_14423,N_14158);
or U15692 (N_15692,N_14365,N_14353);
xnor U15693 (N_15693,N_14198,N_14899);
xnor U15694 (N_15694,N_14953,N_14459);
or U15695 (N_15695,N_14201,N_14239);
xor U15696 (N_15696,N_14758,N_14065);
nand U15697 (N_15697,N_14798,N_14719);
nor U15698 (N_15698,N_14726,N_14410);
and U15699 (N_15699,N_14269,N_14054);
xor U15700 (N_15700,N_14711,N_14388);
and U15701 (N_15701,N_14542,N_14803);
nor U15702 (N_15702,N_14999,N_14398);
and U15703 (N_15703,N_14250,N_14182);
and U15704 (N_15704,N_14587,N_14541);
and U15705 (N_15705,N_14657,N_14320);
and U15706 (N_15706,N_14246,N_14755);
xnor U15707 (N_15707,N_14023,N_14657);
xor U15708 (N_15708,N_14404,N_14513);
or U15709 (N_15709,N_14418,N_14267);
xor U15710 (N_15710,N_14582,N_14688);
nand U15711 (N_15711,N_14055,N_14360);
nor U15712 (N_15712,N_14721,N_14509);
xnor U15713 (N_15713,N_14613,N_14151);
or U15714 (N_15714,N_14442,N_14263);
nand U15715 (N_15715,N_14355,N_14247);
xor U15716 (N_15716,N_14176,N_14381);
or U15717 (N_15717,N_14937,N_14636);
nor U15718 (N_15718,N_14011,N_14835);
nand U15719 (N_15719,N_14450,N_14537);
nand U15720 (N_15720,N_14720,N_14323);
xnor U15721 (N_15721,N_14327,N_14162);
nor U15722 (N_15722,N_14635,N_14070);
or U15723 (N_15723,N_14728,N_14922);
nand U15724 (N_15724,N_14854,N_14278);
xnor U15725 (N_15725,N_14431,N_14065);
nand U15726 (N_15726,N_14962,N_14387);
xnor U15727 (N_15727,N_14174,N_14902);
nand U15728 (N_15728,N_14434,N_14944);
xnor U15729 (N_15729,N_14891,N_14069);
nor U15730 (N_15730,N_14287,N_14535);
nand U15731 (N_15731,N_14012,N_14820);
and U15732 (N_15732,N_14142,N_14499);
or U15733 (N_15733,N_14500,N_14020);
nand U15734 (N_15734,N_14916,N_14788);
nand U15735 (N_15735,N_14707,N_14320);
xor U15736 (N_15736,N_14718,N_14595);
nor U15737 (N_15737,N_14724,N_14005);
nor U15738 (N_15738,N_14780,N_14200);
nor U15739 (N_15739,N_14340,N_14019);
or U15740 (N_15740,N_14786,N_14315);
nand U15741 (N_15741,N_14146,N_14839);
xnor U15742 (N_15742,N_14532,N_14636);
nand U15743 (N_15743,N_14731,N_14635);
xor U15744 (N_15744,N_14010,N_14679);
and U15745 (N_15745,N_14240,N_14340);
and U15746 (N_15746,N_14517,N_14142);
or U15747 (N_15747,N_14295,N_14404);
or U15748 (N_15748,N_14526,N_14065);
nand U15749 (N_15749,N_14498,N_14266);
nand U15750 (N_15750,N_14925,N_14260);
and U15751 (N_15751,N_14116,N_14831);
nor U15752 (N_15752,N_14717,N_14984);
and U15753 (N_15753,N_14433,N_14858);
nor U15754 (N_15754,N_14511,N_14072);
or U15755 (N_15755,N_14626,N_14550);
nor U15756 (N_15756,N_14420,N_14595);
and U15757 (N_15757,N_14398,N_14068);
or U15758 (N_15758,N_14679,N_14762);
xor U15759 (N_15759,N_14720,N_14964);
or U15760 (N_15760,N_14732,N_14464);
or U15761 (N_15761,N_14152,N_14413);
nand U15762 (N_15762,N_14639,N_14992);
nor U15763 (N_15763,N_14306,N_14653);
nand U15764 (N_15764,N_14302,N_14791);
or U15765 (N_15765,N_14520,N_14773);
and U15766 (N_15766,N_14046,N_14643);
nor U15767 (N_15767,N_14855,N_14944);
nand U15768 (N_15768,N_14459,N_14393);
or U15769 (N_15769,N_14178,N_14266);
nor U15770 (N_15770,N_14961,N_14856);
nand U15771 (N_15771,N_14698,N_14319);
xor U15772 (N_15772,N_14692,N_14417);
xor U15773 (N_15773,N_14573,N_14012);
nand U15774 (N_15774,N_14175,N_14771);
or U15775 (N_15775,N_14621,N_14587);
and U15776 (N_15776,N_14774,N_14183);
xnor U15777 (N_15777,N_14534,N_14523);
nand U15778 (N_15778,N_14052,N_14983);
nor U15779 (N_15779,N_14670,N_14034);
nor U15780 (N_15780,N_14189,N_14066);
xor U15781 (N_15781,N_14551,N_14007);
nand U15782 (N_15782,N_14689,N_14734);
nor U15783 (N_15783,N_14882,N_14309);
nor U15784 (N_15784,N_14709,N_14225);
and U15785 (N_15785,N_14563,N_14656);
nor U15786 (N_15786,N_14067,N_14523);
and U15787 (N_15787,N_14873,N_14225);
nand U15788 (N_15788,N_14870,N_14978);
and U15789 (N_15789,N_14074,N_14310);
and U15790 (N_15790,N_14269,N_14322);
nand U15791 (N_15791,N_14762,N_14196);
and U15792 (N_15792,N_14161,N_14177);
nor U15793 (N_15793,N_14972,N_14378);
xnor U15794 (N_15794,N_14416,N_14734);
nor U15795 (N_15795,N_14530,N_14679);
nand U15796 (N_15796,N_14673,N_14482);
nand U15797 (N_15797,N_14733,N_14618);
nor U15798 (N_15798,N_14444,N_14760);
nor U15799 (N_15799,N_14902,N_14305);
nand U15800 (N_15800,N_14344,N_14561);
nor U15801 (N_15801,N_14575,N_14802);
xor U15802 (N_15802,N_14146,N_14193);
nor U15803 (N_15803,N_14423,N_14095);
nor U15804 (N_15804,N_14949,N_14639);
or U15805 (N_15805,N_14414,N_14924);
nor U15806 (N_15806,N_14012,N_14107);
or U15807 (N_15807,N_14723,N_14910);
and U15808 (N_15808,N_14176,N_14924);
or U15809 (N_15809,N_14827,N_14949);
nor U15810 (N_15810,N_14114,N_14241);
nand U15811 (N_15811,N_14333,N_14431);
or U15812 (N_15812,N_14575,N_14794);
or U15813 (N_15813,N_14080,N_14497);
nand U15814 (N_15814,N_14639,N_14140);
or U15815 (N_15815,N_14068,N_14905);
nor U15816 (N_15816,N_14584,N_14644);
or U15817 (N_15817,N_14944,N_14333);
nor U15818 (N_15818,N_14027,N_14337);
nand U15819 (N_15819,N_14946,N_14232);
nand U15820 (N_15820,N_14119,N_14444);
or U15821 (N_15821,N_14232,N_14981);
nand U15822 (N_15822,N_14791,N_14360);
and U15823 (N_15823,N_14268,N_14297);
xor U15824 (N_15824,N_14686,N_14917);
and U15825 (N_15825,N_14545,N_14600);
nor U15826 (N_15826,N_14423,N_14549);
or U15827 (N_15827,N_14449,N_14688);
nand U15828 (N_15828,N_14139,N_14220);
xor U15829 (N_15829,N_14590,N_14127);
nand U15830 (N_15830,N_14645,N_14982);
nor U15831 (N_15831,N_14525,N_14334);
or U15832 (N_15832,N_14069,N_14360);
nand U15833 (N_15833,N_14959,N_14257);
nand U15834 (N_15834,N_14426,N_14583);
and U15835 (N_15835,N_14349,N_14844);
nand U15836 (N_15836,N_14866,N_14811);
nand U15837 (N_15837,N_14730,N_14150);
xor U15838 (N_15838,N_14132,N_14699);
xnor U15839 (N_15839,N_14734,N_14087);
and U15840 (N_15840,N_14925,N_14198);
nor U15841 (N_15841,N_14191,N_14904);
or U15842 (N_15842,N_14077,N_14944);
xnor U15843 (N_15843,N_14391,N_14329);
and U15844 (N_15844,N_14203,N_14830);
and U15845 (N_15845,N_14776,N_14783);
and U15846 (N_15846,N_14807,N_14157);
or U15847 (N_15847,N_14338,N_14376);
or U15848 (N_15848,N_14066,N_14302);
nor U15849 (N_15849,N_14421,N_14332);
xnor U15850 (N_15850,N_14765,N_14083);
nand U15851 (N_15851,N_14669,N_14873);
nor U15852 (N_15852,N_14884,N_14076);
xnor U15853 (N_15853,N_14254,N_14138);
and U15854 (N_15854,N_14876,N_14175);
and U15855 (N_15855,N_14517,N_14667);
or U15856 (N_15856,N_14912,N_14375);
xor U15857 (N_15857,N_14618,N_14275);
or U15858 (N_15858,N_14819,N_14760);
and U15859 (N_15859,N_14626,N_14792);
nand U15860 (N_15860,N_14893,N_14132);
nor U15861 (N_15861,N_14576,N_14223);
xor U15862 (N_15862,N_14541,N_14058);
and U15863 (N_15863,N_14394,N_14883);
and U15864 (N_15864,N_14923,N_14318);
nor U15865 (N_15865,N_14202,N_14228);
nor U15866 (N_15866,N_14755,N_14154);
and U15867 (N_15867,N_14494,N_14742);
nor U15868 (N_15868,N_14212,N_14064);
nor U15869 (N_15869,N_14059,N_14120);
xnor U15870 (N_15870,N_14798,N_14284);
nand U15871 (N_15871,N_14583,N_14824);
xnor U15872 (N_15872,N_14143,N_14139);
or U15873 (N_15873,N_14479,N_14498);
nor U15874 (N_15874,N_14418,N_14124);
nand U15875 (N_15875,N_14371,N_14639);
and U15876 (N_15876,N_14270,N_14488);
or U15877 (N_15877,N_14598,N_14751);
or U15878 (N_15878,N_14505,N_14561);
nand U15879 (N_15879,N_14163,N_14529);
or U15880 (N_15880,N_14625,N_14280);
nor U15881 (N_15881,N_14580,N_14564);
nand U15882 (N_15882,N_14910,N_14659);
or U15883 (N_15883,N_14382,N_14186);
or U15884 (N_15884,N_14030,N_14097);
and U15885 (N_15885,N_14060,N_14025);
nand U15886 (N_15886,N_14411,N_14662);
or U15887 (N_15887,N_14060,N_14002);
or U15888 (N_15888,N_14405,N_14777);
or U15889 (N_15889,N_14741,N_14131);
nand U15890 (N_15890,N_14399,N_14556);
xor U15891 (N_15891,N_14140,N_14264);
and U15892 (N_15892,N_14791,N_14930);
nand U15893 (N_15893,N_14338,N_14092);
xnor U15894 (N_15894,N_14304,N_14195);
or U15895 (N_15895,N_14350,N_14830);
nor U15896 (N_15896,N_14940,N_14733);
nor U15897 (N_15897,N_14250,N_14828);
nand U15898 (N_15898,N_14552,N_14868);
or U15899 (N_15899,N_14580,N_14735);
nand U15900 (N_15900,N_14119,N_14589);
xor U15901 (N_15901,N_14206,N_14770);
nand U15902 (N_15902,N_14391,N_14990);
nor U15903 (N_15903,N_14853,N_14921);
nand U15904 (N_15904,N_14267,N_14718);
nand U15905 (N_15905,N_14529,N_14953);
or U15906 (N_15906,N_14804,N_14523);
and U15907 (N_15907,N_14250,N_14468);
and U15908 (N_15908,N_14186,N_14468);
nand U15909 (N_15909,N_14864,N_14332);
xor U15910 (N_15910,N_14793,N_14726);
or U15911 (N_15911,N_14398,N_14441);
xnor U15912 (N_15912,N_14455,N_14566);
nor U15913 (N_15913,N_14393,N_14926);
and U15914 (N_15914,N_14416,N_14443);
or U15915 (N_15915,N_14125,N_14652);
or U15916 (N_15916,N_14427,N_14815);
xnor U15917 (N_15917,N_14601,N_14396);
and U15918 (N_15918,N_14442,N_14402);
nand U15919 (N_15919,N_14197,N_14405);
and U15920 (N_15920,N_14014,N_14413);
nor U15921 (N_15921,N_14259,N_14094);
nand U15922 (N_15922,N_14125,N_14537);
nand U15923 (N_15923,N_14854,N_14008);
nor U15924 (N_15924,N_14316,N_14271);
and U15925 (N_15925,N_14038,N_14955);
nand U15926 (N_15926,N_14844,N_14737);
xor U15927 (N_15927,N_14882,N_14989);
and U15928 (N_15928,N_14212,N_14249);
xnor U15929 (N_15929,N_14179,N_14788);
and U15930 (N_15930,N_14304,N_14936);
and U15931 (N_15931,N_14032,N_14180);
xnor U15932 (N_15932,N_14693,N_14694);
xor U15933 (N_15933,N_14184,N_14160);
or U15934 (N_15934,N_14034,N_14735);
nand U15935 (N_15935,N_14898,N_14549);
or U15936 (N_15936,N_14610,N_14334);
nand U15937 (N_15937,N_14440,N_14740);
nor U15938 (N_15938,N_14344,N_14002);
or U15939 (N_15939,N_14006,N_14759);
xor U15940 (N_15940,N_14770,N_14859);
nand U15941 (N_15941,N_14206,N_14626);
nor U15942 (N_15942,N_14602,N_14158);
nor U15943 (N_15943,N_14704,N_14679);
and U15944 (N_15944,N_14730,N_14634);
or U15945 (N_15945,N_14433,N_14095);
or U15946 (N_15946,N_14356,N_14902);
xnor U15947 (N_15947,N_14627,N_14015);
xor U15948 (N_15948,N_14174,N_14004);
nand U15949 (N_15949,N_14478,N_14042);
nand U15950 (N_15950,N_14852,N_14436);
nand U15951 (N_15951,N_14922,N_14362);
nand U15952 (N_15952,N_14184,N_14201);
nand U15953 (N_15953,N_14946,N_14268);
or U15954 (N_15954,N_14765,N_14719);
xor U15955 (N_15955,N_14576,N_14048);
and U15956 (N_15956,N_14910,N_14610);
and U15957 (N_15957,N_14562,N_14215);
nand U15958 (N_15958,N_14614,N_14433);
or U15959 (N_15959,N_14346,N_14757);
nor U15960 (N_15960,N_14878,N_14346);
xor U15961 (N_15961,N_14788,N_14804);
and U15962 (N_15962,N_14722,N_14447);
and U15963 (N_15963,N_14267,N_14469);
and U15964 (N_15964,N_14758,N_14851);
or U15965 (N_15965,N_14169,N_14357);
nand U15966 (N_15966,N_14749,N_14994);
nand U15967 (N_15967,N_14567,N_14695);
nand U15968 (N_15968,N_14419,N_14066);
and U15969 (N_15969,N_14782,N_14966);
or U15970 (N_15970,N_14589,N_14346);
or U15971 (N_15971,N_14809,N_14797);
and U15972 (N_15972,N_14011,N_14639);
nor U15973 (N_15973,N_14941,N_14221);
and U15974 (N_15974,N_14583,N_14581);
and U15975 (N_15975,N_14865,N_14629);
xnor U15976 (N_15976,N_14823,N_14481);
nor U15977 (N_15977,N_14022,N_14420);
nand U15978 (N_15978,N_14177,N_14932);
nand U15979 (N_15979,N_14584,N_14356);
or U15980 (N_15980,N_14455,N_14940);
nor U15981 (N_15981,N_14744,N_14502);
nand U15982 (N_15982,N_14424,N_14865);
nand U15983 (N_15983,N_14418,N_14299);
or U15984 (N_15984,N_14174,N_14231);
or U15985 (N_15985,N_14393,N_14041);
nand U15986 (N_15986,N_14959,N_14024);
xnor U15987 (N_15987,N_14761,N_14628);
xnor U15988 (N_15988,N_14070,N_14871);
or U15989 (N_15989,N_14852,N_14487);
nor U15990 (N_15990,N_14911,N_14868);
or U15991 (N_15991,N_14317,N_14308);
and U15992 (N_15992,N_14566,N_14301);
nor U15993 (N_15993,N_14023,N_14746);
nand U15994 (N_15994,N_14792,N_14056);
xnor U15995 (N_15995,N_14979,N_14872);
or U15996 (N_15996,N_14716,N_14342);
xnor U15997 (N_15997,N_14845,N_14077);
xnor U15998 (N_15998,N_14851,N_14583);
xor U15999 (N_15999,N_14481,N_14557);
nor U16000 (N_16000,N_15810,N_15575);
nor U16001 (N_16001,N_15966,N_15827);
nor U16002 (N_16002,N_15985,N_15024);
or U16003 (N_16003,N_15833,N_15113);
or U16004 (N_16004,N_15892,N_15094);
and U16005 (N_16005,N_15283,N_15862);
or U16006 (N_16006,N_15793,N_15357);
nor U16007 (N_16007,N_15176,N_15642);
nor U16008 (N_16008,N_15019,N_15585);
and U16009 (N_16009,N_15114,N_15180);
nor U16010 (N_16010,N_15297,N_15930);
and U16011 (N_16011,N_15962,N_15660);
nor U16012 (N_16012,N_15223,N_15516);
or U16013 (N_16013,N_15543,N_15956);
or U16014 (N_16014,N_15060,N_15397);
nand U16015 (N_16015,N_15971,N_15277);
nor U16016 (N_16016,N_15493,N_15133);
or U16017 (N_16017,N_15068,N_15931);
nand U16018 (N_16018,N_15257,N_15684);
nor U16019 (N_16019,N_15441,N_15529);
xnor U16020 (N_16020,N_15664,N_15540);
and U16021 (N_16021,N_15320,N_15579);
nand U16022 (N_16022,N_15851,N_15759);
nor U16023 (N_16023,N_15295,N_15779);
xnor U16024 (N_16024,N_15783,N_15146);
or U16025 (N_16025,N_15795,N_15322);
xor U16026 (N_16026,N_15937,N_15134);
and U16027 (N_16027,N_15603,N_15940);
and U16028 (N_16028,N_15195,N_15991);
nor U16029 (N_16029,N_15392,N_15200);
xnor U16030 (N_16030,N_15785,N_15190);
nand U16031 (N_16031,N_15222,N_15770);
and U16032 (N_16032,N_15828,N_15040);
and U16033 (N_16033,N_15550,N_15921);
nor U16034 (N_16034,N_15254,N_15748);
xor U16035 (N_16035,N_15228,N_15883);
or U16036 (N_16036,N_15062,N_15431);
nor U16037 (N_16037,N_15207,N_15172);
nor U16038 (N_16038,N_15396,N_15382);
nand U16039 (N_16039,N_15141,N_15570);
or U16040 (N_16040,N_15405,N_15671);
nand U16041 (N_16041,N_15789,N_15632);
or U16042 (N_16042,N_15074,N_15026);
nor U16043 (N_16043,N_15319,N_15048);
or U16044 (N_16044,N_15161,N_15410);
nand U16045 (N_16045,N_15373,N_15363);
xor U16046 (N_16046,N_15121,N_15333);
nand U16047 (N_16047,N_15029,N_15343);
nor U16048 (N_16048,N_15238,N_15303);
nor U16049 (N_16049,N_15519,N_15174);
nand U16050 (N_16050,N_15292,N_15525);
nor U16051 (N_16051,N_15701,N_15666);
nand U16052 (N_16052,N_15943,N_15699);
or U16053 (N_16053,N_15577,N_15305);
xor U16054 (N_16054,N_15476,N_15751);
or U16055 (N_16055,N_15462,N_15559);
xor U16056 (N_16056,N_15980,N_15852);
or U16057 (N_16057,N_15855,N_15453);
nor U16058 (N_16058,N_15039,N_15872);
and U16059 (N_16059,N_15440,N_15831);
nand U16060 (N_16060,N_15022,N_15734);
xor U16061 (N_16061,N_15140,N_15918);
nor U16062 (N_16062,N_15767,N_15717);
xnor U16063 (N_16063,N_15327,N_15778);
and U16064 (N_16064,N_15683,N_15188);
and U16065 (N_16065,N_15128,N_15239);
nor U16066 (N_16066,N_15983,N_15732);
xnor U16067 (N_16067,N_15994,N_15663);
nand U16068 (N_16068,N_15435,N_15091);
or U16069 (N_16069,N_15159,N_15950);
or U16070 (N_16070,N_15093,N_15424);
or U16071 (N_16071,N_15466,N_15706);
xnor U16072 (N_16072,N_15420,N_15438);
or U16073 (N_16073,N_15953,N_15434);
xor U16074 (N_16074,N_15809,N_15982);
and U16075 (N_16075,N_15873,N_15471);
and U16076 (N_16076,N_15457,N_15120);
xor U16077 (N_16077,N_15447,N_15201);
nand U16078 (N_16078,N_15170,N_15451);
xnor U16079 (N_16079,N_15766,N_15848);
nand U16080 (N_16080,N_15426,N_15595);
nor U16081 (N_16081,N_15191,N_15563);
xnor U16082 (N_16082,N_15513,N_15482);
nand U16083 (N_16083,N_15057,N_15667);
nor U16084 (N_16084,N_15535,N_15693);
nand U16085 (N_16085,N_15947,N_15477);
and U16086 (N_16086,N_15847,N_15437);
nor U16087 (N_16087,N_15959,N_15499);
and U16088 (N_16088,N_15731,N_15206);
xor U16089 (N_16089,N_15713,N_15934);
and U16090 (N_16090,N_15129,N_15596);
and U16091 (N_16091,N_15491,N_15227);
nor U16092 (N_16092,N_15386,N_15063);
nand U16093 (N_16093,N_15811,N_15349);
or U16094 (N_16094,N_15259,N_15557);
nor U16095 (N_16095,N_15560,N_15240);
or U16096 (N_16096,N_15647,N_15745);
nand U16097 (N_16097,N_15696,N_15924);
or U16098 (N_16098,N_15309,N_15163);
nand U16099 (N_16099,N_15593,N_15271);
nor U16100 (N_16100,N_15840,N_15744);
nor U16101 (N_16101,N_15286,N_15876);
or U16102 (N_16102,N_15193,N_15630);
and U16103 (N_16103,N_15474,N_15698);
and U16104 (N_16104,N_15756,N_15584);
and U16105 (N_16105,N_15674,N_15034);
nor U16106 (N_16106,N_15411,N_15680);
nor U16107 (N_16107,N_15878,N_15501);
nor U16108 (N_16108,N_15043,N_15012);
and U16109 (N_16109,N_15657,N_15013);
or U16110 (N_16110,N_15742,N_15650);
xnor U16111 (N_16111,N_15002,N_15459);
nand U16112 (N_16112,N_15419,N_15167);
or U16113 (N_16113,N_15443,N_15375);
nand U16114 (N_16114,N_15325,N_15211);
or U16115 (N_16115,N_15308,N_15486);
and U16116 (N_16116,N_15097,N_15110);
and U16117 (N_16117,N_15275,N_15977);
xnor U16118 (N_16118,N_15107,N_15638);
xnor U16119 (N_16119,N_15629,N_15580);
nand U16120 (N_16120,N_15866,N_15072);
xor U16121 (N_16121,N_15716,N_15694);
nand U16122 (N_16122,N_15331,N_15210);
and U16123 (N_16123,N_15960,N_15626);
nor U16124 (N_16124,N_15221,N_15708);
xor U16125 (N_16125,N_15186,N_15747);
nand U16126 (N_16126,N_15669,N_15566);
and U16127 (N_16127,N_15164,N_15341);
xor U16128 (N_16128,N_15602,N_15056);
nand U16129 (N_16129,N_15010,N_15591);
nand U16130 (N_16130,N_15350,N_15217);
and U16131 (N_16131,N_15888,N_15504);
nor U16132 (N_16132,N_15661,N_15733);
nor U16133 (N_16133,N_15260,N_15065);
xor U16134 (N_16134,N_15025,N_15433);
or U16135 (N_16135,N_15372,N_15364);
nor U16136 (N_16136,N_15864,N_15242);
nor U16137 (N_16137,N_15967,N_15534);
nand U16138 (N_16138,N_15998,N_15573);
nor U16139 (N_16139,N_15352,N_15954);
nor U16140 (N_16140,N_15802,N_15762);
xnor U16141 (N_16141,N_15345,N_15760);
nor U16142 (N_16142,N_15533,N_15138);
and U16143 (N_16143,N_15387,N_15711);
nand U16144 (N_16144,N_15631,N_15722);
nor U16145 (N_16145,N_15023,N_15205);
or U16146 (N_16146,N_15016,N_15735);
or U16147 (N_16147,N_15938,N_15229);
xnor U16148 (N_16148,N_15512,N_15393);
nand U16149 (N_16149,N_15886,N_15358);
nand U16150 (N_16150,N_15807,N_15402);
nand U16151 (N_16151,N_15598,N_15902);
and U16152 (N_16152,N_15692,N_15755);
xnor U16153 (N_16153,N_15185,N_15498);
xor U16154 (N_16154,N_15652,N_15332);
xnor U16155 (N_16155,N_15678,N_15119);
xor U16156 (N_16156,N_15670,N_15957);
nor U16157 (N_16157,N_15703,N_15542);
or U16158 (N_16158,N_15316,N_15475);
or U16159 (N_16159,N_15881,N_15028);
nand U16160 (N_16160,N_15224,N_15280);
xor U16161 (N_16161,N_15098,N_15900);
nor U16162 (N_16162,N_15503,N_15797);
nor U16163 (N_16163,N_15727,N_15418);
nand U16164 (N_16164,N_15030,N_15311);
nand U16165 (N_16165,N_15355,N_15523);
nor U16166 (N_16166,N_15569,N_15656);
xnor U16167 (N_16167,N_15874,N_15806);
nand U16168 (N_16168,N_15484,N_15600);
xor U16169 (N_16169,N_15117,N_15945);
nand U16170 (N_16170,N_15863,N_15007);
or U16171 (N_16171,N_15335,N_15995);
nor U16172 (N_16172,N_15815,N_15859);
and U16173 (N_16173,N_15099,N_15623);
or U16174 (N_16174,N_15215,N_15880);
xnor U16175 (N_16175,N_15158,N_15336);
nand U16176 (N_16176,N_15446,N_15052);
and U16177 (N_16177,N_15775,N_15171);
nor U16178 (N_16178,N_15112,N_15380);
nor U16179 (N_16179,N_15932,N_15123);
xor U16180 (N_16180,N_15665,N_15076);
and U16181 (N_16181,N_15232,N_15624);
or U16182 (N_16182,N_15160,N_15988);
or U16183 (N_16183,N_15871,N_15248);
or U16184 (N_16184,N_15317,N_15611);
nand U16185 (N_16185,N_15262,N_15891);
nand U16186 (N_16186,N_15515,N_15588);
or U16187 (N_16187,N_15821,N_15547);
and U16188 (N_16188,N_15237,N_15782);
xnor U16189 (N_16189,N_15524,N_15581);
xnor U16190 (N_16190,N_15147,N_15055);
nor U16191 (N_16191,N_15323,N_15483);
nor U16192 (N_16192,N_15673,N_15772);
nand U16193 (N_16193,N_15278,N_15737);
or U16194 (N_16194,N_15620,N_15979);
or U16195 (N_16195,N_15691,N_15688);
xnor U16196 (N_16196,N_15145,N_15870);
and U16197 (N_16197,N_15686,N_15935);
nor U16198 (N_16198,N_15685,N_15369);
nor U16199 (N_16199,N_15951,N_15599);
nand U16200 (N_16200,N_15730,N_15230);
or U16201 (N_16201,N_15106,N_15721);
xor U16202 (N_16202,N_15077,N_15939);
nand U16203 (N_16203,N_15090,N_15495);
xnor U16204 (N_16204,N_15249,N_15073);
or U16205 (N_16205,N_15389,N_15291);
xnor U16206 (N_16206,N_15294,N_15777);
or U16207 (N_16207,N_15901,N_15036);
or U16208 (N_16208,N_15468,N_15787);
or U16209 (N_16209,N_15272,N_15489);
nor U16210 (N_16210,N_15178,N_15554);
xnor U16211 (N_16211,N_15427,N_15911);
and U16212 (N_16212,N_15752,N_15083);
nand U16213 (N_16213,N_15344,N_15627);
or U16214 (N_16214,N_15315,N_15899);
and U16215 (N_16215,N_15398,N_15823);
nand U16216 (N_16216,N_15470,N_15460);
or U16217 (N_16217,N_15909,N_15754);
xnor U16218 (N_16218,N_15067,N_15092);
xnor U16219 (N_16219,N_15682,N_15545);
nor U16220 (N_16220,N_15808,N_15508);
and U16221 (N_16221,N_15480,N_15154);
nor U16222 (N_16222,N_15781,N_15820);
xor U16223 (N_16223,N_15606,N_15976);
xnor U16224 (N_16224,N_15571,N_15908);
nor U16225 (N_16225,N_15890,N_15725);
nor U16226 (N_16226,N_15984,N_15514);
and U16227 (N_16227,N_15084,N_15773);
or U16228 (N_16228,N_15607,N_15915);
or U16229 (N_16229,N_15768,N_15788);
nor U16230 (N_16230,N_15150,N_15613);
or U16231 (N_16231,N_15182,N_15000);
and U16232 (N_16232,N_15845,N_15391);
or U16233 (N_16233,N_15875,N_15075);
and U16234 (N_16234,N_15517,N_15949);
xor U16235 (N_16235,N_15409,N_15882);
nand U16236 (N_16236,N_15465,N_15485);
nor U16237 (N_16237,N_15033,N_15394);
and U16238 (N_16238,N_15149,N_15049);
xnor U16239 (N_16239,N_15739,N_15774);
nand U16240 (N_16240,N_15096,N_15812);
or U16241 (N_16241,N_15518,N_15109);
nor U16242 (N_16242,N_15687,N_15556);
nor U16243 (N_16243,N_15038,N_15996);
or U16244 (N_16244,N_15253,N_15108);
nor U16245 (N_16245,N_15798,N_15124);
nand U16246 (N_16246,N_15233,N_15676);
xnor U16247 (N_16247,N_15078,N_15439);
nor U16248 (N_16248,N_15893,N_15849);
or U16249 (N_16249,N_15836,N_15044);
nor U16250 (N_16250,N_15247,N_15987);
nand U16251 (N_16251,N_15252,N_15689);
nand U16252 (N_16252,N_15758,N_15008);
or U16253 (N_16253,N_15461,N_15913);
or U16254 (N_16254,N_15640,N_15964);
nand U16255 (N_16255,N_15400,N_15243);
and U16256 (N_16256,N_15919,N_15487);
nor U16257 (N_16257,N_15235,N_15791);
xnor U16258 (N_16258,N_15655,N_15609);
and U16259 (N_16259,N_15646,N_15274);
xor U16260 (N_16260,N_15157,N_15047);
nor U16261 (N_16261,N_15526,N_15511);
nand U16262 (N_16262,N_15003,N_15648);
nand U16263 (N_16263,N_15366,N_15144);
xor U16264 (N_16264,N_15269,N_15497);
and U16265 (N_16265,N_15383,N_15955);
or U16266 (N_16266,N_15381,N_15572);
xor U16267 (N_16267,N_15822,N_15565);
and U16268 (N_16268,N_15786,N_15856);
or U16269 (N_16269,N_15738,N_15702);
and U16270 (N_16270,N_15250,N_15050);
and U16271 (N_16271,N_15801,N_15895);
xor U16272 (N_16272,N_15225,N_15763);
nor U16273 (N_16273,N_15729,N_15928);
nor U16274 (N_16274,N_15961,N_15819);
xor U16275 (N_16275,N_15152,N_15081);
nand U16276 (N_16276,N_15654,N_15679);
nand U16277 (N_16277,N_15799,N_15379);
and U16278 (N_16278,N_15992,N_15522);
nand U16279 (N_16279,N_15463,N_15339);
or U16280 (N_16280,N_15415,N_15792);
xor U16281 (N_16281,N_15946,N_15187);
and U16282 (N_16282,N_15346,N_15496);
or U16283 (N_16283,N_15284,N_15153);
nor U16284 (N_16284,N_15726,N_15189);
xor U16285 (N_16285,N_15009,N_15813);
and U16286 (N_16286,N_15436,N_15920);
or U16287 (N_16287,N_15804,N_15532);
xnor U16288 (N_16288,N_15697,N_15213);
or U16289 (N_16289,N_15425,N_15860);
or U16290 (N_16290,N_15625,N_15118);
xnor U16291 (N_16291,N_15968,N_15502);
and U16292 (N_16292,N_15192,N_15743);
nor U16293 (N_16293,N_15850,N_15528);
nand U16294 (N_16294,N_15263,N_15413);
xor U16295 (N_16295,N_15347,N_15478);
nor U16296 (N_16296,N_15279,N_15132);
and U16297 (N_16297,N_15989,N_15651);
xnor U16298 (N_16298,N_15212,N_15423);
nor U16299 (N_16299,N_15111,N_15844);
xor U16300 (N_16300,N_15973,N_15724);
or U16301 (N_16301,N_15906,N_15923);
xor U16302 (N_16302,N_15450,N_15184);
and U16303 (N_16303,N_15634,N_15728);
or U16304 (N_16304,N_15455,N_15965);
xnor U16305 (N_16305,N_15941,N_15066);
xor U16306 (N_16306,N_15367,N_15531);
nor U16307 (N_16307,N_15203,N_15059);
xnor U16308 (N_16308,N_15835,N_15668);
and U16309 (N_16309,N_15417,N_15558);
or U16310 (N_16310,N_15958,N_15199);
nand U16311 (N_16311,N_15970,N_15115);
nand U16312 (N_16312,N_15270,N_15690);
and U16313 (N_16313,N_15538,N_15925);
or U16314 (N_16314,N_15204,N_15162);
xor U16315 (N_16315,N_15614,N_15469);
or U16316 (N_16316,N_15749,N_15710);
xor U16317 (N_16317,N_15544,N_15061);
and U16318 (N_16318,N_15948,N_15136);
nor U16319 (N_16319,N_15541,N_15301);
nand U16320 (N_16320,N_15408,N_15374);
xnor U16321 (N_16321,N_15905,N_15753);
or U16322 (N_16322,N_15549,N_15619);
or U16323 (N_16323,N_15234,N_15045);
or U16324 (N_16324,N_15390,N_15800);
xnor U16325 (N_16325,N_15288,N_15137);
nand U16326 (N_16326,N_15621,N_15826);
and U16327 (N_16327,N_15618,N_15776);
nor U16328 (N_16328,N_15330,N_15633);
xor U16329 (N_16329,N_15551,N_15889);
nor U16330 (N_16330,N_15494,N_15407);
nand U16331 (N_16331,N_15617,N_15298);
or U16332 (N_16332,N_15219,N_15395);
xnor U16333 (N_16333,N_15289,N_15361);
nor U16334 (N_16334,N_15658,N_15546);
and U16335 (N_16335,N_15582,N_15885);
nand U16336 (N_16336,N_15490,N_15051);
and U16337 (N_16337,N_15371,N_15377);
xnor U16338 (N_16338,N_15643,N_15592);
and U16339 (N_16339,N_15429,N_15765);
or U16340 (N_16340,N_15231,N_15853);
or U16341 (N_16341,N_15761,N_15805);
nand U16342 (N_16342,N_15780,N_15127);
and U16343 (N_16343,N_15649,N_15824);
xnor U16344 (N_16344,N_15256,N_15677);
and U16345 (N_16345,N_15903,N_15017);
xnor U16346 (N_16346,N_15927,N_15004);
or U16347 (N_16347,N_15929,N_15884);
and U16348 (N_16348,N_15116,N_15448);
xor U16349 (N_16349,N_15404,N_15299);
or U16350 (N_16350,N_15421,N_15432);
nor U16351 (N_16351,N_15936,N_15583);
and U16352 (N_16352,N_15981,N_15281);
nand U16353 (N_16353,N_15993,N_15353);
or U16354 (N_16354,N_15790,N_15027);
xnor U16355 (N_16355,N_15302,N_15181);
xor U16356 (N_16356,N_15574,N_15403);
or U16357 (N_16357,N_15198,N_15841);
or U16358 (N_16358,N_15509,N_15507);
and U16359 (N_16359,N_15169,N_15832);
nand U16360 (N_16360,N_15926,N_15715);
nand U16361 (N_16361,N_15368,N_15675);
nor U16362 (N_16362,N_15362,N_15088);
xor U16363 (N_16363,N_15071,N_15268);
nand U16364 (N_16364,N_15709,N_15218);
nor U16365 (N_16365,N_15458,N_15287);
and U16366 (N_16366,N_15342,N_15351);
and U16367 (N_16367,N_15539,N_15142);
and U16368 (N_16368,N_15834,N_15456);
nand U16369 (N_16369,N_15401,N_15628);
nand U16370 (N_16370,N_15865,N_15718);
nand U16371 (N_16371,N_15527,N_15705);
xnor U16372 (N_16372,N_15015,N_15058);
or U16373 (N_16373,N_15814,N_15135);
and U16374 (N_16374,N_15416,N_15086);
and U16375 (N_16375,N_15276,N_15131);
or U16376 (N_16376,N_15894,N_15794);
nand U16377 (N_16377,N_15869,N_15264);
and U16378 (N_16378,N_15481,N_15255);
and U16379 (N_16379,N_15720,N_15681);
nor U16380 (N_16380,N_15321,N_15467);
xnor U16381 (N_16381,N_15719,N_15285);
or U16382 (N_16382,N_15179,N_15590);
and U16383 (N_16383,N_15442,N_15054);
or U16384 (N_16384,N_15796,N_15839);
or U16385 (N_16385,N_15561,N_15488);
nand U16386 (N_16386,N_15473,N_15359);
nor U16387 (N_16387,N_15334,N_15356);
nand U16388 (N_16388,N_15552,N_15102);
or U16389 (N_16389,N_15576,N_15293);
or U16390 (N_16390,N_15125,N_15521);
nand U16391 (N_16391,N_15032,N_15622);
nor U16392 (N_16392,N_15639,N_15986);
and U16393 (N_16393,N_15662,N_15388);
or U16394 (N_16394,N_15300,N_15143);
or U16395 (N_16395,N_15035,N_15079);
nand U16396 (N_16396,N_15974,N_15644);
nor U16397 (N_16397,N_15340,N_15616);
nor U16398 (N_16398,N_15328,N_15520);
nand U16399 (N_16399,N_15422,N_15296);
and U16400 (N_16400,N_15216,N_15479);
and U16401 (N_16401,N_15548,N_15879);
xnor U16402 (N_16402,N_15376,N_15365);
xnor U16403 (N_16403,N_15586,N_15750);
and U16404 (N_16404,N_15868,N_15636);
xnor U16405 (N_16405,N_15011,N_15578);
or U16406 (N_16406,N_15612,N_15241);
nor U16407 (N_16407,N_15555,N_15492);
nand U16408 (N_16408,N_15830,N_15904);
xnor U16409 (N_16409,N_15452,N_15313);
nor U16410 (N_16410,N_15020,N_15635);
or U16411 (N_16411,N_15445,N_15916);
nand U16412 (N_16412,N_15089,N_15910);
nand U16413 (N_16413,N_15952,N_15933);
xnor U16414 (N_16414,N_15312,N_15505);
nor U16415 (N_16415,N_15095,N_15087);
nor U16416 (N_16416,N_15304,N_15173);
nand U16417 (N_16417,N_15196,N_15208);
xnor U16418 (N_16418,N_15615,N_15378);
nand U16419 (N_16419,N_15069,N_15282);
nand U16420 (N_16420,N_15053,N_15867);
and U16421 (N_16421,N_15168,N_15412);
and U16422 (N_16422,N_15177,N_15318);
nand U16423 (N_16423,N_15449,N_15506);
nand U16424 (N_16424,N_15897,N_15803);
and U16425 (N_16425,N_15202,N_15246);
xor U16426 (N_16426,N_15338,N_15907);
nor U16427 (N_16427,N_15816,N_15741);
nand U16428 (N_16428,N_15553,N_15014);
nand U16429 (N_16429,N_15194,N_15444);
xor U16430 (N_16430,N_15290,N_15912);
nand U16431 (N_16431,N_15597,N_15082);
nand U16432 (N_16432,N_15963,N_15641);
nand U16433 (N_16433,N_15637,N_15704);
or U16434 (N_16434,N_15354,N_15001);
nor U16435 (N_16435,N_15605,N_15126);
and U16436 (N_16436,N_15251,N_15064);
nand U16437 (N_16437,N_15103,N_15018);
or U16438 (N_16438,N_15307,N_15944);
xnor U16439 (N_16439,N_15324,N_15672);
or U16440 (N_16440,N_15037,N_15165);
or U16441 (N_16441,N_15975,N_15080);
nor U16442 (N_16442,N_15784,N_15370);
xor U16443 (N_16443,N_15854,N_15837);
nand U16444 (N_16444,N_15454,N_15843);
nor U16445 (N_16445,N_15645,N_15046);
nand U16446 (N_16446,N_15700,N_15536);
xnor U16447 (N_16447,N_15414,N_15155);
and U16448 (N_16448,N_15430,N_15156);
xnor U16449 (N_16449,N_15978,N_15510);
or U16450 (N_16450,N_15385,N_15608);
and U16451 (N_16451,N_15214,N_15151);
nand U16452 (N_16452,N_15348,N_15942);
xor U16453 (N_16453,N_15070,N_15031);
nand U16454 (N_16454,N_15306,N_15610);
nor U16455 (N_16455,N_15530,N_15042);
nand U16456 (N_16456,N_15723,N_15266);
nand U16457 (N_16457,N_15148,N_15922);
or U16458 (N_16458,N_15537,N_15261);
and U16459 (N_16459,N_15898,N_15707);
nor U16460 (N_16460,N_15990,N_15384);
and U16461 (N_16461,N_15314,N_15587);
nand U16462 (N_16462,N_15653,N_15175);
xnor U16463 (N_16463,N_15825,N_15265);
nand U16464 (N_16464,N_15769,N_15562);
xnor U16465 (N_16465,N_15464,N_15166);
nand U16466 (N_16466,N_15972,N_15740);
nor U16467 (N_16467,N_15326,N_15746);
and U16468 (N_16468,N_15564,N_15267);
nand U16469 (N_16469,N_15122,N_15568);
and U16470 (N_16470,N_15818,N_15245);
nand U16471 (N_16471,N_15428,N_15310);
xnor U16472 (N_16472,N_15258,N_15838);
nand U16473 (N_16473,N_15917,N_15846);
xor U16474 (N_16474,N_15659,N_15105);
nor U16475 (N_16475,N_15472,N_15757);
xor U16476 (N_16476,N_15604,N_15914);
nor U16477 (N_16477,N_15197,N_15183);
nor U16478 (N_16478,N_15273,N_15500);
or U16479 (N_16479,N_15236,N_15130);
xnor U16480 (N_16480,N_15005,N_15329);
nor U16481 (N_16481,N_15771,N_15220);
or U16482 (N_16482,N_15567,N_15764);
xor U16483 (N_16483,N_15887,N_15006);
or U16484 (N_16484,N_15085,N_15861);
xor U16485 (N_16485,N_15817,N_15858);
or U16486 (N_16486,N_15041,N_15857);
and U16487 (N_16487,N_15021,N_15842);
and U16488 (N_16488,N_15226,N_15209);
or U16489 (N_16489,N_15896,N_15589);
or U16490 (N_16490,N_15594,N_15714);
nor U16491 (N_16491,N_15101,N_15337);
xor U16492 (N_16492,N_15100,N_15399);
and U16493 (N_16493,N_15969,N_15601);
or U16494 (N_16494,N_15360,N_15695);
nand U16495 (N_16495,N_15104,N_15999);
xnor U16496 (N_16496,N_15406,N_15829);
and U16497 (N_16497,N_15877,N_15244);
or U16498 (N_16498,N_15736,N_15997);
and U16499 (N_16499,N_15712,N_15139);
or U16500 (N_16500,N_15344,N_15406);
or U16501 (N_16501,N_15324,N_15298);
and U16502 (N_16502,N_15414,N_15578);
xor U16503 (N_16503,N_15644,N_15696);
and U16504 (N_16504,N_15466,N_15124);
nor U16505 (N_16505,N_15898,N_15103);
xor U16506 (N_16506,N_15368,N_15639);
and U16507 (N_16507,N_15582,N_15588);
or U16508 (N_16508,N_15363,N_15842);
xor U16509 (N_16509,N_15669,N_15217);
xnor U16510 (N_16510,N_15795,N_15456);
or U16511 (N_16511,N_15750,N_15543);
nand U16512 (N_16512,N_15697,N_15776);
xnor U16513 (N_16513,N_15868,N_15433);
nand U16514 (N_16514,N_15485,N_15706);
nor U16515 (N_16515,N_15656,N_15187);
and U16516 (N_16516,N_15943,N_15878);
or U16517 (N_16517,N_15449,N_15840);
or U16518 (N_16518,N_15375,N_15194);
or U16519 (N_16519,N_15544,N_15996);
nand U16520 (N_16520,N_15446,N_15931);
xor U16521 (N_16521,N_15274,N_15559);
and U16522 (N_16522,N_15525,N_15328);
xor U16523 (N_16523,N_15536,N_15972);
or U16524 (N_16524,N_15424,N_15389);
xor U16525 (N_16525,N_15640,N_15592);
nand U16526 (N_16526,N_15055,N_15377);
or U16527 (N_16527,N_15117,N_15664);
or U16528 (N_16528,N_15132,N_15054);
nor U16529 (N_16529,N_15890,N_15308);
xnor U16530 (N_16530,N_15023,N_15497);
xor U16531 (N_16531,N_15013,N_15088);
xnor U16532 (N_16532,N_15152,N_15585);
or U16533 (N_16533,N_15351,N_15366);
xnor U16534 (N_16534,N_15331,N_15175);
xor U16535 (N_16535,N_15850,N_15513);
nor U16536 (N_16536,N_15505,N_15927);
and U16537 (N_16537,N_15325,N_15658);
nor U16538 (N_16538,N_15749,N_15271);
and U16539 (N_16539,N_15771,N_15236);
or U16540 (N_16540,N_15461,N_15331);
nand U16541 (N_16541,N_15795,N_15428);
nand U16542 (N_16542,N_15247,N_15785);
nor U16543 (N_16543,N_15835,N_15788);
nor U16544 (N_16544,N_15508,N_15369);
and U16545 (N_16545,N_15421,N_15980);
and U16546 (N_16546,N_15194,N_15775);
and U16547 (N_16547,N_15622,N_15109);
nand U16548 (N_16548,N_15080,N_15173);
xnor U16549 (N_16549,N_15259,N_15264);
nor U16550 (N_16550,N_15710,N_15356);
nand U16551 (N_16551,N_15134,N_15154);
and U16552 (N_16552,N_15043,N_15119);
or U16553 (N_16553,N_15187,N_15976);
nand U16554 (N_16554,N_15342,N_15402);
and U16555 (N_16555,N_15097,N_15952);
nand U16556 (N_16556,N_15660,N_15228);
xor U16557 (N_16557,N_15694,N_15223);
xnor U16558 (N_16558,N_15177,N_15636);
nand U16559 (N_16559,N_15464,N_15719);
or U16560 (N_16560,N_15615,N_15412);
or U16561 (N_16561,N_15869,N_15638);
nand U16562 (N_16562,N_15237,N_15655);
or U16563 (N_16563,N_15617,N_15708);
nand U16564 (N_16564,N_15134,N_15432);
xnor U16565 (N_16565,N_15049,N_15745);
xnor U16566 (N_16566,N_15558,N_15964);
or U16567 (N_16567,N_15656,N_15277);
xor U16568 (N_16568,N_15657,N_15311);
or U16569 (N_16569,N_15676,N_15542);
and U16570 (N_16570,N_15080,N_15619);
nor U16571 (N_16571,N_15224,N_15994);
and U16572 (N_16572,N_15537,N_15615);
xnor U16573 (N_16573,N_15282,N_15228);
nand U16574 (N_16574,N_15285,N_15626);
and U16575 (N_16575,N_15983,N_15330);
and U16576 (N_16576,N_15960,N_15412);
and U16577 (N_16577,N_15250,N_15578);
nand U16578 (N_16578,N_15600,N_15824);
nor U16579 (N_16579,N_15296,N_15379);
nand U16580 (N_16580,N_15543,N_15479);
or U16581 (N_16581,N_15462,N_15409);
and U16582 (N_16582,N_15550,N_15095);
nand U16583 (N_16583,N_15178,N_15860);
nor U16584 (N_16584,N_15932,N_15530);
or U16585 (N_16585,N_15608,N_15676);
nand U16586 (N_16586,N_15219,N_15078);
xor U16587 (N_16587,N_15782,N_15801);
nor U16588 (N_16588,N_15028,N_15680);
or U16589 (N_16589,N_15272,N_15690);
xor U16590 (N_16590,N_15153,N_15143);
xnor U16591 (N_16591,N_15899,N_15599);
nand U16592 (N_16592,N_15724,N_15974);
and U16593 (N_16593,N_15779,N_15009);
nand U16594 (N_16594,N_15874,N_15537);
xor U16595 (N_16595,N_15860,N_15941);
xnor U16596 (N_16596,N_15602,N_15003);
and U16597 (N_16597,N_15085,N_15908);
nor U16598 (N_16598,N_15699,N_15320);
or U16599 (N_16599,N_15524,N_15632);
nand U16600 (N_16600,N_15006,N_15845);
and U16601 (N_16601,N_15108,N_15638);
xor U16602 (N_16602,N_15232,N_15396);
and U16603 (N_16603,N_15892,N_15797);
xnor U16604 (N_16604,N_15976,N_15055);
nor U16605 (N_16605,N_15241,N_15619);
or U16606 (N_16606,N_15662,N_15990);
and U16607 (N_16607,N_15276,N_15966);
xor U16608 (N_16608,N_15724,N_15060);
and U16609 (N_16609,N_15078,N_15199);
nor U16610 (N_16610,N_15482,N_15104);
or U16611 (N_16611,N_15030,N_15559);
and U16612 (N_16612,N_15010,N_15380);
nor U16613 (N_16613,N_15932,N_15323);
nand U16614 (N_16614,N_15923,N_15036);
or U16615 (N_16615,N_15420,N_15878);
or U16616 (N_16616,N_15466,N_15591);
or U16617 (N_16617,N_15556,N_15951);
xor U16618 (N_16618,N_15161,N_15379);
or U16619 (N_16619,N_15680,N_15841);
nand U16620 (N_16620,N_15330,N_15708);
nand U16621 (N_16621,N_15303,N_15762);
and U16622 (N_16622,N_15223,N_15395);
nor U16623 (N_16623,N_15907,N_15160);
nand U16624 (N_16624,N_15908,N_15068);
and U16625 (N_16625,N_15686,N_15550);
nand U16626 (N_16626,N_15633,N_15817);
xor U16627 (N_16627,N_15632,N_15799);
and U16628 (N_16628,N_15707,N_15546);
xnor U16629 (N_16629,N_15983,N_15800);
nand U16630 (N_16630,N_15041,N_15714);
and U16631 (N_16631,N_15296,N_15692);
or U16632 (N_16632,N_15848,N_15924);
nor U16633 (N_16633,N_15701,N_15359);
xor U16634 (N_16634,N_15646,N_15044);
nor U16635 (N_16635,N_15205,N_15745);
and U16636 (N_16636,N_15523,N_15721);
xor U16637 (N_16637,N_15124,N_15856);
nand U16638 (N_16638,N_15699,N_15930);
xor U16639 (N_16639,N_15900,N_15651);
nand U16640 (N_16640,N_15175,N_15631);
or U16641 (N_16641,N_15343,N_15812);
or U16642 (N_16642,N_15524,N_15019);
and U16643 (N_16643,N_15757,N_15628);
or U16644 (N_16644,N_15722,N_15589);
nand U16645 (N_16645,N_15707,N_15025);
and U16646 (N_16646,N_15064,N_15542);
nand U16647 (N_16647,N_15536,N_15958);
nand U16648 (N_16648,N_15708,N_15977);
or U16649 (N_16649,N_15837,N_15312);
nand U16650 (N_16650,N_15940,N_15592);
nand U16651 (N_16651,N_15764,N_15704);
xor U16652 (N_16652,N_15496,N_15609);
nand U16653 (N_16653,N_15697,N_15337);
nand U16654 (N_16654,N_15958,N_15085);
nand U16655 (N_16655,N_15639,N_15276);
nand U16656 (N_16656,N_15985,N_15065);
or U16657 (N_16657,N_15267,N_15918);
nand U16658 (N_16658,N_15685,N_15538);
nor U16659 (N_16659,N_15537,N_15090);
nor U16660 (N_16660,N_15652,N_15956);
xnor U16661 (N_16661,N_15586,N_15420);
nor U16662 (N_16662,N_15670,N_15245);
and U16663 (N_16663,N_15344,N_15715);
xor U16664 (N_16664,N_15528,N_15068);
and U16665 (N_16665,N_15954,N_15163);
nand U16666 (N_16666,N_15657,N_15620);
xor U16667 (N_16667,N_15201,N_15685);
nor U16668 (N_16668,N_15448,N_15354);
xor U16669 (N_16669,N_15215,N_15036);
or U16670 (N_16670,N_15126,N_15358);
or U16671 (N_16671,N_15730,N_15116);
xor U16672 (N_16672,N_15471,N_15246);
nand U16673 (N_16673,N_15482,N_15100);
xor U16674 (N_16674,N_15838,N_15313);
nand U16675 (N_16675,N_15258,N_15242);
and U16676 (N_16676,N_15995,N_15199);
xnor U16677 (N_16677,N_15735,N_15832);
and U16678 (N_16678,N_15499,N_15168);
nor U16679 (N_16679,N_15393,N_15895);
xnor U16680 (N_16680,N_15361,N_15435);
nor U16681 (N_16681,N_15355,N_15416);
xor U16682 (N_16682,N_15236,N_15362);
and U16683 (N_16683,N_15065,N_15477);
nor U16684 (N_16684,N_15159,N_15368);
or U16685 (N_16685,N_15715,N_15813);
or U16686 (N_16686,N_15850,N_15562);
nand U16687 (N_16687,N_15278,N_15378);
nand U16688 (N_16688,N_15357,N_15260);
nand U16689 (N_16689,N_15761,N_15736);
nor U16690 (N_16690,N_15668,N_15207);
xor U16691 (N_16691,N_15857,N_15360);
nand U16692 (N_16692,N_15874,N_15218);
xor U16693 (N_16693,N_15586,N_15852);
and U16694 (N_16694,N_15057,N_15829);
nor U16695 (N_16695,N_15200,N_15417);
or U16696 (N_16696,N_15745,N_15980);
nand U16697 (N_16697,N_15145,N_15755);
xor U16698 (N_16698,N_15044,N_15585);
and U16699 (N_16699,N_15849,N_15328);
nand U16700 (N_16700,N_15153,N_15502);
or U16701 (N_16701,N_15356,N_15118);
xor U16702 (N_16702,N_15703,N_15149);
nor U16703 (N_16703,N_15653,N_15447);
nor U16704 (N_16704,N_15402,N_15772);
xnor U16705 (N_16705,N_15884,N_15220);
nor U16706 (N_16706,N_15855,N_15779);
nor U16707 (N_16707,N_15668,N_15739);
or U16708 (N_16708,N_15677,N_15521);
and U16709 (N_16709,N_15408,N_15353);
or U16710 (N_16710,N_15000,N_15821);
or U16711 (N_16711,N_15661,N_15991);
or U16712 (N_16712,N_15445,N_15299);
nor U16713 (N_16713,N_15885,N_15502);
nand U16714 (N_16714,N_15931,N_15143);
or U16715 (N_16715,N_15703,N_15191);
and U16716 (N_16716,N_15357,N_15121);
xor U16717 (N_16717,N_15667,N_15622);
nor U16718 (N_16718,N_15276,N_15700);
or U16719 (N_16719,N_15076,N_15044);
or U16720 (N_16720,N_15299,N_15886);
nand U16721 (N_16721,N_15546,N_15030);
or U16722 (N_16722,N_15561,N_15812);
or U16723 (N_16723,N_15329,N_15598);
or U16724 (N_16724,N_15449,N_15717);
xnor U16725 (N_16725,N_15954,N_15845);
nand U16726 (N_16726,N_15287,N_15292);
or U16727 (N_16727,N_15896,N_15492);
xor U16728 (N_16728,N_15813,N_15064);
or U16729 (N_16729,N_15868,N_15322);
or U16730 (N_16730,N_15855,N_15140);
nor U16731 (N_16731,N_15174,N_15091);
nor U16732 (N_16732,N_15113,N_15986);
or U16733 (N_16733,N_15375,N_15553);
or U16734 (N_16734,N_15748,N_15525);
or U16735 (N_16735,N_15848,N_15024);
and U16736 (N_16736,N_15141,N_15251);
nor U16737 (N_16737,N_15875,N_15567);
nand U16738 (N_16738,N_15494,N_15195);
xor U16739 (N_16739,N_15989,N_15963);
or U16740 (N_16740,N_15578,N_15014);
xnor U16741 (N_16741,N_15938,N_15672);
nand U16742 (N_16742,N_15917,N_15571);
or U16743 (N_16743,N_15380,N_15647);
xor U16744 (N_16744,N_15941,N_15661);
nor U16745 (N_16745,N_15512,N_15435);
and U16746 (N_16746,N_15784,N_15813);
nor U16747 (N_16747,N_15789,N_15275);
and U16748 (N_16748,N_15764,N_15758);
or U16749 (N_16749,N_15337,N_15890);
and U16750 (N_16750,N_15007,N_15063);
nor U16751 (N_16751,N_15721,N_15657);
nor U16752 (N_16752,N_15294,N_15915);
and U16753 (N_16753,N_15002,N_15026);
nor U16754 (N_16754,N_15369,N_15233);
and U16755 (N_16755,N_15848,N_15202);
or U16756 (N_16756,N_15909,N_15885);
nor U16757 (N_16757,N_15709,N_15949);
nor U16758 (N_16758,N_15638,N_15338);
or U16759 (N_16759,N_15666,N_15793);
and U16760 (N_16760,N_15555,N_15664);
and U16761 (N_16761,N_15905,N_15214);
nor U16762 (N_16762,N_15501,N_15741);
or U16763 (N_16763,N_15578,N_15773);
nand U16764 (N_16764,N_15632,N_15292);
or U16765 (N_16765,N_15704,N_15468);
or U16766 (N_16766,N_15662,N_15287);
or U16767 (N_16767,N_15237,N_15109);
nor U16768 (N_16768,N_15621,N_15731);
or U16769 (N_16769,N_15391,N_15394);
nor U16770 (N_16770,N_15325,N_15452);
nor U16771 (N_16771,N_15129,N_15223);
nor U16772 (N_16772,N_15489,N_15202);
or U16773 (N_16773,N_15550,N_15409);
xor U16774 (N_16774,N_15810,N_15377);
nand U16775 (N_16775,N_15869,N_15198);
or U16776 (N_16776,N_15829,N_15677);
nor U16777 (N_16777,N_15379,N_15158);
and U16778 (N_16778,N_15234,N_15410);
or U16779 (N_16779,N_15165,N_15200);
and U16780 (N_16780,N_15207,N_15670);
and U16781 (N_16781,N_15633,N_15945);
xnor U16782 (N_16782,N_15108,N_15382);
nor U16783 (N_16783,N_15298,N_15870);
or U16784 (N_16784,N_15122,N_15790);
xor U16785 (N_16785,N_15028,N_15319);
or U16786 (N_16786,N_15104,N_15053);
nand U16787 (N_16787,N_15949,N_15270);
or U16788 (N_16788,N_15689,N_15149);
xnor U16789 (N_16789,N_15392,N_15409);
xor U16790 (N_16790,N_15758,N_15965);
nor U16791 (N_16791,N_15955,N_15119);
nand U16792 (N_16792,N_15918,N_15161);
or U16793 (N_16793,N_15283,N_15772);
and U16794 (N_16794,N_15199,N_15667);
nor U16795 (N_16795,N_15790,N_15964);
nand U16796 (N_16796,N_15717,N_15517);
xnor U16797 (N_16797,N_15406,N_15341);
or U16798 (N_16798,N_15919,N_15506);
nor U16799 (N_16799,N_15714,N_15311);
xor U16800 (N_16800,N_15902,N_15728);
xor U16801 (N_16801,N_15859,N_15280);
xnor U16802 (N_16802,N_15139,N_15181);
xnor U16803 (N_16803,N_15066,N_15867);
or U16804 (N_16804,N_15850,N_15675);
xnor U16805 (N_16805,N_15379,N_15210);
nor U16806 (N_16806,N_15069,N_15061);
nand U16807 (N_16807,N_15262,N_15525);
xor U16808 (N_16808,N_15899,N_15338);
xor U16809 (N_16809,N_15184,N_15487);
nor U16810 (N_16810,N_15294,N_15942);
nor U16811 (N_16811,N_15401,N_15331);
or U16812 (N_16812,N_15676,N_15749);
xor U16813 (N_16813,N_15870,N_15233);
or U16814 (N_16814,N_15535,N_15138);
or U16815 (N_16815,N_15365,N_15293);
xor U16816 (N_16816,N_15982,N_15297);
and U16817 (N_16817,N_15804,N_15272);
nand U16818 (N_16818,N_15810,N_15058);
nand U16819 (N_16819,N_15568,N_15349);
or U16820 (N_16820,N_15438,N_15534);
nand U16821 (N_16821,N_15741,N_15092);
or U16822 (N_16822,N_15605,N_15015);
or U16823 (N_16823,N_15349,N_15615);
nor U16824 (N_16824,N_15974,N_15265);
and U16825 (N_16825,N_15773,N_15279);
or U16826 (N_16826,N_15302,N_15243);
and U16827 (N_16827,N_15210,N_15408);
nor U16828 (N_16828,N_15713,N_15321);
xor U16829 (N_16829,N_15162,N_15679);
xnor U16830 (N_16830,N_15084,N_15759);
nand U16831 (N_16831,N_15597,N_15814);
xnor U16832 (N_16832,N_15248,N_15320);
nand U16833 (N_16833,N_15069,N_15355);
nand U16834 (N_16834,N_15050,N_15660);
nor U16835 (N_16835,N_15423,N_15833);
or U16836 (N_16836,N_15537,N_15735);
or U16837 (N_16837,N_15416,N_15336);
nand U16838 (N_16838,N_15433,N_15601);
xnor U16839 (N_16839,N_15149,N_15297);
nand U16840 (N_16840,N_15716,N_15672);
xnor U16841 (N_16841,N_15940,N_15926);
nor U16842 (N_16842,N_15901,N_15710);
xnor U16843 (N_16843,N_15046,N_15663);
and U16844 (N_16844,N_15498,N_15753);
nor U16845 (N_16845,N_15355,N_15178);
or U16846 (N_16846,N_15531,N_15732);
xnor U16847 (N_16847,N_15159,N_15156);
nand U16848 (N_16848,N_15382,N_15692);
or U16849 (N_16849,N_15025,N_15558);
nand U16850 (N_16850,N_15793,N_15621);
and U16851 (N_16851,N_15022,N_15593);
xor U16852 (N_16852,N_15304,N_15774);
or U16853 (N_16853,N_15652,N_15498);
xnor U16854 (N_16854,N_15595,N_15324);
nor U16855 (N_16855,N_15441,N_15705);
and U16856 (N_16856,N_15993,N_15603);
nor U16857 (N_16857,N_15345,N_15306);
nand U16858 (N_16858,N_15882,N_15108);
nor U16859 (N_16859,N_15554,N_15979);
or U16860 (N_16860,N_15333,N_15403);
and U16861 (N_16861,N_15060,N_15424);
nand U16862 (N_16862,N_15202,N_15803);
nor U16863 (N_16863,N_15696,N_15111);
nor U16864 (N_16864,N_15497,N_15405);
xnor U16865 (N_16865,N_15798,N_15503);
xnor U16866 (N_16866,N_15363,N_15411);
nor U16867 (N_16867,N_15628,N_15551);
nor U16868 (N_16868,N_15370,N_15861);
xnor U16869 (N_16869,N_15091,N_15241);
nand U16870 (N_16870,N_15222,N_15876);
nand U16871 (N_16871,N_15103,N_15400);
nor U16872 (N_16872,N_15226,N_15269);
nor U16873 (N_16873,N_15748,N_15841);
or U16874 (N_16874,N_15583,N_15421);
nor U16875 (N_16875,N_15680,N_15494);
nand U16876 (N_16876,N_15952,N_15627);
nor U16877 (N_16877,N_15088,N_15477);
xor U16878 (N_16878,N_15840,N_15629);
xor U16879 (N_16879,N_15956,N_15561);
and U16880 (N_16880,N_15325,N_15499);
nand U16881 (N_16881,N_15095,N_15125);
nand U16882 (N_16882,N_15121,N_15108);
xnor U16883 (N_16883,N_15430,N_15542);
or U16884 (N_16884,N_15699,N_15534);
or U16885 (N_16885,N_15161,N_15701);
nand U16886 (N_16886,N_15560,N_15419);
and U16887 (N_16887,N_15891,N_15511);
nand U16888 (N_16888,N_15850,N_15558);
or U16889 (N_16889,N_15495,N_15532);
xor U16890 (N_16890,N_15930,N_15898);
or U16891 (N_16891,N_15376,N_15015);
nand U16892 (N_16892,N_15392,N_15551);
nand U16893 (N_16893,N_15550,N_15080);
and U16894 (N_16894,N_15716,N_15836);
or U16895 (N_16895,N_15552,N_15925);
nand U16896 (N_16896,N_15932,N_15238);
nand U16897 (N_16897,N_15378,N_15486);
nor U16898 (N_16898,N_15743,N_15724);
and U16899 (N_16899,N_15194,N_15033);
nand U16900 (N_16900,N_15415,N_15315);
nor U16901 (N_16901,N_15094,N_15680);
nand U16902 (N_16902,N_15634,N_15512);
or U16903 (N_16903,N_15049,N_15122);
nor U16904 (N_16904,N_15961,N_15998);
nand U16905 (N_16905,N_15116,N_15213);
and U16906 (N_16906,N_15995,N_15761);
or U16907 (N_16907,N_15831,N_15320);
or U16908 (N_16908,N_15927,N_15406);
or U16909 (N_16909,N_15565,N_15875);
nor U16910 (N_16910,N_15446,N_15973);
nor U16911 (N_16911,N_15967,N_15116);
nand U16912 (N_16912,N_15993,N_15717);
or U16913 (N_16913,N_15752,N_15874);
nand U16914 (N_16914,N_15939,N_15568);
nor U16915 (N_16915,N_15419,N_15509);
or U16916 (N_16916,N_15194,N_15979);
or U16917 (N_16917,N_15451,N_15464);
and U16918 (N_16918,N_15271,N_15546);
or U16919 (N_16919,N_15944,N_15854);
and U16920 (N_16920,N_15459,N_15662);
nand U16921 (N_16921,N_15329,N_15613);
and U16922 (N_16922,N_15651,N_15872);
nor U16923 (N_16923,N_15808,N_15703);
or U16924 (N_16924,N_15464,N_15387);
nand U16925 (N_16925,N_15619,N_15650);
xnor U16926 (N_16926,N_15761,N_15871);
xor U16927 (N_16927,N_15974,N_15650);
and U16928 (N_16928,N_15198,N_15960);
nand U16929 (N_16929,N_15697,N_15745);
or U16930 (N_16930,N_15198,N_15272);
and U16931 (N_16931,N_15348,N_15007);
and U16932 (N_16932,N_15743,N_15270);
xnor U16933 (N_16933,N_15028,N_15519);
and U16934 (N_16934,N_15641,N_15783);
and U16935 (N_16935,N_15689,N_15986);
nor U16936 (N_16936,N_15412,N_15384);
xnor U16937 (N_16937,N_15647,N_15066);
nor U16938 (N_16938,N_15925,N_15172);
nand U16939 (N_16939,N_15822,N_15485);
nand U16940 (N_16940,N_15945,N_15121);
nor U16941 (N_16941,N_15881,N_15843);
xnor U16942 (N_16942,N_15625,N_15622);
nor U16943 (N_16943,N_15044,N_15249);
and U16944 (N_16944,N_15414,N_15113);
and U16945 (N_16945,N_15937,N_15292);
and U16946 (N_16946,N_15263,N_15254);
nor U16947 (N_16947,N_15040,N_15496);
and U16948 (N_16948,N_15018,N_15695);
and U16949 (N_16949,N_15229,N_15760);
nand U16950 (N_16950,N_15325,N_15765);
xnor U16951 (N_16951,N_15680,N_15632);
xor U16952 (N_16952,N_15204,N_15107);
xnor U16953 (N_16953,N_15583,N_15525);
xor U16954 (N_16954,N_15512,N_15949);
nand U16955 (N_16955,N_15651,N_15158);
and U16956 (N_16956,N_15684,N_15270);
and U16957 (N_16957,N_15921,N_15672);
nor U16958 (N_16958,N_15677,N_15134);
nor U16959 (N_16959,N_15962,N_15953);
nand U16960 (N_16960,N_15305,N_15219);
xnor U16961 (N_16961,N_15373,N_15314);
or U16962 (N_16962,N_15046,N_15903);
nor U16963 (N_16963,N_15175,N_15253);
nand U16964 (N_16964,N_15183,N_15729);
nor U16965 (N_16965,N_15339,N_15510);
or U16966 (N_16966,N_15462,N_15021);
nand U16967 (N_16967,N_15397,N_15473);
xnor U16968 (N_16968,N_15075,N_15220);
and U16969 (N_16969,N_15722,N_15800);
or U16970 (N_16970,N_15962,N_15832);
and U16971 (N_16971,N_15073,N_15695);
xnor U16972 (N_16972,N_15589,N_15723);
nor U16973 (N_16973,N_15211,N_15615);
nor U16974 (N_16974,N_15115,N_15367);
nor U16975 (N_16975,N_15712,N_15604);
xor U16976 (N_16976,N_15749,N_15157);
nor U16977 (N_16977,N_15033,N_15116);
xor U16978 (N_16978,N_15994,N_15024);
and U16979 (N_16979,N_15495,N_15924);
and U16980 (N_16980,N_15460,N_15877);
or U16981 (N_16981,N_15247,N_15563);
and U16982 (N_16982,N_15944,N_15058);
and U16983 (N_16983,N_15953,N_15289);
xor U16984 (N_16984,N_15145,N_15491);
nand U16985 (N_16985,N_15241,N_15181);
nand U16986 (N_16986,N_15079,N_15382);
nor U16987 (N_16987,N_15464,N_15115);
nor U16988 (N_16988,N_15023,N_15728);
xnor U16989 (N_16989,N_15004,N_15537);
and U16990 (N_16990,N_15136,N_15346);
nor U16991 (N_16991,N_15101,N_15072);
xnor U16992 (N_16992,N_15848,N_15951);
nor U16993 (N_16993,N_15104,N_15175);
and U16994 (N_16994,N_15741,N_15209);
nor U16995 (N_16995,N_15582,N_15520);
nor U16996 (N_16996,N_15821,N_15707);
and U16997 (N_16997,N_15887,N_15132);
and U16998 (N_16998,N_15032,N_15859);
nand U16999 (N_16999,N_15771,N_15282);
or U17000 (N_17000,N_16649,N_16712);
nor U17001 (N_17001,N_16382,N_16290);
nor U17002 (N_17002,N_16367,N_16495);
nand U17003 (N_17003,N_16178,N_16188);
nor U17004 (N_17004,N_16944,N_16650);
xnor U17005 (N_17005,N_16301,N_16221);
and U17006 (N_17006,N_16017,N_16139);
and U17007 (N_17007,N_16880,N_16566);
and U17008 (N_17008,N_16969,N_16397);
or U17009 (N_17009,N_16774,N_16304);
nor U17010 (N_17010,N_16825,N_16204);
nand U17011 (N_17011,N_16269,N_16048);
or U17012 (N_17012,N_16603,N_16016);
nand U17013 (N_17013,N_16350,N_16279);
nor U17014 (N_17014,N_16995,N_16539);
and U17015 (N_17015,N_16059,N_16779);
nor U17016 (N_17016,N_16552,N_16896);
nor U17017 (N_17017,N_16671,N_16079);
and U17018 (N_17018,N_16064,N_16713);
nor U17019 (N_17019,N_16311,N_16445);
xnor U17020 (N_17020,N_16665,N_16427);
and U17021 (N_17021,N_16353,N_16099);
nor U17022 (N_17022,N_16676,N_16717);
and U17023 (N_17023,N_16610,N_16894);
nor U17024 (N_17024,N_16757,N_16878);
nand U17025 (N_17025,N_16722,N_16366);
xnor U17026 (N_17026,N_16956,N_16897);
or U17027 (N_17027,N_16881,N_16669);
or U17028 (N_17028,N_16883,N_16563);
or U17029 (N_17029,N_16947,N_16836);
or U17030 (N_17030,N_16497,N_16689);
or U17031 (N_17031,N_16082,N_16095);
nor U17032 (N_17032,N_16511,N_16483);
nand U17033 (N_17033,N_16124,N_16625);
and U17034 (N_17034,N_16485,N_16159);
xor U17035 (N_17035,N_16818,N_16474);
nand U17036 (N_17036,N_16443,N_16068);
or U17037 (N_17037,N_16044,N_16027);
and U17038 (N_17038,N_16292,N_16582);
nand U17039 (N_17039,N_16823,N_16903);
nor U17040 (N_17040,N_16820,N_16954);
nor U17041 (N_17041,N_16280,N_16130);
and U17042 (N_17042,N_16272,N_16096);
nor U17043 (N_17043,N_16386,N_16058);
nor U17044 (N_17044,N_16614,N_16715);
and U17045 (N_17045,N_16472,N_16150);
or U17046 (N_17046,N_16385,N_16329);
xnor U17047 (N_17047,N_16812,N_16768);
and U17048 (N_17048,N_16803,N_16977);
nand U17049 (N_17049,N_16583,N_16761);
or U17050 (N_17050,N_16586,N_16617);
and U17051 (N_17051,N_16448,N_16576);
or U17052 (N_17052,N_16487,N_16642);
or U17053 (N_17053,N_16160,N_16305);
xor U17054 (N_17054,N_16358,N_16673);
nor U17055 (N_17055,N_16006,N_16907);
nor U17056 (N_17056,N_16704,N_16293);
and U17057 (N_17057,N_16807,N_16515);
or U17058 (N_17058,N_16966,N_16257);
or U17059 (N_17059,N_16478,N_16022);
and U17060 (N_17060,N_16776,N_16904);
nor U17061 (N_17061,N_16446,N_16653);
nand U17062 (N_17062,N_16297,N_16683);
or U17063 (N_17063,N_16402,N_16932);
nor U17064 (N_17064,N_16055,N_16876);
or U17065 (N_17065,N_16363,N_16602);
nand U17066 (N_17066,N_16543,N_16937);
xnor U17067 (N_17067,N_16503,N_16829);
and U17068 (N_17068,N_16524,N_16664);
nand U17069 (N_17069,N_16251,N_16789);
nor U17070 (N_17070,N_16200,N_16192);
nand U17071 (N_17071,N_16201,N_16855);
xor U17072 (N_17072,N_16077,N_16113);
xor U17073 (N_17073,N_16641,N_16435);
xnor U17074 (N_17074,N_16481,N_16107);
nor U17075 (N_17075,N_16737,N_16249);
nor U17076 (N_17076,N_16444,N_16615);
nor U17077 (N_17077,N_16106,N_16853);
xor U17078 (N_17078,N_16644,N_16152);
xnor U17079 (N_17079,N_16607,N_16281);
xnor U17080 (N_17080,N_16415,N_16943);
nor U17081 (N_17081,N_16174,N_16838);
nand U17082 (N_17082,N_16869,N_16473);
xnor U17083 (N_17083,N_16529,N_16655);
nand U17084 (N_17084,N_16199,N_16639);
xnor U17085 (N_17085,N_16828,N_16758);
and U17086 (N_17086,N_16522,N_16449);
nand U17087 (N_17087,N_16800,N_16731);
xor U17088 (N_17088,N_16754,N_16685);
nand U17089 (N_17089,N_16792,N_16383);
or U17090 (N_17090,N_16327,N_16310);
or U17091 (N_17091,N_16764,N_16008);
nor U17092 (N_17092,N_16087,N_16451);
nor U17093 (N_17093,N_16744,N_16002);
or U17094 (N_17094,N_16811,N_16061);
nand U17095 (N_17095,N_16624,N_16674);
and U17096 (N_17096,N_16875,N_16960);
and U17097 (N_17097,N_16765,N_16700);
xnor U17098 (N_17098,N_16354,N_16729);
nor U17099 (N_17099,N_16025,N_16767);
and U17100 (N_17100,N_16718,N_16805);
or U17101 (N_17101,N_16546,N_16787);
nor U17102 (N_17102,N_16179,N_16384);
nand U17103 (N_17103,N_16074,N_16263);
and U17104 (N_17104,N_16306,N_16231);
nor U17105 (N_17105,N_16927,N_16637);
nand U17106 (N_17106,N_16373,N_16066);
nor U17107 (N_17107,N_16330,N_16821);
and U17108 (N_17108,N_16234,N_16548);
and U17109 (N_17109,N_16185,N_16656);
xnor U17110 (N_17110,N_16010,N_16030);
nand U17111 (N_17111,N_16773,N_16781);
or U17112 (N_17112,N_16813,N_16312);
and U17113 (N_17113,N_16042,N_16227);
nor U17114 (N_17114,N_16997,N_16344);
and U17115 (N_17115,N_16100,N_16756);
xor U17116 (N_17116,N_16748,N_16725);
or U17117 (N_17117,N_16162,N_16906);
or U17118 (N_17118,N_16108,N_16867);
xnor U17119 (N_17119,N_16392,N_16950);
nor U17120 (N_17120,N_16168,N_16378);
xor U17121 (N_17121,N_16158,N_16532);
nand U17122 (N_17122,N_16254,N_16086);
nor U17123 (N_17123,N_16403,N_16600);
nor U17124 (N_17124,N_16206,N_16952);
nor U17125 (N_17125,N_16136,N_16464);
and U17126 (N_17126,N_16351,N_16049);
and U17127 (N_17127,N_16544,N_16238);
xnor U17128 (N_17128,N_16479,N_16628);
nand U17129 (N_17129,N_16870,N_16285);
nor U17130 (N_17130,N_16347,N_16418);
or U17131 (N_17131,N_16265,N_16413);
or U17132 (N_17132,N_16015,N_16597);
nor U17133 (N_17133,N_16612,N_16393);
xor U17134 (N_17134,N_16680,N_16535);
and U17135 (N_17135,N_16173,N_16577);
nand U17136 (N_17136,N_16195,N_16315);
nand U17137 (N_17137,N_16341,N_16357);
nor U17138 (N_17138,N_16573,N_16459);
xor U17139 (N_17139,N_16585,N_16250);
nand U17140 (N_17140,N_16556,N_16939);
nand U17141 (N_17141,N_16255,N_16802);
and U17142 (N_17142,N_16916,N_16587);
nor U17143 (N_17143,N_16666,N_16203);
and U17144 (N_17144,N_16321,N_16694);
or U17145 (N_17145,N_16619,N_16493);
xor U17146 (N_17146,N_16376,N_16052);
nand U17147 (N_17147,N_16609,N_16958);
and U17148 (N_17148,N_16370,N_16711);
nor U17149 (N_17149,N_16236,N_16699);
or U17150 (N_17150,N_16390,N_16975);
or U17151 (N_17151,N_16430,N_16660);
or U17152 (N_17152,N_16578,N_16986);
nand U17153 (N_17153,N_16364,N_16243);
or U17154 (N_17154,N_16572,N_16885);
nor U17155 (N_17155,N_16678,N_16252);
nand U17156 (N_17156,N_16194,N_16494);
nor U17157 (N_17157,N_16581,N_16702);
nor U17158 (N_17158,N_16338,N_16088);
nor U17159 (N_17159,N_16164,N_16147);
or U17160 (N_17160,N_16466,N_16468);
and U17161 (N_17161,N_16736,N_16777);
xor U17162 (N_17162,N_16374,N_16659);
and U17163 (N_17163,N_16191,N_16510);
or U17164 (N_17164,N_16930,N_16187);
nand U17165 (N_17165,N_16300,N_16491);
xor U17166 (N_17166,N_16984,N_16861);
or U17167 (N_17167,N_16873,N_16111);
and U17168 (N_17168,N_16102,N_16240);
or U17169 (N_17169,N_16295,N_16962);
xor U17170 (N_17170,N_16723,N_16830);
and U17171 (N_17171,N_16901,N_16824);
or U17172 (N_17172,N_16965,N_16706);
and U17173 (N_17173,N_16230,N_16193);
and U17174 (N_17174,N_16452,N_16317);
nand U17175 (N_17175,N_16499,N_16224);
and U17176 (N_17176,N_16313,N_16819);
nor U17177 (N_17177,N_16163,N_16527);
nand U17178 (N_17178,N_16133,N_16772);
or U17179 (N_17179,N_16740,N_16925);
and U17180 (N_17180,N_16902,N_16069);
nor U17181 (N_17181,N_16154,N_16766);
and U17182 (N_17182,N_16601,N_16946);
and U17183 (N_17183,N_16616,N_16851);
nand U17184 (N_17184,N_16982,N_16661);
nand U17185 (N_17185,N_16760,N_16116);
nand U17186 (N_17186,N_16438,N_16567);
or U17187 (N_17187,N_16793,N_16126);
xnor U17188 (N_17188,N_16047,N_16604);
or U17189 (N_17189,N_16498,N_16171);
or U17190 (N_17190,N_16410,N_16755);
and U17191 (N_17191,N_16319,N_16198);
or U17192 (N_17192,N_16634,N_16229);
or U17193 (N_17193,N_16225,N_16505);
and U17194 (N_17194,N_16595,N_16273);
nand U17195 (N_17195,N_16613,N_16127);
xor U17196 (N_17196,N_16749,N_16226);
nand U17197 (N_17197,N_16007,N_16037);
nor U17198 (N_17198,N_16233,N_16588);
and U17199 (N_17199,N_16908,N_16148);
or U17200 (N_17200,N_16530,N_16559);
nor U17201 (N_17201,N_16672,N_16092);
or U17202 (N_17202,N_16284,N_16611);
xor U17203 (N_17203,N_16214,N_16541);
nand U17204 (N_17204,N_16020,N_16633);
or U17205 (N_17205,N_16286,N_16425);
or U17206 (N_17206,N_16399,N_16019);
or U17207 (N_17207,N_16120,N_16089);
xnor U17208 (N_17208,N_16892,N_16372);
nor U17209 (N_17209,N_16118,N_16176);
or U17210 (N_17210,N_16888,N_16647);
and U17211 (N_17211,N_16558,N_16913);
nor U17212 (N_17212,N_16643,N_16788);
or U17213 (N_17213,N_16412,N_16938);
nand U17214 (N_17214,N_16112,N_16850);
nor U17215 (N_17215,N_16291,N_16935);
nor U17216 (N_17216,N_16978,N_16218);
xor U17217 (N_17217,N_16463,N_16332);
nor U17218 (N_17218,N_16062,N_16771);
and U17219 (N_17219,N_16097,N_16668);
and U17220 (N_17220,N_16342,N_16245);
nor U17221 (N_17221,N_16844,N_16899);
nand U17222 (N_17222,N_16730,N_16910);
or U17223 (N_17223,N_16887,N_16557);
or U17224 (N_17224,N_16770,N_16627);
nand U17225 (N_17225,N_16554,N_16705);
nand U17226 (N_17226,N_16038,N_16076);
and U17227 (N_17227,N_16323,N_16396);
or U17228 (N_17228,N_16687,N_16457);
or U17229 (N_17229,N_16362,N_16734);
or U17230 (N_17230,N_16985,N_16921);
or U17231 (N_17231,N_16423,N_16307);
xnor U17232 (N_17232,N_16228,N_16436);
nand U17233 (N_17233,N_16667,N_16941);
xnor U17234 (N_17234,N_16398,N_16948);
xor U17235 (N_17235,N_16769,N_16381);
nor U17236 (N_17236,N_16677,N_16889);
or U17237 (N_17237,N_16465,N_16691);
nand U17238 (N_17238,N_16205,N_16798);
nand U17239 (N_17239,N_16138,N_16222);
nand U17240 (N_17240,N_16506,N_16075);
nor U17241 (N_17241,N_16974,N_16041);
xor U17242 (N_17242,N_16365,N_16360);
nor U17243 (N_17243,N_16476,N_16837);
or U17244 (N_17244,N_16964,N_16697);
nor U17245 (N_17245,N_16931,N_16103);
nor U17246 (N_17246,N_16545,N_16128);
xor U17247 (N_17247,N_16743,N_16945);
and U17248 (N_17248,N_16400,N_16936);
and U17249 (N_17249,N_16630,N_16167);
xnor U17250 (N_17250,N_16727,N_16686);
or U17251 (N_17251,N_16859,N_16652);
and U17252 (N_17252,N_16791,N_16657);
and U17253 (N_17253,N_16504,N_16496);
nand U17254 (N_17254,N_16745,N_16900);
or U17255 (N_17255,N_16141,N_16520);
or U17256 (N_17256,N_16453,N_16560);
and U17257 (N_17257,N_16244,N_16267);
nor U17258 (N_17258,N_16967,N_16843);
nor U17259 (N_17259,N_16209,N_16131);
and U17260 (N_17260,N_16161,N_16458);
nand U17261 (N_17261,N_16085,N_16988);
nor U17262 (N_17262,N_16738,N_16114);
and U17263 (N_17263,N_16762,N_16721);
and U17264 (N_17264,N_16303,N_16388);
and U17265 (N_17265,N_16379,N_16051);
nor U17266 (N_17266,N_16441,N_16759);
nor U17267 (N_17267,N_16434,N_16797);
or U17268 (N_17268,N_16346,N_16999);
and U17269 (N_17269,N_16863,N_16924);
nand U17270 (N_17270,N_16929,N_16909);
nor U17271 (N_17271,N_16839,N_16013);
nor U17272 (N_17272,N_16957,N_16153);
xor U17273 (N_17273,N_16884,N_16011);
and U17274 (N_17274,N_16518,N_16345);
and U17275 (N_17275,N_16440,N_16596);
or U17276 (N_17276,N_16816,N_16296);
and U17277 (N_17277,N_16215,N_16632);
and U17278 (N_17278,N_16809,N_16324);
xnor U17279 (N_17279,N_16698,N_16872);
or U17280 (N_17280,N_16814,N_16923);
nor U17281 (N_17281,N_16523,N_16421);
and U17282 (N_17282,N_16822,N_16490);
or U17283 (N_17283,N_16322,N_16395);
nand U17284 (N_17284,N_16288,N_16155);
nand U17285 (N_17285,N_16747,N_16070);
nand U17286 (N_17286,N_16001,N_16220);
nor U17287 (N_17287,N_16886,N_16857);
or U17288 (N_17288,N_16394,N_16253);
xnor U17289 (N_17289,N_16431,N_16963);
nor U17290 (N_17290,N_16592,N_16391);
or U17291 (N_17291,N_16140,N_16094);
nand U17292 (N_17292,N_16484,N_16340);
and U17293 (N_17293,N_16682,N_16651);
or U17294 (N_17294,N_16531,N_16258);
nor U17295 (N_17295,N_16517,N_16003);
xor U17296 (N_17296,N_16259,N_16898);
or U17297 (N_17297,N_16570,N_16123);
nand U17298 (N_17298,N_16693,N_16039);
nor U17299 (N_17299,N_16550,N_16580);
xnor U17300 (N_17300,N_16084,N_16270);
nor U17301 (N_17301,N_16810,N_16842);
xor U17302 (N_17302,N_16419,N_16264);
and U17303 (N_17303,N_16424,N_16149);
nand U17304 (N_17304,N_16890,N_16513);
nand U17305 (N_17305,N_16492,N_16993);
nor U17306 (N_17306,N_16865,N_16420);
nor U17307 (N_17307,N_16670,N_16368);
or U17308 (N_17308,N_16590,N_16182);
and U17309 (N_17309,N_16063,N_16626);
xor U17310 (N_17310,N_16202,N_16638);
nor U17311 (N_17311,N_16034,N_16605);
and U17312 (N_17312,N_16785,N_16328);
xor U17313 (N_17313,N_16598,N_16752);
and U17314 (N_17314,N_16146,N_16794);
nand U17315 (N_17315,N_16282,N_16940);
or U17316 (N_17316,N_16115,N_16623);
and U17317 (N_17317,N_16525,N_16780);
nand U17318 (N_17318,N_16692,N_16060);
or U17319 (N_17319,N_16914,N_16636);
and U17320 (N_17320,N_16043,N_16417);
nor U17321 (N_17321,N_16143,N_16663);
nand U17322 (N_17322,N_16428,N_16467);
nor U17323 (N_17323,N_16833,N_16742);
xnor U17324 (N_17324,N_16858,N_16714);
nor U17325 (N_17325,N_16004,N_16121);
nand U17326 (N_17326,N_16973,N_16336);
nor U17327 (N_17327,N_16509,N_16868);
nor U17328 (N_17328,N_16181,N_16561);
nand U17329 (N_17329,N_16646,N_16389);
or U17330 (N_17330,N_16720,N_16083);
nand U17331 (N_17331,N_16959,N_16500);
and U17332 (N_17332,N_16536,N_16594);
nor U17333 (N_17333,N_16246,N_16056);
or U17334 (N_17334,N_16864,N_16411);
nor U17335 (N_17335,N_16471,N_16211);
nand U17336 (N_17336,N_16408,N_16526);
nand U17337 (N_17337,N_16537,N_16470);
nand U17338 (N_17338,N_16648,N_16790);
or U17339 (N_17339,N_16835,N_16710);
xnor U17340 (N_17340,N_16090,N_16054);
nand U17341 (N_17341,N_16157,N_16186);
nand U17342 (N_17342,N_16401,N_16387);
and U17343 (N_17343,N_16409,N_16309);
nor U17344 (N_17344,N_16169,N_16934);
nor U17345 (N_17345,N_16343,N_16289);
nand U17346 (N_17346,N_16972,N_16568);
and U17347 (N_17347,N_16562,N_16553);
or U17348 (N_17348,N_16407,N_16675);
or U17349 (N_17349,N_16283,N_16050);
and U17350 (N_17350,N_16276,N_16516);
and U17351 (N_17351,N_16569,N_16980);
or U17352 (N_17352,N_16012,N_16369);
and U17353 (N_17353,N_16105,N_16860);
or U17354 (N_17354,N_16912,N_16018);
and U17355 (N_17355,N_16949,N_16450);
or U17356 (N_17356,N_16442,N_16308);
nor U17357 (N_17357,N_16654,N_16455);
nor U17358 (N_17358,N_16156,N_16073);
or U17359 (N_17359,N_16029,N_16356);
or U17360 (N_17360,N_16057,N_16477);
xnor U17361 (N_17361,N_16071,N_16521);
or U17362 (N_17362,N_16922,N_16219);
nand U17363 (N_17363,N_16905,N_16707);
nand U17364 (N_17364,N_16796,N_16429);
nand U17365 (N_17365,N_16662,N_16987);
or U17366 (N_17366,N_16184,N_16801);
xnor U17367 (N_17367,N_16348,N_16278);
and U17368 (N_17368,N_16508,N_16591);
xor U17369 (N_17369,N_16298,N_16845);
xor U17370 (N_17370,N_16528,N_16533);
or U17371 (N_17371,N_16926,N_16658);
and U17372 (N_17372,N_16942,N_16416);
nor U17373 (N_17373,N_16331,N_16237);
or U17374 (N_17374,N_16507,N_16316);
or U17375 (N_17375,N_16728,N_16489);
nor U17376 (N_17376,N_16165,N_16847);
nor U17377 (N_17377,N_16584,N_16684);
nor U17378 (N_17378,N_16726,N_16262);
and U17379 (N_17379,N_16826,N_16294);
and U17380 (N_17380,N_16241,N_16998);
nor U17381 (N_17381,N_16891,N_16832);
nor U17382 (N_17382,N_16551,N_16917);
or U17383 (N_17383,N_16815,N_16799);
or U17384 (N_17384,N_16349,N_16197);
nor U17385 (N_17385,N_16724,N_16996);
nand U17386 (N_17386,N_16314,N_16575);
xor U17387 (N_17387,N_16433,N_16690);
and U17388 (N_17388,N_16239,N_16189);
nand U17389 (N_17389,N_16122,N_16920);
xnor U17390 (N_17390,N_16260,N_16232);
or U17391 (N_17391,N_16117,N_16877);
or U17392 (N_17392,N_16093,N_16166);
xnor U17393 (N_17393,N_16629,N_16579);
nand U17394 (N_17394,N_16422,N_16091);
nor U17395 (N_17395,N_16716,N_16961);
xnor U17396 (N_17396,N_16359,N_16621);
and U17397 (N_17397,N_16751,N_16437);
nor U17398 (N_17398,N_16512,N_16404);
nand U17399 (N_17399,N_16318,N_16024);
xor U17400 (N_17400,N_16928,N_16971);
xnor U17401 (N_17401,N_16361,N_16371);
and U17402 (N_17402,N_16145,N_16299);
nand U17403 (N_17403,N_16196,N_16172);
nor U17404 (N_17404,N_16775,N_16854);
xnor U17405 (N_17405,N_16135,N_16696);
nor U17406 (N_17406,N_16739,N_16134);
or U17407 (N_17407,N_16635,N_16334);
and U17408 (N_17408,N_16849,N_16708);
nor U17409 (N_17409,N_16337,N_16599);
xor U17410 (N_17410,N_16574,N_16514);
nand U17411 (N_17411,N_16709,N_16036);
nor U17412 (N_17412,N_16593,N_16645);
nor U17413 (N_17413,N_16856,N_16979);
nor U17414 (N_17414,N_16033,N_16763);
xnor U17415 (N_17415,N_16439,N_16866);
xor U17416 (N_17416,N_16480,N_16565);
or U17417 (N_17417,N_16778,N_16137);
nand U17418 (N_17418,N_16486,N_16989);
nand U17419 (N_17419,N_16175,N_16983);
and U17420 (N_17420,N_16072,N_16933);
nand U17421 (N_17421,N_16302,N_16538);
xnor U17422 (N_17422,N_16065,N_16848);
xnor U17423 (N_17423,N_16217,N_16101);
xor U17424 (N_17424,N_16000,N_16426);
or U17425 (N_17425,N_16895,N_16735);
and U17426 (N_17426,N_16753,N_16028);
nor U17427 (N_17427,N_16475,N_16242);
nor U17428 (N_17428,N_16414,N_16216);
nor U17429 (N_17429,N_16879,N_16783);
nor U17430 (N_17430,N_16080,N_16271);
and U17431 (N_17431,N_16447,N_16009);
xnor U17432 (N_17432,N_16352,N_16732);
nor U17433 (N_17433,N_16208,N_16032);
xnor U17434 (N_17434,N_16968,N_16031);
xnor U17435 (N_17435,N_16213,N_16547);
nand U17436 (N_17436,N_16461,N_16488);
nor U17437 (N_17437,N_16631,N_16098);
and U17438 (N_17438,N_16786,N_16992);
or U17439 (N_17439,N_16951,N_16874);
nand U17440 (N_17440,N_16119,N_16335);
xnor U17441 (N_17441,N_16882,N_16741);
nand U17442 (N_17442,N_16564,N_16406);
and U17443 (N_17443,N_16795,N_16223);
and U17444 (N_17444,N_16235,N_16784);
or U17445 (N_17445,N_16377,N_16405);
and U17446 (N_17446,N_16571,N_16210);
nand U17447 (N_17447,N_16081,N_16462);
or U17448 (N_17448,N_16750,N_16469);
and U17449 (N_17449,N_16519,N_16502);
nor U17450 (N_17450,N_16893,N_16014);
or U17451 (N_17451,N_16534,N_16981);
nor U17452 (N_17452,N_16261,N_16695);
nand U17453 (N_17453,N_16976,N_16555);
nand U17454 (N_17454,N_16608,N_16460);
nand U17455 (N_17455,N_16970,N_16919);
xor U17456 (N_17456,N_16190,N_16212);
and U17457 (N_17457,N_16681,N_16104);
nor U17458 (N_17458,N_16132,N_16125);
nor U17459 (N_17459,N_16170,N_16746);
nor U17460 (N_17460,N_16180,N_16256);
and U17461 (N_17461,N_16953,N_16268);
xnor U17462 (N_17462,N_16618,N_16325);
and U17463 (N_17463,N_16040,N_16804);
nor U17464 (N_17464,N_16846,N_16021);
xor U17465 (N_17465,N_16109,N_16990);
nand U17466 (N_17466,N_16918,N_16207);
nor U17467 (N_17467,N_16144,N_16827);
xnor U17468 (N_17468,N_16045,N_16871);
nor U17469 (N_17469,N_16078,N_16053);
nor U17470 (N_17470,N_16177,N_16679);
and U17471 (N_17471,N_16142,N_16620);
nor U17472 (N_17472,N_16248,N_16287);
and U17473 (N_17473,N_16955,N_16733);
nor U17474 (N_17474,N_16701,N_16320);
xor U17475 (N_17475,N_16915,N_16274);
xor U17476 (N_17476,N_16542,N_16589);
nand U17477 (N_17477,N_16703,N_16719);
xor U17478 (N_17478,N_16247,N_16991);
xnor U17479 (N_17479,N_16326,N_16540);
or U17480 (N_17480,N_16852,N_16275);
nor U17481 (N_17481,N_16841,N_16482);
and U17482 (N_17482,N_16501,N_16454);
nor U17483 (N_17483,N_16994,N_16549);
nand U17484 (N_17484,N_16046,N_16110);
nor U17485 (N_17485,N_16817,N_16806);
and U17486 (N_17486,N_16606,N_16375);
or U17487 (N_17487,N_16831,N_16151);
and U17488 (N_17488,N_16023,N_16355);
nand U17489 (N_17489,N_16026,N_16834);
or U17490 (N_17490,N_16035,N_16432);
nor U17491 (N_17491,N_16266,N_16862);
nor U17492 (N_17492,N_16911,N_16129);
xnor U17493 (N_17493,N_16277,N_16380);
or U17494 (N_17494,N_16456,N_16067);
and U17495 (N_17495,N_16688,N_16782);
nor U17496 (N_17496,N_16333,N_16339);
nor U17497 (N_17497,N_16640,N_16622);
nand U17498 (N_17498,N_16183,N_16808);
or U17499 (N_17499,N_16840,N_16005);
xor U17500 (N_17500,N_16771,N_16307);
xor U17501 (N_17501,N_16635,N_16935);
nor U17502 (N_17502,N_16948,N_16243);
and U17503 (N_17503,N_16738,N_16625);
and U17504 (N_17504,N_16896,N_16849);
xnor U17505 (N_17505,N_16546,N_16528);
xor U17506 (N_17506,N_16588,N_16578);
or U17507 (N_17507,N_16371,N_16698);
nand U17508 (N_17508,N_16934,N_16684);
nor U17509 (N_17509,N_16270,N_16523);
or U17510 (N_17510,N_16879,N_16994);
nor U17511 (N_17511,N_16773,N_16832);
nand U17512 (N_17512,N_16557,N_16649);
xnor U17513 (N_17513,N_16598,N_16046);
and U17514 (N_17514,N_16490,N_16708);
nor U17515 (N_17515,N_16679,N_16726);
nand U17516 (N_17516,N_16972,N_16464);
and U17517 (N_17517,N_16351,N_16767);
nand U17518 (N_17518,N_16263,N_16375);
nand U17519 (N_17519,N_16032,N_16092);
or U17520 (N_17520,N_16317,N_16951);
xnor U17521 (N_17521,N_16322,N_16371);
and U17522 (N_17522,N_16107,N_16631);
nand U17523 (N_17523,N_16965,N_16072);
xor U17524 (N_17524,N_16485,N_16597);
xnor U17525 (N_17525,N_16733,N_16844);
and U17526 (N_17526,N_16825,N_16812);
nor U17527 (N_17527,N_16185,N_16459);
and U17528 (N_17528,N_16496,N_16878);
nor U17529 (N_17529,N_16125,N_16598);
nor U17530 (N_17530,N_16780,N_16886);
xnor U17531 (N_17531,N_16411,N_16214);
nor U17532 (N_17532,N_16330,N_16843);
xor U17533 (N_17533,N_16771,N_16940);
nor U17534 (N_17534,N_16775,N_16865);
nand U17535 (N_17535,N_16874,N_16500);
nand U17536 (N_17536,N_16835,N_16706);
nor U17537 (N_17537,N_16073,N_16695);
xnor U17538 (N_17538,N_16161,N_16176);
or U17539 (N_17539,N_16448,N_16413);
xnor U17540 (N_17540,N_16962,N_16072);
nand U17541 (N_17541,N_16179,N_16435);
xnor U17542 (N_17542,N_16292,N_16411);
nor U17543 (N_17543,N_16482,N_16925);
or U17544 (N_17544,N_16143,N_16187);
nor U17545 (N_17545,N_16452,N_16528);
xor U17546 (N_17546,N_16679,N_16587);
or U17547 (N_17547,N_16992,N_16948);
xnor U17548 (N_17548,N_16456,N_16705);
or U17549 (N_17549,N_16375,N_16529);
or U17550 (N_17550,N_16870,N_16823);
xnor U17551 (N_17551,N_16950,N_16930);
nand U17552 (N_17552,N_16674,N_16640);
xor U17553 (N_17553,N_16222,N_16788);
and U17554 (N_17554,N_16237,N_16105);
or U17555 (N_17555,N_16204,N_16516);
xor U17556 (N_17556,N_16278,N_16411);
or U17557 (N_17557,N_16683,N_16365);
nor U17558 (N_17558,N_16652,N_16960);
xor U17559 (N_17559,N_16892,N_16524);
nand U17560 (N_17560,N_16251,N_16857);
or U17561 (N_17561,N_16480,N_16349);
nand U17562 (N_17562,N_16690,N_16591);
nor U17563 (N_17563,N_16545,N_16700);
xor U17564 (N_17564,N_16394,N_16573);
and U17565 (N_17565,N_16072,N_16733);
and U17566 (N_17566,N_16919,N_16841);
or U17567 (N_17567,N_16546,N_16266);
xor U17568 (N_17568,N_16267,N_16611);
and U17569 (N_17569,N_16464,N_16099);
nand U17570 (N_17570,N_16724,N_16884);
or U17571 (N_17571,N_16842,N_16965);
and U17572 (N_17572,N_16195,N_16002);
nand U17573 (N_17573,N_16554,N_16966);
nor U17574 (N_17574,N_16533,N_16314);
xnor U17575 (N_17575,N_16440,N_16929);
nand U17576 (N_17576,N_16907,N_16645);
or U17577 (N_17577,N_16241,N_16972);
nor U17578 (N_17578,N_16181,N_16439);
nor U17579 (N_17579,N_16523,N_16274);
xnor U17580 (N_17580,N_16471,N_16071);
and U17581 (N_17581,N_16878,N_16669);
and U17582 (N_17582,N_16919,N_16385);
xnor U17583 (N_17583,N_16022,N_16665);
and U17584 (N_17584,N_16123,N_16155);
or U17585 (N_17585,N_16349,N_16251);
and U17586 (N_17586,N_16707,N_16048);
nor U17587 (N_17587,N_16059,N_16366);
and U17588 (N_17588,N_16579,N_16699);
xnor U17589 (N_17589,N_16333,N_16862);
or U17590 (N_17590,N_16055,N_16668);
xor U17591 (N_17591,N_16890,N_16748);
nand U17592 (N_17592,N_16667,N_16799);
nand U17593 (N_17593,N_16021,N_16558);
and U17594 (N_17594,N_16559,N_16453);
or U17595 (N_17595,N_16056,N_16375);
or U17596 (N_17596,N_16650,N_16486);
or U17597 (N_17597,N_16090,N_16760);
xnor U17598 (N_17598,N_16950,N_16200);
nand U17599 (N_17599,N_16495,N_16382);
nor U17600 (N_17600,N_16345,N_16355);
nand U17601 (N_17601,N_16314,N_16690);
nor U17602 (N_17602,N_16936,N_16432);
nand U17603 (N_17603,N_16465,N_16494);
xor U17604 (N_17604,N_16640,N_16114);
or U17605 (N_17605,N_16439,N_16830);
or U17606 (N_17606,N_16208,N_16491);
or U17607 (N_17607,N_16455,N_16767);
and U17608 (N_17608,N_16300,N_16848);
nor U17609 (N_17609,N_16355,N_16533);
or U17610 (N_17610,N_16700,N_16346);
nand U17611 (N_17611,N_16556,N_16202);
and U17612 (N_17612,N_16706,N_16618);
nor U17613 (N_17613,N_16042,N_16453);
xnor U17614 (N_17614,N_16712,N_16222);
xnor U17615 (N_17615,N_16602,N_16651);
nor U17616 (N_17616,N_16226,N_16576);
nand U17617 (N_17617,N_16863,N_16913);
nor U17618 (N_17618,N_16393,N_16893);
or U17619 (N_17619,N_16739,N_16340);
or U17620 (N_17620,N_16946,N_16025);
nor U17621 (N_17621,N_16853,N_16269);
nor U17622 (N_17622,N_16856,N_16063);
and U17623 (N_17623,N_16652,N_16301);
nand U17624 (N_17624,N_16667,N_16777);
or U17625 (N_17625,N_16158,N_16049);
or U17626 (N_17626,N_16726,N_16731);
or U17627 (N_17627,N_16963,N_16304);
or U17628 (N_17628,N_16981,N_16265);
xnor U17629 (N_17629,N_16239,N_16271);
or U17630 (N_17630,N_16662,N_16839);
and U17631 (N_17631,N_16532,N_16473);
nor U17632 (N_17632,N_16715,N_16534);
and U17633 (N_17633,N_16509,N_16770);
and U17634 (N_17634,N_16091,N_16624);
nor U17635 (N_17635,N_16185,N_16940);
nor U17636 (N_17636,N_16339,N_16382);
nor U17637 (N_17637,N_16252,N_16609);
nand U17638 (N_17638,N_16941,N_16857);
nor U17639 (N_17639,N_16416,N_16229);
nor U17640 (N_17640,N_16590,N_16735);
and U17641 (N_17641,N_16769,N_16754);
nor U17642 (N_17642,N_16805,N_16533);
nor U17643 (N_17643,N_16467,N_16729);
and U17644 (N_17644,N_16699,N_16130);
xor U17645 (N_17645,N_16778,N_16362);
or U17646 (N_17646,N_16495,N_16717);
nor U17647 (N_17647,N_16208,N_16395);
nor U17648 (N_17648,N_16041,N_16019);
nor U17649 (N_17649,N_16004,N_16983);
and U17650 (N_17650,N_16336,N_16475);
xor U17651 (N_17651,N_16142,N_16732);
nor U17652 (N_17652,N_16602,N_16245);
nand U17653 (N_17653,N_16857,N_16339);
nor U17654 (N_17654,N_16550,N_16586);
and U17655 (N_17655,N_16519,N_16744);
nor U17656 (N_17656,N_16272,N_16647);
and U17657 (N_17657,N_16927,N_16173);
nand U17658 (N_17658,N_16417,N_16480);
and U17659 (N_17659,N_16498,N_16195);
nand U17660 (N_17660,N_16616,N_16307);
nor U17661 (N_17661,N_16652,N_16322);
or U17662 (N_17662,N_16359,N_16297);
or U17663 (N_17663,N_16033,N_16597);
and U17664 (N_17664,N_16932,N_16623);
and U17665 (N_17665,N_16227,N_16380);
or U17666 (N_17666,N_16102,N_16621);
and U17667 (N_17667,N_16452,N_16973);
and U17668 (N_17668,N_16815,N_16916);
xnor U17669 (N_17669,N_16028,N_16923);
and U17670 (N_17670,N_16146,N_16718);
xor U17671 (N_17671,N_16559,N_16909);
and U17672 (N_17672,N_16789,N_16783);
nand U17673 (N_17673,N_16535,N_16137);
and U17674 (N_17674,N_16465,N_16353);
xnor U17675 (N_17675,N_16899,N_16805);
and U17676 (N_17676,N_16347,N_16519);
nor U17677 (N_17677,N_16850,N_16970);
xnor U17678 (N_17678,N_16602,N_16083);
and U17679 (N_17679,N_16964,N_16883);
or U17680 (N_17680,N_16129,N_16938);
and U17681 (N_17681,N_16265,N_16751);
and U17682 (N_17682,N_16217,N_16570);
nor U17683 (N_17683,N_16516,N_16825);
nor U17684 (N_17684,N_16423,N_16185);
xor U17685 (N_17685,N_16590,N_16909);
xnor U17686 (N_17686,N_16849,N_16259);
nand U17687 (N_17687,N_16714,N_16482);
xor U17688 (N_17688,N_16040,N_16588);
nand U17689 (N_17689,N_16020,N_16492);
or U17690 (N_17690,N_16618,N_16184);
xnor U17691 (N_17691,N_16240,N_16922);
nand U17692 (N_17692,N_16251,N_16076);
and U17693 (N_17693,N_16328,N_16366);
and U17694 (N_17694,N_16065,N_16699);
nor U17695 (N_17695,N_16983,N_16337);
nand U17696 (N_17696,N_16616,N_16346);
nor U17697 (N_17697,N_16750,N_16652);
and U17698 (N_17698,N_16482,N_16229);
xor U17699 (N_17699,N_16891,N_16281);
or U17700 (N_17700,N_16700,N_16031);
nor U17701 (N_17701,N_16141,N_16381);
nor U17702 (N_17702,N_16518,N_16332);
xnor U17703 (N_17703,N_16055,N_16793);
and U17704 (N_17704,N_16940,N_16595);
xor U17705 (N_17705,N_16856,N_16718);
and U17706 (N_17706,N_16349,N_16156);
or U17707 (N_17707,N_16295,N_16685);
or U17708 (N_17708,N_16920,N_16822);
nor U17709 (N_17709,N_16796,N_16857);
or U17710 (N_17710,N_16087,N_16190);
and U17711 (N_17711,N_16215,N_16212);
and U17712 (N_17712,N_16847,N_16201);
nand U17713 (N_17713,N_16627,N_16706);
xnor U17714 (N_17714,N_16075,N_16004);
nor U17715 (N_17715,N_16578,N_16456);
or U17716 (N_17716,N_16215,N_16592);
nand U17717 (N_17717,N_16681,N_16238);
and U17718 (N_17718,N_16499,N_16129);
nor U17719 (N_17719,N_16900,N_16161);
or U17720 (N_17720,N_16383,N_16923);
nand U17721 (N_17721,N_16091,N_16228);
nor U17722 (N_17722,N_16431,N_16039);
xor U17723 (N_17723,N_16418,N_16462);
and U17724 (N_17724,N_16547,N_16122);
and U17725 (N_17725,N_16862,N_16740);
nor U17726 (N_17726,N_16967,N_16273);
and U17727 (N_17727,N_16884,N_16827);
nor U17728 (N_17728,N_16974,N_16588);
nand U17729 (N_17729,N_16625,N_16641);
xnor U17730 (N_17730,N_16655,N_16201);
xnor U17731 (N_17731,N_16139,N_16043);
nor U17732 (N_17732,N_16406,N_16724);
and U17733 (N_17733,N_16115,N_16633);
and U17734 (N_17734,N_16428,N_16669);
nand U17735 (N_17735,N_16168,N_16590);
xnor U17736 (N_17736,N_16362,N_16922);
nand U17737 (N_17737,N_16070,N_16984);
nand U17738 (N_17738,N_16681,N_16826);
nor U17739 (N_17739,N_16435,N_16228);
xnor U17740 (N_17740,N_16036,N_16012);
nand U17741 (N_17741,N_16261,N_16451);
nor U17742 (N_17742,N_16963,N_16401);
and U17743 (N_17743,N_16438,N_16632);
or U17744 (N_17744,N_16763,N_16118);
nand U17745 (N_17745,N_16476,N_16067);
or U17746 (N_17746,N_16793,N_16727);
nor U17747 (N_17747,N_16750,N_16613);
nand U17748 (N_17748,N_16244,N_16140);
xnor U17749 (N_17749,N_16792,N_16623);
or U17750 (N_17750,N_16366,N_16783);
nand U17751 (N_17751,N_16988,N_16700);
nand U17752 (N_17752,N_16617,N_16598);
xor U17753 (N_17753,N_16652,N_16317);
and U17754 (N_17754,N_16841,N_16510);
and U17755 (N_17755,N_16534,N_16348);
nand U17756 (N_17756,N_16880,N_16063);
or U17757 (N_17757,N_16219,N_16567);
and U17758 (N_17758,N_16153,N_16597);
nor U17759 (N_17759,N_16363,N_16052);
xnor U17760 (N_17760,N_16957,N_16863);
nor U17761 (N_17761,N_16097,N_16990);
or U17762 (N_17762,N_16897,N_16039);
xnor U17763 (N_17763,N_16009,N_16203);
nand U17764 (N_17764,N_16310,N_16611);
or U17765 (N_17765,N_16302,N_16890);
nor U17766 (N_17766,N_16011,N_16863);
xor U17767 (N_17767,N_16252,N_16441);
xnor U17768 (N_17768,N_16814,N_16242);
or U17769 (N_17769,N_16821,N_16241);
and U17770 (N_17770,N_16381,N_16774);
nand U17771 (N_17771,N_16952,N_16071);
nor U17772 (N_17772,N_16584,N_16043);
xor U17773 (N_17773,N_16852,N_16863);
xnor U17774 (N_17774,N_16010,N_16953);
and U17775 (N_17775,N_16041,N_16118);
or U17776 (N_17776,N_16817,N_16122);
and U17777 (N_17777,N_16437,N_16519);
and U17778 (N_17778,N_16101,N_16165);
or U17779 (N_17779,N_16263,N_16311);
and U17780 (N_17780,N_16831,N_16406);
and U17781 (N_17781,N_16602,N_16956);
nand U17782 (N_17782,N_16643,N_16527);
or U17783 (N_17783,N_16308,N_16755);
or U17784 (N_17784,N_16724,N_16843);
nand U17785 (N_17785,N_16312,N_16267);
nor U17786 (N_17786,N_16948,N_16648);
nor U17787 (N_17787,N_16866,N_16237);
xnor U17788 (N_17788,N_16880,N_16188);
or U17789 (N_17789,N_16271,N_16948);
or U17790 (N_17790,N_16025,N_16831);
nor U17791 (N_17791,N_16473,N_16207);
xnor U17792 (N_17792,N_16825,N_16461);
xor U17793 (N_17793,N_16308,N_16089);
or U17794 (N_17794,N_16037,N_16227);
or U17795 (N_17795,N_16962,N_16223);
or U17796 (N_17796,N_16708,N_16031);
or U17797 (N_17797,N_16022,N_16640);
and U17798 (N_17798,N_16911,N_16431);
and U17799 (N_17799,N_16107,N_16121);
nor U17800 (N_17800,N_16960,N_16054);
and U17801 (N_17801,N_16530,N_16020);
or U17802 (N_17802,N_16715,N_16495);
and U17803 (N_17803,N_16006,N_16231);
nand U17804 (N_17804,N_16222,N_16143);
nor U17805 (N_17805,N_16156,N_16259);
xnor U17806 (N_17806,N_16828,N_16878);
nand U17807 (N_17807,N_16880,N_16353);
nor U17808 (N_17808,N_16337,N_16948);
xor U17809 (N_17809,N_16552,N_16086);
nor U17810 (N_17810,N_16503,N_16359);
and U17811 (N_17811,N_16598,N_16829);
xnor U17812 (N_17812,N_16625,N_16285);
nor U17813 (N_17813,N_16772,N_16923);
xor U17814 (N_17814,N_16088,N_16749);
nand U17815 (N_17815,N_16273,N_16316);
or U17816 (N_17816,N_16805,N_16908);
and U17817 (N_17817,N_16373,N_16281);
nor U17818 (N_17818,N_16230,N_16035);
xor U17819 (N_17819,N_16339,N_16238);
nor U17820 (N_17820,N_16341,N_16516);
and U17821 (N_17821,N_16804,N_16897);
and U17822 (N_17822,N_16878,N_16987);
or U17823 (N_17823,N_16664,N_16721);
and U17824 (N_17824,N_16778,N_16881);
xor U17825 (N_17825,N_16996,N_16556);
and U17826 (N_17826,N_16256,N_16037);
xnor U17827 (N_17827,N_16808,N_16856);
or U17828 (N_17828,N_16276,N_16716);
and U17829 (N_17829,N_16190,N_16959);
xor U17830 (N_17830,N_16151,N_16179);
nand U17831 (N_17831,N_16241,N_16355);
or U17832 (N_17832,N_16014,N_16198);
or U17833 (N_17833,N_16467,N_16954);
nor U17834 (N_17834,N_16409,N_16509);
nor U17835 (N_17835,N_16006,N_16617);
and U17836 (N_17836,N_16518,N_16373);
or U17837 (N_17837,N_16363,N_16002);
nand U17838 (N_17838,N_16568,N_16244);
and U17839 (N_17839,N_16763,N_16784);
and U17840 (N_17840,N_16056,N_16432);
xor U17841 (N_17841,N_16259,N_16597);
xnor U17842 (N_17842,N_16667,N_16208);
nand U17843 (N_17843,N_16908,N_16253);
nand U17844 (N_17844,N_16021,N_16811);
nor U17845 (N_17845,N_16537,N_16816);
or U17846 (N_17846,N_16528,N_16470);
nand U17847 (N_17847,N_16950,N_16673);
or U17848 (N_17848,N_16887,N_16006);
nor U17849 (N_17849,N_16372,N_16994);
and U17850 (N_17850,N_16051,N_16824);
nand U17851 (N_17851,N_16476,N_16790);
xnor U17852 (N_17852,N_16106,N_16533);
nand U17853 (N_17853,N_16417,N_16644);
and U17854 (N_17854,N_16788,N_16533);
or U17855 (N_17855,N_16997,N_16833);
or U17856 (N_17856,N_16508,N_16732);
or U17857 (N_17857,N_16633,N_16040);
nand U17858 (N_17858,N_16382,N_16181);
and U17859 (N_17859,N_16911,N_16074);
and U17860 (N_17860,N_16489,N_16344);
and U17861 (N_17861,N_16585,N_16122);
nor U17862 (N_17862,N_16964,N_16054);
nand U17863 (N_17863,N_16144,N_16012);
nor U17864 (N_17864,N_16846,N_16329);
and U17865 (N_17865,N_16081,N_16190);
or U17866 (N_17866,N_16230,N_16796);
or U17867 (N_17867,N_16153,N_16076);
xor U17868 (N_17868,N_16889,N_16264);
xor U17869 (N_17869,N_16448,N_16159);
or U17870 (N_17870,N_16706,N_16837);
or U17871 (N_17871,N_16054,N_16372);
and U17872 (N_17872,N_16232,N_16602);
or U17873 (N_17873,N_16861,N_16435);
nor U17874 (N_17874,N_16664,N_16418);
nand U17875 (N_17875,N_16266,N_16444);
nor U17876 (N_17876,N_16711,N_16117);
nor U17877 (N_17877,N_16030,N_16890);
or U17878 (N_17878,N_16564,N_16150);
xor U17879 (N_17879,N_16734,N_16279);
and U17880 (N_17880,N_16668,N_16566);
nor U17881 (N_17881,N_16837,N_16875);
nand U17882 (N_17882,N_16830,N_16869);
nor U17883 (N_17883,N_16736,N_16557);
xor U17884 (N_17884,N_16469,N_16684);
or U17885 (N_17885,N_16520,N_16471);
nand U17886 (N_17886,N_16122,N_16452);
nor U17887 (N_17887,N_16569,N_16960);
or U17888 (N_17888,N_16127,N_16190);
and U17889 (N_17889,N_16307,N_16413);
and U17890 (N_17890,N_16424,N_16957);
xor U17891 (N_17891,N_16611,N_16959);
nor U17892 (N_17892,N_16508,N_16627);
xnor U17893 (N_17893,N_16164,N_16076);
nand U17894 (N_17894,N_16811,N_16863);
and U17895 (N_17895,N_16033,N_16703);
nand U17896 (N_17896,N_16840,N_16279);
or U17897 (N_17897,N_16140,N_16751);
nand U17898 (N_17898,N_16209,N_16305);
xor U17899 (N_17899,N_16096,N_16668);
nor U17900 (N_17900,N_16440,N_16672);
and U17901 (N_17901,N_16407,N_16131);
nand U17902 (N_17902,N_16143,N_16410);
and U17903 (N_17903,N_16548,N_16374);
xor U17904 (N_17904,N_16120,N_16566);
nor U17905 (N_17905,N_16264,N_16978);
nor U17906 (N_17906,N_16066,N_16748);
or U17907 (N_17907,N_16271,N_16154);
nand U17908 (N_17908,N_16429,N_16096);
and U17909 (N_17909,N_16280,N_16578);
and U17910 (N_17910,N_16489,N_16368);
or U17911 (N_17911,N_16616,N_16657);
xor U17912 (N_17912,N_16029,N_16524);
nor U17913 (N_17913,N_16284,N_16166);
and U17914 (N_17914,N_16913,N_16803);
nor U17915 (N_17915,N_16217,N_16731);
nand U17916 (N_17916,N_16841,N_16668);
xnor U17917 (N_17917,N_16700,N_16278);
xnor U17918 (N_17918,N_16380,N_16137);
or U17919 (N_17919,N_16708,N_16378);
nor U17920 (N_17920,N_16557,N_16073);
nor U17921 (N_17921,N_16346,N_16403);
nand U17922 (N_17922,N_16537,N_16083);
or U17923 (N_17923,N_16500,N_16134);
or U17924 (N_17924,N_16726,N_16116);
nor U17925 (N_17925,N_16955,N_16413);
nor U17926 (N_17926,N_16191,N_16876);
or U17927 (N_17927,N_16260,N_16227);
or U17928 (N_17928,N_16751,N_16958);
and U17929 (N_17929,N_16587,N_16020);
xor U17930 (N_17930,N_16560,N_16340);
xor U17931 (N_17931,N_16581,N_16864);
nor U17932 (N_17932,N_16947,N_16712);
nor U17933 (N_17933,N_16919,N_16326);
nor U17934 (N_17934,N_16458,N_16843);
nand U17935 (N_17935,N_16441,N_16105);
nand U17936 (N_17936,N_16574,N_16016);
nand U17937 (N_17937,N_16563,N_16810);
or U17938 (N_17938,N_16208,N_16766);
nand U17939 (N_17939,N_16868,N_16156);
nand U17940 (N_17940,N_16894,N_16353);
and U17941 (N_17941,N_16116,N_16066);
nand U17942 (N_17942,N_16063,N_16232);
or U17943 (N_17943,N_16728,N_16891);
nand U17944 (N_17944,N_16708,N_16278);
nand U17945 (N_17945,N_16746,N_16169);
and U17946 (N_17946,N_16213,N_16464);
nor U17947 (N_17947,N_16961,N_16588);
nor U17948 (N_17948,N_16506,N_16989);
nand U17949 (N_17949,N_16957,N_16220);
or U17950 (N_17950,N_16340,N_16700);
nand U17951 (N_17951,N_16164,N_16502);
or U17952 (N_17952,N_16170,N_16980);
or U17953 (N_17953,N_16218,N_16671);
nand U17954 (N_17954,N_16120,N_16431);
and U17955 (N_17955,N_16943,N_16272);
or U17956 (N_17956,N_16342,N_16039);
and U17957 (N_17957,N_16112,N_16151);
and U17958 (N_17958,N_16453,N_16654);
or U17959 (N_17959,N_16577,N_16788);
and U17960 (N_17960,N_16111,N_16758);
nor U17961 (N_17961,N_16788,N_16477);
and U17962 (N_17962,N_16219,N_16287);
nor U17963 (N_17963,N_16881,N_16604);
nor U17964 (N_17964,N_16494,N_16424);
nor U17965 (N_17965,N_16057,N_16449);
nand U17966 (N_17966,N_16339,N_16852);
nor U17967 (N_17967,N_16605,N_16858);
or U17968 (N_17968,N_16578,N_16177);
xnor U17969 (N_17969,N_16149,N_16728);
xnor U17970 (N_17970,N_16913,N_16389);
nand U17971 (N_17971,N_16635,N_16916);
xor U17972 (N_17972,N_16593,N_16948);
nor U17973 (N_17973,N_16586,N_16836);
or U17974 (N_17974,N_16040,N_16171);
nor U17975 (N_17975,N_16946,N_16538);
xnor U17976 (N_17976,N_16751,N_16812);
and U17977 (N_17977,N_16413,N_16802);
nor U17978 (N_17978,N_16996,N_16456);
nand U17979 (N_17979,N_16782,N_16062);
or U17980 (N_17980,N_16299,N_16240);
and U17981 (N_17981,N_16937,N_16875);
xor U17982 (N_17982,N_16683,N_16697);
or U17983 (N_17983,N_16474,N_16664);
or U17984 (N_17984,N_16752,N_16274);
or U17985 (N_17985,N_16374,N_16619);
xnor U17986 (N_17986,N_16896,N_16682);
xor U17987 (N_17987,N_16759,N_16288);
xnor U17988 (N_17988,N_16241,N_16036);
nand U17989 (N_17989,N_16422,N_16693);
or U17990 (N_17990,N_16473,N_16162);
nor U17991 (N_17991,N_16446,N_16424);
nand U17992 (N_17992,N_16524,N_16171);
nand U17993 (N_17993,N_16983,N_16671);
and U17994 (N_17994,N_16917,N_16279);
xor U17995 (N_17995,N_16836,N_16519);
or U17996 (N_17996,N_16469,N_16726);
and U17997 (N_17997,N_16194,N_16517);
nand U17998 (N_17998,N_16420,N_16119);
xnor U17999 (N_17999,N_16370,N_16970);
xnor U18000 (N_18000,N_17267,N_17546);
nand U18001 (N_18001,N_17249,N_17523);
and U18002 (N_18002,N_17117,N_17813);
and U18003 (N_18003,N_17162,N_17601);
nand U18004 (N_18004,N_17357,N_17488);
nor U18005 (N_18005,N_17067,N_17078);
nand U18006 (N_18006,N_17230,N_17703);
nor U18007 (N_18007,N_17322,N_17498);
xnor U18008 (N_18008,N_17531,N_17182);
nand U18009 (N_18009,N_17753,N_17847);
nor U18010 (N_18010,N_17671,N_17110);
nand U18011 (N_18011,N_17168,N_17627);
nand U18012 (N_18012,N_17804,N_17572);
xor U18013 (N_18013,N_17347,N_17743);
nor U18014 (N_18014,N_17918,N_17343);
xor U18015 (N_18015,N_17164,N_17401);
or U18016 (N_18016,N_17589,N_17137);
or U18017 (N_18017,N_17537,N_17636);
xor U18018 (N_18018,N_17680,N_17239);
nand U18019 (N_18019,N_17157,N_17900);
and U18020 (N_18020,N_17303,N_17999);
or U18021 (N_18021,N_17118,N_17910);
and U18022 (N_18022,N_17824,N_17694);
xor U18023 (N_18023,N_17613,N_17834);
nor U18024 (N_18024,N_17500,N_17229);
and U18025 (N_18025,N_17646,N_17723);
xnor U18026 (N_18026,N_17425,N_17189);
nand U18027 (N_18027,N_17822,N_17797);
xnor U18028 (N_18028,N_17340,N_17313);
nor U18029 (N_18029,N_17662,N_17849);
and U18030 (N_18030,N_17967,N_17060);
nor U18031 (N_18031,N_17543,N_17045);
xnor U18032 (N_18032,N_17602,N_17669);
xor U18033 (N_18033,N_17148,N_17643);
and U18034 (N_18034,N_17529,N_17936);
and U18035 (N_18035,N_17036,N_17856);
and U18036 (N_18036,N_17028,N_17782);
and U18037 (N_18037,N_17349,N_17776);
nor U18038 (N_18038,N_17520,N_17408);
and U18039 (N_18039,N_17974,N_17098);
and U18040 (N_18040,N_17360,N_17062);
nor U18041 (N_18041,N_17949,N_17605);
and U18042 (N_18042,N_17200,N_17784);
and U18043 (N_18043,N_17468,N_17258);
nand U18044 (N_18044,N_17640,N_17561);
and U18045 (N_18045,N_17113,N_17158);
nand U18046 (N_18046,N_17415,N_17108);
nand U18047 (N_18047,N_17564,N_17751);
or U18048 (N_18048,N_17462,N_17035);
nor U18049 (N_18049,N_17614,N_17735);
xor U18050 (N_18050,N_17376,N_17076);
or U18051 (N_18051,N_17369,N_17480);
nand U18052 (N_18052,N_17173,N_17147);
nand U18053 (N_18053,N_17870,N_17043);
nor U18054 (N_18054,N_17487,N_17263);
or U18055 (N_18055,N_17474,N_17130);
nor U18056 (N_18056,N_17140,N_17455);
and U18057 (N_18057,N_17335,N_17748);
and U18058 (N_18058,N_17009,N_17330);
and U18059 (N_18059,N_17151,N_17407);
or U18060 (N_18060,N_17556,N_17979);
and U18061 (N_18061,N_17737,N_17368);
nor U18062 (N_18062,N_17865,N_17734);
or U18063 (N_18063,N_17334,N_17190);
nand U18064 (N_18064,N_17504,N_17619);
nand U18065 (N_18065,N_17712,N_17270);
nor U18066 (N_18066,N_17121,N_17586);
xor U18067 (N_18067,N_17687,N_17770);
or U18068 (N_18068,N_17551,N_17491);
and U18069 (N_18069,N_17590,N_17582);
nor U18070 (N_18070,N_17005,N_17746);
xnor U18071 (N_18071,N_17309,N_17383);
and U18072 (N_18072,N_17466,N_17559);
nor U18073 (N_18073,N_17167,N_17534);
nand U18074 (N_18074,N_17152,N_17738);
and U18075 (N_18075,N_17153,N_17789);
nor U18076 (N_18076,N_17653,N_17584);
xor U18077 (N_18077,N_17288,N_17896);
or U18078 (N_18078,N_17844,N_17047);
and U18079 (N_18079,N_17616,N_17105);
or U18080 (N_18080,N_17194,N_17717);
xnor U18081 (N_18081,N_17908,N_17509);
nand U18082 (N_18082,N_17704,N_17165);
xor U18083 (N_18083,N_17833,N_17881);
or U18084 (N_18084,N_17545,N_17302);
nor U18085 (N_18085,N_17928,N_17410);
nor U18086 (N_18086,N_17431,N_17926);
and U18087 (N_18087,N_17650,N_17615);
or U18088 (N_18088,N_17413,N_17435);
nor U18089 (N_18089,N_17639,N_17620);
xnor U18090 (N_18090,N_17450,N_17198);
xor U18091 (N_18091,N_17961,N_17317);
nor U18092 (N_18092,N_17075,N_17766);
and U18093 (N_18093,N_17090,N_17433);
and U18094 (N_18094,N_17858,N_17454);
nor U18095 (N_18095,N_17205,N_17094);
xnor U18096 (N_18096,N_17188,N_17467);
and U18097 (N_18097,N_17510,N_17321);
xnor U18098 (N_18098,N_17237,N_17208);
xnor U18099 (N_18099,N_17986,N_17089);
nor U18100 (N_18100,N_17664,N_17852);
and U18101 (N_18101,N_17750,N_17892);
nand U18102 (N_18102,N_17575,N_17247);
xor U18103 (N_18103,N_17866,N_17227);
nor U18104 (N_18104,N_17146,N_17678);
and U18105 (N_18105,N_17314,N_17581);
xnor U18106 (N_18106,N_17412,N_17940);
or U18107 (N_18107,N_17486,N_17539);
or U18108 (N_18108,N_17095,N_17221);
or U18109 (N_18109,N_17711,N_17315);
xnor U18110 (N_18110,N_17283,N_17262);
or U18111 (N_18111,N_17655,N_17884);
xnor U18112 (N_18112,N_17527,N_17732);
or U18113 (N_18113,N_17690,N_17115);
nand U18114 (N_18114,N_17018,N_17481);
xnor U18115 (N_18115,N_17501,N_17722);
xor U18116 (N_18116,N_17661,N_17037);
xor U18117 (N_18117,N_17790,N_17673);
and U18118 (N_18118,N_17981,N_17346);
nor U18119 (N_18119,N_17378,N_17277);
nand U18120 (N_18120,N_17795,N_17055);
nor U18121 (N_18121,N_17811,N_17295);
and U18122 (N_18122,N_17526,N_17938);
nand U18123 (N_18123,N_17914,N_17930);
nand U18124 (N_18124,N_17719,N_17278);
nor U18125 (N_18125,N_17176,N_17959);
and U18126 (N_18126,N_17339,N_17695);
nor U18127 (N_18127,N_17398,N_17550);
nor U18128 (N_18128,N_17853,N_17511);
and U18129 (N_18129,N_17780,N_17571);
nand U18130 (N_18130,N_17003,N_17679);
or U18131 (N_18131,N_17594,N_17882);
nand U18132 (N_18132,N_17876,N_17869);
nand U18133 (N_18133,N_17429,N_17683);
and U18134 (N_18134,N_17902,N_17887);
or U18135 (N_18135,N_17689,N_17864);
or U18136 (N_18136,N_17924,N_17451);
nor U18137 (N_18137,N_17050,N_17178);
xor U18138 (N_18138,N_17666,N_17456);
nor U18139 (N_18139,N_17141,N_17625);
and U18140 (N_18140,N_17651,N_17469);
xor U18141 (N_18141,N_17720,N_17312);
nor U18142 (N_18142,N_17547,N_17079);
xnor U18143 (N_18143,N_17946,N_17769);
nand U18144 (N_18144,N_17327,N_17994);
nor U18145 (N_18145,N_17492,N_17554);
and U18146 (N_18146,N_17187,N_17266);
nor U18147 (N_18147,N_17440,N_17265);
nor U18148 (N_18148,N_17508,N_17161);
and U18149 (N_18149,N_17820,N_17426);
xnor U18150 (N_18150,N_17225,N_17351);
and U18151 (N_18151,N_17296,N_17143);
nor U18152 (N_18152,N_17760,N_17513);
or U18153 (N_18153,N_17496,N_17987);
xor U18154 (N_18154,N_17871,N_17608);
xor U18155 (N_18155,N_17484,N_17406);
nand U18156 (N_18156,N_17246,N_17993);
nor U18157 (N_18157,N_17555,N_17396);
or U18158 (N_18158,N_17169,N_17175);
nor U18159 (N_18159,N_17960,N_17489);
xnor U18160 (N_18160,N_17862,N_17801);
nand U18161 (N_18161,N_17814,N_17920);
xnor U18162 (N_18162,N_17757,N_17805);
nand U18163 (N_18163,N_17775,N_17464);
or U18164 (N_18164,N_17744,N_17494);
nand U18165 (N_18165,N_17260,N_17040);
and U18166 (N_18166,N_17580,N_17294);
nor U18167 (N_18167,N_17767,N_17058);
or U18168 (N_18168,N_17861,N_17837);
nand U18169 (N_18169,N_17326,N_17109);
nor U18170 (N_18170,N_17848,N_17384);
xor U18171 (N_18171,N_17672,N_17973);
or U18172 (N_18172,N_17197,N_17102);
or U18173 (N_18173,N_17595,N_17476);
nor U18174 (N_18174,N_17250,N_17286);
or U18175 (N_18175,N_17016,N_17693);
and U18176 (N_18176,N_17222,N_17097);
nand U18177 (N_18177,N_17761,N_17966);
or U18178 (N_18178,N_17667,N_17032);
xor U18179 (N_18179,N_17710,N_17017);
xnor U18180 (N_18180,N_17691,N_17830);
nand U18181 (N_18181,N_17955,N_17372);
and U18182 (N_18182,N_17170,N_17785);
xnor U18183 (N_18183,N_17898,N_17729);
xnor U18184 (N_18184,N_17195,N_17381);
xnor U18185 (N_18185,N_17086,N_17536);
nor U18186 (N_18186,N_17002,N_17652);
and U18187 (N_18187,N_17251,N_17524);
and U18188 (N_18188,N_17565,N_17942);
nand U18189 (N_18189,N_17127,N_17968);
xnor U18190 (N_18190,N_17587,N_17088);
nor U18191 (N_18191,N_17739,N_17083);
or U18192 (N_18192,N_17518,N_17919);
or U18193 (N_18193,N_17823,N_17688);
xnor U18194 (N_18194,N_17224,N_17399);
nor U18195 (N_18195,N_17240,N_17647);
nand U18196 (N_18196,N_17293,N_17984);
nand U18197 (N_18197,N_17452,N_17160);
nor U18198 (N_18198,N_17423,N_17515);
nand U18199 (N_18199,N_17080,N_17206);
or U18200 (N_18200,N_17634,N_17868);
xor U18201 (N_18201,N_17259,N_17759);
or U18202 (N_18202,N_17180,N_17975);
nand U18203 (N_18203,N_17568,N_17163);
nor U18204 (N_18204,N_17081,N_17891);
nor U18205 (N_18205,N_17773,N_17063);
xnor U18206 (N_18206,N_17375,N_17107);
nand U18207 (N_18207,N_17845,N_17542);
xnor U18208 (N_18208,N_17054,N_17010);
nand U18209 (N_18209,N_17557,N_17535);
nand U18210 (N_18210,N_17799,N_17519);
nand U18211 (N_18211,N_17872,N_17957);
nor U18212 (N_18212,N_17726,N_17389);
or U18213 (N_18213,N_17913,N_17387);
nand U18214 (N_18214,N_17006,N_17216);
nor U18215 (N_18215,N_17740,N_17716);
and U18216 (N_18216,N_17528,N_17779);
and U18217 (N_18217,N_17235,N_17100);
xor U18218 (N_18218,N_17859,N_17364);
xnor U18219 (N_18219,N_17223,N_17829);
nor U18220 (N_18220,N_17457,N_17414);
or U18221 (N_18221,N_17133,N_17320);
and U18222 (N_18222,N_17254,N_17126);
and U18223 (N_18223,N_17391,N_17706);
or U18224 (N_18224,N_17256,N_17226);
nor U18225 (N_18225,N_17019,N_17171);
nor U18226 (N_18226,N_17422,N_17879);
and U18227 (N_18227,N_17308,N_17709);
and U18228 (N_18228,N_17271,N_17405);
or U18229 (N_18229,N_17521,N_17085);
or U18230 (N_18230,N_17569,N_17988);
nand U18231 (N_18231,N_17934,N_17144);
and U18232 (N_18232,N_17380,N_17752);
or U18233 (N_18233,N_17091,N_17566);
nor U18234 (N_18234,N_17485,N_17185);
or U18235 (N_18235,N_17268,N_17635);
or U18236 (N_18236,N_17417,N_17065);
or U18237 (N_18237,N_17660,N_17715);
or U18238 (N_18238,N_17774,N_17418);
nor U18239 (N_18239,N_17214,N_17329);
nand U18240 (N_18240,N_17969,N_17745);
xnor U18241 (N_18241,N_17436,N_17025);
or U18242 (N_18242,N_17393,N_17034);
xor U18243 (N_18243,N_17649,N_17276);
xnor U18244 (N_18244,N_17939,N_17641);
and U18245 (N_18245,N_17525,N_17241);
nor U18246 (N_18246,N_17082,N_17056);
or U18247 (N_18247,N_17576,N_17787);
xnor U18248 (N_18248,N_17819,N_17609);
and U18249 (N_18249,N_17668,N_17765);
and U18250 (N_18250,N_17186,N_17274);
nand U18251 (N_18251,N_17588,N_17430);
xnor U18252 (N_18252,N_17030,N_17356);
nand U18253 (N_18253,N_17307,N_17041);
and U18254 (N_18254,N_17027,N_17842);
or U18255 (N_18255,N_17827,N_17618);
and U18256 (N_18256,N_17976,N_17793);
and U18257 (N_18257,N_17885,N_17832);
or U18258 (N_18258,N_17791,N_17621);
xnor U18259 (N_18259,N_17702,N_17633);
or U18260 (N_18260,N_17337,N_17142);
and U18261 (N_18261,N_17764,N_17867);
nor U18262 (N_18262,N_17438,N_17261);
xor U18263 (N_18263,N_17730,N_17014);
xnor U18264 (N_18264,N_17473,N_17894);
and U18265 (N_18265,N_17623,N_17447);
nor U18266 (N_18266,N_17733,N_17442);
or U18267 (N_18267,N_17597,N_17021);
and U18268 (N_18268,N_17883,N_17166);
nor U18269 (N_18269,N_17465,N_17828);
xnor U18270 (N_18270,N_17434,N_17382);
and U18271 (N_18271,N_17196,N_17232);
and U18272 (N_18272,N_17290,N_17015);
or U18273 (N_18273,N_17593,N_17252);
nor U18274 (N_18274,N_17145,N_17839);
and U18275 (N_18275,N_17659,N_17850);
nor U18276 (N_18276,N_17310,N_17388);
and U18277 (N_18277,N_17400,N_17495);
nand U18278 (N_18278,N_17802,N_17714);
or U18279 (N_18279,N_17600,N_17922);
or U18280 (N_18280,N_17783,N_17724);
nor U18281 (N_18281,N_17111,N_17817);
or U18282 (N_18282,N_17243,N_17656);
nand U18283 (N_18283,N_17132,N_17355);
or U18284 (N_18284,N_17541,N_17207);
xor U18285 (N_18285,N_17156,N_17472);
or U18286 (N_18286,N_17209,N_17777);
and U18287 (N_18287,N_17906,N_17530);
or U18288 (N_18288,N_17681,N_17831);
or U18289 (N_18289,N_17421,N_17004);
nand U18290 (N_18290,N_17101,N_17980);
nand U18291 (N_18291,N_17754,N_17877);
and U18292 (N_18292,N_17461,N_17395);
nand U18293 (N_18293,N_17069,N_17854);
nand U18294 (N_18294,N_17763,N_17299);
and U18295 (N_18295,N_17234,N_17573);
or U18296 (N_18296,N_17319,N_17971);
nor U18297 (N_18297,N_17120,N_17925);
xnor U18298 (N_18298,N_17591,N_17128);
or U18299 (N_18299,N_17963,N_17297);
nor U18300 (N_18300,N_17670,N_17758);
nand U18301 (N_18301,N_17540,N_17624);
nor U18302 (N_18302,N_17708,N_17912);
and U18303 (N_18303,N_17637,N_17345);
xor U18304 (N_18304,N_17444,N_17825);
xor U18305 (N_18305,N_17701,N_17038);
and U18306 (N_18306,N_17077,N_17272);
or U18307 (N_18307,N_17826,N_17617);
xnor U18308 (N_18308,N_17684,N_17013);
nor U18309 (N_18309,N_17370,N_17786);
and U18310 (N_18310,N_17544,N_17449);
nand U18311 (N_18311,N_17731,N_17304);
xnor U18312 (N_18312,N_17439,N_17948);
xor U18313 (N_18313,N_17696,N_17228);
and U18314 (N_18314,N_17736,N_17218);
xor U18315 (N_18315,N_17927,N_17857);
nand U18316 (N_18316,N_17747,N_17236);
xor U18317 (N_18317,N_17563,N_17478);
nor U18318 (N_18318,N_17211,N_17217);
nand U18319 (N_18319,N_17503,N_17007);
nand U18320 (N_18320,N_17585,N_17497);
and U18321 (N_18321,N_17992,N_17771);
nor U18322 (N_18322,N_17233,N_17812);
nand U18323 (N_18323,N_17843,N_17245);
xnor U18324 (N_18324,N_17134,N_17301);
or U18325 (N_18325,N_17199,N_17291);
or U18326 (N_18326,N_17257,N_17470);
or U18327 (N_18327,N_17685,N_17119);
nand U18328 (N_18328,N_17443,N_17741);
xnor U18329 (N_18329,N_17756,N_17306);
and U18330 (N_18330,N_17603,N_17982);
nand U18331 (N_18331,N_17096,N_17213);
or U18332 (N_18332,N_17950,N_17810);
nor U18333 (N_18333,N_17516,N_17445);
nand U18334 (N_18334,N_17428,N_17798);
and U18335 (N_18335,N_17366,N_17264);
or U18336 (N_18336,N_17064,N_17713);
nor U18337 (N_18337,N_17816,N_17371);
nand U18338 (N_18338,N_17570,N_17807);
and U18339 (N_18339,N_17012,N_17344);
nand U18340 (N_18340,N_17042,N_17172);
or U18341 (N_18341,N_17772,N_17598);
and U18342 (N_18342,N_17579,N_17219);
nand U18343 (N_18343,N_17386,N_17895);
or U18344 (N_18344,N_17354,N_17522);
or U18345 (N_18345,N_17796,N_17644);
xnor U18346 (N_18346,N_17983,N_17359);
xnor U18347 (N_18347,N_17289,N_17944);
nor U18348 (N_18348,N_17749,N_17998);
xnor U18349 (N_18349,N_17562,N_17338);
or U18350 (N_18350,N_17970,N_17803);
xnor U18351 (N_18351,N_17350,N_17174);
or U18352 (N_18352,N_17626,N_17933);
xor U18353 (N_18353,N_17697,N_17284);
xnor U18354 (N_18354,N_17073,N_17092);
xnor U18355 (N_18355,N_17978,N_17332);
or U18356 (N_18356,N_17532,N_17604);
nand U18357 (N_18357,N_17553,N_17855);
or U18358 (N_18358,N_17475,N_17253);
nand U18359 (N_18359,N_17840,N_17479);
nor U18360 (N_18360,N_17996,N_17700);
xnor U18361 (N_18361,N_17070,N_17682);
xor U18362 (N_18362,N_17916,N_17483);
nor U18363 (N_18363,N_17788,N_17139);
nand U18364 (N_18364,N_17074,N_17596);
nand U18365 (N_18365,N_17642,N_17202);
xnor U18366 (N_18366,N_17538,N_17285);
and U18367 (N_18367,N_17499,N_17808);
or U18368 (N_18368,N_17020,N_17698);
and U18369 (N_18369,N_17610,N_17448);
nand U18370 (N_18370,N_17907,N_17792);
or U18371 (N_18371,N_17287,N_17203);
nand U18372 (N_18372,N_17273,N_17402);
nor U18373 (N_18373,N_17215,N_17676);
xnor U18374 (N_18374,N_17155,N_17397);
xor U18375 (N_18375,N_17567,N_17985);
or U18376 (N_18376,N_17149,N_17705);
and U18377 (N_18377,N_17026,N_17201);
xor U18378 (N_18378,N_17929,N_17836);
xnor U18379 (N_18379,N_17099,N_17958);
or U18380 (N_18380,N_17622,N_17901);
or U18381 (N_18381,N_17358,N_17577);
or U18382 (N_18382,N_17956,N_17353);
nand U18383 (N_18383,N_17193,N_17923);
and U18384 (N_18384,N_17333,N_17116);
or U18385 (N_18385,N_17658,N_17059);
or U18386 (N_18386,N_17718,N_17599);
nand U18387 (N_18387,N_17248,N_17851);
or U18388 (N_18388,N_17821,N_17493);
or U18389 (N_18389,N_17392,N_17977);
nand U18390 (N_18390,N_17046,N_17437);
or U18391 (N_18391,N_17815,N_17061);
nor U18392 (N_18392,N_17052,N_17305);
or U18393 (N_18393,N_17583,N_17951);
or U18394 (N_18394,N_17742,N_17361);
nand U18395 (N_18395,N_17725,N_17889);
and U18396 (N_18396,N_17441,N_17794);
nor U18397 (N_18397,N_17051,N_17336);
nor U18398 (N_18398,N_17915,N_17558);
and U18399 (N_18399,N_17179,N_17403);
nor U18400 (N_18400,N_17692,N_17125);
xor U18401 (N_18401,N_17048,N_17878);
or U18402 (N_18402,N_17331,N_17404);
nor U18403 (N_18403,N_17686,N_17023);
nand U18404 (N_18404,N_17282,N_17707);
nand U18405 (N_18405,N_17220,N_17606);
nand U18406 (N_18406,N_17904,N_17275);
and U18407 (N_18407,N_17755,N_17818);
and U18408 (N_18408,N_17533,N_17031);
and U18409 (N_18409,N_17458,N_17029);
xnor U18410 (N_18410,N_17394,N_17093);
or U18411 (N_18411,N_17778,N_17954);
and U18412 (N_18412,N_17654,N_17781);
xor U18413 (N_18413,N_17578,N_17962);
nand U18414 (N_18414,N_17379,N_17548);
xor U18415 (N_18415,N_17880,N_17630);
nor U18416 (N_18416,N_17039,N_17298);
and U18417 (N_18417,N_17318,N_17066);
nor U18418 (N_18418,N_17104,N_17665);
nand U18419 (N_18419,N_17935,N_17033);
nand U18420 (N_18420,N_17941,N_17446);
and U18421 (N_18421,N_17057,N_17860);
and U18422 (N_18422,N_17212,N_17242);
and U18423 (N_18423,N_17341,N_17044);
xor U18424 (N_18424,N_17184,N_17838);
nor U18425 (N_18425,N_17420,N_17611);
and U18426 (N_18426,N_17863,N_17835);
xnor U18427 (N_18427,N_17874,N_17875);
or U18428 (N_18428,N_17997,N_17903);
nand U18429 (N_18429,N_17727,N_17995);
or U18430 (N_18430,N_17324,N_17323);
xnor U18431 (N_18431,N_17238,N_17460);
or U18432 (N_18432,N_17964,N_17138);
nand U18433 (N_18433,N_17490,N_17352);
nand U18434 (N_18434,N_17129,N_17106);
xor U18435 (N_18435,N_17846,N_17365);
xor U18436 (N_18436,N_17677,N_17008);
xor U18437 (N_18437,N_17560,N_17416);
and U18438 (N_18438,N_17432,N_17292);
or U18439 (N_18439,N_17932,N_17279);
and U18440 (N_18440,N_17592,N_17183);
and U18441 (N_18441,N_17103,N_17965);
nand U18442 (N_18442,N_17873,N_17150);
nand U18443 (N_18443,N_17663,N_17897);
xor U18444 (N_18444,N_17482,N_17419);
nand U18445 (N_18445,N_17943,N_17362);
nor U18446 (N_18446,N_17068,N_17629);
nor U18447 (N_18447,N_17348,N_17886);
or U18448 (N_18448,N_17311,N_17280);
nor U18449 (N_18449,N_17638,N_17953);
nor U18450 (N_18450,N_17053,N_17325);
or U18451 (N_18451,N_17363,N_17989);
and U18452 (N_18452,N_17390,N_17244);
nand U18453 (N_18453,N_17024,N_17385);
xnor U18454 (N_18454,N_17409,N_17945);
and U18455 (N_18455,N_17124,N_17506);
xnor U18456 (N_18456,N_17952,N_17931);
or U18457 (N_18457,N_17000,N_17181);
and U18458 (N_18458,N_17947,N_17502);
nor U18459 (N_18459,N_17154,N_17512);
nand U18460 (N_18460,N_17367,N_17657);
and U18461 (N_18461,N_17762,N_17888);
and U18462 (N_18462,N_17768,N_17072);
and U18463 (N_18463,N_17574,N_17177);
nor U18464 (N_18464,N_17123,N_17800);
nor U18465 (N_18465,N_17841,N_17374);
xor U18466 (N_18466,N_17552,N_17377);
or U18467 (N_18467,N_17809,N_17159);
or U18468 (N_18468,N_17991,N_17049);
xnor U18469 (N_18469,N_17972,N_17463);
or U18470 (N_18470,N_17607,N_17674);
xnor U18471 (N_18471,N_17427,N_17549);
and U18472 (N_18472,N_17675,N_17122);
nand U18473 (N_18473,N_17632,N_17631);
nor U18474 (N_18474,N_17453,N_17281);
and U18475 (N_18475,N_17911,N_17909);
nor U18476 (N_18476,N_17131,N_17191);
and U18477 (N_18477,N_17648,N_17917);
nand U18478 (N_18478,N_17001,N_17505);
nor U18479 (N_18479,N_17011,N_17514);
nor U18480 (N_18480,N_17890,N_17328);
or U18481 (N_18481,N_17300,N_17990);
xor U18482 (N_18482,N_17806,N_17192);
xnor U18483 (N_18483,N_17612,N_17905);
xnor U18484 (N_18484,N_17136,N_17899);
nand U18485 (N_18485,N_17645,N_17424);
and U18486 (N_18486,N_17699,N_17921);
nand U18487 (N_18487,N_17507,N_17255);
nor U18488 (N_18488,N_17269,N_17721);
or U18489 (N_18489,N_17893,N_17114);
xor U18490 (N_18490,N_17071,N_17728);
nor U18491 (N_18491,N_17517,N_17084);
and U18492 (N_18492,N_17411,N_17231);
or U18493 (N_18493,N_17342,N_17628);
and U18494 (N_18494,N_17373,N_17477);
nand U18495 (N_18495,N_17135,N_17471);
or U18496 (N_18496,N_17316,N_17210);
nand U18497 (N_18497,N_17937,N_17204);
and U18498 (N_18498,N_17112,N_17459);
nand U18499 (N_18499,N_17087,N_17022);
nand U18500 (N_18500,N_17017,N_17753);
nor U18501 (N_18501,N_17460,N_17401);
nor U18502 (N_18502,N_17637,N_17617);
and U18503 (N_18503,N_17716,N_17076);
xnor U18504 (N_18504,N_17837,N_17630);
or U18505 (N_18505,N_17701,N_17966);
xnor U18506 (N_18506,N_17466,N_17942);
xor U18507 (N_18507,N_17636,N_17445);
or U18508 (N_18508,N_17009,N_17226);
nor U18509 (N_18509,N_17045,N_17273);
and U18510 (N_18510,N_17961,N_17839);
xnor U18511 (N_18511,N_17027,N_17220);
or U18512 (N_18512,N_17065,N_17968);
nand U18513 (N_18513,N_17399,N_17558);
xor U18514 (N_18514,N_17976,N_17577);
xnor U18515 (N_18515,N_17774,N_17830);
nand U18516 (N_18516,N_17151,N_17537);
and U18517 (N_18517,N_17830,N_17919);
nor U18518 (N_18518,N_17156,N_17053);
xnor U18519 (N_18519,N_17614,N_17737);
nand U18520 (N_18520,N_17563,N_17549);
nor U18521 (N_18521,N_17602,N_17830);
or U18522 (N_18522,N_17396,N_17708);
and U18523 (N_18523,N_17855,N_17401);
and U18524 (N_18524,N_17208,N_17968);
xor U18525 (N_18525,N_17903,N_17020);
nand U18526 (N_18526,N_17381,N_17853);
and U18527 (N_18527,N_17853,N_17095);
nor U18528 (N_18528,N_17641,N_17986);
nand U18529 (N_18529,N_17839,N_17569);
xnor U18530 (N_18530,N_17865,N_17665);
nand U18531 (N_18531,N_17075,N_17417);
and U18532 (N_18532,N_17961,N_17620);
or U18533 (N_18533,N_17666,N_17779);
nand U18534 (N_18534,N_17132,N_17803);
xor U18535 (N_18535,N_17915,N_17846);
nand U18536 (N_18536,N_17760,N_17661);
xor U18537 (N_18537,N_17000,N_17530);
nand U18538 (N_18538,N_17595,N_17132);
or U18539 (N_18539,N_17970,N_17037);
xor U18540 (N_18540,N_17075,N_17507);
nor U18541 (N_18541,N_17082,N_17907);
nand U18542 (N_18542,N_17618,N_17589);
and U18543 (N_18543,N_17921,N_17160);
nor U18544 (N_18544,N_17607,N_17072);
or U18545 (N_18545,N_17654,N_17996);
xor U18546 (N_18546,N_17206,N_17742);
nand U18547 (N_18547,N_17270,N_17567);
nand U18548 (N_18548,N_17740,N_17135);
nand U18549 (N_18549,N_17465,N_17870);
or U18550 (N_18550,N_17660,N_17801);
nor U18551 (N_18551,N_17980,N_17095);
nor U18552 (N_18552,N_17096,N_17991);
or U18553 (N_18553,N_17388,N_17598);
or U18554 (N_18554,N_17744,N_17774);
and U18555 (N_18555,N_17819,N_17797);
nand U18556 (N_18556,N_17369,N_17093);
and U18557 (N_18557,N_17578,N_17733);
nand U18558 (N_18558,N_17836,N_17732);
and U18559 (N_18559,N_17714,N_17938);
nand U18560 (N_18560,N_17358,N_17719);
nand U18561 (N_18561,N_17178,N_17905);
xor U18562 (N_18562,N_17716,N_17927);
nand U18563 (N_18563,N_17544,N_17645);
or U18564 (N_18564,N_17476,N_17606);
nand U18565 (N_18565,N_17586,N_17124);
and U18566 (N_18566,N_17514,N_17182);
nand U18567 (N_18567,N_17786,N_17500);
and U18568 (N_18568,N_17104,N_17889);
nor U18569 (N_18569,N_17415,N_17156);
nor U18570 (N_18570,N_17977,N_17742);
and U18571 (N_18571,N_17760,N_17433);
xnor U18572 (N_18572,N_17150,N_17708);
or U18573 (N_18573,N_17984,N_17987);
nor U18574 (N_18574,N_17314,N_17889);
xor U18575 (N_18575,N_17130,N_17949);
xnor U18576 (N_18576,N_17077,N_17872);
xor U18577 (N_18577,N_17669,N_17926);
and U18578 (N_18578,N_17120,N_17082);
nor U18579 (N_18579,N_17893,N_17375);
nand U18580 (N_18580,N_17931,N_17882);
or U18581 (N_18581,N_17196,N_17087);
nand U18582 (N_18582,N_17565,N_17382);
xor U18583 (N_18583,N_17454,N_17145);
and U18584 (N_18584,N_17135,N_17940);
nand U18585 (N_18585,N_17562,N_17801);
nor U18586 (N_18586,N_17826,N_17446);
or U18587 (N_18587,N_17585,N_17293);
or U18588 (N_18588,N_17341,N_17370);
nor U18589 (N_18589,N_17239,N_17270);
or U18590 (N_18590,N_17043,N_17012);
or U18591 (N_18591,N_17844,N_17623);
nor U18592 (N_18592,N_17699,N_17273);
and U18593 (N_18593,N_17996,N_17265);
xnor U18594 (N_18594,N_17037,N_17220);
and U18595 (N_18595,N_17300,N_17597);
nand U18596 (N_18596,N_17442,N_17873);
nand U18597 (N_18597,N_17872,N_17294);
or U18598 (N_18598,N_17442,N_17251);
and U18599 (N_18599,N_17336,N_17241);
and U18600 (N_18600,N_17448,N_17193);
nor U18601 (N_18601,N_17992,N_17825);
nand U18602 (N_18602,N_17011,N_17625);
nor U18603 (N_18603,N_17333,N_17327);
or U18604 (N_18604,N_17262,N_17560);
nand U18605 (N_18605,N_17481,N_17345);
xor U18606 (N_18606,N_17101,N_17582);
and U18607 (N_18607,N_17376,N_17339);
xor U18608 (N_18608,N_17940,N_17146);
nand U18609 (N_18609,N_17912,N_17137);
xnor U18610 (N_18610,N_17940,N_17487);
nor U18611 (N_18611,N_17719,N_17334);
or U18612 (N_18612,N_17931,N_17517);
and U18613 (N_18613,N_17469,N_17755);
or U18614 (N_18614,N_17438,N_17383);
or U18615 (N_18615,N_17842,N_17349);
nor U18616 (N_18616,N_17160,N_17655);
or U18617 (N_18617,N_17333,N_17551);
and U18618 (N_18618,N_17679,N_17096);
nand U18619 (N_18619,N_17607,N_17071);
nor U18620 (N_18620,N_17122,N_17488);
nor U18621 (N_18621,N_17856,N_17762);
or U18622 (N_18622,N_17732,N_17825);
or U18623 (N_18623,N_17205,N_17815);
xor U18624 (N_18624,N_17958,N_17997);
nand U18625 (N_18625,N_17369,N_17359);
nand U18626 (N_18626,N_17980,N_17163);
nor U18627 (N_18627,N_17810,N_17150);
and U18628 (N_18628,N_17020,N_17074);
nor U18629 (N_18629,N_17089,N_17780);
nor U18630 (N_18630,N_17402,N_17569);
nor U18631 (N_18631,N_17196,N_17880);
xnor U18632 (N_18632,N_17991,N_17269);
nand U18633 (N_18633,N_17326,N_17857);
nand U18634 (N_18634,N_17667,N_17664);
xor U18635 (N_18635,N_17203,N_17159);
nor U18636 (N_18636,N_17308,N_17181);
nand U18637 (N_18637,N_17859,N_17635);
or U18638 (N_18638,N_17753,N_17697);
and U18639 (N_18639,N_17368,N_17654);
or U18640 (N_18640,N_17241,N_17988);
xor U18641 (N_18641,N_17476,N_17661);
nand U18642 (N_18642,N_17053,N_17932);
nand U18643 (N_18643,N_17646,N_17690);
xnor U18644 (N_18644,N_17726,N_17179);
nand U18645 (N_18645,N_17226,N_17337);
xnor U18646 (N_18646,N_17842,N_17326);
nand U18647 (N_18647,N_17701,N_17164);
xnor U18648 (N_18648,N_17211,N_17679);
nand U18649 (N_18649,N_17614,N_17484);
nor U18650 (N_18650,N_17593,N_17732);
nor U18651 (N_18651,N_17518,N_17411);
xnor U18652 (N_18652,N_17240,N_17277);
xor U18653 (N_18653,N_17630,N_17294);
or U18654 (N_18654,N_17620,N_17083);
xor U18655 (N_18655,N_17610,N_17780);
and U18656 (N_18656,N_17260,N_17958);
or U18657 (N_18657,N_17377,N_17551);
xnor U18658 (N_18658,N_17904,N_17000);
nor U18659 (N_18659,N_17362,N_17609);
and U18660 (N_18660,N_17985,N_17430);
nor U18661 (N_18661,N_17675,N_17862);
nor U18662 (N_18662,N_17768,N_17965);
xor U18663 (N_18663,N_17627,N_17150);
or U18664 (N_18664,N_17806,N_17853);
nand U18665 (N_18665,N_17546,N_17584);
and U18666 (N_18666,N_17300,N_17027);
nand U18667 (N_18667,N_17948,N_17691);
nor U18668 (N_18668,N_17368,N_17135);
and U18669 (N_18669,N_17193,N_17397);
or U18670 (N_18670,N_17839,N_17438);
nand U18671 (N_18671,N_17650,N_17868);
nor U18672 (N_18672,N_17471,N_17122);
xnor U18673 (N_18673,N_17696,N_17377);
nor U18674 (N_18674,N_17559,N_17475);
or U18675 (N_18675,N_17629,N_17656);
or U18676 (N_18676,N_17753,N_17877);
nand U18677 (N_18677,N_17688,N_17461);
nor U18678 (N_18678,N_17772,N_17337);
nand U18679 (N_18679,N_17510,N_17067);
xnor U18680 (N_18680,N_17704,N_17864);
or U18681 (N_18681,N_17433,N_17600);
nor U18682 (N_18682,N_17944,N_17705);
nand U18683 (N_18683,N_17797,N_17581);
or U18684 (N_18684,N_17687,N_17931);
and U18685 (N_18685,N_17106,N_17795);
xor U18686 (N_18686,N_17352,N_17972);
nor U18687 (N_18687,N_17388,N_17350);
or U18688 (N_18688,N_17272,N_17590);
and U18689 (N_18689,N_17936,N_17482);
or U18690 (N_18690,N_17086,N_17651);
nand U18691 (N_18691,N_17258,N_17273);
or U18692 (N_18692,N_17766,N_17235);
nand U18693 (N_18693,N_17819,N_17599);
and U18694 (N_18694,N_17963,N_17309);
nand U18695 (N_18695,N_17553,N_17294);
nor U18696 (N_18696,N_17290,N_17258);
or U18697 (N_18697,N_17612,N_17327);
nor U18698 (N_18698,N_17224,N_17843);
or U18699 (N_18699,N_17573,N_17166);
nor U18700 (N_18700,N_17471,N_17999);
xor U18701 (N_18701,N_17251,N_17026);
nor U18702 (N_18702,N_17097,N_17707);
nand U18703 (N_18703,N_17837,N_17200);
nand U18704 (N_18704,N_17706,N_17555);
nor U18705 (N_18705,N_17190,N_17604);
xor U18706 (N_18706,N_17525,N_17972);
or U18707 (N_18707,N_17006,N_17679);
or U18708 (N_18708,N_17390,N_17192);
or U18709 (N_18709,N_17193,N_17560);
xor U18710 (N_18710,N_17648,N_17902);
nand U18711 (N_18711,N_17181,N_17998);
and U18712 (N_18712,N_17580,N_17634);
and U18713 (N_18713,N_17081,N_17976);
nor U18714 (N_18714,N_17687,N_17362);
xnor U18715 (N_18715,N_17610,N_17814);
or U18716 (N_18716,N_17253,N_17641);
xor U18717 (N_18717,N_17759,N_17738);
nor U18718 (N_18718,N_17284,N_17112);
nor U18719 (N_18719,N_17251,N_17101);
or U18720 (N_18720,N_17741,N_17651);
and U18721 (N_18721,N_17927,N_17849);
nor U18722 (N_18722,N_17973,N_17038);
nand U18723 (N_18723,N_17357,N_17222);
nor U18724 (N_18724,N_17450,N_17265);
nand U18725 (N_18725,N_17015,N_17983);
nor U18726 (N_18726,N_17712,N_17873);
nand U18727 (N_18727,N_17372,N_17172);
and U18728 (N_18728,N_17443,N_17339);
and U18729 (N_18729,N_17459,N_17224);
or U18730 (N_18730,N_17062,N_17110);
or U18731 (N_18731,N_17643,N_17348);
or U18732 (N_18732,N_17306,N_17344);
nand U18733 (N_18733,N_17960,N_17395);
xnor U18734 (N_18734,N_17092,N_17191);
nor U18735 (N_18735,N_17260,N_17525);
nor U18736 (N_18736,N_17227,N_17161);
and U18737 (N_18737,N_17046,N_17148);
xor U18738 (N_18738,N_17401,N_17391);
nand U18739 (N_18739,N_17562,N_17862);
xor U18740 (N_18740,N_17495,N_17801);
xor U18741 (N_18741,N_17437,N_17149);
and U18742 (N_18742,N_17544,N_17361);
or U18743 (N_18743,N_17468,N_17789);
and U18744 (N_18744,N_17885,N_17921);
nor U18745 (N_18745,N_17376,N_17406);
xor U18746 (N_18746,N_17339,N_17085);
nor U18747 (N_18747,N_17771,N_17116);
xor U18748 (N_18748,N_17624,N_17750);
nor U18749 (N_18749,N_17951,N_17533);
nor U18750 (N_18750,N_17867,N_17616);
xnor U18751 (N_18751,N_17981,N_17877);
nand U18752 (N_18752,N_17131,N_17433);
and U18753 (N_18753,N_17784,N_17431);
or U18754 (N_18754,N_17919,N_17266);
nor U18755 (N_18755,N_17279,N_17907);
or U18756 (N_18756,N_17023,N_17750);
nor U18757 (N_18757,N_17100,N_17110);
nor U18758 (N_18758,N_17799,N_17399);
or U18759 (N_18759,N_17350,N_17484);
nand U18760 (N_18760,N_17187,N_17104);
xor U18761 (N_18761,N_17027,N_17228);
or U18762 (N_18762,N_17662,N_17014);
xnor U18763 (N_18763,N_17163,N_17579);
nand U18764 (N_18764,N_17426,N_17521);
nor U18765 (N_18765,N_17085,N_17867);
or U18766 (N_18766,N_17966,N_17559);
nor U18767 (N_18767,N_17688,N_17179);
xnor U18768 (N_18768,N_17581,N_17599);
nor U18769 (N_18769,N_17054,N_17898);
and U18770 (N_18770,N_17133,N_17560);
xor U18771 (N_18771,N_17769,N_17207);
xor U18772 (N_18772,N_17940,N_17268);
and U18773 (N_18773,N_17554,N_17698);
nand U18774 (N_18774,N_17567,N_17177);
nand U18775 (N_18775,N_17571,N_17686);
or U18776 (N_18776,N_17829,N_17686);
nor U18777 (N_18777,N_17535,N_17979);
nor U18778 (N_18778,N_17065,N_17087);
and U18779 (N_18779,N_17135,N_17375);
or U18780 (N_18780,N_17798,N_17668);
or U18781 (N_18781,N_17431,N_17992);
nand U18782 (N_18782,N_17033,N_17533);
nor U18783 (N_18783,N_17383,N_17331);
or U18784 (N_18784,N_17649,N_17337);
nor U18785 (N_18785,N_17611,N_17026);
nand U18786 (N_18786,N_17011,N_17912);
and U18787 (N_18787,N_17611,N_17560);
nand U18788 (N_18788,N_17656,N_17441);
and U18789 (N_18789,N_17378,N_17282);
nand U18790 (N_18790,N_17918,N_17629);
nor U18791 (N_18791,N_17976,N_17454);
and U18792 (N_18792,N_17482,N_17247);
xor U18793 (N_18793,N_17066,N_17111);
nor U18794 (N_18794,N_17368,N_17733);
or U18795 (N_18795,N_17421,N_17834);
nand U18796 (N_18796,N_17618,N_17067);
nor U18797 (N_18797,N_17142,N_17364);
or U18798 (N_18798,N_17995,N_17239);
or U18799 (N_18799,N_17263,N_17175);
or U18800 (N_18800,N_17259,N_17185);
and U18801 (N_18801,N_17871,N_17392);
nand U18802 (N_18802,N_17921,N_17579);
and U18803 (N_18803,N_17015,N_17682);
nand U18804 (N_18804,N_17111,N_17337);
and U18805 (N_18805,N_17550,N_17455);
and U18806 (N_18806,N_17566,N_17450);
nor U18807 (N_18807,N_17114,N_17259);
xor U18808 (N_18808,N_17104,N_17459);
nand U18809 (N_18809,N_17898,N_17829);
nand U18810 (N_18810,N_17022,N_17897);
nor U18811 (N_18811,N_17067,N_17430);
nand U18812 (N_18812,N_17839,N_17481);
nand U18813 (N_18813,N_17852,N_17177);
or U18814 (N_18814,N_17763,N_17347);
and U18815 (N_18815,N_17834,N_17625);
nor U18816 (N_18816,N_17284,N_17059);
xnor U18817 (N_18817,N_17107,N_17285);
and U18818 (N_18818,N_17993,N_17442);
and U18819 (N_18819,N_17028,N_17708);
and U18820 (N_18820,N_17898,N_17926);
nor U18821 (N_18821,N_17720,N_17798);
and U18822 (N_18822,N_17105,N_17783);
xor U18823 (N_18823,N_17928,N_17990);
xor U18824 (N_18824,N_17986,N_17744);
nand U18825 (N_18825,N_17119,N_17704);
and U18826 (N_18826,N_17703,N_17369);
nand U18827 (N_18827,N_17129,N_17209);
or U18828 (N_18828,N_17145,N_17154);
or U18829 (N_18829,N_17305,N_17769);
xnor U18830 (N_18830,N_17832,N_17482);
nand U18831 (N_18831,N_17156,N_17104);
xnor U18832 (N_18832,N_17892,N_17288);
xnor U18833 (N_18833,N_17255,N_17730);
nand U18834 (N_18834,N_17003,N_17680);
xnor U18835 (N_18835,N_17483,N_17615);
nor U18836 (N_18836,N_17940,N_17234);
nand U18837 (N_18837,N_17023,N_17275);
nand U18838 (N_18838,N_17143,N_17052);
xnor U18839 (N_18839,N_17023,N_17092);
and U18840 (N_18840,N_17234,N_17091);
or U18841 (N_18841,N_17504,N_17690);
or U18842 (N_18842,N_17189,N_17809);
xnor U18843 (N_18843,N_17304,N_17597);
nor U18844 (N_18844,N_17451,N_17062);
xor U18845 (N_18845,N_17242,N_17114);
and U18846 (N_18846,N_17149,N_17559);
nand U18847 (N_18847,N_17457,N_17538);
and U18848 (N_18848,N_17156,N_17484);
xnor U18849 (N_18849,N_17823,N_17340);
nand U18850 (N_18850,N_17475,N_17802);
nand U18851 (N_18851,N_17565,N_17300);
nand U18852 (N_18852,N_17426,N_17670);
nand U18853 (N_18853,N_17902,N_17721);
and U18854 (N_18854,N_17261,N_17866);
and U18855 (N_18855,N_17104,N_17638);
or U18856 (N_18856,N_17743,N_17431);
nand U18857 (N_18857,N_17897,N_17351);
xor U18858 (N_18858,N_17913,N_17763);
or U18859 (N_18859,N_17116,N_17650);
nor U18860 (N_18860,N_17003,N_17777);
or U18861 (N_18861,N_17970,N_17681);
and U18862 (N_18862,N_17411,N_17457);
nor U18863 (N_18863,N_17520,N_17418);
xor U18864 (N_18864,N_17436,N_17189);
nor U18865 (N_18865,N_17422,N_17193);
nor U18866 (N_18866,N_17414,N_17347);
nor U18867 (N_18867,N_17310,N_17109);
or U18868 (N_18868,N_17782,N_17429);
or U18869 (N_18869,N_17550,N_17883);
or U18870 (N_18870,N_17356,N_17324);
and U18871 (N_18871,N_17260,N_17572);
nand U18872 (N_18872,N_17355,N_17716);
and U18873 (N_18873,N_17890,N_17055);
or U18874 (N_18874,N_17299,N_17803);
nand U18875 (N_18875,N_17484,N_17557);
or U18876 (N_18876,N_17347,N_17041);
nand U18877 (N_18877,N_17309,N_17607);
nand U18878 (N_18878,N_17899,N_17078);
or U18879 (N_18879,N_17566,N_17811);
or U18880 (N_18880,N_17349,N_17381);
and U18881 (N_18881,N_17280,N_17971);
or U18882 (N_18882,N_17553,N_17075);
nor U18883 (N_18883,N_17468,N_17278);
or U18884 (N_18884,N_17079,N_17719);
xnor U18885 (N_18885,N_17379,N_17857);
nand U18886 (N_18886,N_17949,N_17248);
and U18887 (N_18887,N_17569,N_17868);
xor U18888 (N_18888,N_17664,N_17038);
nand U18889 (N_18889,N_17587,N_17760);
or U18890 (N_18890,N_17346,N_17418);
nand U18891 (N_18891,N_17291,N_17966);
nand U18892 (N_18892,N_17676,N_17321);
and U18893 (N_18893,N_17118,N_17162);
xor U18894 (N_18894,N_17092,N_17050);
nor U18895 (N_18895,N_17974,N_17342);
or U18896 (N_18896,N_17405,N_17154);
nor U18897 (N_18897,N_17497,N_17610);
or U18898 (N_18898,N_17996,N_17916);
and U18899 (N_18899,N_17740,N_17156);
nand U18900 (N_18900,N_17856,N_17026);
or U18901 (N_18901,N_17487,N_17908);
and U18902 (N_18902,N_17984,N_17083);
nor U18903 (N_18903,N_17770,N_17659);
and U18904 (N_18904,N_17103,N_17803);
nand U18905 (N_18905,N_17610,N_17722);
nor U18906 (N_18906,N_17775,N_17004);
xnor U18907 (N_18907,N_17014,N_17509);
and U18908 (N_18908,N_17701,N_17163);
or U18909 (N_18909,N_17281,N_17689);
xor U18910 (N_18910,N_17564,N_17640);
nor U18911 (N_18911,N_17413,N_17148);
or U18912 (N_18912,N_17304,N_17365);
nand U18913 (N_18913,N_17208,N_17771);
or U18914 (N_18914,N_17462,N_17537);
nor U18915 (N_18915,N_17933,N_17214);
nor U18916 (N_18916,N_17408,N_17107);
nor U18917 (N_18917,N_17919,N_17358);
xor U18918 (N_18918,N_17891,N_17315);
and U18919 (N_18919,N_17021,N_17363);
or U18920 (N_18920,N_17028,N_17050);
and U18921 (N_18921,N_17817,N_17657);
nand U18922 (N_18922,N_17028,N_17944);
or U18923 (N_18923,N_17339,N_17566);
xnor U18924 (N_18924,N_17873,N_17454);
nor U18925 (N_18925,N_17508,N_17335);
or U18926 (N_18926,N_17368,N_17306);
nor U18927 (N_18927,N_17543,N_17924);
xnor U18928 (N_18928,N_17183,N_17938);
and U18929 (N_18929,N_17506,N_17999);
or U18930 (N_18930,N_17428,N_17480);
nor U18931 (N_18931,N_17524,N_17441);
nand U18932 (N_18932,N_17473,N_17655);
or U18933 (N_18933,N_17296,N_17124);
nor U18934 (N_18934,N_17321,N_17872);
and U18935 (N_18935,N_17095,N_17741);
and U18936 (N_18936,N_17250,N_17747);
xnor U18937 (N_18937,N_17281,N_17489);
and U18938 (N_18938,N_17900,N_17518);
nand U18939 (N_18939,N_17120,N_17604);
and U18940 (N_18940,N_17961,N_17145);
or U18941 (N_18941,N_17607,N_17184);
and U18942 (N_18942,N_17983,N_17977);
xnor U18943 (N_18943,N_17274,N_17973);
and U18944 (N_18944,N_17447,N_17887);
or U18945 (N_18945,N_17651,N_17841);
xor U18946 (N_18946,N_17233,N_17895);
or U18947 (N_18947,N_17348,N_17271);
nand U18948 (N_18948,N_17041,N_17781);
and U18949 (N_18949,N_17717,N_17589);
xnor U18950 (N_18950,N_17594,N_17486);
xor U18951 (N_18951,N_17775,N_17118);
and U18952 (N_18952,N_17481,N_17081);
or U18953 (N_18953,N_17450,N_17057);
and U18954 (N_18954,N_17544,N_17937);
and U18955 (N_18955,N_17532,N_17411);
nor U18956 (N_18956,N_17733,N_17418);
nor U18957 (N_18957,N_17113,N_17765);
nor U18958 (N_18958,N_17853,N_17746);
nor U18959 (N_18959,N_17867,N_17791);
xor U18960 (N_18960,N_17155,N_17009);
nand U18961 (N_18961,N_17467,N_17319);
xor U18962 (N_18962,N_17402,N_17870);
and U18963 (N_18963,N_17260,N_17327);
or U18964 (N_18964,N_17944,N_17085);
nor U18965 (N_18965,N_17667,N_17606);
or U18966 (N_18966,N_17043,N_17707);
nor U18967 (N_18967,N_17878,N_17766);
nor U18968 (N_18968,N_17574,N_17860);
or U18969 (N_18969,N_17883,N_17087);
xor U18970 (N_18970,N_17052,N_17878);
nand U18971 (N_18971,N_17170,N_17810);
and U18972 (N_18972,N_17713,N_17343);
nand U18973 (N_18973,N_17061,N_17891);
nand U18974 (N_18974,N_17423,N_17876);
or U18975 (N_18975,N_17927,N_17066);
and U18976 (N_18976,N_17513,N_17433);
xnor U18977 (N_18977,N_17993,N_17602);
nor U18978 (N_18978,N_17629,N_17464);
and U18979 (N_18979,N_17425,N_17129);
nor U18980 (N_18980,N_17250,N_17151);
or U18981 (N_18981,N_17806,N_17811);
nor U18982 (N_18982,N_17731,N_17237);
and U18983 (N_18983,N_17216,N_17967);
and U18984 (N_18984,N_17673,N_17687);
or U18985 (N_18985,N_17088,N_17123);
nand U18986 (N_18986,N_17944,N_17556);
nand U18987 (N_18987,N_17233,N_17366);
or U18988 (N_18988,N_17751,N_17965);
nand U18989 (N_18989,N_17333,N_17320);
xnor U18990 (N_18990,N_17576,N_17616);
or U18991 (N_18991,N_17369,N_17339);
and U18992 (N_18992,N_17231,N_17643);
nor U18993 (N_18993,N_17822,N_17140);
xor U18994 (N_18994,N_17234,N_17739);
and U18995 (N_18995,N_17217,N_17843);
nor U18996 (N_18996,N_17161,N_17613);
and U18997 (N_18997,N_17100,N_17886);
nand U18998 (N_18998,N_17105,N_17178);
nand U18999 (N_18999,N_17039,N_17801);
nor U19000 (N_19000,N_18120,N_18811);
xor U19001 (N_19001,N_18662,N_18507);
or U19002 (N_19002,N_18384,N_18223);
nor U19003 (N_19003,N_18670,N_18289);
or U19004 (N_19004,N_18126,N_18537);
xnor U19005 (N_19005,N_18855,N_18242);
and U19006 (N_19006,N_18191,N_18912);
and U19007 (N_19007,N_18571,N_18613);
or U19008 (N_19008,N_18689,N_18598);
and U19009 (N_19009,N_18683,N_18486);
and U19010 (N_19010,N_18018,N_18642);
nor U19011 (N_19011,N_18247,N_18631);
nand U19012 (N_19012,N_18359,N_18806);
nand U19013 (N_19013,N_18434,N_18625);
nand U19014 (N_19014,N_18213,N_18583);
nand U19015 (N_19015,N_18827,N_18337);
and U19016 (N_19016,N_18921,N_18224);
nor U19017 (N_19017,N_18814,N_18996);
or U19018 (N_19018,N_18742,N_18065);
nand U19019 (N_19019,N_18719,N_18254);
and U19020 (N_19020,N_18380,N_18973);
xnor U19021 (N_19021,N_18949,N_18676);
and U19022 (N_19022,N_18350,N_18512);
nand U19023 (N_19023,N_18734,N_18250);
nand U19024 (N_19024,N_18659,N_18011);
nor U19025 (N_19025,N_18101,N_18252);
or U19026 (N_19026,N_18978,N_18294);
xnor U19027 (N_19027,N_18748,N_18958);
and U19028 (N_19028,N_18131,N_18758);
or U19029 (N_19029,N_18189,N_18526);
and U19030 (N_19030,N_18000,N_18162);
nor U19031 (N_19031,N_18439,N_18248);
nor U19032 (N_19032,N_18013,N_18096);
nand U19033 (N_19033,N_18136,N_18995);
nand U19034 (N_19034,N_18559,N_18493);
nor U19035 (N_19035,N_18737,N_18186);
and U19036 (N_19036,N_18297,N_18857);
and U19037 (N_19037,N_18030,N_18938);
or U19038 (N_19038,N_18476,N_18954);
nor U19039 (N_19039,N_18933,N_18302);
or U19040 (N_19040,N_18951,N_18528);
xor U19041 (N_19041,N_18455,N_18948);
nor U19042 (N_19042,N_18316,N_18522);
nand U19043 (N_19043,N_18220,N_18338);
or U19044 (N_19044,N_18044,N_18356);
and U19045 (N_19045,N_18744,N_18892);
nor U19046 (N_19046,N_18703,N_18490);
nand U19047 (N_19047,N_18881,N_18728);
or U19048 (N_19048,N_18424,N_18389);
nand U19049 (N_19049,N_18756,N_18622);
and U19050 (N_19050,N_18779,N_18755);
xor U19051 (N_19051,N_18792,N_18176);
nor U19052 (N_19052,N_18460,N_18679);
xor U19053 (N_19053,N_18397,N_18109);
or U19054 (N_19054,N_18075,N_18130);
nand U19055 (N_19055,N_18898,N_18196);
nor U19056 (N_19056,N_18444,N_18385);
or U19057 (N_19057,N_18374,N_18909);
xor U19058 (N_19058,N_18729,N_18407);
nand U19059 (N_19059,N_18172,N_18435);
xor U19060 (N_19060,N_18055,N_18817);
xor U19061 (N_19061,N_18104,N_18969);
or U19062 (N_19062,N_18227,N_18416);
xnor U19063 (N_19063,N_18040,N_18853);
nand U19064 (N_19064,N_18209,N_18941);
nor U19065 (N_19065,N_18849,N_18253);
nor U19066 (N_19066,N_18669,N_18680);
xor U19067 (N_19067,N_18555,N_18873);
and U19068 (N_19068,N_18860,N_18922);
or U19069 (N_19069,N_18970,N_18709);
nor U19070 (N_19070,N_18276,N_18904);
nor U19071 (N_19071,N_18212,N_18009);
xnor U19072 (N_19072,N_18574,N_18475);
and U19073 (N_19073,N_18449,N_18417);
or U19074 (N_19074,N_18829,N_18210);
or U19075 (N_19075,N_18722,N_18980);
and U19076 (N_19076,N_18428,N_18221);
nand U19077 (N_19077,N_18433,N_18815);
nor U19078 (N_19078,N_18119,N_18666);
and U19079 (N_19079,N_18095,N_18751);
xnor U19080 (N_19080,N_18968,N_18916);
or U19081 (N_19081,N_18685,N_18557);
or U19082 (N_19082,N_18149,N_18137);
xor U19083 (N_19083,N_18919,N_18003);
xnor U19084 (N_19084,N_18905,N_18303);
and U19085 (N_19085,N_18931,N_18777);
nand U19086 (N_19086,N_18262,N_18151);
or U19087 (N_19087,N_18646,N_18183);
nor U19088 (N_19088,N_18170,N_18627);
or U19089 (N_19089,N_18844,N_18200);
xor U19090 (N_19090,N_18267,N_18166);
or U19091 (N_19091,N_18298,N_18266);
or U19092 (N_19092,N_18379,N_18010);
nor U19093 (N_19093,N_18828,N_18481);
nand U19094 (N_19094,N_18606,N_18317);
and U19095 (N_19095,N_18309,N_18208);
or U19096 (N_19096,N_18002,N_18611);
nand U19097 (N_19097,N_18390,N_18341);
nor U19098 (N_19098,N_18937,N_18988);
or U19099 (N_19099,N_18184,N_18896);
xnor U19100 (N_19100,N_18783,N_18713);
or U19101 (N_19101,N_18863,N_18715);
and U19102 (N_19102,N_18071,N_18875);
or U19103 (N_19103,N_18647,N_18408);
and U19104 (N_19104,N_18946,N_18843);
xnor U19105 (N_19105,N_18764,N_18488);
nor U19106 (N_19106,N_18445,N_18738);
or U19107 (N_19107,N_18834,N_18865);
nand U19108 (N_19108,N_18947,N_18020);
nand U19109 (N_19109,N_18577,N_18567);
nor U19110 (N_19110,N_18401,N_18619);
nor U19111 (N_19111,N_18634,N_18185);
and U19112 (N_19112,N_18100,N_18017);
and U19113 (N_19113,N_18610,N_18386);
nand U19114 (N_19114,N_18382,N_18469);
nor U19115 (N_19115,N_18903,N_18285);
nor U19116 (N_19116,N_18004,N_18496);
nand U19117 (N_19117,N_18305,N_18824);
xnor U19118 (N_19118,N_18510,N_18960);
or U19119 (N_19119,N_18993,N_18800);
nand U19120 (N_19120,N_18812,N_18957);
and U19121 (N_19121,N_18315,N_18048);
xnor U19122 (N_19122,N_18695,N_18110);
xor U19123 (N_19123,N_18655,N_18246);
nor U19124 (N_19124,N_18731,N_18335);
xnor U19125 (N_19125,N_18842,N_18106);
nand U19126 (N_19126,N_18556,N_18767);
nand U19127 (N_19127,N_18098,N_18187);
nand U19128 (N_19128,N_18886,N_18160);
nand U19129 (N_19129,N_18866,N_18026);
and U19130 (N_19130,N_18603,N_18550);
nor U19131 (N_19131,N_18042,N_18362);
or U19132 (N_19132,N_18083,N_18754);
nand U19133 (N_19133,N_18545,N_18453);
or U19134 (N_19134,N_18641,N_18236);
xnor U19135 (N_19135,N_18950,N_18161);
xor U19136 (N_19136,N_18601,N_18699);
or U19137 (N_19137,N_18736,N_18513);
nand U19138 (N_19138,N_18923,N_18205);
or U19139 (N_19139,N_18412,N_18821);
xor U19140 (N_19140,N_18668,N_18838);
nor U19141 (N_19141,N_18217,N_18678);
xor U19142 (N_19142,N_18192,N_18776);
xor U19143 (N_19143,N_18897,N_18354);
xnor U19144 (N_19144,N_18256,N_18630);
or U19145 (N_19145,N_18918,N_18539);
nand U19146 (N_19146,N_18893,N_18122);
xor U19147 (N_19147,N_18039,N_18971);
and U19148 (N_19148,N_18399,N_18464);
nor U19149 (N_19149,N_18050,N_18264);
xor U19150 (N_19150,N_18334,N_18753);
nor U19151 (N_19151,N_18222,N_18259);
xnor U19152 (N_19152,N_18494,N_18770);
xnor U19153 (N_19153,N_18007,N_18295);
or U19154 (N_19154,N_18984,N_18740);
and U19155 (N_19155,N_18752,N_18629);
nand U19156 (N_19156,N_18330,N_18311);
and U19157 (N_19157,N_18956,N_18281);
and U19158 (N_19158,N_18099,N_18308);
xor U19159 (N_19159,N_18690,N_18602);
nand U19160 (N_19160,N_18965,N_18203);
and U19161 (N_19161,N_18219,N_18381);
nand U19162 (N_19162,N_18563,N_18405);
nor U19163 (N_19163,N_18426,N_18833);
xnor U19164 (N_19164,N_18066,N_18070);
nor U19165 (N_19165,N_18310,N_18600);
nand U19166 (N_19166,N_18480,N_18499);
and U19167 (N_19167,N_18218,N_18440);
xor U19168 (N_19168,N_18299,N_18019);
xnor U19169 (N_19169,N_18796,N_18643);
xnor U19170 (N_19170,N_18194,N_18874);
and U19171 (N_19171,N_18051,N_18135);
xor U19172 (N_19172,N_18179,N_18979);
nor U19173 (N_19173,N_18421,N_18193);
xor U19174 (N_19174,N_18608,N_18472);
xnor U19175 (N_19175,N_18663,N_18422);
xor U19176 (N_19176,N_18997,N_18073);
and U19177 (N_19177,N_18465,N_18762);
and U19178 (N_19178,N_18794,N_18702);
nor U19179 (N_19179,N_18558,N_18708);
and U19180 (N_19180,N_18547,N_18721);
and U19181 (N_19181,N_18269,N_18594);
and U19182 (N_19182,N_18793,N_18944);
and U19183 (N_19183,N_18432,N_18573);
nand U19184 (N_19184,N_18133,N_18759);
nand U19185 (N_19185,N_18928,N_18816);
or U19186 (N_19186,N_18998,N_18532);
nand U19187 (N_19187,N_18458,N_18967);
nor U19188 (N_19188,N_18901,N_18983);
and U19189 (N_19189,N_18845,N_18324);
or U19190 (N_19190,N_18060,N_18204);
nor U19191 (N_19191,N_18199,N_18607);
and U19192 (N_19192,N_18275,N_18406);
or U19193 (N_19193,N_18312,N_18357);
xor U19194 (N_19194,N_18700,N_18624);
or U19195 (N_19195,N_18609,N_18163);
xor U19196 (N_19196,N_18047,N_18841);
and U19197 (N_19197,N_18032,N_18878);
xnor U19198 (N_19198,N_18372,N_18913);
nand U19199 (N_19199,N_18470,N_18115);
nor U19200 (N_19200,N_18329,N_18502);
nand U19201 (N_19201,N_18791,N_18053);
xor U19202 (N_19202,N_18045,N_18370);
and U19203 (N_19203,N_18977,N_18024);
and U19204 (N_19204,N_18087,N_18533);
nor U19205 (N_19205,N_18705,N_18962);
and U19206 (N_19206,N_18945,N_18462);
nand U19207 (N_19207,N_18143,N_18771);
nor U19208 (N_19208,N_18725,N_18798);
or U19209 (N_19209,N_18414,N_18012);
nand U19210 (N_19210,N_18714,N_18684);
nor U19211 (N_19211,N_18438,N_18727);
and U19212 (N_19212,N_18241,N_18819);
or U19213 (N_19213,N_18626,N_18884);
xor U19214 (N_19214,N_18207,N_18640);
and U19215 (N_19215,N_18278,N_18079);
and U19216 (N_19216,N_18076,N_18368);
and U19217 (N_19217,N_18720,N_18615);
or U19218 (N_19218,N_18255,N_18046);
nor U19219 (N_19219,N_18711,N_18645);
nor U19220 (N_19220,N_18342,N_18105);
nor U19221 (N_19221,N_18768,N_18775);
xnor U19222 (N_19222,N_18282,N_18346);
nor U19223 (N_19223,N_18038,N_18743);
or U19224 (N_19224,N_18936,N_18336);
nand U19225 (N_19225,N_18323,N_18840);
nand U19226 (N_19226,N_18760,N_18457);
nor U19227 (N_19227,N_18672,N_18847);
and U19228 (N_19228,N_18301,N_18769);
and U19229 (N_19229,N_18590,N_18831);
or U19230 (N_19230,N_18077,N_18925);
nor U19231 (N_19231,N_18034,N_18345);
nand U19232 (N_19232,N_18581,N_18400);
xor U19233 (N_19233,N_18987,N_18850);
nand U19234 (N_19234,N_18569,N_18333);
or U19235 (N_19235,N_18072,N_18484);
and U19236 (N_19236,N_18786,N_18326);
xnor U19237 (N_19237,N_18803,N_18063);
xor U19238 (N_19238,N_18261,N_18249);
or U19239 (N_19239,N_18461,N_18570);
xnor U19240 (N_19240,N_18652,N_18534);
and U19241 (N_19241,N_18154,N_18491);
xor U19242 (N_19242,N_18851,N_18092);
or U19243 (N_19243,N_18891,N_18704);
nor U19244 (N_19244,N_18041,N_18902);
nand U19245 (N_19245,N_18351,N_18466);
xor U19246 (N_19246,N_18353,N_18932);
nand U19247 (N_19247,N_18366,N_18450);
or U19248 (N_19248,N_18848,N_18393);
or U19249 (N_19249,N_18674,N_18809);
xor U19250 (N_19250,N_18430,N_18781);
xor U19251 (N_19251,N_18516,N_18313);
nor U19252 (N_19252,N_18656,N_18061);
xor U19253 (N_19253,N_18832,N_18930);
nor U19254 (N_19254,N_18085,N_18067);
or U19255 (N_19255,N_18177,N_18623);
or U19256 (N_19256,N_18358,N_18520);
and U19257 (N_19257,N_18963,N_18653);
nor U19258 (N_19258,N_18612,N_18530);
xor U19259 (N_19259,N_18173,N_18485);
nand U19260 (N_19260,N_18052,N_18344);
and U19261 (N_19261,N_18155,N_18395);
xor U19262 (N_19262,N_18495,N_18054);
nor U19263 (N_19263,N_18686,N_18211);
nand U19264 (N_19264,N_18637,N_18468);
or U19265 (N_19265,N_18911,N_18283);
or U19266 (N_19266,N_18089,N_18926);
nand U19267 (N_19267,N_18976,N_18745);
nand U19268 (N_19268,N_18023,N_18907);
xor U19269 (N_19269,N_18387,N_18942);
nor U19270 (N_19270,N_18235,N_18867);
and U19271 (N_19271,N_18314,N_18215);
or U19272 (N_19272,N_18291,N_18638);
nand U19273 (N_19273,N_18810,N_18139);
xnor U19274 (N_19274,N_18290,N_18882);
nor U19275 (N_19275,N_18142,N_18028);
nor U19276 (N_19276,N_18578,N_18566);
nor U19277 (N_19277,N_18887,N_18492);
and U19278 (N_19278,N_18031,N_18665);
or U19279 (N_19279,N_18425,N_18503);
nand U19280 (N_19280,N_18562,N_18989);
nand U19281 (N_19281,N_18726,N_18826);
xor U19282 (N_19282,N_18015,N_18489);
nor U19283 (N_19283,N_18103,N_18535);
or U19284 (N_19284,N_18088,N_18304);
xor U19285 (N_19285,N_18251,N_18735);
or U19286 (N_19286,N_18917,N_18145);
and U19287 (N_19287,N_18616,N_18361);
xor U19288 (N_19288,N_18339,N_18182);
nand U19289 (N_19289,N_18620,N_18858);
nor U19290 (N_19290,N_18146,N_18772);
xor U19291 (N_19291,N_18148,N_18966);
or U19292 (N_19292,N_18328,N_18140);
or U19293 (N_19293,N_18093,N_18724);
nor U19294 (N_19294,N_18195,N_18546);
nand U19295 (N_19295,N_18431,N_18080);
and U19296 (N_19296,N_18201,N_18746);
nand U19297 (N_19297,N_18953,N_18749);
nor U19298 (N_19298,N_18514,N_18320);
and U19299 (N_19299,N_18447,N_18349);
xor U19300 (N_19300,N_18765,N_18774);
and U19301 (N_19301,N_18138,N_18293);
nor U19302 (N_19302,N_18270,N_18006);
nand U19303 (N_19303,N_18591,N_18885);
or U19304 (N_19304,N_18257,N_18644);
nand U19305 (N_19305,N_18097,N_18132);
or U19306 (N_19306,N_18994,N_18228);
nor U19307 (N_19307,N_18197,N_18820);
and U19308 (N_19308,N_18376,N_18016);
nand U19309 (N_19309,N_18823,N_18234);
nor U19310 (N_19310,N_18561,N_18542);
or U19311 (N_19311,N_18575,N_18157);
nor U19312 (N_19312,N_18959,N_18322);
xor U19313 (N_19313,N_18274,N_18165);
xnor U19314 (N_19314,N_18279,N_18604);
or U19315 (N_19315,N_18058,N_18617);
or U19316 (N_19316,N_18605,N_18411);
nor U19317 (N_19317,N_18784,N_18409);
nand U19318 (N_19318,N_18799,N_18156);
xnor U19319 (N_19319,N_18924,N_18862);
xor U19320 (N_19320,N_18579,N_18785);
nor U19321 (N_19321,N_18914,N_18482);
or U19322 (N_19322,N_18467,N_18498);
nand U19323 (N_19323,N_18021,N_18548);
nand U19324 (N_19324,N_18108,N_18568);
nor U19325 (N_19325,N_18580,N_18231);
and U19326 (N_19326,N_18692,N_18635);
nand U19327 (N_19327,N_18152,N_18391);
nor U19328 (N_19328,N_18446,N_18168);
or U19329 (N_19329,N_18084,N_18029);
nor U19330 (N_19330,N_18899,N_18325);
xor U19331 (N_19331,N_18505,N_18694);
nor U19332 (N_19332,N_18375,N_18852);
nor U19333 (N_19333,N_18750,N_18477);
nand U19334 (N_19334,N_18332,N_18258);
nor U19335 (N_19335,N_18529,N_18801);
or U19336 (N_19336,N_18373,N_18141);
nor U19337 (N_19337,N_18651,N_18111);
and U19338 (N_19338,N_18908,N_18473);
nor U19339 (N_19339,N_18518,N_18697);
and U19340 (N_19340,N_18365,N_18733);
or U19341 (N_19341,N_18500,N_18369);
nor U19342 (N_19342,N_18915,N_18519);
xnor U19343 (N_19343,N_18036,N_18701);
nor U19344 (N_19344,N_18363,N_18982);
or U19345 (N_19345,N_18698,N_18732);
nor U19346 (N_19346,N_18463,N_18716);
xor U19347 (N_19347,N_18273,N_18091);
or U19348 (N_19348,N_18658,N_18232);
and U19349 (N_19349,N_18596,N_18747);
xnor U19350 (N_19350,N_18509,N_18990);
and U19351 (N_19351,N_18069,N_18240);
and U19352 (N_19352,N_18022,N_18565);
or U19353 (N_19353,N_18420,N_18167);
nand U19354 (N_19354,N_18836,N_18551);
xor U19355 (N_19355,N_18288,N_18696);
nor U19356 (N_19356,N_18286,N_18981);
nor U19357 (N_19357,N_18582,N_18306);
or U19358 (N_19358,N_18964,N_18846);
nor U19359 (N_19359,N_18377,N_18150);
nand U19360 (N_19360,N_18147,N_18371);
nor U19361 (N_19361,N_18654,N_18129);
nor U19362 (N_19362,N_18413,N_18861);
and U19363 (N_19363,N_18991,N_18388);
nand U19364 (N_19364,N_18198,N_18564);
nor U19365 (N_19365,N_18107,N_18807);
xnor U19366 (N_19366,N_18174,N_18307);
xor U19367 (N_19367,N_18049,N_18524);
xor U19368 (N_19368,N_18585,N_18718);
nor U19369 (N_19369,N_18790,N_18515);
nor U19370 (N_19370,N_18789,N_18035);
xnor U19371 (N_19371,N_18830,N_18593);
xor U19372 (N_19372,N_18804,N_18825);
nand U19373 (N_19373,N_18487,N_18835);
or U19374 (N_19374,N_18206,N_18549);
xor U19375 (N_19375,N_18364,N_18415);
xnor U19376 (N_19376,N_18128,N_18025);
nor U19377 (N_19377,N_18442,N_18870);
nand U19378 (N_19378,N_18175,N_18787);
xnor U19379 (N_19379,N_18854,N_18268);
xnor U19380 (N_19380,N_18554,N_18321);
and U19381 (N_19381,N_18531,N_18394);
and U19382 (N_19382,N_18327,N_18889);
and U19383 (N_19383,N_18864,N_18943);
nand U19384 (N_19384,N_18114,N_18527);
and U19385 (N_19385,N_18523,N_18113);
or U19386 (N_19386,N_18974,N_18043);
xor U19387 (N_19387,N_18584,N_18673);
or U19388 (N_19388,N_18525,N_18717);
and U19389 (N_19389,N_18739,N_18214);
or U19390 (N_19390,N_18544,N_18202);
xnor U19391 (N_19391,N_18890,N_18125);
and U19392 (N_19392,N_18871,N_18014);
nor U19393 (N_19393,N_18795,N_18934);
xnor U19394 (N_19394,N_18378,N_18216);
xor U19395 (N_19395,N_18868,N_18396);
or U19396 (N_19396,N_18005,N_18972);
or U19397 (N_19397,N_18621,N_18418);
xor U19398 (N_19398,N_18894,N_18280);
nand U19399 (N_19399,N_18506,N_18284);
nor U19400 (N_19400,N_18521,N_18340);
xor U19401 (N_19401,N_18986,N_18094);
nor U19402 (N_19402,N_18188,N_18360);
nand U19403 (N_19403,N_18682,N_18263);
nor U19404 (N_19404,N_18419,N_18062);
nor U19405 (N_19405,N_18888,N_18300);
xor U19406 (N_19406,N_18730,N_18452);
xnor U19407 (N_19407,N_18741,N_18118);
nor U19408 (N_19408,N_18780,N_18144);
or U19409 (N_19409,N_18560,N_18906);
or U19410 (N_19410,N_18437,N_18123);
and U19411 (N_19411,N_18955,N_18459);
nor U19412 (N_19412,N_18260,N_18027);
nand U19413 (N_19413,N_18008,N_18633);
nor U19414 (N_19414,N_18710,N_18347);
nor U19415 (N_19415,N_18552,N_18927);
nand U19416 (N_19416,N_18999,N_18757);
and U19417 (N_19417,N_18181,N_18859);
nor U19418 (N_19418,N_18504,N_18723);
nand U19419 (N_19419,N_18876,N_18478);
or U19420 (N_19420,N_18802,N_18245);
or U19421 (N_19421,N_18636,N_18667);
or U19422 (N_19422,N_18536,N_18436);
nor U19423 (N_19423,N_18766,N_18383);
and U19424 (N_19424,N_18985,N_18805);
and U19425 (N_19425,N_18423,N_18576);
nor U19426 (N_19426,N_18427,N_18001);
xor U19427 (N_19427,N_18056,N_18343);
nand U19428 (N_19428,N_18112,N_18117);
or U19429 (N_19429,N_18675,N_18586);
nor U19430 (N_19430,N_18102,N_18657);
nand U19431 (N_19431,N_18230,N_18319);
nand U19432 (N_19432,N_18517,N_18090);
nor U19433 (N_19433,N_18920,N_18033);
nand U19434 (N_19434,N_18410,N_18880);
xor U19435 (N_19435,N_18180,N_18454);
nand U19436 (N_19436,N_18479,N_18226);
xor U19437 (N_19437,N_18082,N_18677);
and U19438 (N_19438,N_18074,N_18238);
or U19439 (N_19439,N_18158,N_18788);
or U19440 (N_19440,N_18225,N_18511);
nor U19441 (N_19441,N_18153,N_18543);
or U19442 (N_19442,N_18895,N_18441);
xnor U19443 (N_19443,N_18271,N_18078);
nand U19444 (N_19444,N_18929,N_18761);
xor U19445 (N_19445,N_18121,N_18331);
or U19446 (N_19446,N_18296,N_18367);
and U19447 (N_19447,N_18900,N_18272);
or U19448 (N_19448,N_18244,N_18592);
and U19449 (N_19449,N_18639,N_18839);
and U19450 (N_19450,N_18508,N_18681);
nand U19451 (N_19451,N_18691,N_18939);
xnor U19452 (N_19452,N_18233,N_18037);
xnor U19453 (N_19453,N_18239,N_18541);
nand U19454 (N_19454,N_18352,N_18649);
and U19455 (N_19455,N_18497,N_18355);
nand U19456 (N_19456,N_18597,N_18782);
nor U19457 (N_19457,N_18553,N_18237);
xor U19458 (N_19458,N_18057,N_18822);
and U19459 (N_19459,N_18402,N_18287);
nor U19460 (N_19460,N_18595,N_18773);
or U19461 (N_19461,N_18589,N_18572);
nor U19462 (N_19462,N_18872,N_18116);
xnor U19463 (N_19463,N_18628,N_18975);
nor U19464 (N_19464,N_18171,N_18650);
nor U19465 (N_19465,N_18159,N_18632);
nand U19466 (N_19466,N_18952,N_18178);
and U19467 (N_19467,N_18538,N_18808);
and U19468 (N_19468,N_18471,N_18660);
nor U19469 (N_19469,N_18614,N_18540);
or U19470 (N_19470,N_18059,N_18134);
or U19471 (N_19471,N_18856,N_18869);
xor U19472 (N_19472,N_18501,N_18813);
xor U19473 (N_19473,N_18243,N_18587);
nor U19474 (N_19474,N_18818,N_18277);
nand U19475 (N_19475,N_18797,N_18483);
or U19476 (N_19476,N_18127,N_18706);
nor U19477 (N_19477,N_18687,N_18671);
or U19478 (N_19478,N_18664,N_18618);
and U19479 (N_19479,N_18265,N_18429);
nand U19480 (N_19480,N_18992,N_18599);
xnor U19481 (N_19481,N_18693,N_18474);
nor U19482 (N_19482,N_18961,N_18164);
nor U19483 (N_19483,N_18935,N_18910);
nand U19484 (N_19484,N_18778,N_18837);
xor U19485 (N_19485,N_18124,N_18229);
and U19486 (N_19486,N_18068,N_18064);
nand U19487 (N_19487,N_18883,N_18879);
xnor U19488 (N_19488,N_18318,N_18292);
nor U19489 (N_19489,N_18081,N_18688);
or U19490 (N_19490,N_18448,N_18588);
nor U19491 (N_19491,N_18456,N_18763);
nor U19492 (N_19492,N_18648,N_18451);
and U19493 (N_19493,N_18443,N_18661);
nand U19494 (N_19494,N_18190,N_18403);
xor U19495 (N_19495,N_18348,N_18940);
nand U19496 (N_19496,N_18404,N_18712);
or U19497 (N_19497,N_18169,N_18086);
or U19498 (N_19498,N_18707,N_18398);
xor U19499 (N_19499,N_18877,N_18392);
xor U19500 (N_19500,N_18585,N_18342);
or U19501 (N_19501,N_18442,N_18435);
nor U19502 (N_19502,N_18420,N_18423);
xor U19503 (N_19503,N_18988,N_18378);
or U19504 (N_19504,N_18150,N_18004);
nand U19505 (N_19505,N_18600,N_18813);
and U19506 (N_19506,N_18834,N_18290);
nor U19507 (N_19507,N_18641,N_18703);
nand U19508 (N_19508,N_18646,N_18528);
xnor U19509 (N_19509,N_18761,N_18770);
or U19510 (N_19510,N_18928,N_18237);
nand U19511 (N_19511,N_18070,N_18971);
and U19512 (N_19512,N_18202,N_18955);
nand U19513 (N_19513,N_18369,N_18235);
nand U19514 (N_19514,N_18479,N_18315);
nand U19515 (N_19515,N_18859,N_18741);
and U19516 (N_19516,N_18607,N_18593);
xor U19517 (N_19517,N_18909,N_18872);
xnor U19518 (N_19518,N_18682,N_18560);
or U19519 (N_19519,N_18618,N_18505);
nor U19520 (N_19520,N_18484,N_18509);
xnor U19521 (N_19521,N_18125,N_18202);
or U19522 (N_19522,N_18100,N_18350);
nand U19523 (N_19523,N_18952,N_18265);
or U19524 (N_19524,N_18408,N_18368);
nor U19525 (N_19525,N_18740,N_18294);
and U19526 (N_19526,N_18211,N_18013);
and U19527 (N_19527,N_18788,N_18581);
nand U19528 (N_19528,N_18759,N_18753);
nor U19529 (N_19529,N_18589,N_18910);
xor U19530 (N_19530,N_18324,N_18304);
nand U19531 (N_19531,N_18826,N_18308);
and U19532 (N_19532,N_18545,N_18867);
xnor U19533 (N_19533,N_18981,N_18772);
nor U19534 (N_19534,N_18513,N_18514);
or U19535 (N_19535,N_18179,N_18384);
xor U19536 (N_19536,N_18259,N_18832);
nor U19537 (N_19537,N_18610,N_18936);
nor U19538 (N_19538,N_18183,N_18392);
nand U19539 (N_19539,N_18801,N_18845);
nand U19540 (N_19540,N_18583,N_18934);
and U19541 (N_19541,N_18560,N_18109);
nand U19542 (N_19542,N_18600,N_18710);
nand U19543 (N_19543,N_18887,N_18055);
or U19544 (N_19544,N_18161,N_18913);
and U19545 (N_19545,N_18839,N_18444);
or U19546 (N_19546,N_18836,N_18045);
xnor U19547 (N_19547,N_18688,N_18138);
or U19548 (N_19548,N_18718,N_18715);
nand U19549 (N_19549,N_18136,N_18536);
xor U19550 (N_19550,N_18531,N_18571);
and U19551 (N_19551,N_18591,N_18258);
nor U19552 (N_19552,N_18246,N_18622);
and U19553 (N_19553,N_18285,N_18337);
nand U19554 (N_19554,N_18218,N_18144);
xnor U19555 (N_19555,N_18824,N_18796);
nand U19556 (N_19556,N_18029,N_18260);
and U19557 (N_19557,N_18451,N_18755);
or U19558 (N_19558,N_18212,N_18743);
xor U19559 (N_19559,N_18409,N_18306);
and U19560 (N_19560,N_18770,N_18184);
nand U19561 (N_19561,N_18471,N_18193);
nand U19562 (N_19562,N_18254,N_18489);
or U19563 (N_19563,N_18134,N_18378);
xor U19564 (N_19564,N_18380,N_18502);
nor U19565 (N_19565,N_18441,N_18475);
nand U19566 (N_19566,N_18742,N_18166);
and U19567 (N_19567,N_18016,N_18250);
or U19568 (N_19568,N_18606,N_18960);
xnor U19569 (N_19569,N_18896,N_18035);
nor U19570 (N_19570,N_18352,N_18548);
nor U19571 (N_19571,N_18363,N_18258);
xor U19572 (N_19572,N_18406,N_18283);
xor U19573 (N_19573,N_18460,N_18730);
and U19574 (N_19574,N_18120,N_18879);
nor U19575 (N_19575,N_18088,N_18840);
and U19576 (N_19576,N_18428,N_18940);
or U19577 (N_19577,N_18400,N_18454);
xor U19578 (N_19578,N_18896,N_18915);
and U19579 (N_19579,N_18508,N_18000);
xnor U19580 (N_19580,N_18045,N_18456);
or U19581 (N_19581,N_18488,N_18149);
and U19582 (N_19582,N_18388,N_18171);
nand U19583 (N_19583,N_18791,N_18649);
nand U19584 (N_19584,N_18890,N_18528);
xnor U19585 (N_19585,N_18386,N_18088);
nor U19586 (N_19586,N_18272,N_18885);
xor U19587 (N_19587,N_18505,N_18785);
nand U19588 (N_19588,N_18583,N_18023);
or U19589 (N_19589,N_18835,N_18163);
and U19590 (N_19590,N_18443,N_18874);
or U19591 (N_19591,N_18584,N_18435);
xnor U19592 (N_19592,N_18738,N_18237);
nor U19593 (N_19593,N_18295,N_18628);
or U19594 (N_19594,N_18555,N_18415);
nor U19595 (N_19595,N_18797,N_18916);
and U19596 (N_19596,N_18029,N_18598);
or U19597 (N_19597,N_18149,N_18835);
nand U19598 (N_19598,N_18651,N_18114);
nand U19599 (N_19599,N_18862,N_18417);
or U19600 (N_19600,N_18050,N_18147);
and U19601 (N_19601,N_18025,N_18797);
xnor U19602 (N_19602,N_18850,N_18455);
and U19603 (N_19603,N_18933,N_18660);
or U19604 (N_19604,N_18918,N_18586);
nor U19605 (N_19605,N_18314,N_18845);
and U19606 (N_19606,N_18780,N_18948);
nor U19607 (N_19607,N_18159,N_18542);
or U19608 (N_19608,N_18932,N_18694);
and U19609 (N_19609,N_18396,N_18855);
and U19610 (N_19610,N_18574,N_18889);
nand U19611 (N_19611,N_18398,N_18040);
xor U19612 (N_19612,N_18667,N_18243);
and U19613 (N_19613,N_18356,N_18912);
nor U19614 (N_19614,N_18815,N_18713);
xnor U19615 (N_19615,N_18673,N_18066);
xnor U19616 (N_19616,N_18966,N_18383);
and U19617 (N_19617,N_18327,N_18536);
or U19618 (N_19618,N_18351,N_18919);
nand U19619 (N_19619,N_18866,N_18711);
nand U19620 (N_19620,N_18326,N_18144);
nor U19621 (N_19621,N_18374,N_18352);
nand U19622 (N_19622,N_18017,N_18865);
nor U19623 (N_19623,N_18122,N_18146);
or U19624 (N_19624,N_18795,N_18039);
xnor U19625 (N_19625,N_18936,N_18496);
nor U19626 (N_19626,N_18543,N_18523);
xnor U19627 (N_19627,N_18476,N_18421);
and U19628 (N_19628,N_18412,N_18481);
xnor U19629 (N_19629,N_18267,N_18606);
xnor U19630 (N_19630,N_18548,N_18291);
xor U19631 (N_19631,N_18911,N_18618);
nand U19632 (N_19632,N_18018,N_18189);
and U19633 (N_19633,N_18830,N_18992);
nor U19634 (N_19634,N_18516,N_18018);
or U19635 (N_19635,N_18239,N_18198);
nand U19636 (N_19636,N_18799,N_18939);
nor U19637 (N_19637,N_18460,N_18627);
or U19638 (N_19638,N_18424,N_18222);
nand U19639 (N_19639,N_18127,N_18602);
nor U19640 (N_19640,N_18455,N_18719);
xor U19641 (N_19641,N_18645,N_18697);
or U19642 (N_19642,N_18937,N_18964);
or U19643 (N_19643,N_18296,N_18520);
nand U19644 (N_19644,N_18491,N_18192);
xnor U19645 (N_19645,N_18525,N_18400);
or U19646 (N_19646,N_18907,N_18394);
xor U19647 (N_19647,N_18536,N_18427);
or U19648 (N_19648,N_18731,N_18229);
or U19649 (N_19649,N_18688,N_18579);
nand U19650 (N_19650,N_18144,N_18415);
or U19651 (N_19651,N_18243,N_18846);
or U19652 (N_19652,N_18850,N_18956);
xor U19653 (N_19653,N_18280,N_18547);
nand U19654 (N_19654,N_18822,N_18465);
or U19655 (N_19655,N_18017,N_18686);
or U19656 (N_19656,N_18875,N_18280);
xor U19657 (N_19657,N_18422,N_18429);
nand U19658 (N_19658,N_18843,N_18848);
and U19659 (N_19659,N_18366,N_18520);
or U19660 (N_19660,N_18573,N_18455);
nand U19661 (N_19661,N_18075,N_18915);
and U19662 (N_19662,N_18401,N_18736);
and U19663 (N_19663,N_18028,N_18957);
and U19664 (N_19664,N_18084,N_18069);
xor U19665 (N_19665,N_18893,N_18455);
and U19666 (N_19666,N_18450,N_18687);
nor U19667 (N_19667,N_18309,N_18934);
nand U19668 (N_19668,N_18121,N_18663);
nand U19669 (N_19669,N_18145,N_18959);
and U19670 (N_19670,N_18357,N_18757);
or U19671 (N_19671,N_18857,N_18993);
or U19672 (N_19672,N_18615,N_18043);
nand U19673 (N_19673,N_18394,N_18569);
nor U19674 (N_19674,N_18220,N_18646);
nor U19675 (N_19675,N_18088,N_18868);
xor U19676 (N_19676,N_18555,N_18768);
and U19677 (N_19677,N_18386,N_18613);
nor U19678 (N_19678,N_18744,N_18876);
and U19679 (N_19679,N_18769,N_18866);
nor U19680 (N_19680,N_18533,N_18125);
and U19681 (N_19681,N_18996,N_18660);
nor U19682 (N_19682,N_18032,N_18280);
nand U19683 (N_19683,N_18136,N_18641);
xor U19684 (N_19684,N_18590,N_18808);
nand U19685 (N_19685,N_18937,N_18565);
nand U19686 (N_19686,N_18683,N_18693);
nand U19687 (N_19687,N_18134,N_18582);
and U19688 (N_19688,N_18765,N_18119);
xnor U19689 (N_19689,N_18616,N_18440);
xor U19690 (N_19690,N_18916,N_18298);
xnor U19691 (N_19691,N_18232,N_18806);
and U19692 (N_19692,N_18788,N_18012);
nor U19693 (N_19693,N_18404,N_18321);
nor U19694 (N_19694,N_18664,N_18104);
xor U19695 (N_19695,N_18225,N_18316);
and U19696 (N_19696,N_18799,N_18435);
xnor U19697 (N_19697,N_18361,N_18440);
nand U19698 (N_19698,N_18454,N_18328);
or U19699 (N_19699,N_18798,N_18051);
nor U19700 (N_19700,N_18173,N_18104);
xnor U19701 (N_19701,N_18054,N_18880);
nor U19702 (N_19702,N_18144,N_18762);
nand U19703 (N_19703,N_18342,N_18736);
or U19704 (N_19704,N_18019,N_18291);
xnor U19705 (N_19705,N_18581,N_18648);
nand U19706 (N_19706,N_18922,N_18504);
xnor U19707 (N_19707,N_18890,N_18984);
xor U19708 (N_19708,N_18036,N_18080);
and U19709 (N_19709,N_18759,N_18421);
or U19710 (N_19710,N_18480,N_18910);
nor U19711 (N_19711,N_18003,N_18845);
or U19712 (N_19712,N_18061,N_18675);
or U19713 (N_19713,N_18233,N_18382);
or U19714 (N_19714,N_18812,N_18269);
and U19715 (N_19715,N_18926,N_18030);
xnor U19716 (N_19716,N_18690,N_18583);
and U19717 (N_19717,N_18119,N_18507);
nand U19718 (N_19718,N_18128,N_18057);
nor U19719 (N_19719,N_18046,N_18965);
xor U19720 (N_19720,N_18774,N_18490);
xor U19721 (N_19721,N_18412,N_18315);
xor U19722 (N_19722,N_18220,N_18593);
and U19723 (N_19723,N_18323,N_18097);
nand U19724 (N_19724,N_18400,N_18556);
xor U19725 (N_19725,N_18027,N_18791);
and U19726 (N_19726,N_18317,N_18668);
nor U19727 (N_19727,N_18506,N_18420);
and U19728 (N_19728,N_18850,N_18147);
nor U19729 (N_19729,N_18813,N_18550);
and U19730 (N_19730,N_18278,N_18745);
or U19731 (N_19731,N_18131,N_18386);
xor U19732 (N_19732,N_18749,N_18983);
nand U19733 (N_19733,N_18710,N_18668);
and U19734 (N_19734,N_18639,N_18049);
nand U19735 (N_19735,N_18150,N_18484);
nand U19736 (N_19736,N_18291,N_18320);
or U19737 (N_19737,N_18969,N_18827);
or U19738 (N_19738,N_18011,N_18528);
and U19739 (N_19739,N_18342,N_18313);
nand U19740 (N_19740,N_18707,N_18596);
or U19741 (N_19741,N_18131,N_18658);
xor U19742 (N_19742,N_18722,N_18011);
and U19743 (N_19743,N_18564,N_18353);
nand U19744 (N_19744,N_18032,N_18284);
nand U19745 (N_19745,N_18975,N_18438);
or U19746 (N_19746,N_18324,N_18446);
nand U19747 (N_19747,N_18187,N_18079);
nand U19748 (N_19748,N_18474,N_18467);
or U19749 (N_19749,N_18907,N_18098);
and U19750 (N_19750,N_18480,N_18746);
and U19751 (N_19751,N_18622,N_18816);
xor U19752 (N_19752,N_18284,N_18126);
or U19753 (N_19753,N_18207,N_18203);
nor U19754 (N_19754,N_18342,N_18874);
xnor U19755 (N_19755,N_18110,N_18568);
and U19756 (N_19756,N_18957,N_18148);
xor U19757 (N_19757,N_18326,N_18566);
and U19758 (N_19758,N_18973,N_18427);
and U19759 (N_19759,N_18655,N_18896);
nor U19760 (N_19760,N_18348,N_18284);
xor U19761 (N_19761,N_18044,N_18952);
nor U19762 (N_19762,N_18951,N_18944);
nand U19763 (N_19763,N_18503,N_18613);
or U19764 (N_19764,N_18960,N_18907);
and U19765 (N_19765,N_18928,N_18145);
xor U19766 (N_19766,N_18945,N_18808);
or U19767 (N_19767,N_18011,N_18170);
xnor U19768 (N_19768,N_18892,N_18853);
and U19769 (N_19769,N_18595,N_18092);
nor U19770 (N_19770,N_18488,N_18337);
xor U19771 (N_19771,N_18274,N_18917);
nor U19772 (N_19772,N_18631,N_18453);
or U19773 (N_19773,N_18703,N_18185);
and U19774 (N_19774,N_18288,N_18758);
nor U19775 (N_19775,N_18333,N_18782);
nor U19776 (N_19776,N_18021,N_18098);
or U19777 (N_19777,N_18978,N_18523);
and U19778 (N_19778,N_18293,N_18466);
or U19779 (N_19779,N_18030,N_18325);
xor U19780 (N_19780,N_18157,N_18011);
nand U19781 (N_19781,N_18672,N_18815);
nand U19782 (N_19782,N_18912,N_18110);
nand U19783 (N_19783,N_18983,N_18390);
nand U19784 (N_19784,N_18875,N_18657);
or U19785 (N_19785,N_18975,N_18550);
nand U19786 (N_19786,N_18921,N_18115);
nand U19787 (N_19787,N_18850,N_18944);
nor U19788 (N_19788,N_18265,N_18177);
or U19789 (N_19789,N_18659,N_18649);
xnor U19790 (N_19790,N_18858,N_18277);
nor U19791 (N_19791,N_18252,N_18201);
nor U19792 (N_19792,N_18665,N_18343);
nand U19793 (N_19793,N_18945,N_18190);
nor U19794 (N_19794,N_18157,N_18417);
nor U19795 (N_19795,N_18333,N_18116);
and U19796 (N_19796,N_18531,N_18936);
nor U19797 (N_19797,N_18235,N_18491);
or U19798 (N_19798,N_18546,N_18470);
nand U19799 (N_19799,N_18658,N_18285);
and U19800 (N_19800,N_18166,N_18045);
xnor U19801 (N_19801,N_18105,N_18944);
or U19802 (N_19802,N_18125,N_18208);
nand U19803 (N_19803,N_18865,N_18718);
nand U19804 (N_19804,N_18548,N_18141);
nor U19805 (N_19805,N_18575,N_18872);
or U19806 (N_19806,N_18612,N_18497);
nor U19807 (N_19807,N_18636,N_18927);
nor U19808 (N_19808,N_18043,N_18198);
nand U19809 (N_19809,N_18206,N_18246);
or U19810 (N_19810,N_18431,N_18759);
nand U19811 (N_19811,N_18113,N_18830);
or U19812 (N_19812,N_18030,N_18997);
nor U19813 (N_19813,N_18692,N_18426);
xor U19814 (N_19814,N_18358,N_18477);
and U19815 (N_19815,N_18569,N_18230);
nand U19816 (N_19816,N_18454,N_18634);
nand U19817 (N_19817,N_18016,N_18127);
nand U19818 (N_19818,N_18831,N_18167);
and U19819 (N_19819,N_18214,N_18288);
or U19820 (N_19820,N_18661,N_18604);
and U19821 (N_19821,N_18508,N_18033);
nor U19822 (N_19822,N_18258,N_18282);
or U19823 (N_19823,N_18591,N_18589);
nand U19824 (N_19824,N_18047,N_18164);
xor U19825 (N_19825,N_18922,N_18750);
or U19826 (N_19826,N_18302,N_18350);
nand U19827 (N_19827,N_18809,N_18449);
xnor U19828 (N_19828,N_18037,N_18882);
xnor U19829 (N_19829,N_18357,N_18217);
xnor U19830 (N_19830,N_18882,N_18451);
or U19831 (N_19831,N_18982,N_18633);
nor U19832 (N_19832,N_18232,N_18654);
nand U19833 (N_19833,N_18425,N_18056);
and U19834 (N_19834,N_18979,N_18874);
or U19835 (N_19835,N_18869,N_18094);
nor U19836 (N_19836,N_18573,N_18020);
xnor U19837 (N_19837,N_18083,N_18446);
nor U19838 (N_19838,N_18802,N_18764);
or U19839 (N_19839,N_18891,N_18883);
and U19840 (N_19840,N_18171,N_18353);
or U19841 (N_19841,N_18385,N_18503);
or U19842 (N_19842,N_18132,N_18380);
and U19843 (N_19843,N_18411,N_18904);
xor U19844 (N_19844,N_18691,N_18025);
nor U19845 (N_19845,N_18025,N_18226);
xnor U19846 (N_19846,N_18978,N_18620);
nor U19847 (N_19847,N_18929,N_18132);
or U19848 (N_19848,N_18875,N_18357);
or U19849 (N_19849,N_18112,N_18377);
xnor U19850 (N_19850,N_18749,N_18909);
xor U19851 (N_19851,N_18676,N_18539);
or U19852 (N_19852,N_18633,N_18142);
nand U19853 (N_19853,N_18355,N_18658);
nand U19854 (N_19854,N_18748,N_18835);
or U19855 (N_19855,N_18418,N_18466);
nand U19856 (N_19856,N_18959,N_18143);
and U19857 (N_19857,N_18652,N_18307);
and U19858 (N_19858,N_18306,N_18038);
xnor U19859 (N_19859,N_18837,N_18802);
nand U19860 (N_19860,N_18026,N_18913);
and U19861 (N_19861,N_18847,N_18816);
nor U19862 (N_19862,N_18812,N_18183);
nand U19863 (N_19863,N_18047,N_18801);
xor U19864 (N_19864,N_18280,N_18698);
or U19865 (N_19865,N_18736,N_18945);
or U19866 (N_19866,N_18444,N_18325);
and U19867 (N_19867,N_18073,N_18582);
nand U19868 (N_19868,N_18209,N_18043);
and U19869 (N_19869,N_18480,N_18246);
or U19870 (N_19870,N_18947,N_18694);
and U19871 (N_19871,N_18136,N_18935);
and U19872 (N_19872,N_18603,N_18748);
nand U19873 (N_19873,N_18444,N_18724);
nor U19874 (N_19874,N_18285,N_18597);
or U19875 (N_19875,N_18156,N_18781);
nand U19876 (N_19876,N_18113,N_18390);
nor U19877 (N_19877,N_18631,N_18004);
xnor U19878 (N_19878,N_18457,N_18655);
and U19879 (N_19879,N_18063,N_18506);
xor U19880 (N_19880,N_18658,N_18334);
xor U19881 (N_19881,N_18582,N_18659);
nand U19882 (N_19882,N_18111,N_18872);
or U19883 (N_19883,N_18947,N_18910);
or U19884 (N_19884,N_18553,N_18848);
nor U19885 (N_19885,N_18239,N_18571);
nor U19886 (N_19886,N_18003,N_18599);
or U19887 (N_19887,N_18195,N_18576);
or U19888 (N_19888,N_18136,N_18372);
xor U19889 (N_19889,N_18228,N_18950);
nand U19890 (N_19890,N_18572,N_18363);
nor U19891 (N_19891,N_18315,N_18586);
nor U19892 (N_19892,N_18209,N_18689);
nor U19893 (N_19893,N_18464,N_18449);
nand U19894 (N_19894,N_18664,N_18951);
nand U19895 (N_19895,N_18996,N_18436);
and U19896 (N_19896,N_18641,N_18343);
or U19897 (N_19897,N_18885,N_18061);
nor U19898 (N_19898,N_18124,N_18890);
xor U19899 (N_19899,N_18514,N_18847);
xnor U19900 (N_19900,N_18523,N_18609);
or U19901 (N_19901,N_18101,N_18186);
xnor U19902 (N_19902,N_18657,N_18939);
xor U19903 (N_19903,N_18091,N_18191);
or U19904 (N_19904,N_18831,N_18088);
nand U19905 (N_19905,N_18494,N_18882);
xnor U19906 (N_19906,N_18092,N_18640);
or U19907 (N_19907,N_18345,N_18825);
or U19908 (N_19908,N_18572,N_18209);
xor U19909 (N_19909,N_18134,N_18597);
and U19910 (N_19910,N_18478,N_18506);
nor U19911 (N_19911,N_18532,N_18465);
and U19912 (N_19912,N_18531,N_18069);
nand U19913 (N_19913,N_18617,N_18975);
nor U19914 (N_19914,N_18984,N_18865);
nand U19915 (N_19915,N_18219,N_18957);
xor U19916 (N_19916,N_18130,N_18516);
or U19917 (N_19917,N_18025,N_18638);
nand U19918 (N_19918,N_18289,N_18566);
nor U19919 (N_19919,N_18168,N_18338);
xnor U19920 (N_19920,N_18974,N_18373);
nor U19921 (N_19921,N_18206,N_18929);
or U19922 (N_19922,N_18275,N_18483);
and U19923 (N_19923,N_18984,N_18794);
and U19924 (N_19924,N_18502,N_18779);
or U19925 (N_19925,N_18553,N_18813);
or U19926 (N_19926,N_18486,N_18231);
nor U19927 (N_19927,N_18263,N_18867);
xor U19928 (N_19928,N_18159,N_18605);
and U19929 (N_19929,N_18966,N_18105);
and U19930 (N_19930,N_18192,N_18840);
or U19931 (N_19931,N_18695,N_18160);
xor U19932 (N_19932,N_18893,N_18862);
xor U19933 (N_19933,N_18441,N_18523);
xor U19934 (N_19934,N_18156,N_18749);
nand U19935 (N_19935,N_18954,N_18325);
nand U19936 (N_19936,N_18574,N_18379);
and U19937 (N_19937,N_18046,N_18553);
xnor U19938 (N_19938,N_18545,N_18059);
xor U19939 (N_19939,N_18853,N_18049);
nand U19940 (N_19940,N_18887,N_18545);
nor U19941 (N_19941,N_18764,N_18029);
or U19942 (N_19942,N_18318,N_18495);
nand U19943 (N_19943,N_18374,N_18858);
or U19944 (N_19944,N_18221,N_18462);
nand U19945 (N_19945,N_18094,N_18991);
nor U19946 (N_19946,N_18119,N_18133);
nor U19947 (N_19947,N_18366,N_18646);
nor U19948 (N_19948,N_18956,N_18503);
nand U19949 (N_19949,N_18618,N_18051);
nand U19950 (N_19950,N_18474,N_18566);
and U19951 (N_19951,N_18266,N_18666);
xor U19952 (N_19952,N_18815,N_18527);
nand U19953 (N_19953,N_18204,N_18940);
or U19954 (N_19954,N_18462,N_18510);
and U19955 (N_19955,N_18926,N_18203);
or U19956 (N_19956,N_18838,N_18452);
nand U19957 (N_19957,N_18469,N_18388);
and U19958 (N_19958,N_18492,N_18856);
or U19959 (N_19959,N_18741,N_18013);
and U19960 (N_19960,N_18848,N_18325);
and U19961 (N_19961,N_18680,N_18192);
and U19962 (N_19962,N_18365,N_18482);
xnor U19963 (N_19963,N_18146,N_18530);
xor U19964 (N_19964,N_18822,N_18027);
nand U19965 (N_19965,N_18561,N_18046);
and U19966 (N_19966,N_18615,N_18032);
nand U19967 (N_19967,N_18198,N_18263);
xor U19968 (N_19968,N_18484,N_18352);
or U19969 (N_19969,N_18813,N_18045);
or U19970 (N_19970,N_18508,N_18802);
or U19971 (N_19971,N_18025,N_18237);
and U19972 (N_19972,N_18485,N_18362);
xor U19973 (N_19973,N_18629,N_18894);
xor U19974 (N_19974,N_18710,N_18103);
xor U19975 (N_19975,N_18471,N_18815);
nor U19976 (N_19976,N_18308,N_18720);
and U19977 (N_19977,N_18391,N_18379);
or U19978 (N_19978,N_18981,N_18328);
or U19979 (N_19979,N_18376,N_18940);
and U19980 (N_19980,N_18567,N_18058);
or U19981 (N_19981,N_18860,N_18172);
xor U19982 (N_19982,N_18762,N_18915);
nand U19983 (N_19983,N_18433,N_18332);
and U19984 (N_19984,N_18716,N_18413);
nand U19985 (N_19985,N_18345,N_18511);
xnor U19986 (N_19986,N_18942,N_18028);
and U19987 (N_19987,N_18113,N_18697);
nor U19988 (N_19988,N_18084,N_18090);
or U19989 (N_19989,N_18515,N_18020);
and U19990 (N_19990,N_18611,N_18968);
or U19991 (N_19991,N_18079,N_18436);
nand U19992 (N_19992,N_18489,N_18385);
nand U19993 (N_19993,N_18652,N_18588);
nor U19994 (N_19994,N_18341,N_18752);
or U19995 (N_19995,N_18807,N_18922);
nor U19996 (N_19996,N_18953,N_18238);
and U19997 (N_19997,N_18945,N_18637);
nor U19998 (N_19998,N_18422,N_18570);
nand U19999 (N_19999,N_18851,N_18899);
nand U20000 (N_20000,N_19154,N_19414);
and U20001 (N_20001,N_19254,N_19468);
nand U20002 (N_20002,N_19309,N_19239);
or U20003 (N_20003,N_19068,N_19578);
or U20004 (N_20004,N_19881,N_19998);
nand U20005 (N_20005,N_19766,N_19838);
nor U20006 (N_20006,N_19776,N_19315);
xnor U20007 (N_20007,N_19408,N_19509);
nand U20008 (N_20008,N_19188,N_19111);
nand U20009 (N_20009,N_19301,N_19859);
xor U20010 (N_20010,N_19931,N_19382);
and U20011 (N_20011,N_19769,N_19522);
and U20012 (N_20012,N_19010,N_19991);
and U20013 (N_20013,N_19675,N_19950);
nor U20014 (N_20014,N_19302,N_19822);
nand U20015 (N_20015,N_19780,N_19595);
and U20016 (N_20016,N_19586,N_19189);
and U20017 (N_20017,N_19872,N_19243);
nor U20018 (N_20018,N_19056,N_19972);
xnor U20019 (N_20019,N_19582,N_19963);
and U20020 (N_20020,N_19303,N_19373);
or U20021 (N_20021,N_19794,N_19916);
nand U20022 (N_20022,N_19561,N_19423);
or U20023 (N_20023,N_19037,N_19692);
nor U20024 (N_20024,N_19957,N_19014);
nor U20025 (N_20025,N_19394,N_19133);
and U20026 (N_20026,N_19678,N_19238);
xor U20027 (N_20027,N_19223,N_19273);
and U20028 (N_20028,N_19244,N_19287);
xnor U20029 (N_20029,N_19230,N_19554);
or U20030 (N_20030,N_19547,N_19869);
xor U20031 (N_20031,N_19713,N_19300);
and U20032 (N_20032,N_19528,N_19719);
or U20033 (N_20033,N_19623,N_19220);
xor U20034 (N_20034,N_19562,N_19613);
xor U20035 (N_20035,N_19319,N_19824);
nor U20036 (N_20036,N_19217,N_19514);
or U20037 (N_20037,N_19695,N_19874);
xor U20038 (N_20038,N_19158,N_19674);
nor U20039 (N_20039,N_19877,N_19240);
nand U20040 (N_20040,N_19176,N_19521);
nand U20041 (N_20041,N_19927,N_19344);
or U20042 (N_20042,N_19529,N_19199);
nand U20043 (N_20043,N_19702,N_19140);
nor U20044 (N_20044,N_19117,N_19572);
nor U20045 (N_20045,N_19345,N_19211);
and U20046 (N_20046,N_19632,N_19180);
xor U20047 (N_20047,N_19648,N_19918);
or U20048 (N_20048,N_19857,N_19323);
or U20049 (N_20049,N_19488,N_19668);
nand U20050 (N_20050,N_19749,N_19608);
nand U20051 (N_20051,N_19272,N_19215);
and U20052 (N_20052,N_19296,N_19544);
nor U20053 (N_20053,N_19427,N_19185);
or U20054 (N_20054,N_19486,N_19086);
xor U20055 (N_20055,N_19641,N_19246);
xnor U20056 (N_20056,N_19019,N_19042);
nor U20057 (N_20057,N_19842,N_19059);
xor U20058 (N_20058,N_19393,N_19699);
xnor U20059 (N_20059,N_19729,N_19625);
nand U20060 (N_20060,N_19288,N_19966);
nand U20061 (N_20061,N_19754,N_19866);
and U20062 (N_20062,N_19809,N_19581);
and U20063 (N_20063,N_19232,N_19577);
nand U20064 (N_20064,N_19829,N_19525);
nand U20065 (N_20065,N_19849,N_19642);
xnor U20066 (N_20066,N_19862,N_19790);
or U20067 (N_20067,N_19880,N_19186);
nor U20068 (N_20068,N_19083,N_19763);
nand U20069 (N_20069,N_19173,N_19707);
nand U20070 (N_20070,N_19747,N_19367);
or U20071 (N_20071,N_19314,N_19353);
and U20072 (N_20072,N_19843,N_19928);
nand U20073 (N_20073,N_19257,N_19597);
nor U20074 (N_20074,N_19316,N_19920);
xor U20075 (N_20075,N_19654,N_19557);
and U20076 (N_20076,N_19429,N_19099);
nor U20077 (N_20077,N_19580,N_19762);
nor U20078 (N_20078,N_19310,N_19725);
nand U20079 (N_20079,N_19819,N_19341);
and U20080 (N_20080,N_19233,N_19500);
or U20081 (N_20081,N_19934,N_19018);
nand U20082 (N_20082,N_19566,N_19498);
or U20083 (N_20083,N_19221,N_19552);
nor U20084 (N_20084,N_19941,N_19493);
xnor U20085 (N_20085,N_19046,N_19385);
xor U20086 (N_20086,N_19801,N_19386);
nand U20087 (N_20087,N_19737,N_19067);
or U20088 (N_20088,N_19646,N_19813);
xnor U20089 (N_20089,N_19171,N_19962);
and U20090 (N_20090,N_19779,N_19938);
nand U20091 (N_20091,N_19636,N_19555);
and U20092 (N_20092,N_19628,N_19282);
nor U20093 (N_20093,N_19279,N_19759);
and U20094 (N_20094,N_19698,N_19893);
nor U20095 (N_20095,N_19292,N_19760);
nor U20096 (N_20096,N_19494,N_19569);
xnor U20097 (N_20097,N_19376,N_19953);
xnor U20098 (N_20098,N_19935,N_19103);
nand U20099 (N_20099,N_19085,N_19601);
nand U20100 (N_20100,N_19850,N_19480);
xnor U20101 (N_20101,N_19281,N_19722);
or U20102 (N_20102,N_19216,N_19976);
nor U20103 (N_20103,N_19756,N_19047);
and U20104 (N_20104,N_19491,N_19207);
xnor U20105 (N_20105,N_19676,N_19050);
nand U20106 (N_20106,N_19734,N_19073);
nor U20107 (N_20107,N_19327,N_19040);
nand U20108 (N_20108,N_19968,N_19691);
xnor U20109 (N_20109,N_19411,N_19637);
xor U20110 (N_20110,N_19999,N_19477);
xor U20111 (N_20111,N_19510,N_19959);
nand U20112 (N_20112,N_19121,N_19481);
nand U20113 (N_20113,N_19131,N_19432);
nor U20114 (N_20114,N_19590,N_19655);
or U20115 (N_20115,N_19157,N_19504);
or U20116 (N_20116,N_19114,N_19129);
and U20117 (N_20117,N_19271,N_19030);
xor U20118 (N_20118,N_19191,N_19816);
nand U20119 (N_20119,N_19192,N_19716);
nand U20120 (N_20120,N_19396,N_19090);
or U20121 (N_20121,N_19937,N_19008);
nand U20122 (N_20122,N_19553,N_19791);
and U20123 (N_20123,N_19029,N_19075);
nor U20124 (N_20124,N_19727,N_19783);
xnor U20125 (N_20125,N_19600,N_19952);
nand U20126 (N_20126,N_19563,N_19820);
or U20127 (N_20127,N_19827,N_19084);
nand U20128 (N_20128,N_19908,N_19712);
xor U20129 (N_20129,N_19418,N_19096);
nor U20130 (N_20130,N_19583,N_19492);
nand U20131 (N_20131,N_19017,N_19197);
or U20132 (N_20132,N_19592,N_19457);
xor U20133 (N_20133,N_19259,N_19139);
and U20134 (N_20134,N_19253,N_19422);
xnor U20135 (N_20135,N_19120,N_19036);
xor U20136 (N_20136,N_19177,N_19377);
nand U20137 (N_20137,N_19439,N_19770);
nand U20138 (N_20138,N_19359,N_19960);
or U20139 (N_20139,N_19093,N_19921);
xnor U20140 (N_20140,N_19907,N_19440);
and U20141 (N_20141,N_19404,N_19144);
xor U20142 (N_20142,N_19902,N_19889);
xnor U20143 (N_20143,N_19104,N_19946);
nor U20144 (N_20144,N_19992,N_19571);
xor U20145 (N_20145,N_19389,N_19058);
and U20146 (N_20146,N_19564,N_19967);
and U20147 (N_20147,N_19003,N_19265);
or U20148 (N_20148,N_19996,N_19403);
and U20149 (N_20149,N_19318,N_19064);
or U20150 (N_20150,N_19011,N_19392);
or U20151 (N_20151,N_19679,N_19627);
xnor U20152 (N_20152,N_19884,N_19169);
nor U20153 (N_20153,N_19735,N_19844);
or U20154 (N_20154,N_19665,N_19026);
nand U20155 (N_20155,N_19610,N_19693);
xnor U20156 (N_20156,N_19619,N_19971);
xnor U20157 (N_20157,N_19497,N_19080);
xor U20158 (N_20158,N_19081,N_19306);
and U20159 (N_20159,N_19800,N_19645);
and U20160 (N_20160,N_19771,N_19823);
and U20161 (N_20161,N_19669,N_19043);
nand U20162 (N_20162,N_19644,N_19974);
or U20163 (N_20163,N_19774,N_19864);
xnor U20164 (N_20164,N_19052,N_19746);
nor U20165 (N_20165,N_19087,N_19156);
nor U20166 (N_20166,N_19295,N_19406);
nor U20167 (N_20167,N_19615,N_19773);
and U20168 (N_20168,N_19540,N_19179);
and U20169 (N_20169,N_19175,N_19170);
or U20170 (N_20170,N_19245,N_19242);
or U20171 (N_20171,N_19039,N_19055);
xnor U20172 (N_20172,N_19092,N_19095);
nand U20173 (N_20173,N_19778,N_19706);
nor U20174 (N_20174,N_19975,N_19425);
xor U20175 (N_20175,N_19984,N_19347);
xnor U20176 (N_20176,N_19442,N_19714);
nor U20177 (N_20177,N_19621,N_19127);
nand U20178 (N_20178,N_19351,N_19049);
and U20179 (N_20179,N_19155,N_19740);
nor U20180 (N_20180,N_19202,N_19579);
nand U20181 (N_20181,N_19153,N_19689);
and U20182 (N_20182,N_19431,N_19006);
xor U20183 (N_20183,N_19333,N_19079);
and U20184 (N_20184,N_19210,N_19062);
or U20185 (N_20185,N_19659,N_19501);
nand U20186 (N_20186,N_19417,N_19410);
xnor U20187 (N_20187,N_19035,N_19730);
xnor U20188 (N_20188,N_19428,N_19275);
and U20189 (N_20189,N_19970,N_19409);
xor U20190 (N_20190,N_19704,N_19291);
nor U20191 (N_20191,N_19321,N_19513);
nor U20192 (N_20192,N_19383,N_19784);
xnor U20193 (N_20193,N_19936,N_19366);
nor U20194 (N_20194,N_19728,N_19053);
nand U20195 (N_20195,N_19997,N_19841);
nor U20196 (N_20196,N_19524,N_19939);
nand U20197 (N_20197,N_19196,N_19463);
xor U20198 (N_20198,N_19370,N_19435);
xnor U20199 (N_20199,N_19867,N_19584);
nor U20200 (N_20200,N_19368,N_19201);
or U20201 (N_20201,N_19982,N_19596);
nor U20202 (N_20202,N_19923,N_19551);
or U20203 (N_20203,N_19206,N_19005);
and U20204 (N_20204,N_19150,N_19865);
xnor U20205 (N_20205,N_19748,N_19395);
or U20206 (N_20206,N_19940,N_19467);
and U20207 (N_20207,N_19890,N_19237);
xor U20208 (N_20208,N_19136,N_19828);
xor U20209 (N_20209,N_19187,N_19038);
xor U20210 (N_20210,N_19836,N_19671);
or U20211 (N_20211,N_19720,N_19012);
nand U20212 (N_20212,N_19799,N_19231);
or U20213 (N_20213,N_19147,N_19878);
or U20214 (N_20214,N_19349,N_19797);
nand U20215 (N_20215,N_19885,N_19482);
nor U20216 (N_20216,N_19032,N_19961);
or U20217 (N_20217,N_19496,N_19919);
xor U20218 (N_20218,N_19328,N_19560);
nor U20219 (N_20219,N_19276,N_19299);
xor U20220 (N_20220,N_19834,N_19015);
nor U20221 (N_20221,N_19786,N_19002);
nor U20222 (N_20222,N_19362,N_19110);
nand U20223 (N_20223,N_19490,N_19887);
nand U20224 (N_20224,N_19516,N_19335);
nand U20225 (N_20225,N_19757,N_19883);
and U20226 (N_20226,N_19682,N_19915);
nand U20227 (N_20227,N_19474,N_19174);
and U20228 (N_20228,N_19777,N_19643);
and U20229 (N_20229,N_19806,N_19218);
nand U20230 (N_20230,N_19534,N_19565);
nor U20231 (N_20231,N_19891,N_19313);
nor U20232 (N_20232,N_19744,N_19280);
xnor U20233 (N_20233,N_19751,N_19639);
and U20234 (N_20234,N_19726,N_19863);
xnor U20235 (N_20235,N_19476,N_19649);
and U20236 (N_20236,N_19954,N_19585);
xor U20237 (N_20237,N_19687,N_19629);
xor U20238 (N_20238,N_19266,N_19614);
nor U20239 (N_20239,N_19985,N_19663);
nor U20240 (N_20240,N_19401,N_19441);
xor U20241 (N_20241,N_19159,N_19402);
xnor U20242 (N_20242,N_19262,N_19261);
or U20243 (N_20243,N_19978,N_19149);
xnor U20244 (N_20244,N_19145,N_19804);
nand U20245 (N_20245,N_19124,N_19882);
nand U20246 (N_20246,N_19944,N_19853);
xnor U20247 (N_20247,N_19361,N_19696);
nand U20248 (N_20248,N_19826,N_19694);
or U20249 (N_20249,N_19214,N_19478);
nor U20250 (N_20250,N_19647,N_19977);
and U20251 (N_20251,N_19115,N_19100);
xnor U20252 (N_20252,N_19473,N_19788);
or U20253 (N_20253,N_19852,N_19503);
or U20254 (N_20254,N_19447,N_19371);
and U20255 (N_20255,N_19567,N_19453);
nand U20256 (N_20256,N_19297,N_19098);
and U20257 (N_20257,N_19624,N_19166);
and U20258 (N_20258,N_19742,N_19988);
nor U20259 (N_20259,N_19004,N_19876);
xnor U20260 (N_20260,N_19250,N_19072);
and U20261 (N_20261,N_19690,N_19357);
nor U20262 (N_20262,N_19130,N_19556);
or U20263 (N_20263,N_19445,N_19286);
nand U20264 (N_20264,N_19023,N_19617);
nor U20265 (N_20265,N_19559,N_19143);
xnor U20266 (N_20266,N_19113,N_19071);
nand U20267 (N_20267,N_19616,N_19116);
nand U20268 (N_20268,N_19449,N_19465);
nand U20269 (N_20269,N_19810,N_19903);
and U20270 (N_20270,N_19917,N_19650);
or U20271 (N_20271,N_19451,N_19020);
and U20272 (N_20272,N_19336,N_19229);
and U20273 (N_20273,N_19724,N_19125);
nand U20274 (N_20274,N_19994,N_19929);
xnor U20275 (N_20275,N_19270,N_19993);
nand U20276 (N_20276,N_19350,N_19733);
nor U20277 (N_20277,N_19673,N_19094);
nor U20278 (N_20278,N_19677,N_19811);
and U20279 (N_20279,N_19980,N_19956);
xor U20280 (N_20280,N_19979,N_19343);
nor U20281 (N_20281,N_19594,N_19717);
nand U20282 (N_20282,N_19886,N_19833);
or U20283 (N_20283,N_19308,N_19048);
xnor U20284 (N_20284,N_19798,N_19205);
and U20285 (N_20285,N_19485,N_19575);
or U20286 (N_20286,N_19054,N_19045);
and U20287 (N_20287,N_19651,N_19711);
nand U20288 (N_20288,N_19190,N_19587);
and U20289 (N_20289,N_19815,N_19424);
xor U20290 (N_20290,N_19028,N_19164);
nand U20291 (N_20291,N_19892,N_19543);
or U20292 (N_20292,N_19787,N_19024);
xor U20293 (N_20293,N_19860,N_19546);
nand U20294 (N_20294,N_19375,N_19443);
or U20295 (N_20295,N_19986,N_19945);
nand U20296 (N_20296,N_19142,N_19568);
xor U20297 (N_20297,N_19895,N_19334);
xnor U20298 (N_20298,N_19235,N_19227);
or U20299 (N_20299,N_19989,N_19470);
nand U20300 (N_20300,N_19298,N_19458);
nand U20301 (N_20301,N_19203,N_19549);
xnor U20302 (N_20302,N_19352,N_19835);
xnor U20303 (N_20303,N_19538,N_19965);
nor U20304 (N_20304,N_19796,N_19123);
or U20305 (N_20305,N_19000,N_19576);
and U20306 (N_20306,N_19499,N_19495);
xnor U20307 (N_20307,N_19413,N_19364);
xnor U20308 (N_20308,N_19195,N_19452);
and U20309 (N_20309,N_19700,N_19021);
nor U20310 (N_20310,N_19948,N_19660);
or U20311 (N_20311,N_19795,N_19515);
or U20312 (N_20312,N_19633,N_19102);
nor U20313 (N_20313,N_19412,N_19317);
or U20314 (N_20314,N_19661,N_19511);
xnor U20315 (N_20315,N_19620,N_19926);
xor U20316 (N_20316,N_19340,N_19708);
xnor U20317 (N_20317,N_19063,N_19263);
and U20318 (N_20318,N_19471,N_19162);
or U20319 (N_20319,N_19911,N_19082);
or U20320 (N_20320,N_19839,N_19074);
and U20321 (N_20321,N_19635,N_19922);
and U20322 (N_20322,N_19964,N_19854);
or U20323 (N_20323,N_19830,N_19683);
xnor U20324 (N_20324,N_19378,N_19430);
or U20325 (N_20325,N_19475,N_19066);
nand U20326 (N_20326,N_19523,N_19208);
and U20327 (N_20327,N_19752,N_19894);
nand U20328 (N_20328,N_19775,N_19840);
nand U20329 (N_20329,N_19598,N_19924);
nand U20330 (N_20330,N_19051,N_19723);
xor U20331 (N_20331,N_19322,N_19606);
nand U20332 (N_20332,N_19466,N_19033);
or U20333 (N_20333,N_19535,N_19420);
or U20334 (N_20334,N_19767,N_19384);
nor U20335 (N_20335,N_19252,N_19832);
or U20336 (N_20336,N_19812,N_19947);
or U20337 (N_20337,N_19932,N_19871);
nand U20338 (N_20338,N_19851,N_19264);
nand U20339 (N_20339,N_19731,N_19355);
or U20340 (N_20340,N_19548,N_19027);
nand U20341 (N_20341,N_19198,N_19137);
nand U20342 (N_20342,N_19520,N_19070);
nor U20343 (N_20343,N_19900,N_19405);
nor U20344 (N_20344,N_19283,N_19888);
xor U20345 (N_20345,N_19837,N_19387);
nand U20346 (N_20346,N_19326,N_19348);
nand U20347 (N_20347,N_19680,N_19667);
xor U20348 (N_20348,N_19653,N_19284);
and U20349 (N_20349,N_19134,N_19101);
xor U20350 (N_20350,N_19141,N_19305);
nand U20351 (N_20351,N_19391,N_19304);
nand U20352 (N_20352,N_19901,N_19703);
nor U20353 (N_20353,N_19255,N_19460);
xor U20354 (N_20354,N_19446,N_19438);
nand U20355 (N_20355,N_19588,N_19570);
and U20356 (N_20356,N_19664,N_19289);
nand U20357 (N_20357,N_19789,N_19705);
nand U20358 (N_20358,N_19455,N_19541);
nor U20359 (N_20359,N_19507,N_19818);
nor U20360 (N_20360,N_19505,N_19331);
nand U20361 (N_20361,N_19533,N_19831);
nand U20362 (N_20362,N_19126,N_19802);
nand U20363 (N_20363,N_19224,N_19433);
xor U20364 (N_20364,N_19656,N_19905);
or U20365 (N_20365,N_19715,N_19290);
and U20366 (N_20366,N_19013,N_19088);
and U20367 (N_20367,N_19226,N_19861);
and U20368 (N_20368,N_19407,N_19904);
nand U20369 (N_20369,N_19181,N_19397);
or U20370 (N_20370,N_19077,N_19573);
nand U20371 (N_20371,N_19057,N_19163);
nand U20372 (N_20372,N_19128,N_19631);
and U20373 (N_20373,N_19419,N_19256);
nand U20374 (N_20374,N_19845,N_19324);
nand U20375 (N_20375,N_19542,N_19607);
or U20376 (N_20376,N_19078,N_19846);
or U20377 (N_20377,N_19269,N_19897);
nand U20378 (N_20378,N_19372,N_19400);
or U20379 (N_20379,N_19739,N_19898);
and U20380 (N_20380,N_19416,N_19109);
xor U20381 (N_20381,N_19168,N_19479);
nand U20382 (N_20382,N_19545,N_19450);
nor U20383 (N_20383,N_19951,N_19868);
and U20384 (N_20384,N_19518,N_19219);
nand U20385 (N_20385,N_19076,N_19686);
nand U20386 (N_20386,N_19765,N_19112);
nand U20387 (N_20387,N_19670,N_19914);
or U20388 (N_20388,N_19681,N_19634);
nor U20389 (N_20389,N_19856,N_19360);
nand U20390 (N_20390,N_19151,N_19436);
nand U20391 (N_20391,N_19750,N_19987);
or U20392 (N_20392,N_19658,N_19574);
nand U20393 (N_20393,N_19380,N_19990);
nor U20394 (N_20394,N_19278,N_19148);
nor U20395 (N_20395,N_19178,N_19146);
xnor U20396 (N_20396,N_19605,N_19875);
and U20397 (N_20397,N_19374,N_19462);
or U20398 (N_20398,N_19065,N_19906);
nand U20399 (N_20399,N_19817,N_19709);
or U20400 (N_20400,N_19983,N_19484);
nand U20401 (N_20401,N_19307,N_19294);
and U20402 (N_20402,N_19710,N_19459);
or U20403 (N_20403,N_19517,N_19933);
nand U20404 (N_20404,N_19225,N_19666);
xor U20405 (N_20405,N_19356,N_19388);
nor U20406 (N_20406,N_19167,N_19685);
or U20407 (N_20407,N_19069,N_19558);
nand U20408 (N_20408,N_19909,N_19132);
xnor U20409 (N_20409,N_19122,N_19949);
xnor U20410 (N_20410,N_19955,N_19506);
xnor U20411 (N_20411,N_19593,N_19236);
or U20412 (N_20412,N_19193,N_19325);
nor U20413 (N_20413,N_19358,N_19119);
and U20414 (N_20414,N_19089,N_19138);
nor U20415 (N_20415,N_19009,N_19622);
and U20416 (N_20416,N_19807,N_19461);
xnor U20417 (N_20417,N_19061,N_19415);
and U20418 (N_20418,N_19204,N_19808);
or U20419 (N_20419,N_19531,N_19022);
or U20420 (N_20420,N_19684,N_19031);
xnor U20421 (N_20421,N_19354,N_19662);
and U20422 (N_20422,N_19489,N_19539);
or U20423 (N_20423,N_19638,N_19161);
and U20424 (N_20424,N_19738,N_19320);
nand U20425 (N_20425,N_19258,N_19034);
xnor U20426 (N_20426,N_19526,N_19721);
xor U20427 (N_20427,N_19234,N_19532);
nand U20428 (N_20428,N_19483,N_19814);
or U20429 (N_20429,N_19041,N_19228);
xor U20430 (N_20430,N_19172,N_19925);
xnor U20431 (N_20431,N_19611,N_19339);
nand U20432 (N_20432,N_19285,N_19332);
xnor U20433 (N_20433,N_19761,N_19688);
nand U20434 (N_20434,N_19603,N_19741);
nor U20435 (N_20435,N_19312,N_19626);
nand U20436 (N_20436,N_19589,N_19672);
nand U20437 (N_20437,N_19274,N_19222);
or U20438 (N_20438,N_19848,N_19247);
and U20439 (N_20439,N_19912,N_19241);
xnor U20440 (N_20440,N_19160,N_19330);
and U20441 (N_20441,N_19910,N_19530);
nor U20442 (N_20442,N_19456,N_19652);
xnor U20443 (N_20443,N_19260,N_19896);
xnor U20444 (N_20444,N_19399,N_19943);
xnor U20445 (N_20445,N_19311,N_19899);
and U20446 (N_20446,N_19398,N_19758);
nand U20447 (N_20447,N_19793,N_19942);
and U20448 (N_20448,N_19591,N_19434);
or U20449 (N_20449,N_19873,N_19200);
nand U20450 (N_20450,N_19487,N_19165);
nand U20451 (N_20451,N_19248,N_19855);
xor U20452 (N_20452,N_19701,N_19437);
nand U20453 (N_20453,N_19697,N_19502);
or U20454 (N_20454,N_19426,N_19105);
or U20455 (N_20455,N_19379,N_19753);
nand U20456 (N_20456,N_19277,N_19184);
nand U20457 (N_20457,N_19421,N_19369);
and U20458 (N_20458,N_19007,N_19772);
or U20459 (N_20459,N_19390,N_19512);
nand U20460 (N_20460,N_19870,N_19792);
nand U20461 (N_20461,N_19930,N_19657);
or U20462 (N_20462,N_19448,N_19293);
or U20463 (N_20463,N_19609,N_19183);
and U20464 (N_20464,N_19097,N_19550);
xnor U20465 (N_20465,N_19847,N_19016);
or U20466 (N_20466,N_19755,N_19958);
and U20467 (N_20467,N_19106,N_19381);
nand U20468 (N_20468,N_19182,N_19805);
xnor U20469 (N_20469,N_19267,N_19969);
nor U20470 (N_20470,N_19337,N_19821);
nor U20471 (N_20471,N_19212,N_19858);
or U20472 (N_20472,N_19508,N_19044);
and U20473 (N_20473,N_19537,N_19251);
nand U20474 (N_20474,N_19444,N_19768);
nor U20475 (N_20475,N_19599,N_19060);
or U20476 (N_20476,N_19365,N_19743);
nor U20477 (N_20477,N_19527,N_19329);
or U20478 (N_20478,N_19194,N_19879);
or U20479 (N_20479,N_19249,N_19732);
or U20480 (N_20480,N_19825,N_19107);
xnor U20481 (N_20481,N_19640,N_19618);
xor U20482 (N_20482,N_19764,N_19472);
and U20483 (N_20483,N_19519,N_19342);
nand U20484 (N_20484,N_19782,N_19454);
nand U20485 (N_20485,N_19108,N_19736);
and U20486 (N_20486,N_19209,N_19338);
nor U20487 (N_20487,N_19152,N_19630);
or U20488 (N_20488,N_19604,N_19913);
nor U20489 (N_20489,N_19745,N_19973);
xnor U20490 (N_20490,N_19464,N_19981);
nand U20491 (N_20491,N_19781,N_19612);
nand U20492 (N_20492,N_19536,N_19346);
or U20493 (N_20493,N_19363,N_19469);
and U20494 (N_20494,N_19803,N_19091);
and U20495 (N_20495,N_19268,N_19135);
xor U20496 (N_20496,N_19025,N_19118);
nor U20497 (N_20497,N_19001,N_19995);
and U20498 (N_20498,N_19785,N_19213);
nor U20499 (N_20499,N_19718,N_19602);
nor U20500 (N_20500,N_19452,N_19959);
and U20501 (N_20501,N_19212,N_19129);
nand U20502 (N_20502,N_19108,N_19827);
xor U20503 (N_20503,N_19416,N_19540);
nand U20504 (N_20504,N_19505,N_19907);
nor U20505 (N_20505,N_19756,N_19031);
or U20506 (N_20506,N_19587,N_19956);
nand U20507 (N_20507,N_19856,N_19892);
nor U20508 (N_20508,N_19791,N_19245);
xnor U20509 (N_20509,N_19903,N_19104);
and U20510 (N_20510,N_19105,N_19078);
and U20511 (N_20511,N_19244,N_19105);
nor U20512 (N_20512,N_19488,N_19013);
or U20513 (N_20513,N_19265,N_19691);
nor U20514 (N_20514,N_19113,N_19047);
and U20515 (N_20515,N_19179,N_19573);
xnor U20516 (N_20516,N_19901,N_19931);
and U20517 (N_20517,N_19771,N_19274);
or U20518 (N_20518,N_19185,N_19245);
or U20519 (N_20519,N_19877,N_19136);
nand U20520 (N_20520,N_19953,N_19618);
xor U20521 (N_20521,N_19490,N_19400);
xor U20522 (N_20522,N_19538,N_19899);
or U20523 (N_20523,N_19110,N_19886);
xor U20524 (N_20524,N_19679,N_19856);
nand U20525 (N_20525,N_19042,N_19441);
xnor U20526 (N_20526,N_19623,N_19795);
or U20527 (N_20527,N_19846,N_19213);
or U20528 (N_20528,N_19027,N_19413);
or U20529 (N_20529,N_19822,N_19237);
nand U20530 (N_20530,N_19028,N_19135);
or U20531 (N_20531,N_19272,N_19721);
or U20532 (N_20532,N_19992,N_19153);
and U20533 (N_20533,N_19536,N_19510);
or U20534 (N_20534,N_19264,N_19758);
and U20535 (N_20535,N_19224,N_19096);
nand U20536 (N_20536,N_19215,N_19632);
and U20537 (N_20537,N_19016,N_19409);
nand U20538 (N_20538,N_19043,N_19477);
or U20539 (N_20539,N_19434,N_19229);
nor U20540 (N_20540,N_19844,N_19722);
and U20541 (N_20541,N_19061,N_19052);
nand U20542 (N_20542,N_19972,N_19136);
nor U20543 (N_20543,N_19824,N_19353);
nor U20544 (N_20544,N_19695,N_19977);
and U20545 (N_20545,N_19143,N_19642);
xor U20546 (N_20546,N_19971,N_19263);
nand U20547 (N_20547,N_19776,N_19048);
xnor U20548 (N_20548,N_19954,N_19483);
nand U20549 (N_20549,N_19646,N_19613);
and U20550 (N_20550,N_19453,N_19883);
xor U20551 (N_20551,N_19206,N_19410);
xor U20552 (N_20552,N_19226,N_19960);
xnor U20553 (N_20553,N_19726,N_19076);
nand U20554 (N_20554,N_19059,N_19383);
and U20555 (N_20555,N_19346,N_19525);
and U20556 (N_20556,N_19551,N_19276);
or U20557 (N_20557,N_19760,N_19279);
or U20558 (N_20558,N_19431,N_19513);
nor U20559 (N_20559,N_19407,N_19668);
xnor U20560 (N_20560,N_19633,N_19218);
xnor U20561 (N_20561,N_19761,N_19225);
nor U20562 (N_20562,N_19238,N_19485);
or U20563 (N_20563,N_19490,N_19001);
nand U20564 (N_20564,N_19052,N_19170);
nor U20565 (N_20565,N_19547,N_19836);
nor U20566 (N_20566,N_19601,N_19062);
and U20567 (N_20567,N_19195,N_19011);
nand U20568 (N_20568,N_19930,N_19150);
or U20569 (N_20569,N_19673,N_19905);
nor U20570 (N_20570,N_19685,N_19356);
xnor U20571 (N_20571,N_19246,N_19082);
nand U20572 (N_20572,N_19581,N_19225);
nor U20573 (N_20573,N_19274,N_19365);
and U20574 (N_20574,N_19951,N_19746);
nor U20575 (N_20575,N_19115,N_19405);
or U20576 (N_20576,N_19123,N_19537);
nor U20577 (N_20577,N_19814,N_19545);
nand U20578 (N_20578,N_19845,N_19461);
xor U20579 (N_20579,N_19115,N_19584);
or U20580 (N_20580,N_19764,N_19443);
or U20581 (N_20581,N_19156,N_19265);
or U20582 (N_20582,N_19638,N_19194);
nor U20583 (N_20583,N_19877,N_19869);
or U20584 (N_20584,N_19179,N_19863);
and U20585 (N_20585,N_19715,N_19981);
nand U20586 (N_20586,N_19972,N_19873);
and U20587 (N_20587,N_19940,N_19376);
and U20588 (N_20588,N_19093,N_19455);
and U20589 (N_20589,N_19352,N_19361);
and U20590 (N_20590,N_19112,N_19414);
or U20591 (N_20591,N_19629,N_19061);
xor U20592 (N_20592,N_19802,N_19580);
xnor U20593 (N_20593,N_19367,N_19334);
or U20594 (N_20594,N_19266,N_19608);
or U20595 (N_20595,N_19888,N_19776);
or U20596 (N_20596,N_19717,N_19341);
and U20597 (N_20597,N_19179,N_19774);
or U20598 (N_20598,N_19076,N_19816);
nand U20599 (N_20599,N_19583,N_19062);
xor U20600 (N_20600,N_19047,N_19312);
nand U20601 (N_20601,N_19421,N_19194);
or U20602 (N_20602,N_19553,N_19345);
xor U20603 (N_20603,N_19339,N_19552);
and U20604 (N_20604,N_19478,N_19746);
nor U20605 (N_20605,N_19058,N_19334);
or U20606 (N_20606,N_19697,N_19264);
nand U20607 (N_20607,N_19654,N_19997);
xnor U20608 (N_20608,N_19461,N_19706);
and U20609 (N_20609,N_19627,N_19880);
or U20610 (N_20610,N_19578,N_19604);
nand U20611 (N_20611,N_19290,N_19078);
and U20612 (N_20612,N_19258,N_19977);
and U20613 (N_20613,N_19126,N_19085);
and U20614 (N_20614,N_19902,N_19952);
xor U20615 (N_20615,N_19693,N_19435);
nor U20616 (N_20616,N_19878,N_19881);
xnor U20617 (N_20617,N_19217,N_19037);
nor U20618 (N_20618,N_19277,N_19010);
nand U20619 (N_20619,N_19325,N_19406);
and U20620 (N_20620,N_19651,N_19224);
xor U20621 (N_20621,N_19140,N_19089);
xor U20622 (N_20622,N_19643,N_19562);
or U20623 (N_20623,N_19992,N_19956);
and U20624 (N_20624,N_19510,N_19388);
and U20625 (N_20625,N_19019,N_19577);
and U20626 (N_20626,N_19455,N_19098);
nand U20627 (N_20627,N_19033,N_19860);
or U20628 (N_20628,N_19245,N_19516);
and U20629 (N_20629,N_19418,N_19289);
or U20630 (N_20630,N_19889,N_19527);
nor U20631 (N_20631,N_19969,N_19873);
xnor U20632 (N_20632,N_19515,N_19658);
nor U20633 (N_20633,N_19130,N_19199);
or U20634 (N_20634,N_19888,N_19631);
nand U20635 (N_20635,N_19810,N_19782);
nand U20636 (N_20636,N_19505,N_19663);
nand U20637 (N_20637,N_19091,N_19480);
xor U20638 (N_20638,N_19174,N_19984);
xnor U20639 (N_20639,N_19339,N_19599);
and U20640 (N_20640,N_19285,N_19019);
nor U20641 (N_20641,N_19961,N_19439);
xnor U20642 (N_20642,N_19999,N_19497);
nand U20643 (N_20643,N_19451,N_19547);
xnor U20644 (N_20644,N_19884,N_19303);
and U20645 (N_20645,N_19243,N_19330);
nor U20646 (N_20646,N_19221,N_19162);
or U20647 (N_20647,N_19121,N_19382);
xor U20648 (N_20648,N_19280,N_19021);
nor U20649 (N_20649,N_19072,N_19777);
nand U20650 (N_20650,N_19572,N_19394);
nand U20651 (N_20651,N_19374,N_19749);
nor U20652 (N_20652,N_19151,N_19282);
nor U20653 (N_20653,N_19538,N_19286);
or U20654 (N_20654,N_19668,N_19630);
or U20655 (N_20655,N_19834,N_19459);
or U20656 (N_20656,N_19675,N_19725);
nand U20657 (N_20657,N_19066,N_19326);
nand U20658 (N_20658,N_19872,N_19057);
nor U20659 (N_20659,N_19530,N_19153);
or U20660 (N_20660,N_19541,N_19011);
and U20661 (N_20661,N_19103,N_19060);
nor U20662 (N_20662,N_19079,N_19761);
and U20663 (N_20663,N_19626,N_19402);
and U20664 (N_20664,N_19918,N_19232);
nor U20665 (N_20665,N_19090,N_19140);
nor U20666 (N_20666,N_19036,N_19953);
nand U20667 (N_20667,N_19832,N_19046);
xnor U20668 (N_20668,N_19653,N_19110);
or U20669 (N_20669,N_19096,N_19704);
nand U20670 (N_20670,N_19060,N_19820);
nor U20671 (N_20671,N_19963,N_19631);
and U20672 (N_20672,N_19786,N_19822);
or U20673 (N_20673,N_19091,N_19235);
nand U20674 (N_20674,N_19712,N_19592);
and U20675 (N_20675,N_19339,N_19539);
xnor U20676 (N_20676,N_19756,N_19568);
xnor U20677 (N_20677,N_19328,N_19845);
and U20678 (N_20678,N_19715,N_19582);
or U20679 (N_20679,N_19585,N_19207);
and U20680 (N_20680,N_19010,N_19331);
nor U20681 (N_20681,N_19942,N_19980);
nand U20682 (N_20682,N_19096,N_19420);
nor U20683 (N_20683,N_19617,N_19132);
xnor U20684 (N_20684,N_19208,N_19356);
and U20685 (N_20685,N_19928,N_19109);
nor U20686 (N_20686,N_19319,N_19822);
and U20687 (N_20687,N_19621,N_19491);
or U20688 (N_20688,N_19005,N_19914);
xnor U20689 (N_20689,N_19247,N_19679);
nand U20690 (N_20690,N_19357,N_19774);
nand U20691 (N_20691,N_19396,N_19610);
nand U20692 (N_20692,N_19248,N_19140);
or U20693 (N_20693,N_19883,N_19761);
xnor U20694 (N_20694,N_19806,N_19498);
or U20695 (N_20695,N_19809,N_19681);
xor U20696 (N_20696,N_19732,N_19153);
xnor U20697 (N_20697,N_19787,N_19367);
nor U20698 (N_20698,N_19974,N_19827);
nor U20699 (N_20699,N_19110,N_19134);
xnor U20700 (N_20700,N_19272,N_19107);
xor U20701 (N_20701,N_19440,N_19938);
nor U20702 (N_20702,N_19111,N_19662);
nand U20703 (N_20703,N_19341,N_19484);
or U20704 (N_20704,N_19837,N_19060);
or U20705 (N_20705,N_19997,N_19912);
xnor U20706 (N_20706,N_19292,N_19397);
nand U20707 (N_20707,N_19115,N_19759);
nand U20708 (N_20708,N_19056,N_19365);
nand U20709 (N_20709,N_19579,N_19334);
nor U20710 (N_20710,N_19606,N_19366);
nand U20711 (N_20711,N_19583,N_19762);
nand U20712 (N_20712,N_19486,N_19302);
nand U20713 (N_20713,N_19429,N_19340);
nor U20714 (N_20714,N_19207,N_19675);
xor U20715 (N_20715,N_19991,N_19658);
nand U20716 (N_20716,N_19427,N_19542);
or U20717 (N_20717,N_19652,N_19035);
nand U20718 (N_20718,N_19832,N_19586);
nor U20719 (N_20719,N_19771,N_19077);
and U20720 (N_20720,N_19761,N_19438);
and U20721 (N_20721,N_19269,N_19688);
nor U20722 (N_20722,N_19206,N_19483);
xnor U20723 (N_20723,N_19281,N_19569);
and U20724 (N_20724,N_19668,N_19376);
and U20725 (N_20725,N_19768,N_19046);
nand U20726 (N_20726,N_19182,N_19780);
nand U20727 (N_20727,N_19518,N_19480);
and U20728 (N_20728,N_19351,N_19663);
and U20729 (N_20729,N_19638,N_19213);
and U20730 (N_20730,N_19836,N_19752);
or U20731 (N_20731,N_19804,N_19533);
or U20732 (N_20732,N_19920,N_19709);
and U20733 (N_20733,N_19010,N_19956);
nand U20734 (N_20734,N_19941,N_19602);
nand U20735 (N_20735,N_19826,N_19489);
and U20736 (N_20736,N_19598,N_19178);
xnor U20737 (N_20737,N_19422,N_19760);
and U20738 (N_20738,N_19754,N_19406);
or U20739 (N_20739,N_19591,N_19099);
or U20740 (N_20740,N_19019,N_19766);
and U20741 (N_20741,N_19416,N_19007);
xnor U20742 (N_20742,N_19461,N_19925);
or U20743 (N_20743,N_19276,N_19968);
and U20744 (N_20744,N_19021,N_19296);
xor U20745 (N_20745,N_19550,N_19171);
xnor U20746 (N_20746,N_19517,N_19668);
nor U20747 (N_20747,N_19890,N_19802);
and U20748 (N_20748,N_19960,N_19955);
nor U20749 (N_20749,N_19437,N_19569);
xnor U20750 (N_20750,N_19722,N_19492);
xor U20751 (N_20751,N_19945,N_19305);
and U20752 (N_20752,N_19336,N_19989);
xor U20753 (N_20753,N_19819,N_19610);
and U20754 (N_20754,N_19495,N_19393);
or U20755 (N_20755,N_19550,N_19695);
nor U20756 (N_20756,N_19752,N_19292);
and U20757 (N_20757,N_19157,N_19120);
xnor U20758 (N_20758,N_19114,N_19531);
and U20759 (N_20759,N_19018,N_19596);
or U20760 (N_20760,N_19620,N_19260);
nor U20761 (N_20761,N_19197,N_19566);
or U20762 (N_20762,N_19112,N_19245);
xnor U20763 (N_20763,N_19750,N_19961);
xor U20764 (N_20764,N_19040,N_19046);
xor U20765 (N_20765,N_19768,N_19623);
and U20766 (N_20766,N_19496,N_19316);
and U20767 (N_20767,N_19796,N_19160);
nor U20768 (N_20768,N_19898,N_19335);
nand U20769 (N_20769,N_19359,N_19416);
xor U20770 (N_20770,N_19981,N_19708);
xnor U20771 (N_20771,N_19752,N_19438);
xor U20772 (N_20772,N_19331,N_19305);
nor U20773 (N_20773,N_19151,N_19633);
and U20774 (N_20774,N_19462,N_19577);
nor U20775 (N_20775,N_19158,N_19889);
and U20776 (N_20776,N_19634,N_19274);
nor U20777 (N_20777,N_19880,N_19424);
and U20778 (N_20778,N_19417,N_19443);
xor U20779 (N_20779,N_19745,N_19688);
nor U20780 (N_20780,N_19378,N_19022);
nand U20781 (N_20781,N_19656,N_19647);
xor U20782 (N_20782,N_19304,N_19688);
nor U20783 (N_20783,N_19821,N_19653);
xnor U20784 (N_20784,N_19226,N_19062);
nor U20785 (N_20785,N_19489,N_19715);
nor U20786 (N_20786,N_19934,N_19343);
and U20787 (N_20787,N_19847,N_19446);
and U20788 (N_20788,N_19909,N_19104);
nand U20789 (N_20789,N_19954,N_19777);
xnor U20790 (N_20790,N_19012,N_19919);
xnor U20791 (N_20791,N_19712,N_19720);
nand U20792 (N_20792,N_19298,N_19021);
xnor U20793 (N_20793,N_19825,N_19659);
nand U20794 (N_20794,N_19091,N_19455);
or U20795 (N_20795,N_19665,N_19330);
and U20796 (N_20796,N_19078,N_19427);
or U20797 (N_20797,N_19105,N_19609);
xor U20798 (N_20798,N_19135,N_19918);
nand U20799 (N_20799,N_19178,N_19293);
nor U20800 (N_20800,N_19726,N_19055);
or U20801 (N_20801,N_19834,N_19284);
and U20802 (N_20802,N_19138,N_19920);
or U20803 (N_20803,N_19580,N_19409);
nor U20804 (N_20804,N_19794,N_19503);
nor U20805 (N_20805,N_19238,N_19346);
nor U20806 (N_20806,N_19970,N_19509);
nor U20807 (N_20807,N_19581,N_19769);
xor U20808 (N_20808,N_19790,N_19394);
nand U20809 (N_20809,N_19410,N_19423);
nand U20810 (N_20810,N_19386,N_19484);
xor U20811 (N_20811,N_19718,N_19598);
nand U20812 (N_20812,N_19322,N_19501);
nand U20813 (N_20813,N_19808,N_19093);
and U20814 (N_20814,N_19318,N_19059);
xor U20815 (N_20815,N_19386,N_19612);
or U20816 (N_20816,N_19806,N_19189);
xor U20817 (N_20817,N_19580,N_19706);
nand U20818 (N_20818,N_19073,N_19387);
or U20819 (N_20819,N_19157,N_19193);
or U20820 (N_20820,N_19773,N_19101);
and U20821 (N_20821,N_19102,N_19893);
xor U20822 (N_20822,N_19729,N_19373);
nand U20823 (N_20823,N_19824,N_19554);
or U20824 (N_20824,N_19245,N_19131);
xor U20825 (N_20825,N_19091,N_19645);
or U20826 (N_20826,N_19221,N_19332);
nor U20827 (N_20827,N_19722,N_19666);
and U20828 (N_20828,N_19220,N_19227);
and U20829 (N_20829,N_19256,N_19065);
and U20830 (N_20830,N_19498,N_19743);
or U20831 (N_20831,N_19973,N_19810);
or U20832 (N_20832,N_19132,N_19085);
or U20833 (N_20833,N_19705,N_19525);
nor U20834 (N_20834,N_19646,N_19020);
nor U20835 (N_20835,N_19146,N_19482);
xor U20836 (N_20836,N_19625,N_19111);
nand U20837 (N_20837,N_19155,N_19816);
xnor U20838 (N_20838,N_19576,N_19356);
nand U20839 (N_20839,N_19323,N_19979);
or U20840 (N_20840,N_19466,N_19887);
and U20841 (N_20841,N_19989,N_19759);
or U20842 (N_20842,N_19012,N_19187);
and U20843 (N_20843,N_19457,N_19770);
xnor U20844 (N_20844,N_19887,N_19372);
xnor U20845 (N_20845,N_19735,N_19586);
nand U20846 (N_20846,N_19627,N_19144);
xor U20847 (N_20847,N_19731,N_19507);
nand U20848 (N_20848,N_19101,N_19600);
or U20849 (N_20849,N_19130,N_19645);
nand U20850 (N_20850,N_19244,N_19575);
nand U20851 (N_20851,N_19268,N_19375);
and U20852 (N_20852,N_19978,N_19076);
nor U20853 (N_20853,N_19334,N_19300);
or U20854 (N_20854,N_19696,N_19656);
or U20855 (N_20855,N_19795,N_19593);
and U20856 (N_20856,N_19327,N_19717);
or U20857 (N_20857,N_19717,N_19883);
nor U20858 (N_20858,N_19170,N_19948);
nor U20859 (N_20859,N_19204,N_19741);
or U20860 (N_20860,N_19831,N_19803);
nor U20861 (N_20861,N_19630,N_19280);
or U20862 (N_20862,N_19630,N_19383);
xor U20863 (N_20863,N_19892,N_19678);
nand U20864 (N_20864,N_19782,N_19722);
nand U20865 (N_20865,N_19168,N_19806);
nand U20866 (N_20866,N_19654,N_19878);
or U20867 (N_20867,N_19862,N_19242);
nand U20868 (N_20868,N_19136,N_19312);
or U20869 (N_20869,N_19552,N_19521);
nand U20870 (N_20870,N_19632,N_19904);
nor U20871 (N_20871,N_19348,N_19422);
nand U20872 (N_20872,N_19813,N_19096);
and U20873 (N_20873,N_19975,N_19314);
nor U20874 (N_20874,N_19037,N_19452);
or U20875 (N_20875,N_19836,N_19435);
or U20876 (N_20876,N_19166,N_19812);
and U20877 (N_20877,N_19434,N_19280);
xnor U20878 (N_20878,N_19851,N_19776);
or U20879 (N_20879,N_19005,N_19705);
xnor U20880 (N_20880,N_19178,N_19931);
or U20881 (N_20881,N_19795,N_19191);
and U20882 (N_20882,N_19716,N_19451);
nor U20883 (N_20883,N_19224,N_19669);
and U20884 (N_20884,N_19466,N_19783);
xnor U20885 (N_20885,N_19212,N_19384);
nand U20886 (N_20886,N_19824,N_19032);
nor U20887 (N_20887,N_19169,N_19214);
xor U20888 (N_20888,N_19068,N_19641);
xnor U20889 (N_20889,N_19678,N_19235);
xor U20890 (N_20890,N_19811,N_19128);
xnor U20891 (N_20891,N_19531,N_19658);
nor U20892 (N_20892,N_19688,N_19663);
or U20893 (N_20893,N_19278,N_19617);
and U20894 (N_20894,N_19813,N_19571);
or U20895 (N_20895,N_19332,N_19157);
and U20896 (N_20896,N_19215,N_19610);
xnor U20897 (N_20897,N_19106,N_19063);
xor U20898 (N_20898,N_19620,N_19094);
and U20899 (N_20899,N_19876,N_19895);
and U20900 (N_20900,N_19461,N_19283);
nor U20901 (N_20901,N_19149,N_19703);
xor U20902 (N_20902,N_19610,N_19611);
nand U20903 (N_20903,N_19421,N_19262);
xor U20904 (N_20904,N_19531,N_19816);
xor U20905 (N_20905,N_19410,N_19677);
nand U20906 (N_20906,N_19736,N_19947);
xor U20907 (N_20907,N_19180,N_19900);
nor U20908 (N_20908,N_19161,N_19629);
xnor U20909 (N_20909,N_19157,N_19220);
nor U20910 (N_20910,N_19748,N_19518);
nand U20911 (N_20911,N_19090,N_19590);
or U20912 (N_20912,N_19285,N_19245);
nand U20913 (N_20913,N_19615,N_19482);
or U20914 (N_20914,N_19963,N_19743);
xnor U20915 (N_20915,N_19375,N_19794);
or U20916 (N_20916,N_19133,N_19144);
nand U20917 (N_20917,N_19439,N_19234);
and U20918 (N_20918,N_19190,N_19595);
or U20919 (N_20919,N_19990,N_19626);
and U20920 (N_20920,N_19652,N_19316);
or U20921 (N_20921,N_19582,N_19656);
nand U20922 (N_20922,N_19639,N_19688);
and U20923 (N_20923,N_19663,N_19174);
or U20924 (N_20924,N_19506,N_19139);
nor U20925 (N_20925,N_19524,N_19742);
xor U20926 (N_20926,N_19723,N_19888);
and U20927 (N_20927,N_19942,N_19936);
xnor U20928 (N_20928,N_19882,N_19222);
xor U20929 (N_20929,N_19896,N_19984);
or U20930 (N_20930,N_19311,N_19581);
and U20931 (N_20931,N_19572,N_19335);
nand U20932 (N_20932,N_19070,N_19112);
nand U20933 (N_20933,N_19923,N_19410);
nor U20934 (N_20934,N_19701,N_19299);
and U20935 (N_20935,N_19896,N_19899);
nand U20936 (N_20936,N_19489,N_19700);
or U20937 (N_20937,N_19617,N_19044);
nor U20938 (N_20938,N_19719,N_19284);
nor U20939 (N_20939,N_19744,N_19463);
xor U20940 (N_20940,N_19553,N_19626);
nor U20941 (N_20941,N_19500,N_19522);
nor U20942 (N_20942,N_19158,N_19278);
and U20943 (N_20943,N_19312,N_19570);
and U20944 (N_20944,N_19941,N_19232);
xnor U20945 (N_20945,N_19442,N_19664);
nand U20946 (N_20946,N_19185,N_19679);
and U20947 (N_20947,N_19827,N_19063);
or U20948 (N_20948,N_19578,N_19522);
nor U20949 (N_20949,N_19238,N_19825);
nor U20950 (N_20950,N_19685,N_19296);
or U20951 (N_20951,N_19295,N_19539);
nor U20952 (N_20952,N_19361,N_19051);
or U20953 (N_20953,N_19590,N_19248);
or U20954 (N_20954,N_19462,N_19380);
or U20955 (N_20955,N_19742,N_19018);
nor U20956 (N_20956,N_19405,N_19869);
or U20957 (N_20957,N_19710,N_19005);
nor U20958 (N_20958,N_19179,N_19529);
xor U20959 (N_20959,N_19234,N_19332);
or U20960 (N_20960,N_19683,N_19189);
nand U20961 (N_20961,N_19324,N_19828);
and U20962 (N_20962,N_19707,N_19215);
or U20963 (N_20963,N_19595,N_19922);
xnor U20964 (N_20964,N_19615,N_19527);
and U20965 (N_20965,N_19195,N_19016);
nor U20966 (N_20966,N_19275,N_19988);
nor U20967 (N_20967,N_19932,N_19459);
or U20968 (N_20968,N_19641,N_19865);
nor U20969 (N_20969,N_19514,N_19526);
xnor U20970 (N_20970,N_19515,N_19350);
or U20971 (N_20971,N_19054,N_19182);
xnor U20972 (N_20972,N_19707,N_19907);
nor U20973 (N_20973,N_19625,N_19028);
nand U20974 (N_20974,N_19084,N_19539);
xnor U20975 (N_20975,N_19187,N_19441);
nand U20976 (N_20976,N_19361,N_19180);
nor U20977 (N_20977,N_19396,N_19351);
xnor U20978 (N_20978,N_19506,N_19905);
or U20979 (N_20979,N_19655,N_19830);
xor U20980 (N_20980,N_19858,N_19042);
xnor U20981 (N_20981,N_19670,N_19351);
nand U20982 (N_20982,N_19770,N_19649);
xnor U20983 (N_20983,N_19263,N_19913);
nor U20984 (N_20984,N_19013,N_19320);
nand U20985 (N_20985,N_19078,N_19793);
and U20986 (N_20986,N_19285,N_19231);
and U20987 (N_20987,N_19934,N_19794);
nand U20988 (N_20988,N_19454,N_19083);
and U20989 (N_20989,N_19508,N_19307);
or U20990 (N_20990,N_19987,N_19923);
and U20991 (N_20991,N_19654,N_19581);
and U20992 (N_20992,N_19324,N_19806);
or U20993 (N_20993,N_19130,N_19338);
and U20994 (N_20994,N_19894,N_19074);
and U20995 (N_20995,N_19282,N_19422);
nor U20996 (N_20996,N_19231,N_19827);
nand U20997 (N_20997,N_19214,N_19706);
or U20998 (N_20998,N_19627,N_19505);
xnor U20999 (N_20999,N_19619,N_19917);
or U21000 (N_21000,N_20321,N_20466);
xor U21001 (N_21001,N_20939,N_20996);
or U21002 (N_21002,N_20176,N_20608);
nand U21003 (N_21003,N_20428,N_20850);
nor U21004 (N_21004,N_20730,N_20600);
nand U21005 (N_21005,N_20742,N_20698);
xor U21006 (N_21006,N_20822,N_20301);
nand U21007 (N_21007,N_20292,N_20553);
nor U21008 (N_21008,N_20255,N_20672);
and U21009 (N_21009,N_20219,N_20794);
or U21010 (N_21010,N_20015,N_20772);
and U21011 (N_21011,N_20193,N_20477);
and U21012 (N_21012,N_20530,N_20297);
nor U21013 (N_21013,N_20699,N_20796);
xnor U21014 (N_21014,N_20688,N_20873);
and U21015 (N_21015,N_20327,N_20966);
or U21016 (N_21016,N_20992,N_20941);
xor U21017 (N_21017,N_20729,N_20037);
xor U21018 (N_21018,N_20066,N_20564);
and U21019 (N_21019,N_20005,N_20731);
nand U21020 (N_21020,N_20139,N_20159);
xnor U21021 (N_21021,N_20481,N_20618);
nor U21022 (N_21022,N_20187,N_20231);
and U21023 (N_21023,N_20432,N_20505);
nand U21024 (N_21024,N_20899,N_20583);
xor U21025 (N_21025,N_20640,N_20419);
xor U21026 (N_21026,N_20149,N_20323);
or U21027 (N_21027,N_20767,N_20749);
xor U21028 (N_21028,N_20874,N_20174);
or U21029 (N_21029,N_20011,N_20085);
and U21030 (N_21030,N_20702,N_20467);
or U21031 (N_21031,N_20524,N_20629);
or U21032 (N_21032,N_20907,N_20832);
xnor U21033 (N_21033,N_20570,N_20389);
or U21034 (N_21034,N_20230,N_20778);
or U21035 (N_21035,N_20398,N_20995);
nor U21036 (N_21036,N_20980,N_20185);
nand U21037 (N_21037,N_20058,N_20240);
nor U21038 (N_21038,N_20844,N_20206);
nor U21039 (N_21039,N_20764,N_20334);
xor U21040 (N_21040,N_20599,N_20726);
and U21041 (N_21041,N_20829,N_20962);
nand U21042 (N_21042,N_20133,N_20735);
nor U21043 (N_21043,N_20320,N_20302);
xnor U21044 (N_21044,N_20578,N_20346);
xnor U21045 (N_21045,N_20169,N_20867);
nand U21046 (N_21046,N_20342,N_20399);
and U21047 (N_21047,N_20619,N_20353);
and U21048 (N_21048,N_20606,N_20792);
xnor U21049 (N_21049,N_20090,N_20465);
and U21050 (N_21050,N_20961,N_20827);
nor U21051 (N_21051,N_20331,N_20842);
nand U21052 (N_21052,N_20910,N_20486);
nand U21053 (N_21053,N_20359,N_20442);
xor U21054 (N_21054,N_20551,N_20179);
and U21055 (N_21055,N_20934,N_20659);
nand U21056 (N_21056,N_20237,N_20709);
nor U21057 (N_21057,N_20492,N_20958);
nand U21058 (N_21058,N_20009,N_20110);
xnor U21059 (N_21059,N_20135,N_20851);
and U21060 (N_21060,N_20682,N_20663);
nand U21061 (N_21061,N_20040,N_20417);
or U21062 (N_21062,N_20859,N_20100);
and U21063 (N_21063,N_20126,N_20340);
and U21064 (N_21064,N_20454,N_20054);
nor U21065 (N_21065,N_20523,N_20987);
and U21066 (N_21066,N_20444,N_20164);
xor U21067 (N_21067,N_20386,N_20194);
and U21068 (N_21068,N_20871,N_20025);
xnor U21069 (N_21069,N_20434,N_20865);
xor U21070 (N_21070,N_20991,N_20002);
and U21071 (N_21071,N_20338,N_20294);
xnor U21072 (N_21072,N_20122,N_20036);
nor U21073 (N_21073,N_20830,N_20216);
xnor U21074 (N_21074,N_20213,N_20579);
and U21075 (N_21075,N_20623,N_20568);
and U21076 (N_21076,N_20445,N_20979);
xnor U21077 (N_21077,N_20718,N_20636);
nor U21078 (N_21078,N_20549,N_20300);
nor U21079 (N_21079,N_20032,N_20339);
or U21080 (N_21080,N_20312,N_20086);
and U21081 (N_21081,N_20499,N_20106);
and U21082 (N_21082,N_20746,N_20348);
and U21083 (N_21083,N_20437,N_20156);
nor U21084 (N_21084,N_20379,N_20113);
or U21085 (N_21085,N_20968,N_20614);
and U21086 (N_21086,N_20083,N_20686);
xor U21087 (N_21087,N_20581,N_20155);
nand U21088 (N_21088,N_20819,N_20502);
xnor U21089 (N_21089,N_20922,N_20175);
and U21090 (N_21090,N_20960,N_20522);
or U21091 (N_21091,N_20453,N_20092);
and U21092 (N_21092,N_20247,N_20217);
nor U21093 (N_21093,N_20949,N_20006);
and U21094 (N_21094,N_20520,N_20864);
and U21095 (N_21095,N_20265,N_20809);
nor U21096 (N_21096,N_20261,N_20412);
nand U21097 (N_21097,N_20021,N_20970);
and U21098 (N_21098,N_20147,N_20203);
nor U21099 (N_21099,N_20138,N_20236);
nor U21100 (N_21100,N_20634,N_20983);
nand U21101 (N_21101,N_20103,N_20542);
nor U21102 (N_21102,N_20439,N_20343);
nor U21103 (N_21103,N_20798,N_20114);
xnor U21104 (N_21104,N_20161,N_20836);
nand U21105 (N_21105,N_20993,N_20413);
xnor U21106 (N_21106,N_20986,N_20436);
xnor U21107 (N_21107,N_20531,N_20763);
or U21108 (N_21108,N_20567,N_20330);
or U21109 (N_21109,N_20226,N_20532);
xor U21110 (N_21110,N_20503,N_20047);
nor U21111 (N_21111,N_20953,N_20184);
nor U21112 (N_21112,N_20645,N_20109);
or U21113 (N_21113,N_20306,N_20335);
nand U21114 (N_21114,N_20325,N_20501);
nor U21115 (N_21115,N_20890,N_20653);
nand U21116 (N_21116,N_20266,N_20616);
xnor U21117 (N_21117,N_20029,N_20031);
nor U21118 (N_21118,N_20153,N_20264);
nor U21119 (N_21119,N_20635,N_20038);
or U21120 (N_21120,N_20136,N_20391);
and U21121 (N_21121,N_20057,N_20761);
and U21122 (N_21122,N_20811,N_20356);
nor U21123 (N_21123,N_20725,N_20456);
xor U21124 (N_21124,N_20202,N_20768);
nand U21125 (N_21125,N_20372,N_20738);
xnor U21126 (N_21126,N_20207,N_20183);
or U21127 (N_21127,N_20607,N_20282);
nor U21128 (N_21128,N_20807,N_20494);
nor U21129 (N_21129,N_20198,N_20420);
or U21130 (N_21130,N_20368,N_20493);
or U21131 (N_21131,N_20740,N_20234);
and U21132 (N_21132,N_20878,N_20592);
nor U21133 (N_21133,N_20246,N_20518);
and U21134 (N_21134,N_20228,N_20162);
or U21135 (N_21135,N_20209,N_20943);
or U21136 (N_21136,N_20068,N_20818);
xor U21137 (N_21137,N_20181,N_20951);
and U21138 (N_21138,N_20963,N_20509);
nand U21139 (N_21139,N_20401,N_20008);
or U21140 (N_21140,N_20733,N_20506);
and U21141 (N_21141,N_20920,N_20650);
and U21142 (N_21142,N_20096,N_20797);
nor U21143 (N_21143,N_20559,N_20075);
nor U21144 (N_21144,N_20393,N_20957);
nand U21145 (N_21145,N_20762,N_20076);
and U21146 (N_21146,N_20846,N_20383);
nor U21147 (N_21147,N_20081,N_20329);
or U21148 (N_21148,N_20690,N_20596);
nand U21149 (N_21149,N_20351,N_20286);
xnor U21150 (N_21150,N_20847,N_20728);
nand U21151 (N_21151,N_20357,N_20214);
nor U21152 (N_21152,N_20938,N_20710);
or U21153 (N_21153,N_20295,N_20558);
or U21154 (N_21154,N_20367,N_20802);
nor U21155 (N_21155,N_20358,N_20223);
and U21156 (N_21156,N_20681,N_20831);
and U21157 (N_21157,N_20491,N_20188);
nor U21158 (N_21158,N_20272,N_20575);
and U21159 (N_21159,N_20259,N_20345);
and U21160 (N_21160,N_20269,N_20648);
xnor U21161 (N_21161,N_20414,N_20862);
nand U21162 (N_21162,N_20540,N_20630);
nand U21163 (N_21163,N_20459,N_20022);
or U21164 (N_21164,N_20661,N_20803);
xor U21165 (N_21165,N_20571,N_20249);
and U21166 (N_21166,N_20257,N_20416);
or U21167 (N_21167,N_20318,N_20780);
nor U21168 (N_21168,N_20157,N_20902);
nor U21169 (N_21169,N_20990,N_20786);
nand U21170 (N_21170,N_20598,N_20756);
nor U21171 (N_21171,N_20039,N_20489);
nand U21172 (N_21172,N_20839,N_20869);
xnor U21173 (N_21173,N_20285,N_20123);
and U21174 (N_21174,N_20547,N_20984);
nand U21175 (N_21175,N_20546,N_20651);
nor U21176 (N_21176,N_20378,N_20003);
nand U21177 (N_21177,N_20887,N_20077);
nor U21178 (N_21178,N_20160,N_20909);
xnor U21179 (N_21179,N_20468,N_20543);
nor U21180 (N_21180,N_20557,N_20163);
and U21181 (N_21181,N_20610,N_20349);
nor U21182 (N_21182,N_20152,N_20994);
or U21183 (N_21183,N_20253,N_20643);
or U21184 (N_21184,N_20521,N_20460);
nor U21185 (N_21185,N_20171,N_20055);
and U21186 (N_21186,N_20609,N_20576);
or U21187 (N_21187,N_20470,N_20069);
nor U21188 (N_21188,N_20158,N_20143);
and U21189 (N_21189,N_20314,N_20215);
xor U21190 (N_21190,N_20999,N_20433);
nand U21191 (N_21191,N_20224,N_20438);
xnor U21192 (N_21192,N_20712,N_20552);
or U21193 (N_21193,N_20475,N_20748);
and U21194 (N_21194,N_20324,N_20063);
xor U21195 (N_21195,N_20913,N_20923);
or U21196 (N_21196,N_20988,N_20586);
nand U21197 (N_21197,N_20125,N_20424);
nand U21198 (N_21198,N_20151,N_20646);
and U21199 (N_21199,N_20944,N_20402);
and U21200 (N_21200,N_20976,N_20471);
xnor U21201 (N_21201,N_20895,N_20685);
nor U21202 (N_21202,N_20917,N_20997);
nor U21203 (N_21203,N_20880,N_20779);
and U21204 (N_21204,N_20601,N_20930);
or U21205 (N_21205,N_20916,N_20554);
and U21206 (N_21206,N_20277,N_20482);
nand U21207 (N_21207,N_20099,N_20450);
nand U21208 (N_21208,N_20095,N_20817);
or U21209 (N_21209,N_20409,N_20637);
or U21210 (N_21210,N_20507,N_20755);
nor U21211 (N_21211,N_20573,N_20590);
xnor U21212 (N_21212,N_20026,N_20361);
and U21213 (N_21213,N_20906,N_20799);
nor U21214 (N_21214,N_20189,N_20727);
or U21215 (N_21215,N_20644,N_20411);
and U21216 (N_21216,N_20977,N_20824);
nor U21217 (N_21217,N_20239,N_20204);
nand U21218 (N_21218,N_20448,N_20254);
xor U21219 (N_21219,N_20404,N_20737);
nor U21220 (N_21220,N_20469,N_20550);
or U21221 (N_21221,N_20537,N_20132);
or U21222 (N_21222,N_20900,N_20805);
and U21223 (N_21223,N_20130,N_20855);
or U21224 (N_21224,N_20860,N_20921);
nor U21225 (N_21225,N_20782,N_20381);
nand U21226 (N_21226,N_20056,N_20064);
xor U21227 (N_21227,N_20192,N_20734);
or U21228 (N_21228,N_20889,N_20043);
and U21229 (N_21229,N_20362,N_20928);
xnor U21230 (N_21230,N_20671,N_20875);
and U21231 (N_21231,N_20177,N_20089);
nor U21232 (N_21232,N_20197,N_20510);
xnor U21233 (N_21233,N_20408,N_20049);
or U21234 (N_21234,N_20248,N_20476);
nor U21235 (N_21235,N_20369,N_20828);
and U21236 (N_21236,N_20677,N_20182);
nor U21237 (N_21237,N_20858,N_20708);
or U21238 (N_21238,N_20561,N_20884);
or U21239 (N_21239,N_20473,N_20915);
nor U21240 (N_21240,N_20891,N_20933);
or U21241 (N_21241,N_20441,N_20388);
or U21242 (N_21242,N_20757,N_20879);
nor U21243 (N_21243,N_20816,N_20597);
nand U21244 (N_21244,N_20680,N_20704);
and U21245 (N_21245,N_20059,N_20539);
nor U21246 (N_21246,N_20825,N_20079);
nand U21247 (N_21247,N_20484,N_20418);
and U21248 (N_21248,N_20898,N_20497);
and U21249 (N_21249,N_20082,N_20569);
and U21250 (N_21250,N_20380,N_20341);
or U21251 (N_21251,N_20654,N_20914);
or U21252 (N_21252,N_20784,N_20632);
nand U21253 (N_21253,N_20766,N_20812);
and U21254 (N_21254,N_20528,N_20691);
nand U21255 (N_21255,N_20973,N_20344);
nor U21256 (N_21256,N_20487,N_20225);
or U21257 (N_21257,N_20200,N_20694);
and U21258 (N_21258,N_20304,N_20229);
or U21259 (N_21259,N_20050,N_20897);
nor U21260 (N_21260,N_20422,N_20942);
or U21261 (N_21261,N_20087,N_20752);
nand U21262 (N_21262,N_20769,N_20041);
and U21263 (N_21263,N_20291,N_20876);
nand U21264 (N_21264,N_20676,N_20689);
and U21265 (N_21265,N_20795,N_20387);
nand U21266 (N_21266,N_20080,N_20117);
nor U21267 (N_21267,N_20227,N_20745);
and U21268 (N_21268,N_20364,N_20791);
nand U21269 (N_21269,N_20978,N_20626);
nand U21270 (N_21270,N_20919,N_20585);
and U21271 (N_21271,N_20741,N_20771);
and U21272 (N_21272,N_20102,N_20668);
and U21273 (N_21273,N_20326,N_20777);
nor U21274 (N_21274,N_20319,N_20273);
nor U21275 (N_21275,N_20131,N_20244);
nand U21276 (N_21276,N_20017,N_20696);
or U21277 (N_21277,N_20211,N_20027);
or U21278 (N_21278,N_20396,N_20800);
nor U21279 (N_21279,N_20426,N_20360);
and U21280 (N_21280,N_20870,N_20395);
nor U21281 (N_21281,N_20695,N_20628);
and U21282 (N_21282,N_20885,N_20736);
nor U21283 (N_21283,N_20883,N_20400);
xor U21284 (N_21284,N_20703,N_20739);
and U21285 (N_21285,N_20462,N_20390);
nor U21286 (N_21286,N_20834,N_20370);
and U21287 (N_21287,N_20508,N_20621);
nor U21288 (N_21288,N_20714,N_20589);
nand U21289 (N_21289,N_20972,N_20515);
or U21290 (N_21290,N_20406,N_20974);
xor U21291 (N_21291,N_20290,N_20280);
nor U21292 (N_21292,N_20425,N_20529);
nand U21293 (N_21293,N_20602,N_20713);
and U21294 (N_21294,N_20955,N_20101);
and U21295 (N_21295,N_20905,N_20283);
nor U21296 (N_21296,N_20810,N_20641);
nor U21297 (N_21297,N_20371,N_20104);
or U21298 (N_21298,N_20514,N_20299);
xnor U21299 (N_21299,N_20513,N_20337);
nor U21300 (N_21300,N_20721,N_20724);
nor U21301 (N_21301,N_20580,N_20052);
nor U21302 (N_21302,N_20093,N_20144);
and U21303 (N_21303,N_20750,N_20118);
or U21304 (N_21304,N_20279,N_20000);
nor U21305 (N_21305,N_20111,N_20649);
nor U21306 (N_21306,N_20045,N_20806);
nor U21307 (N_21307,N_20281,N_20952);
xor U21308 (N_21308,N_20071,N_20271);
xnor U21309 (N_21309,N_20669,N_20815);
xor U21310 (N_21310,N_20877,N_20019);
and U21311 (N_21311,N_20781,N_20936);
nand U21312 (N_21312,N_20010,N_20566);
nor U21313 (N_21313,N_20754,N_20872);
nand U21314 (N_21314,N_20480,N_20853);
and U21315 (N_21315,N_20275,N_20582);
nor U21316 (N_21316,N_20073,N_20046);
nand U21317 (N_21317,N_20033,N_20051);
xnor U21318 (N_21318,N_20533,N_20956);
nand U21319 (N_21319,N_20655,N_20720);
or U21320 (N_21320,N_20289,N_20317);
nand U21321 (N_21321,N_20773,N_20954);
nand U21322 (N_21322,N_20455,N_20284);
or U21323 (N_21323,N_20925,N_20336);
and U21324 (N_21324,N_20770,N_20250);
nor U21325 (N_21325,N_20555,N_20427);
xor U21326 (N_21326,N_20121,N_20541);
nor U21327 (N_21327,N_20094,N_20904);
or U21328 (N_21328,N_20967,N_20293);
nand U21329 (N_21329,N_20821,N_20969);
xnor U21330 (N_21330,N_20622,N_20201);
and U21331 (N_21331,N_20205,N_20852);
and U21332 (N_21332,N_20534,N_20701);
nand U21333 (N_21333,N_20804,N_20751);
nand U21334 (N_21334,N_20382,N_20421);
or U21335 (N_21335,N_20447,N_20732);
or U21336 (N_21336,N_20927,N_20423);
and U21337 (N_21337,N_20747,N_20683);
nor U21338 (N_21338,N_20516,N_20405);
and U21339 (N_21339,N_20882,N_20170);
xnor U21340 (N_21340,N_20394,N_20788);
or U21341 (N_21341,N_20451,N_20793);
and U21342 (N_21342,N_20260,N_20268);
and U21343 (N_21343,N_20893,N_20191);
or U21344 (N_21344,N_20233,N_20526);
and U21345 (N_21345,N_20307,N_20373);
nand U21346 (N_21346,N_20212,N_20243);
nor U21347 (N_21347,N_20670,N_20097);
xnor U21348 (N_21348,N_20311,N_20020);
and U21349 (N_21349,N_20474,N_20431);
and U21350 (N_21350,N_20166,N_20638);
nand U21351 (N_21351,N_20127,N_20947);
or U21352 (N_21352,N_20857,N_20775);
nand U21353 (N_21353,N_20587,N_20856);
nand U21354 (N_21354,N_20107,N_20639);
or U21355 (N_21355,N_20758,N_20065);
nor U21356 (N_21356,N_20971,N_20262);
xnor U21357 (N_21357,N_20556,N_20863);
xor U21358 (N_21358,N_20430,N_20625);
or U21359 (N_21359,N_20940,N_20888);
or U21360 (N_21360,N_20678,N_20222);
and U21361 (N_21361,N_20035,N_20098);
nor U21362 (N_21362,N_20563,N_20004);
or U21363 (N_21363,N_20753,N_20042);
and U21364 (N_21364,N_20245,N_20403);
nor U21365 (N_21365,N_20841,N_20605);
and U21366 (N_21366,N_20415,N_20146);
xnor U21367 (N_21367,N_20313,N_20538);
or U21368 (N_21368,N_20479,N_20823);
nor U21369 (N_21369,N_20363,N_20692);
nand U21370 (N_21370,N_20196,N_20744);
nor U21371 (N_21371,N_20464,N_20584);
or U21372 (N_21372,N_20208,N_20776);
or U21373 (N_21373,N_20911,N_20124);
xnor U21374 (N_21374,N_20478,N_20642);
xor U21375 (N_21375,N_20760,N_20572);
and U21376 (N_21376,N_20588,N_20140);
xor U21377 (N_21377,N_20931,N_20165);
nand U21378 (N_21378,N_20717,N_20410);
nand U21379 (N_21379,N_20835,N_20658);
xnor U21380 (N_21380,N_20615,N_20813);
or U21381 (N_21381,N_20034,N_20315);
or U21382 (N_21382,N_20016,N_20964);
or U21383 (N_21383,N_20544,N_20377);
and U21384 (N_21384,N_20705,N_20119);
nor U21385 (N_21385,N_20088,N_20950);
xnor U21386 (N_21386,N_20785,N_20808);
xor U21387 (N_21387,N_20693,N_20662);
and U21388 (N_21388,N_20886,N_20854);
and U21389 (N_21389,N_20376,N_20684);
nand U21390 (N_21390,N_20332,N_20134);
or U21391 (N_21391,N_20665,N_20903);
nand U21392 (N_21392,N_20959,N_20759);
xor U21393 (N_21393,N_20715,N_20894);
xor U21394 (N_21394,N_20723,N_20627);
nor U21395 (N_21395,N_20633,N_20631);
and U21396 (N_21396,N_20595,N_20276);
xor U21397 (N_21397,N_20504,N_20154);
or U21398 (N_21398,N_20707,N_20826);
xor U21399 (N_21399,N_20845,N_20374);
xnor U21400 (N_21400,N_20485,N_20789);
nor U21401 (N_21401,N_20697,N_20490);
or U21402 (N_21402,N_20861,N_20355);
xnor U21403 (N_21403,N_20574,N_20765);
or U21404 (N_21404,N_20912,N_20365);
nor U21405 (N_21405,N_20001,N_20221);
xor U21406 (N_21406,N_20981,N_20141);
nor U21407 (N_21407,N_20446,N_20366);
or U21408 (N_21408,N_20199,N_20354);
and U21409 (N_21409,N_20242,N_20932);
nor U21410 (N_21410,N_20392,N_20652);
nor U21411 (N_21411,N_20060,N_20500);
xor U21412 (N_21412,N_20310,N_20946);
xnor U21413 (N_21413,N_20180,N_20989);
nand U21414 (N_21414,N_20620,N_20743);
nand U21415 (N_21415,N_20129,N_20790);
nor U21416 (N_21416,N_20679,N_20975);
and U21417 (N_21417,N_20985,N_20945);
xnor U21418 (N_21418,N_20048,N_20145);
nor U21419 (N_21419,N_20053,N_20116);
or U21420 (N_21420,N_20613,N_20577);
and U21421 (N_21421,N_20591,N_20929);
nand U21422 (N_21422,N_20218,N_20435);
or U21423 (N_21423,N_20078,N_20624);
nand U21424 (N_21424,N_20288,N_20612);
and U21425 (N_21425,N_20287,N_20881);
xnor U21426 (N_21426,N_20687,N_20072);
nor U21427 (N_21427,N_20926,N_20316);
or U21428 (N_21428,N_20309,N_20948);
xnor U21429 (N_21429,N_20148,N_20673);
and U21430 (N_21430,N_20924,N_20023);
and U21431 (N_21431,N_20868,N_20527);
or U21432 (N_21432,N_20560,N_20461);
and U21433 (N_21433,N_20722,N_20562);
or U21434 (N_21434,N_20593,N_20190);
nor U21435 (N_21435,N_20232,N_20173);
nand U21436 (N_21436,N_20472,N_20656);
nand U21437 (N_21437,N_20647,N_20061);
and U21438 (N_21438,N_20303,N_20814);
nor U21439 (N_21439,N_20278,N_20128);
nor U21440 (N_21440,N_20716,N_20167);
xnor U21441 (N_21441,N_20463,N_20112);
and U21442 (N_21442,N_20801,N_20664);
xor U21443 (N_21443,N_20115,N_20700);
xor U21444 (N_21444,N_20308,N_20074);
or U21445 (N_21445,N_20998,N_20711);
xor U21446 (N_21446,N_20525,N_20142);
nor U21447 (N_21447,N_20384,N_20840);
and U21448 (N_21448,N_20512,N_20007);
nand U21449 (N_21449,N_20536,N_20298);
nand U21450 (N_21450,N_20267,N_20440);
xnor U21451 (N_21451,N_20787,N_20168);
or U21452 (N_21452,N_20517,N_20603);
and U21453 (N_21453,N_20675,N_20030);
nand U21454 (N_21454,N_20186,N_20982);
nand U21455 (N_21455,N_20305,N_20347);
or U21456 (N_21456,N_20495,N_20866);
xor U21457 (N_21457,N_20018,N_20296);
nand U21458 (N_21458,N_20833,N_20024);
xnor U21459 (N_21459,N_20918,N_20935);
and U21460 (N_21460,N_20901,N_20235);
nand U21461 (N_21461,N_20496,N_20070);
and U21462 (N_21462,N_20498,N_20848);
nor U21463 (N_21463,N_20238,N_20657);
and U21464 (N_21464,N_20660,N_20706);
and U21465 (N_21465,N_20044,N_20210);
xor U21466 (N_21466,N_20091,N_20062);
and U21467 (N_21467,N_20352,N_20220);
nand U21468 (N_21468,N_20195,N_20838);
or U21469 (N_21469,N_20565,N_20274);
or U21470 (N_21470,N_20594,N_20892);
nor U21471 (N_21471,N_20252,N_20908);
and U21472 (N_21472,N_20013,N_20783);
and U21473 (N_21473,N_20084,N_20849);
or U21474 (N_21474,N_20458,N_20137);
or U21475 (N_21475,N_20178,N_20028);
nor U21476 (N_21476,N_20251,N_20604);
or U21477 (N_21477,N_20256,N_20322);
xnor U21478 (N_21478,N_20443,N_20397);
or U21479 (N_21479,N_20067,N_20241);
xnor U21480 (N_21480,N_20407,N_20483);
xor U21481 (N_21481,N_20452,N_20719);
nor U21482 (N_21482,N_20449,N_20774);
or U21483 (N_21483,N_20511,N_20150);
xnor U21484 (N_21484,N_20012,N_20333);
nand U21485 (N_21485,N_20488,N_20258);
or U21486 (N_21486,N_20350,N_20270);
xor U21487 (N_21487,N_20375,N_20328);
and U21488 (N_21488,N_20617,N_20666);
nor U21489 (N_21489,N_20172,N_20896);
nand U21490 (N_21490,N_20548,N_20611);
or U21491 (N_21491,N_20120,N_20429);
xnor U21492 (N_21492,N_20263,N_20674);
nor U21493 (N_21493,N_20545,N_20108);
nor U21494 (N_21494,N_20667,N_20457);
nand U21495 (N_21495,N_20820,N_20519);
and U21496 (N_21496,N_20105,N_20965);
or U21497 (N_21497,N_20014,N_20843);
nor U21498 (N_21498,N_20535,N_20837);
nand U21499 (N_21499,N_20385,N_20937);
and U21500 (N_21500,N_20826,N_20519);
nor U21501 (N_21501,N_20443,N_20456);
or U21502 (N_21502,N_20984,N_20451);
and U21503 (N_21503,N_20077,N_20881);
and U21504 (N_21504,N_20295,N_20592);
and U21505 (N_21505,N_20161,N_20202);
and U21506 (N_21506,N_20875,N_20149);
xnor U21507 (N_21507,N_20294,N_20387);
nand U21508 (N_21508,N_20793,N_20912);
nand U21509 (N_21509,N_20613,N_20705);
nor U21510 (N_21510,N_20706,N_20923);
nand U21511 (N_21511,N_20240,N_20671);
nor U21512 (N_21512,N_20376,N_20721);
or U21513 (N_21513,N_20398,N_20724);
or U21514 (N_21514,N_20849,N_20346);
nand U21515 (N_21515,N_20787,N_20696);
nand U21516 (N_21516,N_20904,N_20830);
or U21517 (N_21517,N_20910,N_20129);
nor U21518 (N_21518,N_20188,N_20535);
nand U21519 (N_21519,N_20700,N_20425);
nand U21520 (N_21520,N_20652,N_20864);
nand U21521 (N_21521,N_20422,N_20335);
or U21522 (N_21522,N_20533,N_20502);
or U21523 (N_21523,N_20184,N_20028);
or U21524 (N_21524,N_20755,N_20348);
nand U21525 (N_21525,N_20132,N_20341);
nor U21526 (N_21526,N_20863,N_20260);
nand U21527 (N_21527,N_20041,N_20135);
or U21528 (N_21528,N_20419,N_20671);
or U21529 (N_21529,N_20709,N_20716);
xor U21530 (N_21530,N_20183,N_20239);
and U21531 (N_21531,N_20189,N_20883);
xnor U21532 (N_21532,N_20742,N_20626);
nor U21533 (N_21533,N_20142,N_20287);
or U21534 (N_21534,N_20176,N_20849);
xor U21535 (N_21535,N_20881,N_20239);
nand U21536 (N_21536,N_20033,N_20923);
nor U21537 (N_21537,N_20435,N_20170);
and U21538 (N_21538,N_20335,N_20997);
and U21539 (N_21539,N_20416,N_20395);
and U21540 (N_21540,N_20813,N_20602);
xor U21541 (N_21541,N_20346,N_20638);
and U21542 (N_21542,N_20974,N_20133);
and U21543 (N_21543,N_20625,N_20618);
or U21544 (N_21544,N_20376,N_20124);
or U21545 (N_21545,N_20620,N_20532);
nand U21546 (N_21546,N_20095,N_20874);
xor U21547 (N_21547,N_20300,N_20093);
or U21548 (N_21548,N_20260,N_20243);
nor U21549 (N_21549,N_20900,N_20152);
and U21550 (N_21550,N_20984,N_20808);
and U21551 (N_21551,N_20633,N_20416);
nor U21552 (N_21552,N_20140,N_20258);
and U21553 (N_21553,N_20960,N_20622);
or U21554 (N_21554,N_20058,N_20503);
and U21555 (N_21555,N_20327,N_20247);
xor U21556 (N_21556,N_20446,N_20360);
and U21557 (N_21557,N_20061,N_20293);
or U21558 (N_21558,N_20002,N_20920);
and U21559 (N_21559,N_20083,N_20188);
and U21560 (N_21560,N_20378,N_20875);
nor U21561 (N_21561,N_20196,N_20872);
or U21562 (N_21562,N_20807,N_20376);
and U21563 (N_21563,N_20717,N_20738);
nor U21564 (N_21564,N_20226,N_20158);
nor U21565 (N_21565,N_20939,N_20047);
nand U21566 (N_21566,N_20656,N_20192);
nor U21567 (N_21567,N_20237,N_20600);
or U21568 (N_21568,N_20339,N_20374);
nor U21569 (N_21569,N_20627,N_20148);
and U21570 (N_21570,N_20026,N_20836);
and U21571 (N_21571,N_20596,N_20371);
or U21572 (N_21572,N_20717,N_20635);
xor U21573 (N_21573,N_20423,N_20526);
xor U21574 (N_21574,N_20405,N_20503);
xor U21575 (N_21575,N_20303,N_20768);
nor U21576 (N_21576,N_20001,N_20868);
xor U21577 (N_21577,N_20413,N_20651);
or U21578 (N_21578,N_20065,N_20332);
or U21579 (N_21579,N_20728,N_20606);
and U21580 (N_21580,N_20084,N_20068);
or U21581 (N_21581,N_20991,N_20840);
nand U21582 (N_21582,N_20371,N_20009);
nand U21583 (N_21583,N_20035,N_20181);
and U21584 (N_21584,N_20459,N_20439);
nand U21585 (N_21585,N_20057,N_20834);
nor U21586 (N_21586,N_20156,N_20222);
and U21587 (N_21587,N_20764,N_20433);
or U21588 (N_21588,N_20640,N_20354);
and U21589 (N_21589,N_20222,N_20423);
and U21590 (N_21590,N_20643,N_20900);
or U21591 (N_21591,N_20598,N_20759);
xor U21592 (N_21592,N_20918,N_20500);
or U21593 (N_21593,N_20450,N_20918);
xor U21594 (N_21594,N_20368,N_20059);
nor U21595 (N_21595,N_20725,N_20130);
or U21596 (N_21596,N_20876,N_20774);
nor U21597 (N_21597,N_20079,N_20102);
and U21598 (N_21598,N_20422,N_20751);
and U21599 (N_21599,N_20596,N_20357);
or U21600 (N_21600,N_20216,N_20540);
or U21601 (N_21601,N_20973,N_20503);
nand U21602 (N_21602,N_20111,N_20763);
xor U21603 (N_21603,N_20253,N_20287);
and U21604 (N_21604,N_20835,N_20640);
nand U21605 (N_21605,N_20917,N_20756);
and U21606 (N_21606,N_20472,N_20487);
and U21607 (N_21607,N_20586,N_20585);
nor U21608 (N_21608,N_20817,N_20060);
nor U21609 (N_21609,N_20451,N_20996);
nand U21610 (N_21610,N_20871,N_20620);
nor U21611 (N_21611,N_20112,N_20638);
xnor U21612 (N_21612,N_20444,N_20989);
nand U21613 (N_21613,N_20018,N_20130);
and U21614 (N_21614,N_20789,N_20542);
nor U21615 (N_21615,N_20164,N_20379);
nand U21616 (N_21616,N_20316,N_20426);
xor U21617 (N_21617,N_20803,N_20302);
or U21618 (N_21618,N_20137,N_20237);
xor U21619 (N_21619,N_20552,N_20632);
and U21620 (N_21620,N_20720,N_20852);
and U21621 (N_21621,N_20844,N_20684);
and U21622 (N_21622,N_20073,N_20627);
nor U21623 (N_21623,N_20294,N_20483);
nand U21624 (N_21624,N_20779,N_20427);
nand U21625 (N_21625,N_20493,N_20784);
nand U21626 (N_21626,N_20657,N_20720);
nand U21627 (N_21627,N_20617,N_20062);
nor U21628 (N_21628,N_20334,N_20110);
or U21629 (N_21629,N_20446,N_20939);
and U21630 (N_21630,N_20092,N_20080);
or U21631 (N_21631,N_20926,N_20972);
and U21632 (N_21632,N_20149,N_20677);
and U21633 (N_21633,N_20581,N_20056);
nor U21634 (N_21634,N_20075,N_20696);
or U21635 (N_21635,N_20384,N_20793);
and U21636 (N_21636,N_20850,N_20940);
or U21637 (N_21637,N_20231,N_20479);
nand U21638 (N_21638,N_20432,N_20837);
nor U21639 (N_21639,N_20283,N_20873);
xor U21640 (N_21640,N_20485,N_20610);
xnor U21641 (N_21641,N_20020,N_20864);
and U21642 (N_21642,N_20741,N_20739);
and U21643 (N_21643,N_20220,N_20426);
nor U21644 (N_21644,N_20765,N_20716);
and U21645 (N_21645,N_20289,N_20810);
xnor U21646 (N_21646,N_20567,N_20783);
xor U21647 (N_21647,N_20751,N_20826);
and U21648 (N_21648,N_20220,N_20171);
nand U21649 (N_21649,N_20393,N_20429);
or U21650 (N_21650,N_20104,N_20842);
or U21651 (N_21651,N_20471,N_20851);
and U21652 (N_21652,N_20567,N_20043);
or U21653 (N_21653,N_20771,N_20888);
nor U21654 (N_21654,N_20550,N_20564);
or U21655 (N_21655,N_20564,N_20327);
nand U21656 (N_21656,N_20349,N_20168);
xor U21657 (N_21657,N_20176,N_20299);
nand U21658 (N_21658,N_20021,N_20985);
nor U21659 (N_21659,N_20990,N_20525);
nand U21660 (N_21660,N_20499,N_20576);
and U21661 (N_21661,N_20960,N_20551);
nor U21662 (N_21662,N_20576,N_20494);
and U21663 (N_21663,N_20313,N_20091);
nor U21664 (N_21664,N_20016,N_20461);
and U21665 (N_21665,N_20473,N_20519);
nor U21666 (N_21666,N_20756,N_20876);
and U21667 (N_21667,N_20749,N_20386);
nor U21668 (N_21668,N_20689,N_20780);
nand U21669 (N_21669,N_20901,N_20139);
and U21670 (N_21670,N_20356,N_20466);
xnor U21671 (N_21671,N_20260,N_20635);
and U21672 (N_21672,N_20717,N_20959);
xor U21673 (N_21673,N_20644,N_20827);
or U21674 (N_21674,N_20096,N_20511);
nand U21675 (N_21675,N_20579,N_20882);
xnor U21676 (N_21676,N_20282,N_20557);
and U21677 (N_21677,N_20068,N_20971);
or U21678 (N_21678,N_20067,N_20172);
or U21679 (N_21679,N_20021,N_20278);
and U21680 (N_21680,N_20247,N_20481);
or U21681 (N_21681,N_20819,N_20074);
and U21682 (N_21682,N_20663,N_20508);
and U21683 (N_21683,N_20000,N_20934);
nor U21684 (N_21684,N_20222,N_20324);
or U21685 (N_21685,N_20046,N_20565);
or U21686 (N_21686,N_20791,N_20731);
nand U21687 (N_21687,N_20131,N_20663);
nand U21688 (N_21688,N_20648,N_20695);
nand U21689 (N_21689,N_20668,N_20263);
nor U21690 (N_21690,N_20773,N_20749);
nand U21691 (N_21691,N_20434,N_20667);
or U21692 (N_21692,N_20826,N_20571);
and U21693 (N_21693,N_20470,N_20652);
nand U21694 (N_21694,N_20674,N_20348);
nor U21695 (N_21695,N_20968,N_20756);
or U21696 (N_21696,N_20352,N_20418);
and U21697 (N_21697,N_20713,N_20663);
or U21698 (N_21698,N_20654,N_20022);
xor U21699 (N_21699,N_20520,N_20118);
xor U21700 (N_21700,N_20005,N_20223);
nor U21701 (N_21701,N_20069,N_20766);
nor U21702 (N_21702,N_20362,N_20604);
xor U21703 (N_21703,N_20405,N_20385);
or U21704 (N_21704,N_20874,N_20037);
or U21705 (N_21705,N_20410,N_20563);
and U21706 (N_21706,N_20232,N_20856);
or U21707 (N_21707,N_20067,N_20267);
xnor U21708 (N_21708,N_20284,N_20119);
and U21709 (N_21709,N_20634,N_20674);
xnor U21710 (N_21710,N_20940,N_20838);
and U21711 (N_21711,N_20788,N_20712);
nand U21712 (N_21712,N_20259,N_20952);
xnor U21713 (N_21713,N_20503,N_20231);
xor U21714 (N_21714,N_20747,N_20780);
xnor U21715 (N_21715,N_20960,N_20977);
and U21716 (N_21716,N_20105,N_20197);
nor U21717 (N_21717,N_20244,N_20257);
nand U21718 (N_21718,N_20444,N_20735);
and U21719 (N_21719,N_20407,N_20526);
nor U21720 (N_21720,N_20036,N_20121);
nor U21721 (N_21721,N_20453,N_20651);
or U21722 (N_21722,N_20718,N_20142);
and U21723 (N_21723,N_20806,N_20834);
nor U21724 (N_21724,N_20134,N_20382);
or U21725 (N_21725,N_20950,N_20139);
and U21726 (N_21726,N_20285,N_20709);
nand U21727 (N_21727,N_20576,N_20981);
or U21728 (N_21728,N_20374,N_20907);
nor U21729 (N_21729,N_20793,N_20945);
or U21730 (N_21730,N_20397,N_20481);
and U21731 (N_21731,N_20521,N_20420);
or U21732 (N_21732,N_20746,N_20004);
nand U21733 (N_21733,N_20114,N_20945);
or U21734 (N_21734,N_20849,N_20601);
and U21735 (N_21735,N_20571,N_20703);
and U21736 (N_21736,N_20322,N_20100);
or U21737 (N_21737,N_20788,N_20379);
xnor U21738 (N_21738,N_20376,N_20151);
or U21739 (N_21739,N_20725,N_20995);
xnor U21740 (N_21740,N_20989,N_20577);
and U21741 (N_21741,N_20879,N_20827);
and U21742 (N_21742,N_20385,N_20451);
xor U21743 (N_21743,N_20222,N_20503);
nor U21744 (N_21744,N_20959,N_20732);
nor U21745 (N_21745,N_20804,N_20726);
or U21746 (N_21746,N_20445,N_20215);
xnor U21747 (N_21747,N_20158,N_20402);
and U21748 (N_21748,N_20421,N_20987);
and U21749 (N_21749,N_20133,N_20147);
nor U21750 (N_21750,N_20318,N_20171);
or U21751 (N_21751,N_20903,N_20238);
or U21752 (N_21752,N_20592,N_20947);
xnor U21753 (N_21753,N_20700,N_20798);
nor U21754 (N_21754,N_20095,N_20204);
xnor U21755 (N_21755,N_20388,N_20854);
and U21756 (N_21756,N_20305,N_20820);
and U21757 (N_21757,N_20480,N_20628);
nor U21758 (N_21758,N_20908,N_20911);
xnor U21759 (N_21759,N_20381,N_20619);
nand U21760 (N_21760,N_20955,N_20339);
nand U21761 (N_21761,N_20181,N_20917);
nand U21762 (N_21762,N_20102,N_20839);
or U21763 (N_21763,N_20795,N_20871);
or U21764 (N_21764,N_20173,N_20031);
or U21765 (N_21765,N_20655,N_20044);
and U21766 (N_21766,N_20557,N_20159);
and U21767 (N_21767,N_20955,N_20493);
and U21768 (N_21768,N_20326,N_20208);
and U21769 (N_21769,N_20540,N_20886);
nor U21770 (N_21770,N_20759,N_20512);
xor U21771 (N_21771,N_20420,N_20498);
xnor U21772 (N_21772,N_20153,N_20485);
xnor U21773 (N_21773,N_20639,N_20415);
xor U21774 (N_21774,N_20264,N_20218);
nor U21775 (N_21775,N_20815,N_20671);
nor U21776 (N_21776,N_20983,N_20595);
xor U21777 (N_21777,N_20206,N_20905);
and U21778 (N_21778,N_20131,N_20769);
or U21779 (N_21779,N_20520,N_20513);
xor U21780 (N_21780,N_20813,N_20305);
nand U21781 (N_21781,N_20239,N_20887);
and U21782 (N_21782,N_20247,N_20872);
xor U21783 (N_21783,N_20926,N_20352);
nand U21784 (N_21784,N_20929,N_20072);
nand U21785 (N_21785,N_20760,N_20515);
nor U21786 (N_21786,N_20673,N_20873);
nor U21787 (N_21787,N_20788,N_20192);
and U21788 (N_21788,N_20048,N_20310);
nand U21789 (N_21789,N_20112,N_20375);
or U21790 (N_21790,N_20302,N_20493);
xnor U21791 (N_21791,N_20408,N_20757);
nor U21792 (N_21792,N_20525,N_20217);
or U21793 (N_21793,N_20915,N_20158);
xnor U21794 (N_21794,N_20373,N_20414);
and U21795 (N_21795,N_20791,N_20199);
and U21796 (N_21796,N_20925,N_20546);
or U21797 (N_21797,N_20699,N_20628);
nor U21798 (N_21798,N_20683,N_20266);
nor U21799 (N_21799,N_20072,N_20875);
or U21800 (N_21800,N_20098,N_20197);
nand U21801 (N_21801,N_20502,N_20723);
and U21802 (N_21802,N_20828,N_20589);
nor U21803 (N_21803,N_20556,N_20225);
and U21804 (N_21804,N_20376,N_20330);
nand U21805 (N_21805,N_20136,N_20386);
nand U21806 (N_21806,N_20634,N_20131);
or U21807 (N_21807,N_20852,N_20040);
xor U21808 (N_21808,N_20145,N_20512);
and U21809 (N_21809,N_20398,N_20686);
nor U21810 (N_21810,N_20207,N_20593);
nand U21811 (N_21811,N_20210,N_20337);
and U21812 (N_21812,N_20948,N_20739);
xor U21813 (N_21813,N_20474,N_20477);
nor U21814 (N_21814,N_20015,N_20127);
or U21815 (N_21815,N_20718,N_20696);
xnor U21816 (N_21816,N_20119,N_20289);
xnor U21817 (N_21817,N_20154,N_20995);
nand U21818 (N_21818,N_20112,N_20236);
nand U21819 (N_21819,N_20433,N_20196);
nand U21820 (N_21820,N_20747,N_20920);
xor U21821 (N_21821,N_20569,N_20267);
nand U21822 (N_21822,N_20756,N_20717);
or U21823 (N_21823,N_20716,N_20920);
xnor U21824 (N_21824,N_20334,N_20822);
xor U21825 (N_21825,N_20233,N_20707);
nand U21826 (N_21826,N_20220,N_20294);
nor U21827 (N_21827,N_20308,N_20608);
and U21828 (N_21828,N_20089,N_20056);
xnor U21829 (N_21829,N_20924,N_20452);
xor U21830 (N_21830,N_20722,N_20474);
or U21831 (N_21831,N_20893,N_20842);
and U21832 (N_21832,N_20243,N_20482);
nand U21833 (N_21833,N_20669,N_20274);
nor U21834 (N_21834,N_20619,N_20836);
and U21835 (N_21835,N_20109,N_20930);
and U21836 (N_21836,N_20458,N_20525);
nor U21837 (N_21837,N_20006,N_20754);
or U21838 (N_21838,N_20440,N_20620);
nand U21839 (N_21839,N_20783,N_20951);
and U21840 (N_21840,N_20987,N_20247);
and U21841 (N_21841,N_20809,N_20595);
nand U21842 (N_21842,N_20824,N_20616);
and U21843 (N_21843,N_20929,N_20220);
or U21844 (N_21844,N_20968,N_20969);
and U21845 (N_21845,N_20237,N_20994);
or U21846 (N_21846,N_20209,N_20773);
and U21847 (N_21847,N_20229,N_20260);
nand U21848 (N_21848,N_20611,N_20967);
nand U21849 (N_21849,N_20824,N_20002);
xor U21850 (N_21850,N_20754,N_20258);
nand U21851 (N_21851,N_20364,N_20719);
and U21852 (N_21852,N_20507,N_20487);
and U21853 (N_21853,N_20939,N_20273);
nor U21854 (N_21854,N_20078,N_20337);
and U21855 (N_21855,N_20650,N_20133);
or U21856 (N_21856,N_20810,N_20445);
or U21857 (N_21857,N_20630,N_20263);
or U21858 (N_21858,N_20568,N_20418);
or U21859 (N_21859,N_20178,N_20743);
nor U21860 (N_21860,N_20549,N_20588);
and U21861 (N_21861,N_20569,N_20487);
xor U21862 (N_21862,N_20371,N_20702);
xor U21863 (N_21863,N_20928,N_20005);
xnor U21864 (N_21864,N_20326,N_20956);
xnor U21865 (N_21865,N_20208,N_20911);
nor U21866 (N_21866,N_20494,N_20694);
nand U21867 (N_21867,N_20246,N_20297);
and U21868 (N_21868,N_20774,N_20566);
and U21869 (N_21869,N_20579,N_20565);
nor U21870 (N_21870,N_20979,N_20175);
nor U21871 (N_21871,N_20504,N_20824);
nor U21872 (N_21872,N_20357,N_20774);
and U21873 (N_21873,N_20688,N_20135);
nand U21874 (N_21874,N_20660,N_20166);
or U21875 (N_21875,N_20759,N_20719);
xor U21876 (N_21876,N_20535,N_20468);
nand U21877 (N_21877,N_20767,N_20532);
or U21878 (N_21878,N_20946,N_20707);
xnor U21879 (N_21879,N_20588,N_20225);
and U21880 (N_21880,N_20510,N_20486);
and U21881 (N_21881,N_20007,N_20735);
xnor U21882 (N_21882,N_20976,N_20393);
nand U21883 (N_21883,N_20241,N_20598);
nor U21884 (N_21884,N_20572,N_20162);
and U21885 (N_21885,N_20582,N_20903);
nor U21886 (N_21886,N_20750,N_20101);
and U21887 (N_21887,N_20440,N_20637);
nand U21888 (N_21888,N_20188,N_20497);
nor U21889 (N_21889,N_20117,N_20533);
nor U21890 (N_21890,N_20426,N_20530);
xor U21891 (N_21891,N_20594,N_20260);
nand U21892 (N_21892,N_20062,N_20059);
nor U21893 (N_21893,N_20329,N_20506);
or U21894 (N_21894,N_20245,N_20038);
and U21895 (N_21895,N_20568,N_20273);
nand U21896 (N_21896,N_20888,N_20730);
xnor U21897 (N_21897,N_20757,N_20350);
nand U21898 (N_21898,N_20058,N_20659);
or U21899 (N_21899,N_20769,N_20913);
nor U21900 (N_21900,N_20656,N_20784);
and U21901 (N_21901,N_20475,N_20673);
and U21902 (N_21902,N_20524,N_20059);
and U21903 (N_21903,N_20290,N_20461);
and U21904 (N_21904,N_20679,N_20104);
and U21905 (N_21905,N_20258,N_20687);
or U21906 (N_21906,N_20315,N_20280);
and U21907 (N_21907,N_20698,N_20625);
xnor U21908 (N_21908,N_20543,N_20207);
xnor U21909 (N_21909,N_20292,N_20212);
and U21910 (N_21910,N_20792,N_20040);
nor U21911 (N_21911,N_20527,N_20978);
xor U21912 (N_21912,N_20896,N_20161);
xor U21913 (N_21913,N_20868,N_20451);
and U21914 (N_21914,N_20734,N_20869);
nor U21915 (N_21915,N_20138,N_20303);
nand U21916 (N_21916,N_20878,N_20418);
or U21917 (N_21917,N_20493,N_20809);
nor U21918 (N_21918,N_20756,N_20958);
nor U21919 (N_21919,N_20819,N_20473);
xnor U21920 (N_21920,N_20839,N_20579);
nand U21921 (N_21921,N_20711,N_20041);
and U21922 (N_21922,N_20861,N_20308);
nand U21923 (N_21923,N_20021,N_20998);
xor U21924 (N_21924,N_20279,N_20723);
and U21925 (N_21925,N_20634,N_20306);
or U21926 (N_21926,N_20535,N_20746);
or U21927 (N_21927,N_20593,N_20630);
nor U21928 (N_21928,N_20962,N_20570);
nand U21929 (N_21929,N_20568,N_20654);
or U21930 (N_21930,N_20376,N_20348);
nor U21931 (N_21931,N_20642,N_20468);
nand U21932 (N_21932,N_20331,N_20890);
nor U21933 (N_21933,N_20714,N_20111);
and U21934 (N_21934,N_20268,N_20423);
nand U21935 (N_21935,N_20321,N_20200);
and U21936 (N_21936,N_20188,N_20715);
and U21937 (N_21937,N_20427,N_20061);
or U21938 (N_21938,N_20097,N_20908);
xor U21939 (N_21939,N_20876,N_20248);
nand U21940 (N_21940,N_20601,N_20722);
nor U21941 (N_21941,N_20355,N_20110);
and U21942 (N_21942,N_20773,N_20589);
nor U21943 (N_21943,N_20407,N_20372);
xnor U21944 (N_21944,N_20901,N_20851);
xor U21945 (N_21945,N_20458,N_20251);
xor U21946 (N_21946,N_20069,N_20924);
xor U21947 (N_21947,N_20304,N_20015);
nor U21948 (N_21948,N_20390,N_20647);
or U21949 (N_21949,N_20673,N_20689);
or U21950 (N_21950,N_20245,N_20630);
or U21951 (N_21951,N_20515,N_20721);
nand U21952 (N_21952,N_20118,N_20543);
nand U21953 (N_21953,N_20524,N_20073);
nand U21954 (N_21954,N_20871,N_20294);
nor U21955 (N_21955,N_20653,N_20210);
nor U21956 (N_21956,N_20412,N_20540);
xnor U21957 (N_21957,N_20680,N_20255);
nor U21958 (N_21958,N_20450,N_20469);
xor U21959 (N_21959,N_20717,N_20218);
and U21960 (N_21960,N_20951,N_20958);
xor U21961 (N_21961,N_20109,N_20622);
or U21962 (N_21962,N_20726,N_20189);
nor U21963 (N_21963,N_20690,N_20370);
and U21964 (N_21964,N_20170,N_20775);
or U21965 (N_21965,N_20289,N_20086);
and U21966 (N_21966,N_20047,N_20322);
nand U21967 (N_21967,N_20684,N_20478);
or U21968 (N_21968,N_20401,N_20636);
or U21969 (N_21969,N_20025,N_20672);
and U21970 (N_21970,N_20520,N_20991);
nor U21971 (N_21971,N_20916,N_20856);
nor U21972 (N_21972,N_20194,N_20666);
nand U21973 (N_21973,N_20939,N_20179);
nand U21974 (N_21974,N_20185,N_20784);
and U21975 (N_21975,N_20204,N_20230);
nand U21976 (N_21976,N_20031,N_20276);
and U21977 (N_21977,N_20419,N_20606);
xor U21978 (N_21978,N_20751,N_20310);
or U21979 (N_21979,N_20589,N_20945);
nand U21980 (N_21980,N_20636,N_20881);
nand U21981 (N_21981,N_20729,N_20646);
or U21982 (N_21982,N_20889,N_20406);
nand U21983 (N_21983,N_20801,N_20335);
nor U21984 (N_21984,N_20453,N_20765);
xor U21985 (N_21985,N_20217,N_20066);
nor U21986 (N_21986,N_20509,N_20603);
nand U21987 (N_21987,N_20525,N_20047);
nor U21988 (N_21988,N_20970,N_20069);
and U21989 (N_21989,N_20518,N_20359);
xor U21990 (N_21990,N_20796,N_20966);
and U21991 (N_21991,N_20720,N_20548);
and U21992 (N_21992,N_20396,N_20231);
nand U21993 (N_21993,N_20080,N_20437);
nor U21994 (N_21994,N_20300,N_20685);
nor U21995 (N_21995,N_20155,N_20051);
and U21996 (N_21996,N_20968,N_20464);
nor U21997 (N_21997,N_20516,N_20613);
and U21998 (N_21998,N_20690,N_20029);
nor U21999 (N_21999,N_20194,N_20371);
nor U22000 (N_22000,N_21675,N_21846);
or U22001 (N_22001,N_21439,N_21040);
and U22002 (N_22002,N_21505,N_21274);
and U22003 (N_22003,N_21001,N_21171);
or U22004 (N_22004,N_21487,N_21698);
or U22005 (N_22005,N_21045,N_21112);
xor U22006 (N_22006,N_21773,N_21015);
xor U22007 (N_22007,N_21780,N_21845);
nand U22008 (N_22008,N_21939,N_21399);
and U22009 (N_22009,N_21166,N_21793);
nand U22010 (N_22010,N_21071,N_21096);
nand U22011 (N_22011,N_21438,N_21530);
or U22012 (N_22012,N_21694,N_21479);
and U22013 (N_22013,N_21336,N_21656);
xor U22014 (N_22014,N_21492,N_21197);
xor U22015 (N_22015,N_21172,N_21629);
nor U22016 (N_22016,N_21127,N_21181);
nand U22017 (N_22017,N_21450,N_21951);
nand U22018 (N_22018,N_21499,N_21791);
and U22019 (N_22019,N_21583,N_21103);
or U22020 (N_22020,N_21122,N_21940);
nand U22021 (N_22021,N_21260,N_21580);
nand U22022 (N_22022,N_21763,N_21282);
nor U22023 (N_22023,N_21707,N_21472);
nor U22024 (N_22024,N_21524,N_21387);
nor U22025 (N_22025,N_21866,N_21292);
nand U22026 (N_22026,N_21135,N_21139);
or U22027 (N_22027,N_21605,N_21140);
nor U22028 (N_22028,N_21111,N_21288);
nor U22029 (N_22029,N_21654,N_21434);
nor U22030 (N_22030,N_21736,N_21988);
or U22031 (N_22031,N_21941,N_21596);
or U22032 (N_22032,N_21851,N_21673);
or U22033 (N_22033,N_21618,N_21099);
nor U22034 (N_22034,N_21690,N_21655);
and U22035 (N_22035,N_21235,N_21076);
xnor U22036 (N_22036,N_21073,N_21848);
or U22037 (N_22037,N_21511,N_21170);
nand U22038 (N_22038,N_21781,N_21083);
and U22039 (N_22039,N_21110,N_21987);
nand U22040 (N_22040,N_21386,N_21131);
xnor U22041 (N_22041,N_21755,N_21760);
and U22042 (N_22042,N_21508,N_21588);
nor U22043 (N_22043,N_21327,N_21027);
and U22044 (N_22044,N_21776,N_21869);
or U22045 (N_22045,N_21921,N_21772);
nand U22046 (N_22046,N_21735,N_21569);
xnor U22047 (N_22047,N_21651,N_21306);
nand U22048 (N_22048,N_21341,N_21196);
nor U22049 (N_22049,N_21899,N_21437);
and U22050 (N_22050,N_21979,N_21631);
nor U22051 (N_22051,N_21446,N_21659);
and U22052 (N_22052,N_21897,N_21565);
nand U22053 (N_22053,N_21035,N_21346);
nor U22054 (N_22054,N_21643,N_21182);
or U22055 (N_22055,N_21396,N_21029);
and U22056 (N_22056,N_21345,N_21089);
nor U22057 (N_22057,N_21177,N_21774);
or U22058 (N_22058,N_21075,N_21902);
nor U22059 (N_22059,N_21679,N_21536);
or U22060 (N_22060,N_21610,N_21849);
nor U22061 (N_22061,N_21217,N_21710);
or U22062 (N_22062,N_21000,N_21882);
or U22063 (N_22063,N_21028,N_21555);
nand U22064 (N_22064,N_21312,N_21350);
and U22065 (N_22065,N_21043,N_21115);
or U22066 (N_22066,N_21668,N_21372);
xnor U22067 (N_22067,N_21400,N_21314);
nor U22068 (N_22068,N_21389,N_21276);
nor U22069 (N_22069,N_21244,N_21435);
nor U22070 (N_22070,N_21955,N_21245);
nor U22071 (N_22071,N_21861,N_21480);
and U22072 (N_22072,N_21687,N_21008);
xor U22073 (N_22073,N_21419,N_21982);
and U22074 (N_22074,N_21486,N_21325);
and U22075 (N_22075,N_21607,N_21381);
nor U22076 (N_22076,N_21191,N_21677);
xor U22077 (N_22077,N_21534,N_21506);
or U22078 (N_22078,N_21599,N_21269);
or U22079 (N_22079,N_21151,N_21092);
nor U22080 (N_22080,N_21459,N_21440);
or U22081 (N_22081,N_21612,N_21875);
or U22082 (N_22082,N_21109,N_21616);
and U22083 (N_22083,N_21176,N_21717);
xor U22084 (N_22084,N_21259,N_21783);
and U22085 (N_22085,N_21187,N_21518);
or U22086 (N_22086,N_21761,N_21832);
xnor U22087 (N_22087,N_21806,N_21165);
nor U22088 (N_22088,N_21792,N_21582);
nand U22089 (N_22089,N_21065,N_21989);
nor U22090 (N_22090,N_21398,N_21746);
nor U22091 (N_22091,N_21994,N_21993);
xnor U22092 (N_22092,N_21408,N_21658);
nand U22093 (N_22093,N_21461,N_21041);
nand U22094 (N_22094,N_21595,N_21403);
or U22095 (N_22095,N_21887,N_21404);
or U22096 (N_22096,N_21578,N_21996);
and U22097 (N_22097,N_21558,N_21681);
xnor U22098 (N_22098,N_21978,N_21749);
xor U22099 (N_22099,N_21753,N_21010);
or U22100 (N_22100,N_21265,N_21817);
and U22101 (N_22101,N_21488,N_21369);
or U22102 (N_22102,N_21741,N_21152);
nor U22103 (N_22103,N_21708,N_21415);
and U22104 (N_22104,N_21652,N_21380);
and U22105 (N_22105,N_21744,N_21729);
nor U22106 (N_22106,N_21669,N_21934);
nor U22107 (N_22107,N_21769,N_21337);
or U22108 (N_22108,N_21591,N_21164);
nand U22109 (N_22109,N_21782,N_21912);
or U22110 (N_22110,N_21964,N_21302);
nand U22111 (N_22111,N_21348,N_21986);
or U22112 (N_22112,N_21237,N_21836);
nand U22113 (N_22113,N_21295,N_21917);
and U22114 (N_22114,N_21329,N_21503);
or U22115 (N_22115,N_21367,N_21999);
xnor U22116 (N_22116,N_21830,N_21764);
and U22117 (N_22117,N_21829,N_21750);
nor U22118 (N_22118,N_21309,N_21064);
nor U22119 (N_22119,N_21990,N_21510);
or U22120 (N_22120,N_21824,N_21891);
xnor U22121 (N_22121,N_21491,N_21128);
or U22122 (N_22122,N_21519,N_21406);
nor U22123 (N_22123,N_21250,N_21856);
or U22124 (N_22124,N_21920,N_21020);
or U22125 (N_22125,N_21330,N_21827);
or U22126 (N_22126,N_21107,N_21393);
and U22127 (N_22127,N_21496,N_21739);
nor U22128 (N_22128,N_21003,N_21294);
nand U22129 (N_22129,N_21664,N_21696);
or U22130 (N_22130,N_21077,N_21141);
nor U22131 (N_22131,N_21428,N_21397);
nor U22132 (N_22132,N_21030,N_21971);
nor U22133 (N_22133,N_21215,N_21590);
and U22134 (N_22134,N_21100,N_21357);
or U22135 (N_22135,N_21087,N_21896);
and U22136 (N_22136,N_21870,N_21258);
and U22137 (N_22137,N_21156,N_21860);
nand U22138 (N_22138,N_21786,N_21721);
nand U22139 (N_22139,N_21624,N_21936);
or U22140 (N_22140,N_21837,N_21044);
and U22141 (N_22141,N_21646,N_21497);
nor U22142 (N_22142,N_21208,N_21078);
or U22143 (N_22143,N_21642,N_21974);
nand U22144 (N_22144,N_21037,N_21561);
nand U22145 (N_22145,N_21207,N_21129);
nand U22146 (N_22146,N_21961,N_21431);
and U22147 (N_22147,N_21150,N_21685);
or U22148 (N_22148,N_21731,N_21401);
xor U22149 (N_22149,N_21012,N_21257);
nor U22150 (N_22150,N_21952,N_21105);
nor U22151 (N_22151,N_21737,N_21771);
or U22152 (N_22152,N_21745,N_21353);
nor U22153 (N_22153,N_21262,N_21678);
xor U22154 (N_22154,N_21185,N_21436);
and U22155 (N_22155,N_21085,N_21533);
and U22156 (N_22156,N_21236,N_21615);
or U22157 (N_22157,N_21038,N_21842);
and U22158 (N_22158,N_21362,N_21918);
or U22159 (N_22159,N_21722,N_21323);
and U22160 (N_22160,N_21444,N_21297);
xor U22161 (N_22161,N_21514,N_21416);
or U22162 (N_22162,N_21844,N_21680);
xor U22163 (N_22163,N_21532,N_21219);
nand U22164 (N_22164,N_21058,N_21812);
nand U22165 (N_22165,N_21512,N_21146);
xor U22166 (N_22166,N_21481,N_21351);
nor U22167 (N_22167,N_21700,N_21720);
xnor U22168 (N_22168,N_21602,N_21756);
or U22169 (N_22169,N_21795,N_21452);
or U22170 (N_22170,N_21432,N_21854);
nor U22171 (N_22171,N_21959,N_21732);
and U22172 (N_22172,N_21914,N_21116);
nor U22173 (N_22173,N_21778,N_21877);
nor U22174 (N_22174,N_21104,N_21084);
and U22175 (N_22175,N_21332,N_21826);
nand U22176 (N_22176,N_21925,N_21815);
nand U22177 (N_22177,N_21467,N_21261);
nor U22178 (N_22178,N_21963,N_21334);
and U22179 (N_22179,N_21883,N_21935);
or U22180 (N_22180,N_21178,N_21402);
xor U22181 (N_22181,N_21671,N_21316);
or U22182 (N_22182,N_21859,N_21888);
xnor U22183 (N_22183,N_21466,N_21930);
or U22184 (N_22184,N_21377,N_21242);
nor U22185 (N_22185,N_21821,N_21210);
nor U22186 (N_22186,N_21388,N_21179);
or U22187 (N_22187,N_21047,N_21560);
xor U22188 (N_22188,N_21313,N_21973);
or U22189 (N_22189,N_21825,N_21807);
nand U22190 (N_22190,N_21944,N_21095);
xnor U22191 (N_22191,N_21320,N_21279);
or U22192 (N_22192,N_21800,N_21447);
nand U22193 (N_22193,N_21238,N_21291);
nand U22194 (N_22194,N_21338,N_21828);
or U22195 (N_22195,N_21442,N_21542);
nor U22196 (N_22196,N_21123,N_21418);
and U22197 (N_22197,N_21661,N_21233);
nand U22198 (N_22198,N_21991,N_21395);
nand U22199 (N_22199,N_21133,N_21190);
or U22200 (N_22200,N_21676,N_21992);
nor U22201 (N_22201,N_21886,N_21688);
and U22202 (N_22202,N_21553,N_21335);
nand U22203 (N_22203,N_21706,N_21305);
and U22204 (N_22204,N_21134,N_21547);
and U22205 (N_22205,N_21649,N_21384);
nor U22206 (N_22206,N_21787,N_21169);
nand U22207 (N_22207,N_21541,N_21522);
nand U22208 (N_22208,N_21019,N_21922);
and U22209 (N_22209,N_21342,N_21412);
nor U22210 (N_22210,N_21173,N_21153);
and U22211 (N_22211,N_21862,N_21251);
nand U22212 (N_22212,N_21834,N_21485);
nor U22213 (N_22213,N_21878,N_21392);
or U22214 (N_22214,N_21718,N_21711);
and U22215 (N_22215,N_21249,N_21716);
and U22216 (N_22216,N_21502,N_21748);
or U22217 (N_22217,N_21509,N_21126);
nand U22218 (N_22218,N_21998,N_21570);
or U22219 (N_22219,N_21052,N_21034);
or U22220 (N_22220,N_21378,N_21876);
nand U22221 (N_22221,N_21319,N_21523);
or U22222 (N_22222,N_21638,N_21119);
nand U22223 (N_22223,N_21976,N_21552);
nor U22224 (N_22224,N_21054,N_21841);
xor U22225 (N_22225,N_21200,N_21026);
nand U22226 (N_22226,N_21080,N_21061);
nor U22227 (N_22227,N_21589,N_21670);
nand U22228 (N_22228,N_21660,N_21630);
or U22229 (N_22229,N_21002,N_21637);
nand U22230 (N_22230,N_21229,N_21429);
xor U22231 (N_22231,N_21548,N_21082);
or U22232 (N_22232,N_21268,N_21189);
nand U22233 (N_22233,N_21333,N_21066);
and U22234 (N_22234,N_21241,N_21593);
nor U22235 (N_22235,N_21243,N_21340);
and U22236 (N_22236,N_21234,N_21374);
nor U22237 (N_22237,N_21222,N_21929);
or U22238 (N_22238,N_21136,N_21867);
and U22239 (N_22239,N_21407,N_21443);
nor U22240 (N_22240,N_21206,N_21873);
xnor U22241 (N_22241,N_21551,N_21254);
or U22242 (N_22242,N_21013,N_21183);
xnor U22243 (N_22243,N_21272,N_21231);
nand U22244 (N_22244,N_21193,N_21872);
nand U22245 (N_22245,N_21120,N_21124);
nand U22246 (N_22246,N_21451,N_21995);
xor U22247 (N_22247,N_21881,N_21009);
nor U22248 (N_22248,N_21470,N_21142);
or U22249 (N_22249,N_21476,N_21725);
xor U22250 (N_22250,N_21747,N_21069);
nand U22251 (N_22251,N_21050,N_21603);
or U22252 (N_22252,N_21892,N_21803);
nand U22253 (N_22253,N_21568,N_21409);
or U22254 (N_22254,N_21211,N_21063);
nor U22255 (N_22255,N_21563,N_21529);
nor U22256 (N_22256,N_21703,N_21927);
xor U22257 (N_22257,N_21537,N_21702);
xnor U22258 (N_22258,N_21705,N_21811);
xnor U22259 (N_22259,N_21263,N_21494);
xor U22260 (N_22260,N_21360,N_21521);
xor U22261 (N_22261,N_21714,N_21890);
nand U22262 (N_22262,N_21566,N_21347);
nand U22263 (N_22263,N_21801,N_21853);
and U22264 (N_22264,N_21454,N_21311);
xor U22265 (N_22265,N_21144,N_21449);
xor U22266 (N_22266,N_21425,N_21363);
xnor U22267 (N_22267,N_21619,N_21007);
xor U22268 (N_22268,N_21754,N_21270);
and U22269 (N_22269,N_21657,N_21898);
xnor U22270 (N_22270,N_21928,N_21535);
nand U22271 (N_22271,N_21933,N_21184);
xor U22272 (N_22272,N_21086,N_21067);
nor U22273 (N_22273,N_21108,N_21445);
or U22274 (N_22274,N_21968,N_21515);
xor U22275 (N_22275,N_21430,N_21816);
or U22276 (N_22276,N_21271,N_21545);
and U22277 (N_22277,N_21813,N_21018);
or U22278 (N_22278,N_21255,N_21352);
xnor U22279 (N_22279,N_21025,N_21919);
or U22280 (N_22280,N_21033,N_21125);
nand U22281 (N_22281,N_21275,N_21885);
xor U22282 (N_22282,N_21477,N_21611);
nor U22283 (N_22283,N_21057,N_21321);
xor U22284 (N_22284,N_21022,N_21868);
nand U22285 (N_22285,N_21056,N_21239);
or U22286 (N_22286,N_21493,N_21613);
nor U22287 (N_22287,N_21132,N_21594);
xor U22288 (N_22288,N_21137,N_21463);
nor U22289 (N_22289,N_21500,N_21473);
and U22290 (N_22290,N_21310,N_21525);
or U22291 (N_22291,N_21517,N_21383);
xnor U22292 (N_22292,N_21884,N_21970);
nand U22293 (N_22293,N_21354,N_21820);
xor U22294 (N_22294,N_21223,N_21574);
nor U22295 (N_22295,N_21055,N_21364);
or U22296 (N_22296,N_21953,N_21647);
nor U22297 (N_22297,N_21550,N_21621);
nand U22298 (N_22298,N_21201,N_21068);
xnor U22299 (N_22299,N_21290,N_21556);
nand U22300 (N_22300,N_21549,N_21118);
or U22301 (N_22301,N_21584,N_21960);
xnor U22302 (N_22302,N_21014,N_21411);
nand U22303 (N_22303,N_21424,N_21130);
and U22304 (N_22304,N_21833,N_21228);
nand U22305 (N_22305,N_21088,N_21328);
nor U22306 (N_22306,N_21915,N_21965);
nor U22307 (N_22307,N_21246,N_21874);
xnor U22308 (N_22308,N_21462,N_21909);
nor U22309 (N_22309,N_21983,N_21916);
and U22310 (N_22310,N_21997,N_21726);
and U22311 (N_22311,N_21048,N_21662);
xor U22312 (N_22312,N_21689,N_21375);
xor U22313 (N_22313,N_21723,N_21650);
or U22314 (N_22314,N_21379,N_21391);
and U22315 (N_22315,N_21728,N_21456);
xnor U22316 (N_22316,N_21053,N_21091);
or U22317 (N_22317,N_21453,N_21768);
xnor U22318 (N_22318,N_21847,N_21592);
or U22319 (N_22319,N_21543,N_21984);
xor U22320 (N_22320,N_21648,N_21980);
and U22321 (N_22321,N_21317,N_21031);
and U22322 (N_22322,N_21214,N_21281);
nand U22323 (N_22323,N_21308,N_21942);
or U22324 (N_22324,N_21796,N_21343);
and U22325 (N_22325,N_21893,N_21004);
nand U22326 (N_22326,N_21232,N_21433);
or U22327 (N_22327,N_21490,N_21526);
and U22328 (N_22328,N_21699,N_21098);
or U22329 (N_22329,N_21913,N_21017);
nand U22330 (N_22330,N_21175,N_21021);
nor U22331 (N_22331,N_21704,N_21759);
and U22332 (N_22332,N_21455,N_21609);
or U22333 (N_22333,N_21385,N_21641);
nand U22334 (N_22334,N_21969,N_21839);
xor U22335 (N_22335,N_21474,N_21938);
nor U22336 (N_22336,N_21572,N_21227);
nor U22337 (N_22337,N_21784,N_21168);
nand U22338 (N_22338,N_21005,N_21831);
nand U22339 (N_22339,N_21417,N_21225);
nand U22340 (N_22340,N_21079,N_21911);
and U22341 (N_22341,N_21620,N_21538);
nor U22342 (N_22342,N_21039,N_21743);
and U22343 (N_22343,N_21159,N_21908);
nor U22344 (N_22344,N_21220,N_21252);
xor U22345 (N_22345,N_21213,N_21838);
and U22346 (N_22346,N_21701,N_21684);
and U22347 (N_22347,N_21149,N_21577);
nand U22348 (N_22348,N_21634,N_21958);
nand U22349 (N_22349,N_21709,N_21036);
and U22350 (N_22350,N_21777,N_21966);
and U22351 (N_22351,N_21757,N_21277);
nor U22352 (N_22352,N_21427,N_21686);
and U22353 (N_22353,N_21307,N_21835);
nor U22354 (N_22354,N_21484,N_21879);
or U22355 (N_22355,N_21770,N_21138);
nand U22356 (N_22356,N_21198,N_21163);
nand U22357 (N_22357,N_21394,N_21923);
and U22358 (N_22358,N_21516,N_21957);
and U22359 (N_22359,N_21597,N_21426);
or U22360 (N_22360,N_21947,N_21559);
xor U22361 (N_22361,N_21857,N_21247);
or U22362 (N_22362,N_21954,N_21267);
or U22363 (N_22363,N_21625,N_21051);
nor U22364 (N_22364,N_21102,N_21468);
or U22365 (N_22365,N_21587,N_21376);
nand U22366 (N_22366,N_21790,N_21871);
nand U22367 (N_22367,N_21683,N_21483);
nand U22368 (N_22368,N_21300,N_21632);
and U22369 (N_22369,N_21006,N_21301);
or U22370 (N_22370,N_21023,N_21808);
nor U22371 (N_22371,N_21962,N_21864);
and U22372 (N_22372,N_21785,N_21738);
nand U22373 (N_22373,N_21606,N_21799);
xor U22374 (N_22374,N_21950,N_21557);
xor U22375 (N_22375,N_21926,N_21161);
nand U22376 (N_22376,N_21788,N_21576);
nand U22377 (N_22377,N_21667,N_21949);
xnor U22378 (N_22378,N_21666,N_21956);
xor U22379 (N_22379,N_21863,N_21059);
xnor U22380 (N_22380,N_21205,N_21810);
nor U22381 (N_22381,N_21016,N_21901);
xnor U22382 (N_22382,N_21469,N_21212);
nand U22383 (N_22383,N_21818,N_21880);
nand U22384 (N_22384,N_21458,N_21423);
nor U22385 (N_22385,N_21303,N_21633);
and U22386 (N_22386,N_21285,N_21286);
nor U22387 (N_22387,N_21218,N_21216);
and U22388 (N_22388,N_21042,N_21298);
nand U22389 (N_22389,N_21644,N_21324);
or U22390 (N_22390,N_21192,N_21366);
and U22391 (N_22391,N_21062,N_21627);
nand U22392 (N_22392,N_21900,N_21501);
nor U22393 (N_22393,N_21758,N_21948);
xor U22394 (N_22394,N_21157,N_21840);
nor U22395 (N_22395,N_21371,N_21766);
nand U22396 (N_22396,N_21356,N_21697);
and U22397 (N_22397,N_21622,N_21567);
nand U22398 (N_22398,N_21665,N_21167);
or U22399 (N_22399,N_21554,N_21373);
and U22400 (N_22400,N_21283,N_21358);
and U22401 (N_22401,N_21504,N_21287);
nor U22402 (N_22402,N_21284,N_21230);
and U22403 (N_22403,N_21636,N_21730);
nor U22404 (N_22404,N_21145,N_21639);
nand U22405 (N_22405,N_21539,N_21060);
xor U22406 (N_22406,N_21626,N_21361);
nor U22407 (N_22407,N_21489,N_21202);
and U22408 (N_22408,N_21931,N_21289);
nor U22409 (N_22409,N_21405,N_21614);
or U22410 (N_22410,N_21204,N_21465);
nand U22411 (N_22411,N_21413,N_21601);
nor U22412 (N_22412,N_21188,N_21106);
xor U22413 (N_22413,N_21628,N_21221);
nand U22414 (N_22414,N_21011,N_21097);
nor U22415 (N_22415,N_21674,N_21765);
nor U22416 (N_22416,N_21390,N_21719);
or U22417 (N_22417,N_21421,N_21160);
nor U22418 (N_22418,N_21617,N_21148);
and U22419 (N_22419,N_21441,N_21967);
nor U22420 (N_22420,N_21932,N_21762);
or U22421 (N_22421,N_21562,N_21822);
or U22422 (N_22422,N_21315,N_21798);
and U22423 (N_22423,N_21322,N_21571);
nand U22424 (N_22424,N_21304,N_21977);
or U22425 (N_22425,N_21843,N_21645);
or U22426 (N_22426,N_21695,N_21448);
and U22427 (N_22427,N_21653,N_21946);
or U22428 (N_22428,N_21155,N_21471);
nand U22429 (N_22429,N_21672,N_21520);
and U22430 (N_22430,N_21823,N_21850);
xor U22431 (N_22431,N_21802,N_21712);
and U22432 (N_22432,N_21895,N_21349);
and U22433 (N_22433,N_21733,N_21344);
or U22434 (N_22434,N_21478,N_21852);
or U22435 (N_22435,N_21740,N_21414);
or U22436 (N_22436,N_21158,N_21498);
xnor U22437 (N_22437,N_21814,N_21663);
xnor U22438 (N_22438,N_21299,N_21121);
and U22439 (N_22439,N_21635,N_21331);
nor U22440 (N_22440,N_21370,N_21203);
nor U22441 (N_22441,N_21819,N_21904);
xor U22442 (N_22442,N_21046,N_21195);
xnor U22443 (N_22443,N_21117,N_21154);
or U22444 (N_22444,N_21460,N_21804);
xor U22445 (N_22445,N_21248,N_21355);
and U22446 (N_22446,N_21858,N_21180);
nand U22447 (N_22447,N_21495,N_21573);
or U22448 (N_22448,N_21032,N_21420);
and U22449 (N_22449,N_21972,N_21368);
nor U22450 (N_22450,N_21296,N_21608);
nand U22451 (N_22451,N_21585,N_21072);
nand U22452 (N_22452,N_21975,N_21640);
nor U22453 (N_22453,N_21256,N_21779);
nand U22454 (N_22454,N_21093,N_21094);
nor U22455 (N_22455,N_21507,N_21318);
and U22456 (N_22456,N_21855,N_21604);
nand U22457 (N_22457,N_21586,N_21945);
and U22458 (N_22458,N_21422,N_21113);
nand U22459 (N_22459,N_21074,N_21564);
xor U22460 (N_22460,N_21049,N_21905);
xnor U22461 (N_22461,N_21775,N_21894);
nor U22462 (N_22462,N_21194,N_21924);
xnor U22463 (N_22463,N_21147,N_21903);
nor U22464 (N_22464,N_21727,N_21253);
xor U22465 (N_22465,N_21081,N_21513);
xnor U22466 (N_22466,N_21693,N_21365);
or U22467 (N_22467,N_21937,N_21598);
xor U22468 (N_22468,N_21715,N_21174);
and U22469 (N_22469,N_21410,N_21359);
nand U22470 (N_22470,N_21280,N_21546);
and U22471 (N_22471,N_21943,N_21527);
nand U22472 (N_22472,N_21575,N_21691);
or U22473 (N_22473,N_21226,N_21809);
or U22474 (N_22474,N_21865,N_21224);
and U22475 (N_22475,N_21767,N_21579);
and U22476 (N_22476,N_21752,N_21457);
or U22477 (N_22477,N_21906,N_21278);
and U22478 (N_22478,N_21742,N_21464);
nand U22479 (N_22479,N_21794,N_21907);
nand U22480 (N_22480,N_21724,N_21540);
xnor U22481 (N_22481,N_21692,N_21339);
and U22482 (N_22482,N_21266,N_21682);
or U22483 (N_22483,N_21581,N_21382);
xnor U22484 (N_22484,N_21751,N_21475);
xnor U22485 (N_22485,N_21240,N_21985);
nand U22486 (N_22486,N_21531,N_21544);
and U22487 (N_22487,N_21114,N_21101);
xnor U22488 (N_22488,N_21209,N_21789);
nor U22489 (N_22489,N_21600,N_21293);
nor U22490 (N_22490,N_21070,N_21199);
nand U22491 (N_22491,N_21734,N_21090);
nand U22492 (N_22492,N_21889,N_21713);
and U22493 (N_22493,N_21482,N_21264);
nand U22494 (N_22494,N_21186,N_21326);
xnor U22495 (N_22495,N_21981,N_21528);
and U22496 (N_22496,N_21273,N_21910);
nand U22497 (N_22497,N_21797,N_21024);
or U22498 (N_22498,N_21623,N_21805);
nand U22499 (N_22499,N_21143,N_21162);
or U22500 (N_22500,N_21643,N_21150);
nand U22501 (N_22501,N_21276,N_21343);
or U22502 (N_22502,N_21145,N_21500);
nor U22503 (N_22503,N_21949,N_21577);
nor U22504 (N_22504,N_21686,N_21253);
and U22505 (N_22505,N_21350,N_21290);
and U22506 (N_22506,N_21946,N_21593);
nor U22507 (N_22507,N_21174,N_21615);
and U22508 (N_22508,N_21304,N_21306);
nor U22509 (N_22509,N_21715,N_21818);
xnor U22510 (N_22510,N_21076,N_21290);
or U22511 (N_22511,N_21934,N_21744);
nor U22512 (N_22512,N_21959,N_21461);
or U22513 (N_22513,N_21543,N_21634);
and U22514 (N_22514,N_21000,N_21093);
xnor U22515 (N_22515,N_21584,N_21288);
and U22516 (N_22516,N_21968,N_21340);
and U22517 (N_22517,N_21726,N_21911);
nand U22518 (N_22518,N_21997,N_21074);
nand U22519 (N_22519,N_21489,N_21046);
nand U22520 (N_22520,N_21742,N_21001);
and U22521 (N_22521,N_21013,N_21408);
nor U22522 (N_22522,N_21921,N_21136);
or U22523 (N_22523,N_21163,N_21749);
xor U22524 (N_22524,N_21453,N_21017);
nor U22525 (N_22525,N_21966,N_21336);
xor U22526 (N_22526,N_21203,N_21241);
nor U22527 (N_22527,N_21700,N_21255);
nor U22528 (N_22528,N_21646,N_21371);
xor U22529 (N_22529,N_21869,N_21669);
and U22530 (N_22530,N_21963,N_21234);
or U22531 (N_22531,N_21997,N_21834);
xnor U22532 (N_22532,N_21862,N_21645);
nor U22533 (N_22533,N_21549,N_21702);
nor U22534 (N_22534,N_21569,N_21120);
xor U22535 (N_22535,N_21559,N_21673);
nand U22536 (N_22536,N_21635,N_21615);
nor U22537 (N_22537,N_21010,N_21052);
nand U22538 (N_22538,N_21977,N_21205);
and U22539 (N_22539,N_21567,N_21862);
or U22540 (N_22540,N_21258,N_21511);
nor U22541 (N_22541,N_21212,N_21887);
nor U22542 (N_22542,N_21532,N_21078);
and U22543 (N_22543,N_21360,N_21255);
or U22544 (N_22544,N_21616,N_21086);
or U22545 (N_22545,N_21118,N_21851);
nand U22546 (N_22546,N_21669,N_21010);
xor U22547 (N_22547,N_21259,N_21251);
nor U22548 (N_22548,N_21466,N_21457);
nand U22549 (N_22549,N_21395,N_21472);
or U22550 (N_22550,N_21858,N_21561);
and U22551 (N_22551,N_21913,N_21204);
nor U22552 (N_22552,N_21830,N_21947);
nand U22553 (N_22553,N_21997,N_21541);
nor U22554 (N_22554,N_21406,N_21170);
nor U22555 (N_22555,N_21846,N_21416);
xnor U22556 (N_22556,N_21026,N_21690);
nand U22557 (N_22557,N_21095,N_21125);
nor U22558 (N_22558,N_21205,N_21657);
nor U22559 (N_22559,N_21158,N_21487);
xor U22560 (N_22560,N_21828,N_21658);
nand U22561 (N_22561,N_21594,N_21958);
nor U22562 (N_22562,N_21652,N_21911);
and U22563 (N_22563,N_21873,N_21008);
nand U22564 (N_22564,N_21153,N_21818);
nand U22565 (N_22565,N_21009,N_21492);
xnor U22566 (N_22566,N_21532,N_21851);
nand U22567 (N_22567,N_21890,N_21847);
xor U22568 (N_22568,N_21719,N_21439);
or U22569 (N_22569,N_21220,N_21761);
or U22570 (N_22570,N_21687,N_21942);
nand U22571 (N_22571,N_21061,N_21995);
or U22572 (N_22572,N_21109,N_21282);
xnor U22573 (N_22573,N_21141,N_21635);
nand U22574 (N_22574,N_21660,N_21596);
nor U22575 (N_22575,N_21109,N_21239);
nor U22576 (N_22576,N_21944,N_21118);
or U22577 (N_22577,N_21464,N_21769);
and U22578 (N_22578,N_21242,N_21957);
and U22579 (N_22579,N_21716,N_21476);
or U22580 (N_22580,N_21832,N_21342);
xnor U22581 (N_22581,N_21649,N_21061);
xor U22582 (N_22582,N_21056,N_21057);
or U22583 (N_22583,N_21104,N_21208);
or U22584 (N_22584,N_21437,N_21253);
and U22585 (N_22585,N_21947,N_21002);
and U22586 (N_22586,N_21394,N_21453);
nand U22587 (N_22587,N_21527,N_21978);
or U22588 (N_22588,N_21809,N_21593);
xnor U22589 (N_22589,N_21377,N_21316);
and U22590 (N_22590,N_21052,N_21531);
and U22591 (N_22591,N_21164,N_21518);
nand U22592 (N_22592,N_21391,N_21834);
or U22593 (N_22593,N_21759,N_21275);
and U22594 (N_22594,N_21472,N_21051);
xor U22595 (N_22595,N_21474,N_21894);
xnor U22596 (N_22596,N_21108,N_21840);
and U22597 (N_22597,N_21850,N_21489);
nand U22598 (N_22598,N_21634,N_21054);
xnor U22599 (N_22599,N_21690,N_21402);
nor U22600 (N_22600,N_21361,N_21690);
xor U22601 (N_22601,N_21160,N_21712);
xnor U22602 (N_22602,N_21563,N_21642);
or U22603 (N_22603,N_21286,N_21319);
and U22604 (N_22604,N_21265,N_21267);
and U22605 (N_22605,N_21319,N_21957);
nand U22606 (N_22606,N_21329,N_21843);
nand U22607 (N_22607,N_21455,N_21556);
and U22608 (N_22608,N_21283,N_21050);
nor U22609 (N_22609,N_21969,N_21838);
and U22610 (N_22610,N_21185,N_21650);
nor U22611 (N_22611,N_21389,N_21982);
nand U22612 (N_22612,N_21387,N_21810);
xor U22613 (N_22613,N_21525,N_21659);
or U22614 (N_22614,N_21337,N_21306);
nor U22615 (N_22615,N_21961,N_21513);
xor U22616 (N_22616,N_21193,N_21251);
nand U22617 (N_22617,N_21888,N_21980);
nand U22618 (N_22618,N_21015,N_21267);
and U22619 (N_22619,N_21400,N_21089);
and U22620 (N_22620,N_21052,N_21369);
nand U22621 (N_22621,N_21257,N_21769);
and U22622 (N_22622,N_21817,N_21651);
nand U22623 (N_22623,N_21628,N_21258);
nor U22624 (N_22624,N_21092,N_21664);
or U22625 (N_22625,N_21401,N_21252);
nor U22626 (N_22626,N_21791,N_21989);
nor U22627 (N_22627,N_21216,N_21172);
xor U22628 (N_22628,N_21413,N_21884);
nand U22629 (N_22629,N_21388,N_21045);
xnor U22630 (N_22630,N_21667,N_21781);
nand U22631 (N_22631,N_21801,N_21128);
nor U22632 (N_22632,N_21039,N_21144);
and U22633 (N_22633,N_21516,N_21340);
or U22634 (N_22634,N_21141,N_21798);
or U22635 (N_22635,N_21788,N_21418);
or U22636 (N_22636,N_21122,N_21383);
and U22637 (N_22637,N_21294,N_21986);
nor U22638 (N_22638,N_21573,N_21915);
or U22639 (N_22639,N_21139,N_21224);
and U22640 (N_22640,N_21883,N_21070);
xor U22641 (N_22641,N_21226,N_21022);
and U22642 (N_22642,N_21954,N_21174);
or U22643 (N_22643,N_21888,N_21043);
xor U22644 (N_22644,N_21441,N_21717);
xor U22645 (N_22645,N_21466,N_21679);
nor U22646 (N_22646,N_21217,N_21982);
xnor U22647 (N_22647,N_21021,N_21509);
nand U22648 (N_22648,N_21466,N_21223);
or U22649 (N_22649,N_21142,N_21415);
or U22650 (N_22650,N_21723,N_21405);
nor U22651 (N_22651,N_21417,N_21726);
or U22652 (N_22652,N_21538,N_21347);
or U22653 (N_22653,N_21909,N_21549);
xnor U22654 (N_22654,N_21590,N_21715);
and U22655 (N_22655,N_21600,N_21676);
or U22656 (N_22656,N_21849,N_21792);
or U22657 (N_22657,N_21832,N_21266);
xor U22658 (N_22658,N_21036,N_21285);
and U22659 (N_22659,N_21177,N_21306);
nor U22660 (N_22660,N_21086,N_21283);
nor U22661 (N_22661,N_21750,N_21849);
or U22662 (N_22662,N_21197,N_21443);
nand U22663 (N_22663,N_21456,N_21927);
or U22664 (N_22664,N_21629,N_21639);
or U22665 (N_22665,N_21748,N_21464);
nor U22666 (N_22666,N_21267,N_21521);
and U22667 (N_22667,N_21251,N_21194);
nor U22668 (N_22668,N_21441,N_21576);
or U22669 (N_22669,N_21284,N_21180);
nor U22670 (N_22670,N_21478,N_21275);
and U22671 (N_22671,N_21403,N_21290);
and U22672 (N_22672,N_21743,N_21899);
nor U22673 (N_22673,N_21615,N_21783);
nor U22674 (N_22674,N_21646,N_21207);
or U22675 (N_22675,N_21538,N_21067);
xnor U22676 (N_22676,N_21640,N_21747);
nor U22677 (N_22677,N_21623,N_21838);
xnor U22678 (N_22678,N_21807,N_21709);
nor U22679 (N_22679,N_21110,N_21270);
xor U22680 (N_22680,N_21531,N_21818);
and U22681 (N_22681,N_21068,N_21196);
and U22682 (N_22682,N_21675,N_21977);
and U22683 (N_22683,N_21396,N_21461);
nand U22684 (N_22684,N_21764,N_21282);
xor U22685 (N_22685,N_21148,N_21318);
nand U22686 (N_22686,N_21905,N_21876);
or U22687 (N_22687,N_21409,N_21805);
nand U22688 (N_22688,N_21696,N_21508);
and U22689 (N_22689,N_21384,N_21146);
nor U22690 (N_22690,N_21371,N_21499);
xnor U22691 (N_22691,N_21595,N_21519);
nor U22692 (N_22692,N_21236,N_21367);
and U22693 (N_22693,N_21827,N_21439);
or U22694 (N_22694,N_21856,N_21426);
and U22695 (N_22695,N_21732,N_21710);
nand U22696 (N_22696,N_21993,N_21353);
nand U22697 (N_22697,N_21025,N_21584);
xnor U22698 (N_22698,N_21038,N_21096);
xnor U22699 (N_22699,N_21856,N_21818);
xnor U22700 (N_22700,N_21229,N_21228);
nor U22701 (N_22701,N_21810,N_21093);
or U22702 (N_22702,N_21337,N_21589);
nand U22703 (N_22703,N_21902,N_21160);
nand U22704 (N_22704,N_21808,N_21835);
nand U22705 (N_22705,N_21761,N_21511);
or U22706 (N_22706,N_21057,N_21757);
nand U22707 (N_22707,N_21870,N_21433);
or U22708 (N_22708,N_21181,N_21868);
or U22709 (N_22709,N_21448,N_21416);
nand U22710 (N_22710,N_21327,N_21650);
nor U22711 (N_22711,N_21139,N_21489);
nor U22712 (N_22712,N_21492,N_21779);
and U22713 (N_22713,N_21102,N_21029);
xor U22714 (N_22714,N_21904,N_21210);
nor U22715 (N_22715,N_21980,N_21071);
or U22716 (N_22716,N_21309,N_21753);
nor U22717 (N_22717,N_21258,N_21217);
nor U22718 (N_22718,N_21817,N_21267);
or U22719 (N_22719,N_21110,N_21067);
xor U22720 (N_22720,N_21627,N_21890);
nor U22721 (N_22721,N_21263,N_21106);
xnor U22722 (N_22722,N_21316,N_21044);
xor U22723 (N_22723,N_21677,N_21554);
nand U22724 (N_22724,N_21344,N_21271);
or U22725 (N_22725,N_21922,N_21097);
or U22726 (N_22726,N_21839,N_21938);
nand U22727 (N_22727,N_21692,N_21604);
and U22728 (N_22728,N_21172,N_21632);
or U22729 (N_22729,N_21082,N_21468);
xor U22730 (N_22730,N_21059,N_21871);
nor U22731 (N_22731,N_21207,N_21254);
and U22732 (N_22732,N_21809,N_21454);
and U22733 (N_22733,N_21681,N_21106);
nor U22734 (N_22734,N_21822,N_21365);
nor U22735 (N_22735,N_21378,N_21890);
xor U22736 (N_22736,N_21815,N_21435);
or U22737 (N_22737,N_21214,N_21129);
and U22738 (N_22738,N_21600,N_21361);
nor U22739 (N_22739,N_21883,N_21739);
nand U22740 (N_22740,N_21684,N_21422);
xor U22741 (N_22741,N_21572,N_21569);
and U22742 (N_22742,N_21911,N_21470);
and U22743 (N_22743,N_21633,N_21982);
or U22744 (N_22744,N_21479,N_21002);
nor U22745 (N_22745,N_21846,N_21686);
and U22746 (N_22746,N_21385,N_21610);
nand U22747 (N_22747,N_21679,N_21966);
nand U22748 (N_22748,N_21745,N_21322);
nand U22749 (N_22749,N_21985,N_21164);
nand U22750 (N_22750,N_21547,N_21359);
nor U22751 (N_22751,N_21333,N_21829);
xor U22752 (N_22752,N_21903,N_21367);
and U22753 (N_22753,N_21358,N_21397);
or U22754 (N_22754,N_21444,N_21000);
xor U22755 (N_22755,N_21101,N_21697);
or U22756 (N_22756,N_21991,N_21910);
nand U22757 (N_22757,N_21267,N_21674);
xor U22758 (N_22758,N_21954,N_21029);
and U22759 (N_22759,N_21996,N_21826);
nor U22760 (N_22760,N_21889,N_21983);
nor U22761 (N_22761,N_21265,N_21413);
or U22762 (N_22762,N_21507,N_21361);
nand U22763 (N_22763,N_21687,N_21352);
or U22764 (N_22764,N_21563,N_21036);
nor U22765 (N_22765,N_21723,N_21190);
and U22766 (N_22766,N_21495,N_21614);
or U22767 (N_22767,N_21097,N_21161);
nand U22768 (N_22768,N_21360,N_21168);
and U22769 (N_22769,N_21750,N_21031);
and U22770 (N_22770,N_21518,N_21104);
and U22771 (N_22771,N_21957,N_21462);
nor U22772 (N_22772,N_21940,N_21858);
nor U22773 (N_22773,N_21237,N_21135);
or U22774 (N_22774,N_21104,N_21513);
and U22775 (N_22775,N_21549,N_21688);
nand U22776 (N_22776,N_21377,N_21865);
xor U22777 (N_22777,N_21080,N_21029);
xor U22778 (N_22778,N_21304,N_21642);
xnor U22779 (N_22779,N_21320,N_21600);
and U22780 (N_22780,N_21193,N_21106);
xnor U22781 (N_22781,N_21499,N_21119);
or U22782 (N_22782,N_21871,N_21870);
nor U22783 (N_22783,N_21001,N_21966);
nor U22784 (N_22784,N_21116,N_21545);
nand U22785 (N_22785,N_21203,N_21573);
or U22786 (N_22786,N_21702,N_21822);
and U22787 (N_22787,N_21159,N_21707);
xnor U22788 (N_22788,N_21043,N_21338);
xnor U22789 (N_22789,N_21214,N_21137);
xnor U22790 (N_22790,N_21998,N_21223);
nand U22791 (N_22791,N_21841,N_21062);
or U22792 (N_22792,N_21903,N_21365);
nor U22793 (N_22793,N_21432,N_21821);
nand U22794 (N_22794,N_21985,N_21579);
xor U22795 (N_22795,N_21720,N_21132);
xor U22796 (N_22796,N_21139,N_21608);
xnor U22797 (N_22797,N_21668,N_21451);
or U22798 (N_22798,N_21393,N_21955);
nand U22799 (N_22799,N_21071,N_21710);
and U22800 (N_22800,N_21262,N_21723);
or U22801 (N_22801,N_21659,N_21293);
or U22802 (N_22802,N_21019,N_21527);
nand U22803 (N_22803,N_21763,N_21671);
nor U22804 (N_22804,N_21755,N_21345);
and U22805 (N_22805,N_21332,N_21045);
xor U22806 (N_22806,N_21011,N_21838);
or U22807 (N_22807,N_21722,N_21391);
xnor U22808 (N_22808,N_21343,N_21411);
and U22809 (N_22809,N_21064,N_21774);
nand U22810 (N_22810,N_21539,N_21561);
or U22811 (N_22811,N_21546,N_21929);
or U22812 (N_22812,N_21312,N_21481);
nand U22813 (N_22813,N_21321,N_21360);
nand U22814 (N_22814,N_21977,N_21469);
nor U22815 (N_22815,N_21842,N_21071);
nand U22816 (N_22816,N_21618,N_21439);
nor U22817 (N_22817,N_21531,N_21271);
nor U22818 (N_22818,N_21455,N_21760);
or U22819 (N_22819,N_21658,N_21126);
or U22820 (N_22820,N_21135,N_21750);
nand U22821 (N_22821,N_21134,N_21694);
or U22822 (N_22822,N_21631,N_21653);
nor U22823 (N_22823,N_21214,N_21762);
nand U22824 (N_22824,N_21912,N_21282);
or U22825 (N_22825,N_21629,N_21788);
nand U22826 (N_22826,N_21885,N_21929);
nand U22827 (N_22827,N_21346,N_21024);
nand U22828 (N_22828,N_21242,N_21241);
xor U22829 (N_22829,N_21601,N_21304);
xor U22830 (N_22830,N_21836,N_21560);
xnor U22831 (N_22831,N_21738,N_21452);
xor U22832 (N_22832,N_21255,N_21070);
or U22833 (N_22833,N_21421,N_21066);
xnor U22834 (N_22834,N_21652,N_21145);
nand U22835 (N_22835,N_21813,N_21390);
nor U22836 (N_22836,N_21159,N_21894);
xor U22837 (N_22837,N_21766,N_21797);
and U22838 (N_22838,N_21972,N_21307);
xnor U22839 (N_22839,N_21946,N_21154);
and U22840 (N_22840,N_21129,N_21714);
xnor U22841 (N_22841,N_21427,N_21593);
nor U22842 (N_22842,N_21010,N_21769);
nand U22843 (N_22843,N_21390,N_21517);
or U22844 (N_22844,N_21709,N_21441);
nor U22845 (N_22845,N_21616,N_21362);
or U22846 (N_22846,N_21735,N_21945);
xor U22847 (N_22847,N_21344,N_21886);
nand U22848 (N_22848,N_21394,N_21357);
nand U22849 (N_22849,N_21156,N_21966);
xnor U22850 (N_22850,N_21758,N_21539);
nand U22851 (N_22851,N_21805,N_21177);
nand U22852 (N_22852,N_21774,N_21886);
nor U22853 (N_22853,N_21256,N_21076);
nand U22854 (N_22854,N_21781,N_21535);
nor U22855 (N_22855,N_21143,N_21248);
xor U22856 (N_22856,N_21692,N_21300);
and U22857 (N_22857,N_21450,N_21815);
or U22858 (N_22858,N_21352,N_21740);
and U22859 (N_22859,N_21383,N_21926);
and U22860 (N_22860,N_21464,N_21019);
or U22861 (N_22861,N_21972,N_21381);
nor U22862 (N_22862,N_21069,N_21202);
or U22863 (N_22863,N_21324,N_21970);
xnor U22864 (N_22864,N_21449,N_21058);
or U22865 (N_22865,N_21023,N_21529);
nand U22866 (N_22866,N_21777,N_21234);
or U22867 (N_22867,N_21998,N_21619);
xor U22868 (N_22868,N_21352,N_21322);
nand U22869 (N_22869,N_21590,N_21005);
xor U22870 (N_22870,N_21965,N_21973);
nor U22871 (N_22871,N_21909,N_21598);
xor U22872 (N_22872,N_21005,N_21957);
xnor U22873 (N_22873,N_21252,N_21494);
nor U22874 (N_22874,N_21583,N_21253);
and U22875 (N_22875,N_21394,N_21489);
nand U22876 (N_22876,N_21365,N_21341);
and U22877 (N_22877,N_21334,N_21088);
and U22878 (N_22878,N_21389,N_21557);
xnor U22879 (N_22879,N_21808,N_21658);
nand U22880 (N_22880,N_21252,N_21577);
nand U22881 (N_22881,N_21585,N_21296);
nand U22882 (N_22882,N_21135,N_21535);
xor U22883 (N_22883,N_21013,N_21335);
and U22884 (N_22884,N_21386,N_21469);
or U22885 (N_22885,N_21080,N_21613);
xnor U22886 (N_22886,N_21788,N_21779);
or U22887 (N_22887,N_21797,N_21825);
xor U22888 (N_22888,N_21767,N_21499);
xnor U22889 (N_22889,N_21732,N_21359);
xnor U22890 (N_22890,N_21352,N_21961);
or U22891 (N_22891,N_21911,N_21474);
nand U22892 (N_22892,N_21557,N_21928);
and U22893 (N_22893,N_21426,N_21133);
and U22894 (N_22894,N_21520,N_21359);
xor U22895 (N_22895,N_21001,N_21765);
or U22896 (N_22896,N_21229,N_21877);
and U22897 (N_22897,N_21349,N_21312);
and U22898 (N_22898,N_21895,N_21542);
nand U22899 (N_22899,N_21577,N_21983);
xor U22900 (N_22900,N_21804,N_21166);
nand U22901 (N_22901,N_21272,N_21277);
nand U22902 (N_22902,N_21162,N_21613);
nand U22903 (N_22903,N_21345,N_21605);
nor U22904 (N_22904,N_21689,N_21756);
xor U22905 (N_22905,N_21653,N_21277);
or U22906 (N_22906,N_21456,N_21431);
xor U22907 (N_22907,N_21118,N_21389);
or U22908 (N_22908,N_21491,N_21711);
xor U22909 (N_22909,N_21562,N_21627);
or U22910 (N_22910,N_21918,N_21073);
or U22911 (N_22911,N_21572,N_21348);
nor U22912 (N_22912,N_21943,N_21244);
nor U22913 (N_22913,N_21567,N_21023);
nand U22914 (N_22914,N_21302,N_21077);
and U22915 (N_22915,N_21466,N_21036);
nand U22916 (N_22916,N_21056,N_21781);
nand U22917 (N_22917,N_21185,N_21129);
nor U22918 (N_22918,N_21913,N_21873);
or U22919 (N_22919,N_21604,N_21972);
and U22920 (N_22920,N_21379,N_21452);
nor U22921 (N_22921,N_21418,N_21421);
and U22922 (N_22922,N_21886,N_21722);
and U22923 (N_22923,N_21758,N_21227);
and U22924 (N_22924,N_21462,N_21578);
nor U22925 (N_22925,N_21255,N_21619);
nand U22926 (N_22926,N_21637,N_21276);
xor U22927 (N_22927,N_21461,N_21687);
and U22928 (N_22928,N_21549,N_21293);
xnor U22929 (N_22929,N_21771,N_21620);
and U22930 (N_22930,N_21989,N_21190);
nand U22931 (N_22931,N_21540,N_21075);
xnor U22932 (N_22932,N_21972,N_21116);
and U22933 (N_22933,N_21661,N_21431);
and U22934 (N_22934,N_21128,N_21895);
and U22935 (N_22935,N_21209,N_21373);
nor U22936 (N_22936,N_21975,N_21998);
xor U22937 (N_22937,N_21414,N_21230);
xor U22938 (N_22938,N_21761,N_21688);
xnor U22939 (N_22939,N_21549,N_21896);
xor U22940 (N_22940,N_21812,N_21443);
xnor U22941 (N_22941,N_21053,N_21879);
nand U22942 (N_22942,N_21856,N_21351);
and U22943 (N_22943,N_21232,N_21000);
xnor U22944 (N_22944,N_21005,N_21105);
or U22945 (N_22945,N_21630,N_21901);
and U22946 (N_22946,N_21616,N_21729);
or U22947 (N_22947,N_21833,N_21951);
nor U22948 (N_22948,N_21608,N_21607);
xnor U22949 (N_22949,N_21406,N_21455);
nand U22950 (N_22950,N_21207,N_21630);
nor U22951 (N_22951,N_21662,N_21852);
and U22952 (N_22952,N_21109,N_21062);
nor U22953 (N_22953,N_21352,N_21497);
or U22954 (N_22954,N_21569,N_21994);
and U22955 (N_22955,N_21125,N_21222);
or U22956 (N_22956,N_21382,N_21626);
xnor U22957 (N_22957,N_21856,N_21828);
and U22958 (N_22958,N_21120,N_21928);
nor U22959 (N_22959,N_21319,N_21949);
or U22960 (N_22960,N_21337,N_21588);
nand U22961 (N_22961,N_21569,N_21359);
xor U22962 (N_22962,N_21061,N_21920);
xor U22963 (N_22963,N_21347,N_21935);
nand U22964 (N_22964,N_21760,N_21649);
nor U22965 (N_22965,N_21476,N_21880);
and U22966 (N_22966,N_21526,N_21836);
or U22967 (N_22967,N_21628,N_21516);
or U22968 (N_22968,N_21557,N_21703);
xnor U22969 (N_22969,N_21765,N_21770);
nor U22970 (N_22970,N_21132,N_21180);
xor U22971 (N_22971,N_21511,N_21646);
nor U22972 (N_22972,N_21709,N_21310);
and U22973 (N_22973,N_21941,N_21679);
nor U22974 (N_22974,N_21499,N_21752);
and U22975 (N_22975,N_21831,N_21893);
and U22976 (N_22976,N_21514,N_21444);
nor U22977 (N_22977,N_21947,N_21284);
or U22978 (N_22978,N_21566,N_21396);
nand U22979 (N_22979,N_21497,N_21001);
nor U22980 (N_22980,N_21187,N_21383);
nand U22981 (N_22981,N_21259,N_21480);
and U22982 (N_22982,N_21454,N_21650);
or U22983 (N_22983,N_21796,N_21440);
or U22984 (N_22984,N_21983,N_21854);
or U22985 (N_22985,N_21526,N_21261);
xnor U22986 (N_22986,N_21278,N_21415);
and U22987 (N_22987,N_21358,N_21097);
xor U22988 (N_22988,N_21398,N_21048);
nand U22989 (N_22989,N_21390,N_21127);
nor U22990 (N_22990,N_21200,N_21660);
nor U22991 (N_22991,N_21216,N_21483);
or U22992 (N_22992,N_21962,N_21713);
nand U22993 (N_22993,N_21975,N_21475);
and U22994 (N_22994,N_21373,N_21813);
or U22995 (N_22995,N_21973,N_21851);
and U22996 (N_22996,N_21516,N_21110);
and U22997 (N_22997,N_21071,N_21780);
and U22998 (N_22998,N_21848,N_21651);
nor U22999 (N_22999,N_21679,N_21874);
and U23000 (N_23000,N_22159,N_22322);
nor U23001 (N_23001,N_22502,N_22423);
xor U23002 (N_23002,N_22766,N_22475);
xnor U23003 (N_23003,N_22319,N_22468);
or U23004 (N_23004,N_22767,N_22626);
and U23005 (N_23005,N_22980,N_22362);
nand U23006 (N_23006,N_22131,N_22897);
or U23007 (N_23007,N_22261,N_22177);
or U23008 (N_23008,N_22492,N_22915);
and U23009 (N_23009,N_22176,N_22971);
and U23010 (N_23010,N_22305,N_22257);
and U23011 (N_23011,N_22955,N_22228);
nor U23012 (N_23012,N_22393,N_22563);
and U23013 (N_23013,N_22802,N_22372);
nor U23014 (N_23014,N_22841,N_22637);
nand U23015 (N_23015,N_22365,N_22211);
xnor U23016 (N_23016,N_22146,N_22214);
or U23017 (N_23017,N_22594,N_22990);
and U23018 (N_23018,N_22227,N_22989);
and U23019 (N_23019,N_22086,N_22441);
xnor U23020 (N_23020,N_22616,N_22115);
nor U23021 (N_23021,N_22507,N_22470);
nor U23022 (N_23022,N_22660,N_22545);
nor U23023 (N_23023,N_22657,N_22093);
nor U23024 (N_23024,N_22346,N_22341);
and U23025 (N_23025,N_22585,N_22624);
or U23026 (N_23026,N_22930,N_22831);
xor U23027 (N_23027,N_22366,N_22771);
and U23028 (N_23028,N_22705,N_22091);
or U23029 (N_23029,N_22071,N_22128);
nor U23030 (N_23030,N_22108,N_22247);
nor U23031 (N_23031,N_22168,N_22753);
and U23032 (N_23032,N_22076,N_22263);
nand U23033 (N_23033,N_22278,N_22401);
nand U23034 (N_23034,N_22537,N_22813);
nand U23035 (N_23035,N_22758,N_22613);
and U23036 (N_23036,N_22386,N_22924);
nor U23037 (N_23037,N_22495,N_22557);
nand U23038 (N_23038,N_22727,N_22420);
xnor U23039 (N_23039,N_22986,N_22892);
nor U23040 (N_23040,N_22041,N_22796);
nand U23041 (N_23041,N_22325,N_22439);
and U23042 (N_23042,N_22785,N_22044);
nor U23043 (N_23043,N_22260,N_22781);
xor U23044 (N_23044,N_22815,N_22552);
nand U23045 (N_23045,N_22474,N_22419);
nor U23046 (N_23046,N_22623,N_22693);
nor U23047 (N_23047,N_22584,N_22191);
nand U23048 (N_23048,N_22901,N_22060);
xnor U23049 (N_23049,N_22764,N_22374);
nand U23050 (N_23050,N_22772,N_22575);
and U23051 (N_23051,N_22493,N_22605);
and U23052 (N_23052,N_22975,N_22745);
and U23053 (N_23053,N_22588,N_22857);
xnor U23054 (N_23054,N_22996,N_22883);
xor U23055 (N_23055,N_22740,N_22694);
xnor U23056 (N_23056,N_22016,N_22617);
and U23057 (N_23057,N_22377,N_22824);
nand U23058 (N_23058,N_22593,N_22804);
nand U23059 (N_23059,N_22438,N_22382);
and U23060 (N_23060,N_22524,N_22598);
xnor U23061 (N_23061,N_22890,N_22236);
nand U23062 (N_23062,N_22369,N_22483);
xor U23063 (N_23063,N_22416,N_22117);
and U23064 (N_23064,N_22392,N_22183);
xnor U23065 (N_23065,N_22925,N_22821);
xor U23066 (N_23066,N_22097,N_22424);
nand U23067 (N_23067,N_22381,N_22718);
nand U23068 (N_23068,N_22453,N_22048);
nor U23069 (N_23069,N_22042,N_22118);
xnor U23070 (N_23070,N_22875,N_22929);
or U23071 (N_23071,N_22065,N_22982);
nand U23072 (N_23072,N_22978,N_22564);
nor U23073 (N_23073,N_22581,N_22997);
xor U23074 (N_23074,N_22242,N_22210);
xor U23075 (N_23075,N_22167,N_22334);
nor U23076 (N_23076,N_22269,N_22449);
xor U23077 (N_23077,N_22773,N_22948);
nand U23078 (N_23078,N_22787,N_22618);
or U23079 (N_23079,N_22153,N_22685);
nand U23080 (N_23080,N_22390,N_22513);
and U23081 (N_23081,N_22992,N_22414);
or U23082 (N_23082,N_22953,N_22706);
nand U23083 (N_23083,N_22778,N_22239);
or U23084 (N_23084,N_22583,N_22850);
xor U23085 (N_23085,N_22595,N_22232);
and U23086 (N_23086,N_22122,N_22479);
or U23087 (N_23087,N_22505,N_22205);
or U23088 (N_23088,N_22161,N_22387);
or U23089 (N_23089,N_22422,N_22272);
xor U23090 (N_23090,N_22889,N_22163);
nor U23091 (N_23091,N_22789,N_22709);
nand U23092 (N_23092,N_22648,N_22240);
nor U23093 (N_23093,N_22360,N_22107);
xor U23094 (N_23094,N_22763,N_22826);
or U23095 (N_23095,N_22469,N_22208);
or U23096 (N_23096,N_22506,N_22641);
nand U23097 (N_23097,N_22612,N_22794);
and U23098 (N_23098,N_22729,N_22716);
xor U23099 (N_23099,N_22017,N_22528);
nand U23100 (N_23100,N_22994,N_22877);
nand U23101 (N_23101,N_22030,N_22779);
and U23102 (N_23102,N_22212,N_22072);
nand U23103 (N_23103,N_22881,N_22610);
xnor U23104 (N_23104,N_22429,N_22898);
xnor U23105 (N_23105,N_22678,N_22238);
nor U23106 (N_23106,N_22849,N_22103);
or U23107 (N_23107,N_22172,N_22171);
nor U23108 (N_23108,N_22047,N_22486);
nand U23109 (N_23109,N_22330,N_22809);
nand U23110 (N_23110,N_22795,N_22320);
and U23111 (N_23111,N_22525,N_22052);
nor U23112 (N_23112,N_22291,N_22104);
or U23113 (N_23113,N_22001,N_22406);
or U23114 (N_23114,N_22855,N_22150);
or U23115 (N_23115,N_22683,N_22039);
and U23116 (N_23116,N_22943,N_22958);
nand U23117 (N_23117,N_22417,N_22477);
xnor U23118 (N_23118,N_22735,N_22137);
nand U23119 (N_23119,N_22517,N_22918);
nor U23120 (N_23120,N_22088,N_22717);
and U23121 (N_23121,N_22644,N_22113);
nor U23122 (N_23122,N_22669,N_22684);
nor U23123 (N_23123,N_22891,N_22409);
and U23124 (N_23124,N_22286,N_22184);
nor U23125 (N_23125,N_22723,N_22762);
nand U23126 (N_23126,N_22871,N_22018);
or U23127 (N_23127,N_22614,N_22887);
and U23128 (N_23128,N_22218,N_22459);
xor U23129 (N_23129,N_22661,N_22741);
nor U23130 (N_23130,N_22664,N_22932);
nand U23131 (N_23131,N_22731,N_22193);
and U23132 (N_23132,N_22699,N_22124);
nand U23133 (N_23133,N_22285,N_22636);
xor U23134 (N_23134,N_22920,N_22885);
or U23135 (N_23135,N_22970,N_22730);
nor U23136 (N_23136,N_22548,N_22814);
nor U23137 (N_23137,N_22518,N_22457);
and U23138 (N_23138,N_22295,N_22798);
or U23139 (N_23139,N_22913,N_22700);
or U23140 (N_23140,N_22508,N_22127);
xnor U23141 (N_23141,N_22323,N_22421);
nand U23142 (N_23142,N_22155,N_22911);
or U23143 (N_23143,N_22467,N_22586);
nor U23144 (N_23144,N_22848,N_22009);
and U23145 (N_23145,N_22051,N_22573);
nor U23146 (N_23146,N_22682,N_22349);
or U23147 (N_23147,N_22491,N_22570);
nand U23148 (N_23148,N_22345,N_22977);
xor U23149 (N_23149,N_22268,N_22514);
xnor U23150 (N_23150,N_22966,N_22974);
and U23151 (N_23151,N_22547,N_22324);
and U23152 (N_23152,N_22264,N_22830);
nor U23153 (N_23153,N_22602,N_22222);
or U23154 (N_23154,N_22301,N_22357);
or U23155 (N_23155,N_22724,N_22968);
nand U23156 (N_23156,N_22542,N_22946);
nor U23157 (N_23157,N_22936,N_22099);
and U23158 (N_23158,N_22534,N_22756);
xor U23159 (N_23159,N_22645,N_22267);
and U23160 (N_23160,N_22859,N_22769);
xnor U23161 (N_23161,N_22343,N_22904);
nand U23162 (N_23162,N_22375,N_22535);
and U23163 (N_23163,N_22774,N_22659);
nand U23164 (N_23164,N_22793,N_22111);
nor U23165 (N_23165,N_22029,N_22383);
nand U23166 (N_23166,N_22102,N_22998);
nand U23167 (N_23167,N_22510,N_22567);
nand U23168 (N_23168,N_22199,N_22630);
and U23169 (N_23169,N_22942,N_22165);
nand U23170 (N_23170,N_22022,N_22649);
and U23171 (N_23171,N_22728,N_22309);
and U23172 (N_23172,N_22253,N_22750);
or U23173 (N_23173,N_22311,N_22248);
and U23174 (N_23174,N_22187,N_22520);
nand U23175 (N_23175,N_22189,N_22209);
xor U23176 (N_23176,N_22005,N_22845);
nor U23177 (N_23177,N_22355,N_22835);
nor U23178 (N_23178,N_22589,N_22903);
nand U23179 (N_23179,N_22962,N_22504);
nor U23180 (N_23180,N_22204,N_22079);
and U23181 (N_23181,N_22241,N_22270);
nand U23182 (N_23182,N_22021,N_22461);
xor U23183 (N_23183,N_22391,N_22095);
nand U23184 (N_23184,N_22689,N_22080);
xnor U23185 (N_23185,N_22152,N_22344);
nor U23186 (N_23186,N_22299,N_22579);
nand U23187 (N_23187,N_22959,N_22023);
xnor U23188 (N_23188,N_22655,N_22512);
xnor U23189 (N_23189,N_22234,N_22351);
or U23190 (N_23190,N_22237,N_22791);
nand U23191 (N_23191,N_22668,N_22412);
nand U23192 (N_23192,N_22806,N_22100);
nor U23193 (N_23193,N_22577,N_22829);
nor U23194 (N_23194,N_22940,N_22494);
and U23195 (N_23195,N_22621,N_22280);
nand U23196 (N_23196,N_22482,N_22574);
or U23197 (N_23197,N_22003,N_22134);
nand U23198 (N_23198,N_22780,N_22714);
nor U23199 (N_23199,N_22854,N_22591);
or U23200 (N_23200,N_22034,N_22752);
xnor U23201 (N_23201,N_22147,N_22969);
or U23202 (N_23202,N_22279,N_22036);
and U23203 (N_23203,N_22004,N_22761);
nand U23204 (N_23204,N_22526,N_22556);
xnor U23205 (N_23205,N_22129,N_22569);
nand U23206 (N_23206,N_22865,N_22817);
xnor U23207 (N_23207,N_22646,N_22202);
nand U23208 (N_23208,N_22571,N_22909);
or U23209 (N_23209,N_22979,N_22656);
nor U23210 (N_23210,N_22712,N_22873);
and U23211 (N_23211,N_22415,N_22020);
nand U23212 (N_23212,N_22064,N_22175);
and U23213 (N_23213,N_22148,N_22331);
and U23214 (N_23214,N_22775,N_22028);
or U23215 (N_23215,N_22303,N_22370);
xor U23216 (N_23216,N_22460,N_22490);
or U23217 (N_23217,N_22335,N_22398);
and U23218 (N_23218,N_22995,N_22456);
xnor U23219 (N_23219,N_22861,N_22067);
xor U23220 (N_23220,N_22058,N_22462);
nand U23221 (N_23221,N_22266,N_22277);
nor U23222 (N_23222,N_22884,N_22606);
xnor U23223 (N_23223,N_22770,N_22686);
or U23224 (N_23224,N_22927,N_22478);
or U23225 (N_23225,N_22522,N_22224);
xor U23226 (N_23226,N_22213,N_22098);
and U23227 (N_23227,N_22938,N_22704);
and U23228 (N_23228,N_22447,N_22084);
nand U23229 (N_23229,N_22838,N_22035);
nor U23230 (N_23230,N_22484,N_22380);
xor U23231 (N_23231,N_22089,N_22832);
xnor U23232 (N_23232,N_22288,N_22216);
or U23233 (N_23233,N_22307,N_22258);
and U23234 (N_23234,N_22455,N_22869);
or U23235 (N_23235,N_22697,N_22851);
and U23236 (N_23236,N_22519,N_22116);
xnor U23237 (N_23237,N_22905,N_22967);
and U23238 (N_23238,N_22825,N_22054);
nor U23239 (N_23239,N_22452,N_22436);
and U23240 (N_23240,N_22642,N_22059);
xnor U23241 (N_23241,N_22130,N_22434);
and U23242 (N_23242,N_22900,N_22139);
and U23243 (N_23243,N_22874,N_22445);
and U23244 (N_23244,N_22870,N_22866);
xnor U23245 (N_23245,N_22596,N_22354);
nand U23246 (N_23246,N_22653,N_22939);
nor U23247 (N_23247,N_22895,N_22008);
nor U23248 (N_23248,N_22226,N_22867);
nor U23249 (N_23249,N_22050,N_22275);
nor U23250 (N_23250,N_22799,N_22114);
and U23251 (N_23251,N_22919,N_22852);
or U23252 (N_23252,N_22732,N_22533);
or U23253 (N_23253,N_22912,N_22011);
nand U23254 (N_23254,N_22976,N_22444);
xnor U23255 (N_23255,N_22283,N_22294);
xnor U23256 (N_23256,N_22244,N_22543);
nor U23257 (N_23257,N_22120,N_22040);
and U23258 (N_23258,N_22687,N_22411);
nor U23259 (N_23259,N_22092,N_22880);
and U23260 (N_23260,N_22744,N_22371);
and U23261 (N_23261,N_22647,N_22529);
and U23262 (N_23262,N_22639,N_22907);
xor U23263 (N_23263,N_22627,N_22609);
xor U23264 (N_23264,N_22576,N_22466);
and U23265 (N_23265,N_22201,N_22746);
xnor U23266 (N_23266,N_22255,N_22135);
nor U23267 (N_23267,N_22643,N_22549);
nand U23268 (N_23268,N_22726,N_22074);
or U23269 (N_23269,N_22140,N_22014);
xnor U23270 (N_23270,N_22822,N_22332);
or U23271 (N_23271,N_22910,N_22676);
nand U23272 (N_23272,N_22565,N_22496);
nand U23273 (N_23273,N_22551,N_22720);
nand U23274 (N_23274,N_22688,N_22707);
nor U23275 (N_23275,N_22427,N_22908);
or U23276 (N_23276,N_22056,N_22840);
or U23277 (N_23277,N_22776,N_22151);
and U23278 (N_23278,N_22336,N_22158);
nand U23279 (N_23279,N_22801,N_22562);
nand U23280 (N_23280,N_22265,N_22077);
and U23281 (N_23281,N_22431,N_22068);
nand U23282 (N_23282,N_22703,N_22471);
and U23283 (N_23283,N_22680,N_22734);
nand U23284 (N_23284,N_22843,N_22828);
nor U23285 (N_23285,N_22405,N_22677);
nor U23286 (N_23286,N_22473,N_22179);
nor U23287 (N_23287,N_22329,N_22310);
nand U23288 (N_23288,N_22983,N_22634);
xor U23289 (N_23289,N_22950,N_22738);
xor U23290 (N_23290,N_22666,N_22923);
xor U23291 (N_23291,N_22066,N_22464);
nor U23292 (N_23292,N_22608,N_22252);
nor U23293 (N_23293,N_22451,N_22662);
nor U23294 (N_23294,N_22378,N_22742);
or U23295 (N_23295,N_22934,N_22027);
xnor U23296 (N_23296,N_22190,N_22230);
nand U23297 (N_23297,N_22546,N_22715);
nor U23298 (N_23298,N_22757,N_22057);
xor U23299 (N_23299,N_22160,N_22019);
xor U23300 (N_23300,N_22192,N_22157);
nand U23301 (N_23301,N_22797,N_22651);
or U23302 (N_23302,N_22333,N_22396);
nand U23303 (N_23303,N_22635,N_22868);
nand U23304 (N_23304,N_22458,N_22862);
nand U23305 (N_23305,N_22481,N_22926);
nand U23306 (N_23306,N_22864,N_22105);
xor U23307 (N_23307,N_22652,N_22149);
and U23308 (N_23308,N_22364,N_22561);
and U23309 (N_23309,N_22872,N_22245);
or U23310 (N_23310,N_22070,N_22572);
xor U23311 (N_23311,N_22788,N_22296);
and U23312 (N_23312,N_22987,N_22203);
xnor U23313 (N_23313,N_22094,N_22082);
or U23314 (N_23314,N_22297,N_22181);
xor U23315 (N_23315,N_22026,N_22418);
xor U23316 (N_23316,N_22600,N_22225);
or U23317 (N_23317,N_22553,N_22480);
nor U23318 (N_23318,N_22818,N_22413);
nor U23319 (N_23319,N_22917,N_22031);
nand U23320 (N_23320,N_22988,N_22782);
nand U23321 (N_23321,N_22200,N_22816);
and U23322 (N_23322,N_22748,N_22235);
nand U23323 (N_23323,N_22428,N_22006);
nor U23324 (N_23324,N_22404,N_22142);
nand U23325 (N_23325,N_22170,N_22198);
or U23326 (N_23326,N_22856,N_22601);
and U23327 (N_23327,N_22515,N_22132);
nand U23328 (N_23328,N_22388,N_22217);
and U23329 (N_23329,N_22195,N_22672);
nand U23330 (N_23330,N_22592,N_22844);
xor U23331 (N_23331,N_22300,N_22282);
and U23332 (N_23332,N_22555,N_22560);
xor U23333 (N_23333,N_22860,N_22273);
nand U23334 (N_23334,N_22629,N_22043);
nand U23335 (N_23335,N_22085,N_22281);
nand U23336 (N_23336,N_22143,N_22681);
nand U23337 (N_23337,N_22347,N_22024);
nor U23338 (N_23338,N_22069,N_22298);
or U23339 (N_23339,N_22407,N_22038);
or U23340 (N_23340,N_22182,N_22803);
and U23341 (N_23341,N_22931,N_22587);
and U23342 (N_23342,N_22622,N_22509);
or U23343 (N_23343,N_22194,N_22389);
or U23344 (N_23344,N_22985,N_22174);
xnor U23345 (N_23345,N_22500,N_22532);
xnor U23346 (N_23346,N_22373,N_22733);
and U23347 (N_23347,N_22550,N_22765);
nor U23348 (N_23348,N_22454,N_22619);
and U23349 (N_23349,N_22823,N_22442);
or U23350 (N_23350,N_22960,N_22197);
xor U23351 (N_23351,N_22708,N_22376);
or U23352 (N_23352,N_22073,N_22751);
and U23353 (N_23353,N_22807,N_22433);
and U23354 (N_23354,N_22119,N_22719);
nand U23355 (N_23355,N_22081,N_22304);
or U23356 (N_23356,N_22558,N_22790);
nand U23357 (N_23357,N_22002,N_22944);
nand U23358 (N_23358,N_22658,N_22087);
and U23359 (N_23359,N_22246,N_22759);
nor U23360 (N_23360,N_22358,N_22367);
nand U23361 (N_23361,N_22747,N_22498);
or U23362 (N_23362,N_22896,N_22338);
nor U23363 (N_23363,N_22062,N_22952);
nor U23364 (N_23364,N_22692,N_22679);
nor U23365 (N_23365,N_22876,N_22945);
xnor U23366 (N_23366,N_22049,N_22957);
nor U23367 (N_23367,N_22702,N_22604);
or U23368 (N_23368,N_22947,N_22650);
or U23369 (N_23369,N_22568,N_22965);
nor U23370 (N_23370,N_22321,N_22465);
and U23371 (N_23371,N_22410,N_22437);
nor U23372 (N_23372,N_22858,N_22786);
nor U23373 (N_23373,N_22096,N_22126);
or U23374 (N_23374,N_22327,N_22691);
nor U23375 (N_23375,N_22219,N_22951);
and U23376 (N_23376,N_22169,N_22141);
nand U23377 (N_23377,N_22981,N_22274);
nand U23378 (N_23378,N_22670,N_22262);
and U23379 (N_23379,N_22863,N_22013);
and U23380 (N_23380,N_22805,N_22206);
xnor U23381 (N_23381,N_22276,N_22501);
and U23382 (N_23382,N_22725,N_22984);
nand U23383 (N_23383,N_22783,N_22012);
or U23384 (N_23384,N_22611,N_22640);
xor U23385 (N_23385,N_22544,N_22145);
xor U23386 (N_23386,N_22739,N_22937);
nor U23387 (N_23387,N_22136,N_22760);
xnor U23388 (N_23388,N_22882,N_22839);
xor U23389 (N_23389,N_22173,N_22949);
xor U23390 (N_23390,N_22620,N_22736);
or U23391 (N_23391,N_22886,N_22554);
xnor U23392 (N_23392,N_22359,N_22207);
and U23393 (N_23393,N_22254,N_22231);
or U23394 (N_23394,N_22743,N_22921);
and U23395 (N_23395,N_22768,N_22582);
nand U23396 (N_23396,N_22559,N_22340);
xor U23397 (N_23397,N_22314,N_22511);
nor U23398 (N_23398,N_22698,N_22223);
and U23399 (N_23399,N_22671,N_22403);
or U23400 (N_23400,N_22928,N_22394);
xnor U23401 (N_23401,N_22721,N_22308);
nand U23402 (N_23402,N_22633,N_22178);
xnor U23403 (N_23403,N_22902,N_22450);
nor U23404 (N_23404,N_22055,N_22590);
xnor U23405 (N_23405,N_22527,N_22144);
and U23406 (N_23406,N_22337,N_22888);
nor U23407 (N_23407,N_22722,N_22667);
nor U23408 (N_23408,N_22166,N_22833);
or U23409 (N_23409,N_22312,N_22318);
xor U23410 (N_23410,N_22836,N_22138);
and U23411 (N_23411,N_22993,N_22025);
xnor U23412 (N_23412,N_22430,N_22665);
and U23413 (N_23413,N_22538,N_22906);
nor U23414 (N_23414,N_22625,N_22954);
or U23415 (N_23415,N_22063,N_22922);
or U23416 (N_23416,N_22654,N_22353);
or U23417 (N_23417,N_22164,N_22638);
xor U23418 (N_23418,N_22603,N_22315);
nor U23419 (N_23419,N_22597,N_22125);
nand U23420 (N_23420,N_22154,N_22631);
nand U23421 (N_23421,N_22292,N_22083);
or U23422 (N_23422,N_22015,N_22536);
and U23423 (N_23423,N_22488,N_22162);
or U23424 (N_23424,N_22326,N_22271);
xnor U23425 (N_23425,N_22800,N_22348);
nand U23426 (N_23426,N_22489,N_22632);
nor U23427 (N_23427,N_22792,N_22363);
nand U23428 (N_23428,N_22251,N_22425);
and U23429 (N_23429,N_22061,N_22808);
or U23430 (N_23430,N_22221,N_22819);
nor U23431 (N_23431,N_22476,N_22487);
nand U23432 (N_23432,N_22754,N_22010);
or U23433 (N_23433,N_22289,N_22188);
nor U23434 (N_23434,N_22400,N_22810);
or U23435 (N_23435,N_22399,N_22379);
and U23436 (N_23436,N_22110,N_22916);
nand U23437 (N_23437,N_22991,N_22032);
or U23438 (N_23438,N_22385,N_22185);
nor U23439 (N_23439,N_22847,N_22408);
or U23440 (N_23440,N_22499,N_22186);
or U23441 (N_23441,N_22302,N_22287);
and U23442 (N_23442,N_22531,N_22812);
or U23443 (N_23443,N_22133,N_22313);
nor U23444 (N_23444,N_22249,N_22749);
and U23445 (N_23445,N_22395,N_22293);
or U23446 (N_23446,N_22196,N_22316);
or U23447 (N_23447,N_22259,N_22397);
nor U23448 (N_23448,N_22090,N_22899);
nand U23449 (N_23449,N_22834,N_22820);
nor U23450 (N_23450,N_22615,N_22243);
or U23451 (N_23451,N_22432,N_22811);
nor U23452 (N_23452,N_22894,N_22485);
and U23453 (N_23453,N_22463,N_22503);
nor U23454 (N_23454,N_22737,N_22933);
and U23455 (N_23455,N_22256,N_22827);
xor U23456 (N_23456,N_22878,N_22578);
or U23457 (N_23457,N_22000,N_22448);
nand U23458 (N_23458,N_22710,N_22229);
and U23459 (N_23459,N_22446,N_22963);
and U23460 (N_23460,N_22961,N_22690);
nand U23461 (N_23461,N_22007,N_22384);
and U23462 (N_23462,N_22516,N_22673);
xor U23463 (N_23463,N_22443,N_22290);
nor U23464 (N_23464,N_22777,N_22109);
xor U23465 (N_23465,N_22711,N_22053);
and U23466 (N_23466,N_22837,N_22342);
nand U23467 (N_23467,N_22893,N_22033);
nand U23468 (N_23468,N_22101,N_22112);
xnor U23469 (N_23469,N_22607,N_22361);
and U23470 (N_23470,N_22663,N_22156);
nor U23471 (N_23471,N_22580,N_22755);
nand U23472 (N_23472,N_22037,N_22696);
and U23473 (N_23473,N_22914,N_22973);
nand U23474 (N_23474,N_22306,N_22075);
and U23475 (N_23475,N_22356,N_22941);
or U23476 (N_23476,N_22540,N_22972);
nor U23477 (N_23477,N_22846,N_22713);
or U23478 (N_23478,N_22964,N_22853);
xnor U23479 (N_23479,N_22935,N_22566);
nor U23480 (N_23480,N_22180,N_22078);
or U23481 (N_23481,N_22539,N_22628);
or U23482 (N_23482,N_22472,N_22368);
and U23483 (N_23483,N_22339,N_22523);
nor U23484 (N_23484,N_22435,N_22440);
xor U23485 (N_23485,N_22215,N_22328);
nand U23486 (N_23486,N_22599,N_22352);
or U23487 (N_23487,N_22250,N_22045);
or U23488 (N_23488,N_22121,N_22674);
and U23489 (N_23489,N_22497,N_22284);
nor U23490 (N_23490,N_22233,N_22402);
nor U23491 (N_23491,N_22701,N_22350);
or U23492 (N_23492,N_22426,N_22879);
nand U23493 (N_23493,N_22046,N_22106);
or U23494 (N_23494,N_22784,N_22220);
nor U23495 (N_23495,N_22123,N_22675);
xor U23496 (N_23496,N_22521,N_22695);
xor U23497 (N_23497,N_22956,N_22541);
nand U23498 (N_23498,N_22999,N_22317);
and U23499 (N_23499,N_22530,N_22842);
and U23500 (N_23500,N_22047,N_22609);
nand U23501 (N_23501,N_22256,N_22804);
nor U23502 (N_23502,N_22460,N_22083);
xor U23503 (N_23503,N_22141,N_22330);
xor U23504 (N_23504,N_22641,N_22119);
and U23505 (N_23505,N_22844,N_22244);
or U23506 (N_23506,N_22127,N_22788);
nor U23507 (N_23507,N_22580,N_22290);
nor U23508 (N_23508,N_22625,N_22020);
nand U23509 (N_23509,N_22260,N_22793);
nand U23510 (N_23510,N_22429,N_22332);
nand U23511 (N_23511,N_22505,N_22657);
and U23512 (N_23512,N_22463,N_22328);
xnor U23513 (N_23513,N_22512,N_22050);
xor U23514 (N_23514,N_22244,N_22449);
or U23515 (N_23515,N_22666,N_22999);
and U23516 (N_23516,N_22540,N_22234);
and U23517 (N_23517,N_22395,N_22257);
and U23518 (N_23518,N_22905,N_22772);
or U23519 (N_23519,N_22982,N_22304);
nand U23520 (N_23520,N_22689,N_22105);
or U23521 (N_23521,N_22409,N_22159);
and U23522 (N_23522,N_22194,N_22118);
nor U23523 (N_23523,N_22211,N_22650);
xnor U23524 (N_23524,N_22317,N_22758);
and U23525 (N_23525,N_22584,N_22414);
nand U23526 (N_23526,N_22074,N_22663);
xor U23527 (N_23527,N_22672,N_22948);
or U23528 (N_23528,N_22086,N_22841);
xor U23529 (N_23529,N_22795,N_22200);
nor U23530 (N_23530,N_22236,N_22394);
or U23531 (N_23531,N_22391,N_22874);
or U23532 (N_23532,N_22162,N_22917);
nand U23533 (N_23533,N_22979,N_22118);
xnor U23534 (N_23534,N_22963,N_22252);
or U23535 (N_23535,N_22684,N_22196);
or U23536 (N_23536,N_22282,N_22580);
nor U23537 (N_23537,N_22603,N_22167);
and U23538 (N_23538,N_22523,N_22333);
xor U23539 (N_23539,N_22004,N_22144);
nor U23540 (N_23540,N_22678,N_22424);
nand U23541 (N_23541,N_22913,N_22702);
nor U23542 (N_23542,N_22069,N_22810);
nand U23543 (N_23543,N_22113,N_22178);
or U23544 (N_23544,N_22695,N_22569);
nand U23545 (N_23545,N_22538,N_22580);
xnor U23546 (N_23546,N_22430,N_22402);
nand U23547 (N_23547,N_22911,N_22906);
xnor U23548 (N_23548,N_22058,N_22951);
nand U23549 (N_23549,N_22719,N_22969);
nand U23550 (N_23550,N_22510,N_22481);
xor U23551 (N_23551,N_22124,N_22080);
nand U23552 (N_23552,N_22974,N_22364);
xor U23553 (N_23553,N_22992,N_22998);
xnor U23554 (N_23554,N_22360,N_22012);
or U23555 (N_23555,N_22281,N_22193);
or U23556 (N_23556,N_22292,N_22924);
and U23557 (N_23557,N_22877,N_22450);
or U23558 (N_23558,N_22877,N_22520);
or U23559 (N_23559,N_22853,N_22976);
xor U23560 (N_23560,N_22922,N_22193);
or U23561 (N_23561,N_22734,N_22690);
nor U23562 (N_23562,N_22742,N_22514);
nor U23563 (N_23563,N_22722,N_22512);
xor U23564 (N_23564,N_22192,N_22599);
nor U23565 (N_23565,N_22833,N_22379);
nor U23566 (N_23566,N_22356,N_22350);
and U23567 (N_23567,N_22379,N_22574);
xnor U23568 (N_23568,N_22532,N_22432);
nor U23569 (N_23569,N_22905,N_22057);
nor U23570 (N_23570,N_22171,N_22987);
nor U23571 (N_23571,N_22559,N_22174);
and U23572 (N_23572,N_22111,N_22709);
xnor U23573 (N_23573,N_22323,N_22644);
and U23574 (N_23574,N_22606,N_22253);
nand U23575 (N_23575,N_22972,N_22817);
and U23576 (N_23576,N_22067,N_22693);
nor U23577 (N_23577,N_22114,N_22361);
xor U23578 (N_23578,N_22772,N_22685);
xor U23579 (N_23579,N_22700,N_22374);
nor U23580 (N_23580,N_22669,N_22813);
or U23581 (N_23581,N_22856,N_22250);
or U23582 (N_23582,N_22505,N_22225);
xnor U23583 (N_23583,N_22723,N_22628);
nor U23584 (N_23584,N_22348,N_22287);
xor U23585 (N_23585,N_22534,N_22474);
and U23586 (N_23586,N_22453,N_22163);
nor U23587 (N_23587,N_22793,N_22203);
nor U23588 (N_23588,N_22062,N_22643);
xor U23589 (N_23589,N_22101,N_22984);
nand U23590 (N_23590,N_22686,N_22968);
nor U23591 (N_23591,N_22676,N_22918);
and U23592 (N_23592,N_22835,N_22068);
xor U23593 (N_23593,N_22656,N_22377);
xor U23594 (N_23594,N_22456,N_22246);
nand U23595 (N_23595,N_22166,N_22247);
or U23596 (N_23596,N_22451,N_22616);
xor U23597 (N_23597,N_22011,N_22381);
nor U23598 (N_23598,N_22995,N_22889);
xnor U23599 (N_23599,N_22714,N_22474);
or U23600 (N_23600,N_22661,N_22570);
nand U23601 (N_23601,N_22330,N_22814);
xnor U23602 (N_23602,N_22766,N_22848);
and U23603 (N_23603,N_22142,N_22657);
or U23604 (N_23604,N_22770,N_22521);
nor U23605 (N_23605,N_22013,N_22493);
or U23606 (N_23606,N_22301,N_22910);
or U23607 (N_23607,N_22346,N_22245);
xnor U23608 (N_23608,N_22183,N_22599);
and U23609 (N_23609,N_22466,N_22733);
nor U23610 (N_23610,N_22298,N_22283);
xor U23611 (N_23611,N_22573,N_22254);
xnor U23612 (N_23612,N_22837,N_22391);
nand U23613 (N_23613,N_22145,N_22677);
or U23614 (N_23614,N_22535,N_22230);
or U23615 (N_23615,N_22761,N_22756);
nor U23616 (N_23616,N_22264,N_22099);
nand U23617 (N_23617,N_22993,N_22543);
or U23618 (N_23618,N_22181,N_22557);
xor U23619 (N_23619,N_22233,N_22739);
and U23620 (N_23620,N_22660,N_22346);
nand U23621 (N_23621,N_22760,N_22929);
nand U23622 (N_23622,N_22592,N_22121);
nor U23623 (N_23623,N_22511,N_22165);
and U23624 (N_23624,N_22345,N_22799);
nor U23625 (N_23625,N_22962,N_22612);
xor U23626 (N_23626,N_22475,N_22898);
and U23627 (N_23627,N_22691,N_22614);
nand U23628 (N_23628,N_22375,N_22217);
or U23629 (N_23629,N_22487,N_22034);
nor U23630 (N_23630,N_22333,N_22351);
nand U23631 (N_23631,N_22546,N_22088);
nor U23632 (N_23632,N_22475,N_22125);
and U23633 (N_23633,N_22567,N_22371);
xor U23634 (N_23634,N_22218,N_22616);
nor U23635 (N_23635,N_22124,N_22561);
or U23636 (N_23636,N_22393,N_22446);
and U23637 (N_23637,N_22492,N_22499);
and U23638 (N_23638,N_22220,N_22770);
xor U23639 (N_23639,N_22023,N_22150);
and U23640 (N_23640,N_22106,N_22559);
or U23641 (N_23641,N_22752,N_22788);
nor U23642 (N_23642,N_22572,N_22169);
nand U23643 (N_23643,N_22190,N_22617);
or U23644 (N_23644,N_22260,N_22613);
nor U23645 (N_23645,N_22331,N_22096);
or U23646 (N_23646,N_22401,N_22150);
nor U23647 (N_23647,N_22802,N_22610);
or U23648 (N_23648,N_22194,N_22816);
or U23649 (N_23649,N_22272,N_22078);
nand U23650 (N_23650,N_22192,N_22181);
xor U23651 (N_23651,N_22064,N_22038);
nor U23652 (N_23652,N_22505,N_22700);
and U23653 (N_23653,N_22565,N_22378);
xor U23654 (N_23654,N_22769,N_22099);
nor U23655 (N_23655,N_22464,N_22984);
and U23656 (N_23656,N_22534,N_22029);
nor U23657 (N_23657,N_22961,N_22140);
and U23658 (N_23658,N_22136,N_22709);
nor U23659 (N_23659,N_22051,N_22401);
or U23660 (N_23660,N_22289,N_22871);
or U23661 (N_23661,N_22398,N_22922);
nand U23662 (N_23662,N_22363,N_22397);
nand U23663 (N_23663,N_22601,N_22832);
and U23664 (N_23664,N_22532,N_22262);
nor U23665 (N_23665,N_22103,N_22057);
or U23666 (N_23666,N_22122,N_22069);
or U23667 (N_23667,N_22100,N_22946);
or U23668 (N_23668,N_22109,N_22642);
nand U23669 (N_23669,N_22689,N_22387);
xnor U23670 (N_23670,N_22237,N_22197);
nand U23671 (N_23671,N_22838,N_22491);
or U23672 (N_23672,N_22236,N_22685);
or U23673 (N_23673,N_22740,N_22046);
or U23674 (N_23674,N_22386,N_22244);
and U23675 (N_23675,N_22740,N_22438);
or U23676 (N_23676,N_22258,N_22837);
and U23677 (N_23677,N_22126,N_22784);
nor U23678 (N_23678,N_22737,N_22599);
xor U23679 (N_23679,N_22578,N_22593);
nand U23680 (N_23680,N_22789,N_22595);
nand U23681 (N_23681,N_22459,N_22983);
nand U23682 (N_23682,N_22649,N_22139);
or U23683 (N_23683,N_22631,N_22903);
or U23684 (N_23684,N_22526,N_22185);
xnor U23685 (N_23685,N_22268,N_22685);
or U23686 (N_23686,N_22556,N_22663);
nor U23687 (N_23687,N_22309,N_22261);
nor U23688 (N_23688,N_22392,N_22240);
xor U23689 (N_23689,N_22722,N_22578);
or U23690 (N_23690,N_22393,N_22658);
nand U23691 (N_23691,N_22340,N_22250);
and U23692 (N_23692,N_22744,N_22226);
and U23693 (N_23693,N_22310,N_22901);
and U23694 (N_23694,N_22722,N_22870);
nand U23695 (N_23695,N_22019,N_22254);
or U23696 (N_23696,N_22811,N_22991);
xor U23697 (N_23697,N_22021,N_22632);
or U23698 (N_23698,N_22357,N_22404);
nand U23699 (N_23699,N_22897,N_22367);
or U23700 (N_23700,N_22315,N_22600);
nand U23701 (N_23701,N_22031,N_22108);
nor U23702 (N_23702,N_22730,N_22228);
and U23703 (N_23703,N_22732,N_22044);
nand U23704 (N_23704,N_22175,N_22289);
nand U23705 (N_23705,N_22815,N_22496);
and U23706 (N_23706,N_22974,N_22342);
or U23707 (N_23707,N_22785,N_22091);
nand U23708 (N_23708,N_22883,N_22539);
nor U23709 (N_23709,N_22585,N_22856);
and U23710 (N_23710,N_22952,N_22497);
nor U23711 (N_23711,N_22119,N_22262);
xor U23712 (N_23712,N_22958,N_22912);
nand U23713 (N_23713,N_22438,N_22007);
or U23714 (N_23714,N_22015,N_22918);
or U23715 (N_23715,N_22497,N_22294);
nor U23716 (N_23716,N_22521,N_22133);
and U23717 (N_23717,N_22969,N_22500);
or U23718 (N_23718,N_22640,N_22503);
xor U23719 (N_23719,N_22176,N_22830);
and U23720 (N_23720,N_22965,N_22080);
or U23721 (N_23721,N_22478,N_22885);
nand U23722 (N_23722,N_22428,N_22091);
or U23723 (N_23723,N_22840,N_22249);
and U23724 (N_23724,N_22497,N_22915);
xnor U23725 (N_23725,N_22348,N_22100);
or U23726 (N_23726,N_22492,N_22055);
and U23727 (N_23727,N_22180,N_22099);
nor U23728 (N_23728,N_22512,N_22098);
xor U23729 (N_23729,N_22007,N_22470);
nor U23730 (N_23730,N_22902,N_22705);
and U23731 (N_23731,N_22088,N_22762);
nor U23732 (N_23732,N_22275,N_22216);
xor U23733 (N_23733,N_22475,N_22370);
and U23734 (N_23734,N_22974,N_22340);
and U23735 (N_23735,N_22345,N_22754);
and U23736 (N_23736,N_22384,N_22497);
and U23737 (N_23737,N_22050,N_22962);
xnor U23738 (N_23738,N_22402,N_22382);
nand U23739 (N_23739,N_22274,N_22780);
and U23740 (N_23740,N_22640,N_22806);
nor U23741 (N_23741,N_22939,N_22561);
or U23742 (N_23742,N_22474,N_22213);
xnor U23743 (N_23743,N_22174,N_22832);
and U23744 (N_23744,N_22879,N_22237);
nand U23745 (N_23745,N_22725,N_22861);
xor U23746 (N_23746,N_22189,N_22757);
or U23747 (N_23747,N_22600,N_22394);
xor U23748 (N_23748,N_22680,N_22354);
nor U23749 (N_23749,N_22985,N_22871);
and U23750 (N_23750,N_22052,N_22241);
nand U23751 (N_23751,N_22689,N_22135);
and U23752 (N_23752,N_22042,N_22319);
and U23753 (N_23753,N_22766,N_22030);
or U23754 (N_23754,N_22922,N_22114);
xor U23755 (N_23755,N_22700,N_22656);
xnor U23756 (N_23756,N_22183,N_22836);
xor U23757 (N_23757,N_22398,N_22022);
nor U23758 (N_23758,N_22953,N_22791);
xor U23759 (N_23759,N_22778,N_22720);
or U23760 (N_23760,N_22305,N_22279);
and U23761 (N_23761,N_22126,N_22858);
nand U23762 (N_23762,N_22618,N_22139);
and U23763 (N_23763,N_22810,N_22361);
nor U23764 (N_23764,N_22178,N_22139);
and U23765 (N_23765,N_22587,N_22139);
xnor U23766 (N_23766,N_22108,N_22513);
nand U23767 (N_23767,N_22033,N_22928);
nand U23768 (N_23768,N_22427,N_22324);
nor U23769 (N_23769,N_22248,N_22031);
or U23770 (N_23770,N_22114,N_22238);
and U23771 (N_23771,N_22850,N_22636);
and U23772 (N_23772,N_22971,N_22463);
nand U23773 (N_23773,N_22227,N_22110);
nand U23774 (N_23774,N_22779,N_22234);
xor U23775 (N_23775,N_22954,N_22239);
nor U23776 (N_23776,N_22895,N_22088);
or U23777 (N_23777,N_22021,N_22638);
nand U23778 (N_23778,N_22796,N_22042);
xor U23779 (N_23779,N_22497,N_22078);
and U23780 (N_23780,N_22667,N_22702);
or U23781 (N_23781,N_22234,N_22478);
xor U23782 (N_23782,N_22120,N_22016);
or U23783 (N_23783,N_22435,N_22271);
or U23784 (N_23784,N_22376,N_22698);
nor U23785 (N_23785,N_22155,N_22383);
xor U23786 (N_23786,N_22484,N_22653);
nand U23787 (N_23787,N_22815,N_22861);
or U23788 (N_23788,N_22090,N_22825);
nand U23789 (N_23789,N_22744,N_22599);
nand U23790 (N_23790,N_22880,N_22245);
or U23791 (N_23791,N_22243,N_22129);
or U23792 (N_23792,N_22244,N_22145);
or U23793 (N_23793,N_22647,N_22937);
or U23794 (N_23794,N_22673,N_22745);
and U23795 (N_23795,N_22973,N_22390);
nor U23796 (N_23796,N_22274,N_22005);
nor U23797 (N_23797,N_22443,N_22784);
nand U23798 (N_23798,N_22327,N_22345);
or U23799 (N_23799,N_22738,N_22352);
and U23800 (N_23800,N_22413,N_22606);
xnor U23801 (N_23801,N_22057,N_22901);
and U23802 (N_23802,N_22008,N_22894);
xnor U23803 (N_23803,N_22192,N_22934);
xor U23804 (N_23804,N_22284,N_22583);
or U23805 (N_23805,N_22639,N_22846);
nand U23806 (N_23806,N_22868,N_22790);
nor U23807 (N_23807,N_22567,N_22117);
and U23808 (N_23808,N_22317,N_22227);
nor U23809 (N_23809,N_22396,N_22169);
or U23810 (N_23810,N_22391,N_22699);
xor U23811 (N_23811,N_22489,N_22498);
nor U23812 (N_23812,N_22160,N_22407);
or U23813 (N_23813,N_22343,N_22919);
nand U23814 (N_23814,N_22096,N_22356);
nor U23815 (N_23815,N_22684,N_22728);
or U23816 (N_23816,N_22494,N_22345);
or U23817 (N_23817,N_22228,N_22391);
xnor U23818 (N_23818,N_22356,N_22001);
nand U23819 (N_23819,N_22393,N_22831);
nand U23820 (N_23820,N_22024,N_22855);
and U23821 (N_23821,N_22615,N_22452);
and U23822 (N_23822,N_22401,N_22908);
and U23823 (N_23823,N_22232,N_22605);
xor U23824 (N_23824,N_22976,N_22762);
nor U23825 (N_23825,N_22978,N_22609);
xor U23826 (N_23826,N_22869,N_22980);
or U23827 (N_23827,N_22841,N_22792);
nand U23828 (N_23828,N_22174,N_22733);
nor U23829 (N_23829,N_22731,N_22537);
or U23830 (N_23830,N_22169,N_22393);
and U23831 (N_23831,N_22845,N_22629);
xor U23832 (N_23832,N_22786,N_22179);
or U23833 (N_23833,N_22705,N_22393);
nor U23834 (N_23834,N_22306,N_22067);
xnor U23835 (N_23835,N_22865,N_22052);
and U23836 (N_23836,N_22893,N_22513);
and U23837 (N_23837,N_22666,N_22657);
nand U23838 (N_23838,N_22359,N_22512);
nor U23839 (N_23839,N_22440,N_22371);
or U23840 (N_23840,N_22993,N_22502);
or U23841 (N_23841,N_22131,N_22167);
xor U23842 (N_23842,N_22734,N_22745);
nand U23843 (N_23843,N_22458,N_22006);
or U23844 (N_23844,N_22482,N_22532);
nand U23845 (N_23845,N_22701,N_22065);
or U23846 (N_23846,N_22604,N_22190);
or U23847 (N_23847,N_22834,N_22783);
and U23848 (N_23848,N_22942,N_22616);
xnor U23849 (N_23849,N_22350,N_22248);
and U23850 (N_23850,N_22795,N_22417);
nor U23851 (N_23851,N_22973,N_22398);
nand U23852 (N_23852,N_22808,N_22367);
and U23853 (N_23853,N_22200,N_22536);
nand U23854 (N_23854,N_22263,N_22965);
and U23855 (N_23855,N_22938,N_22597);
and U23856 (N_23856,N_22627,N_22408);
nor U23857 (N_23857,N_22573,N_22589);
or U23858 (N_23858,N_22013,N_22114);
xnor U23859 (N_23859,N_22012,N_22884);
or U23860 (N_23860,N_22044,N_22969);
and U23861 (N_23861,N_22593,N_22170);
xnor U23862 (N_23862,N_22743,N_22213);
nor U23863 (N_23863,N_22228,N_22926);
or U23864 (N_23864,N_22763,N_22685);
and U23865 (N_23865,N_22585,N_22704);
nor U23866 (N_23866,N_22705,N_22761);
nor U23867 (N_23867,N_22441,N_22688);
xnor U23868 (N_23868,N_22733,N_22580);
or U23869 (N_23869,N_22210,N_22848);
and U23870 (N_23870,N_22033,N_22439);
xor U23871 (N_23871,N_22795,N_22400);
xnor U23872 (N_23872,N_22381,N_22042);
or U23873 (N_23873,N_22824,N_22464);
xnor U23874 (N_23874,N_22571,N_22126);
xor U23875 (N_23875,N_22374,N_22595);
nand U23876 (N_23876,N_22880,N_22959);
and U23877 (N_23877,N_22075,N_22769);
nand U23878 (N_23878,N_22093,N_22703);
xnor U23879 (N_23879,N_22949,N_22053);
xor U23880 (N_23880,N_22858,N_22400);
and U23881 (N_23881,N_22077,N_22923);
nand U23882 (N_23882,N_22305,N_22253);
or U23883 (N_23883,N_22683,N_22063);
nand U23884 (N_23884,N_22275,N_22619);
and U23885 (N_23885,N_22445,N_22659);
and U23886 (N_23886,N_22001,N_22456);
or U23887 (N_23887,N_22995,N_22871);
xor U23888 (N_23888,N_22311,N_22199);
xnor U23889 (N_23889,N_22066,N_22510);
and U23890 (N_23890,N_22826,N_22897);
xor U23891 (N_23891,N_22575,N_22640);
nand U23892 (N_23892,N_22988,N_22432);
nor U23893 (N_23893,N_22256,N_22888);
and U23894 (N_23894,N_22169,N_22386);
xnor U23895 (N_23895,N_22226,N_22076);
nand U23896 (N_23896,N_22475,N_22567);
or U23897 (N_23897,N_22277,N_22275);
or U23898 (N_23898,N_22734,N_22348);
or U23899 (N_23899,N_22454,N_22471);
nand U23900 (N_23900,N_22254,N_22575);
nand U23901 (N_23901,N_22259,N_22918);
nand U23902 (N_23902,N_22201,N_22848);
nand U23903 (N_23903,N_22517,N_22720);
and U23904 (N_23904,N_22921,N_22916);
and U23905 (N_23905,N_22435,N_22599);
xnor U23906 (N_23906,N_22391,N_22407);
xor U23907 (N_23907,N_22802,N_22962);
nand U23908 (N_23908,N_22763,N_22772);
nor U23909 (N_23909,N_22200,N_22555);
and U23910 (N_23910,N_22649,N_22904);
nor U23911 (N_23911,N_22923,N_22237);
xnor U23912 (N_23912,N_22323,N_22795);
xnor U23913 (N_23913,N_22592,N_22108);
nor U23914 (N_23914,N_22175,N_22946);
and U23915 (N_23915,N_22820,N_22665);
nand U23916 (N_23916,N_22105,N_22328);
xor U23917 (N_23917,N_22834,N_22675);
nor U23918 (N_23918,N_22278,N_22983);
nand U23919 (N_23919,N_22211,N_22859);
nand U23920 (N_23920,N_22295,N_22619);
or U23921 (N_23921,N_22720,N_22530);
nand U23922 (N_23922,N_22643,N_22618);
and U23923 (N_23923,N_22270,N_22495);
xor U23924 (N_23924,N_22659,N_22522);
and U23925 (N_23925,N_22661,N_22506);
and U23926 (N_23926,N_22820,N_22707);
or U23927 (N_23927,N_22637,N_22802);
or U23928 (N_23928,N_22898,N_22124);
and U23929 (N_23929,N_22329,N_22686);
nor U23930 (N_23930,N_22277,N_22910);
xnor U23931 (N_23931,N_22149,N_22055);
and U23932 (N_23932,N_22193,N_22894);
nor U23933 (N_23933,N_22136,N_22938);
nand U23934 (N_23934,N_22425,N_22590);
nor U23935 (N_23935,N_22198,N_22588);
and U23936 (N_23936,N_22037,N_22779);
nor U23937 (N_23937,N_22529,N_22005);
nor U23938 (N_23938,N_22830,N_22429);
and U23939 (N_23939,N_22015,N_22310);
nor U23940 (N_23940,N_22751,N_22163);
nor U23941 (N_23941,N_22332,N_22956);
nor U23942 (N_23942,N_22389,N_22225);
xor U23943 (N_23943,N_22033,N_22175);
and U23944 (N_23944,N_22397,N_22437);
nand U23945 (N_23945,N_22871,N_22128);
xnor U23946 (N_23946,N_22649,N_22603);
or U23947 (N_23947,N_22957,N_22904);
or U23948 (N_23948,N_22645,N_22073);
nor U23949 (N_23949,N_22170,N_22087);
and U23950 (N_23950,N_22840,N_22051);
or U23951 (N_23951,N_22332,N_22333);
nor U23952 (N_23952,N_22688,N_22857);
and U23953 (N_23953,N_22457,N_22264);
xnor U23954 (N_23954,N_22933,N_22383);
and U23955 (N_23955,N_22629,N_22079);
or U23956 (N_23956,N_22257,N_22814);
nor U23957 (N_23957,N_22436,N_22635);
or U23958 (N_23958,N_22519,N_22735);
nor U23959 (N_23959,N_22147,N_22913);
and U23960 (N_23960,N_22910,N_22978);
nor U23961 (N_23961,N_22005,N_22537);
nor U23962 (N_23962,N_22606,N_22554);
and U23963 (N_23963,N_22879,N_22960);
nand U23964 (N_23964,N_22072,N_22166);
and U23965 (N_23965,N_22990,N_22951);
xor U23966 (N_23966,N_22430,N_22455);
xor U23967 (N_23967,N_22006,N_22359);
nand U23968 (N_23968,N_22993,N_22469);
xor U23969 (N_23969,N_22524,N_22678);
nor U23970 (N_23970,N_22632,N_22721);
nand U23971 (N_23971,N_22979,N_22912);
xor U23972 (N_23972,N_22746,N_22172);
and U23973 (N_23973,N_22443,N_22432);
nand U23974 (N_23974,N_22521,N_22509);
nor U23975 (N_23975,N_22696,N_22278);
and U23976 (N_23976,N_22784,N_22828);
nand U23977 (N_23977,N_22459,N_22511);
and U23978 (N_23978,N_22568,N_22941);
nor U23979 (N_23979,N_22820,N_22068);
nand U23980 (N_23980,N_22266,N_22741);
nand U23981 (N_23981,N_22033,N_22409);
and U23982 (N_23982,N_22389,N_22217);
nor U23983 (N_23983,N_22455,N_22140);
nand U23984 (N_23984,N_22520,N_22020);
xor U23985 (N_23985,N_22699,N_22604);
xnor U23986 (N_23986,N_22999,N_22833);
and U23987 (N_23987,N_22461,N_22287);
nor U23988 (N_23988,N_22673,N_22383);
and U23989 (N_23989,N_22826,N_22627);
nand U23990 (N_23990,N_22153,N_22170);
nand U23991 (N_23991,N_22816,N_22182);
and U23992 (N_23992,N_22894,N_22139);
nor U23993 (N_23993,N_22740,N_22962);
and U23994 (N_23994,N_22693,N_22647);
nand U23995 (N_23995,N_22850,N_22745);
or U23996 (N_23996,N_22375,N_22000);
nand U23997 (N_23997,N_22978,N_22121);
nor U23998 (N_23998,N_22085,N_22140);
xnor U23999 (N_23999,N_22094,N_22836);
and U24000 (N_24000,N_23710,N_23187);
xnor U24001 (N_24001,N_23237,N_23361);
and U24002 (N_24002,N_23828,N_23162);
xnor U24003 (N_24003,N_23435,N_23570);
nand U24004 (N_24004,N_23822,N_23697);
and U24005 (N_24005,N_23809,N_23795);
nand U24006 (N_24006,N_23036,N_23636);
nor U24007 (N_24007,N_23356,N_23083);
or U24008 (N_24008,N_23864,N_23902);
nor U24009 (N_24009,N_23528,N_23645);
nor U24010 (N_24010,N_23625,N_23722);
xnor U24011 (N_24011,N_23772,N_23825);
and U24012 (N_24012,N_23583,N_23723);
xor U24013 (N_24013,N_23863,N_23171);
nor U24014 (N_24014,N_23299,N_23285);
xor U24015 (N_24015,N_23151,N_23935);
xnor U24016 (N_24016,N_23951,N_23911);
nor U24017 (N_24017,N_23368,N_23553);
or U24018 (N_24018,N_23531,N_23229);
or U24019 (N_24019,N_23381,N_23076);
or U24020 (N_24020,N_23947,N_23558);
and U24021 (N_24021,N_23526,N_23439);
or U24022 (N_24022,N_23120,N_23525);
xor U24023 (N_24023,N_23853,N_23923);
nor U24024 (N_24024,N_23071,N_23750);
nand U24025 (N_24025,N_23228,N_23728);
nand U24026 (N_24026,N_23634,N_23061);
nand U24027 (N_24027,N_23040,N_23980);
nor U24028 (N_24028,N_23465,N_23388);
nor U24029 (N_24029,N_23940,N_23370);
xnor U24030 (N_24030,N_23939,N_23736);
or U24031 (N_24031,N_23610,N_23340);
nor U24032 (N_24032,N_23762,N_23430);
nand U24033 (N_24033,N_23290,N_23433);
nand U24034 (N_24034,N_23358,N_23894);
xor U24035 (N_24035,N_23956,N_23986);
xor U24036 (N_24036,N_23378,N_23487);
xnor U24037 (N_24037,N_23540,N_23987);
nor U24038 (N_24038,N_23860,N_23932);
nand U24039 (N_24039,N_23605,N_23600);
nor U24040 (N_24040,N_23993,N_23239);
xor U24041 (N_24041,N_23963,N_23738);
or U24042 (N_24042,N_23573,N_23082);
or U24043 (N_24043,N_23387,N_23760);
or U24044 (N_24044,N_23617,N_23431);
xnor U24045 (N_24045,N_23154,N_23359);
or U24046 (N_24046,N_23618,N_23020);
and U24047 (N_24047,N_23885,N_23862);
xnor U24048 (N_24048,N_23308,N_23018);
nor U24049 (N_24049,N_23629,N_23702);
nor U24050 (N_24050,N_23852,N_23635);
nand U24051 (N_24051,N_23765,N_23786);
nor U24052 (N_24052,N_23950,N_23432);
xor U24053 (N_24053,N_23177,N_23596);
or U24054 (N_24054,N_23405,N_23063);
and U24055 (N_24055,N_23633,N_23773);
nand U24056 (N_24056,N_23218,N_23066);
nor U24057 (N_24057,N_23791,N_23444);
xnor U24058 (N_24058,N_23344,N_23812);
xor U24059 (N_24059,N_23555,N_23365);
or U24060 (N_24060,N_23719,N_23623);
nor U24061 (N_24061,N_23478,N_23582);
nand U24062 (N_24062,N_23148,N_23797);
nor U24063 (N_24063,N_23204,N_23622);
and U24064 (N_24064,N_23014,N_23088);
nor U24065 (N_24065,N_23944,N_23805);
and U24066 (N_24066,N_23459,N_23338);
nand U24067 (N_24067,N_23499,N_23657);
nand U24068 (N_24068,N_23630,N_23476);
xnor U24069 (N_24069,N_23469,N_23390);
xor U24070 (N_24070,N_23073,N_23845);
or U24071 (N_24071,N_23671,N_23998);
and U24072 (N_24072,N_23628,N_23116);
and U24073 (N_24073,N_23727,N_23042);
xor U24074 (N_24074,N_23079,N_23699);
nand U24075 (N_24075,N_23690,N_23906);
nor U24076 (N_24076,N_23578,N_23128);
nand U24077 (N_24077,N_23122,N_23245);
or U24078 (N_24078,N_23008,N_23592);
nand U24079 (N_24079,N_23134,N_23886);
xnor U24080 (N_24080,N_23757,N_23114);
or U24081 (N_24081,N_23002,N_23590);
xor U24082 (N_24082,N_23241,N_23734);
xnor U24083 (N_24083,N_23900,N_23268);
xnor U24084 (N_24084,N_23659,N_23203);
or U24085 (N_24085,N_23050,N_23824);
or U24086 (N_24086,N_23047,N_23997);
nand U24087 (N_24087,N_23319,N_23927);
nor U24088 (N_24088,N_23826,N_23137);
and U24089 (N_24089,N_23252,N_23312);
xnor U24090 (N_24090,N_23733,N_23904);
xor U24091 (N_24091,N_23631,N_23856);
nor U24092 (N_24092,N_23747,N_23677);
nand U24093 (N_24093,N_23070,N_23206);
xor U24094 (N_24094,N_23872,N_23039);
or U24095 (N_24095,N_23286,N_23157);
nand U24096 (N_24096,N_23191,N_23649);
xnor U24097 (N_24097,N_23403,N_23059);
and U24098 (N_24098,N_23785,N_23244);
nor U24099 (N_24099,N_23873,N_23982);
nand U24100 (N_24100,N_23011,N_23876);
xor U24101 (N_24101,N_23353,N_23597);
or U24102 (N_24102,N_23505,N_23411);
or U24103 (N_24103,N_23049,N_23816);
nand U24104 (N_24104,N_23491,N_23326);
nand U24105 (N_24105,N_23046,N_23546);
nand U24106 (N_24106,N_23243,N_23043);
xor U24107 (N_24107,N_23003,N_23793);
xor U24108 (N_24108,N_23041,N_23027);
or U24109 (N_24109,N_23075,N_23840);
nand U24110 (N_24110,N_23682,N_23990);
nor U24111 (N_24111,N_23096,N_23751);
or U24112 (N_24112,N_23077,N_23099);
or U24113 (N_24113,N_23847,N_23424);
and U24114 (N_24114,N_23695,N_23908);
or U24115 (N_24115,N_23588,N_23918);
nor U24116 (N_24116,N_23930,N_23305);
xor U24117 (N_24117,N_23668,N_23410);
xnor U24118 (N_24118,N_23521,N_23745);
nand U24119 (N_24119,N_23587,N_23084);
nand U24120 (N_24120,N_23579,N_23145);
and U24121 (N_24121,N_23804,N_23067);
xor U24122 (N_24122,N_23320,N_23779);
xnor U24123 (N_24123,N_23961,N_23953);
or U24124 (N_24124,N_23504,N_23337);
nand U24125 (N_24125,N_23163,N_23194);
or U24126 (N_24126,N_23849,N_23983);
and U24127 (N_24127,N_23179,N_23161);
or U24128 (N_24128,N_23472,N_23445);
nand U24129 (N_24129,N_23141,N_23520);
nand U24130 (N_24130,N_23292,N_23153);
or U24131 (N_24131,N_23341,N_23038);
and U24132 (N_24132,N_23523,N_23580);
xnor U24133 (N_24133,N_23543,N_23352);
xnor U24134 (N_24134,N_23574,N_23720);
nor U24135 (N_24135,N_23730,N_23934);
or U24136 (N_24136,N_23267,N_23530);
and U24137 (N_24137,N_23575,N_23330);
and U24138 (N_24138,N_23484,N_23205);
or U24139 (N_24139,N_23461,N_23185);
or U24140 (N_24140,N_23278,N_23064);
xor U24141 (N_24141,N_23373,N_23781);
xor U24142 (N_24142,N_23182,N_23032);
xnor U24143 (N_24143,N_23264,N_23614);
nand U24144 (N_24144,N_23251,N_23887);
xnor U24145 (N_24145,N_23334,N_23989);
nand U24146 (N_24146,N_23955,N_23113);
nor U24147 (N_24147,N_23829,N_23542);
nand U24148 (N_24148,N_23641,N_23080);
and U24149 (N_24149,N_23089,N_23306);
xnor U24150 (N_24150,N_23313,N_23323);
nor U24151 (N_24151,N_23721,N_23057);
nand U24152 (N_24152,N_23053,N_23767);
or U24153 (N_24153,N_23941,N_23324);
or U24154 (N_24154,N_23518,N_23201);
and U24155 (N_24155,N_23716,N_23207);
or U24156 (N_24156,N_23477,N_23907);
nand U24157 (N_24157,N_23665,N_23310);
xnor U24158 (N_24158,N_23492,N_23425);
xnor U24159 (N_24159,N_23656,N_23176);
and U24160 (N_24160,N_23969,N_23170);
or U24161 (N_24161,N_23679,N_23266);
or U24162 (N_24162,N_23529,N_23115);
nand U24163 (N_24163,N_23369,N_23893);
nand U24164 (N_24164,N_23848,N_23602);
and U24165 (N_24165,N_23945,N_23770);
xor U24166 (N_24166,N_23005,N_23929);
or U24167 (N_24167,N_23235,N_23339);
or U24168 (N_24168,N_23992,N_23220);
xor U24169 (N_24169,N_23263,N_23458);
nor U24170 (N_24170,N_23619,N_23835);
and U24171 (N_24171,N_23783,N_23891);
nor U24172 (N_24172,N_23650,N_23216);
and U24173 (N_24173,N_23644,N_23949);
or U24174 (N_24174,N_23703,N_23627);
and U24175 (N_24175,N_23680,N_23815);
or U24176 (N_24176,N_23468,N_23150);
nand U24177 (N_24177,N_23744,N_23357);
xnor U24178 (N_24178,N_23706,N_23759);
nor U24179 (N_24179,N_23401,N_23565);
and U24180 (N_24180,N_23513,N_23283);
nor U24181 (N_24181,N_23909,N_23265);
xnor U24182 (N_24182,N_23708,N_23867);
nor U24183 (N_24183,N_23015,N_23965);
nand U24184 (N_24184,N_23796,N_23117);
and U24185 (N_24185,N_23282,N_23561);
nor U24186 (N_24186,N_23470,N_23807);
or U24187 (N_24187,N_23475,N_23350);
nor U24188 (N_24188,N_23414,N_23551);
or U24189 (N_24189,N_23924,N_23097);
nand U24190 (N_24190,N_23164,N_23506);
nand U24191 (N_24191,N_23914,N_23510);
nand U24192 (N_24192,N_23557,N_23764);
nor U24193 (N_24193,N_23107,N_23234);
nand U24194 (N_24194,N_23402,N_23545);
xnor U24195 (N_24195,N_23919,N_23156);
xor U24196 (N_24196,N_23763,N_23406);
and U24197 (N_24197,N_23321,N_23654);
nand U24198 (N_24198,N_23496,N_23591);
or U24199 (N_24199,N_23712,N_23422);
xnor U24200 (N_24200,N_23714,N_23776);
or U24201 (N_24201,N_23599,N_23256);
xnor U24202 (N_24202,N_23780,N_23878);
nor U24203 (N_24203,N_23186,N_23547);
xor U24204 (N_24204,N_23869,N_23731);
and U24205 (N_24205,N_23495,N_23322);
and U24206 (N_24206,N_23819,N_23537);
and U24207 (N_24207,N_23771,N_23604);
and U24208 (N_24208,N_23655,N_23007);
or U24209 (N_24209,N_23926,N_23143);
xor U24210 (N_24210,N_23126,N_23407);
nand U24211 (N_24211,N_23823,N_23144);
or U24212 (N_24212,N_23613,N_23742);
nor U24213 (N_24213,N_23977,N_23632);
and U24214 (N_24214,N_23412,N_23442);
nor U24215 (N_24215,N_23087,N_23512);
xor U24216 (N_24216,N_23684,N_23379);
xor U24217 (N_24217,N_23519,N_23960);
nor U24218 (N_24218,N_23219,N_23010);
or U24219 (N_24219,N_23548,N_23846);
or U24220 (N_24220,N_23971,N_23693);
nand U24221 (N_24221,N_23647,N_23328);
nand U24222 (N_24222,N_23500,N_23367);
nor U24223 (N_24223,N_23225,N_23464);
or U24224 (N_24224,N_23090,N_23291);
or U24225 (N_24225,N_23842,N_23777);
nor U24226 (N_24226,N_23384,N_23451);
nor U24227 (N_24227,N_23094,N_23417);
nor U24228 (N_24228,N_23189,N_23917);
xor U24229 (N_24229,N_23851,N_23473);
nor U24230 (N_24230,N_23678,N_23515);
and U24231 (N_24231,N_23025,N_23511);
nor U24232 (N_24232,N_23843,N_23142);
xnor U24233 (N_24233,N_23584,N_23966);
xnor U24234 (N_24234,N_23389,N_23118);
xnor U24235 (N_24235,N_23922,N_23101);
xor U24236 (N_24236,N_23810,N_23952);
and U24237 (N_24237,N_23022,N_23754);
and U24238 (N_24238,N_23503,N_23016);
and U24239 (N_24239,N_23972,N_23131);
nand U24240 (N_24240,N_23300,N_23676);
nand U24241 (N_24241,N_23827,N_23211);
nor U24242 (N_24242,N_23688,N_23769);
or U24243 (N_24243,N_23385,N_23937);
and U24244 (N_24244,N_23253,N_23416);
or U24245 (N_24245,N_23446,N_23355);
xnor U24246 (N_24246,N_23261,N_23569);
nand U24247 (N_24247,N_23844,N_23274);
and U24248 (N_24248,N_23527,N_23399);
nor U24249 (N_24249,N_23741,N_23994);
xor U24250 (N_24250,N_23559,N_23535);
nand U24251 (N_24251,N_23354,N_23607);
and U24252 (N_24252,N_23861,N_23169);
xnor U24253 (N_24253,N_23901,N_23912);
and U24254 (N_24254,N_23766,N_23611);
nor U24255 (N_24255,N_23294,N_23086);
and U24256 (N_24256,N_23098,N_23035);
xor U24257 (N_24257,N_23858,N_23124);
nand U24258 (N_24258,N_23013,N_23288);
and U24259 (N_24259,N_23774,N_23670);
nand U24260 (N_24260,N_23434,N_23105);
nor U24261 (N_24261,N_23441,N_23563);
xor U24262 (N_24262,N_23335,N_23497);
or U24263 (N_24263,N_23889,N_23111);
xnor U24264 (N_24264,N_23467,N_23481);
xor U24265 (N_24265,N_23638,N_23713);
xnor U24266 (N_24266,N_23250,N_23806);
nand U24267 (N_24267,N_23155,N_23874);
or U24268 (N_24268,N_23855,N_23023);
xor U24269 (N_24269,N_23062,N_23593);
nor U24270 (N_24270,N_23740,N_23167);
xor U24271 (N_24271,N_23129,N_23314);
nand U24272 (N_24272,N_23995,N_23209);
nor U24273 (N_24273,N_23637,N_23502);
and U24274 (N_24274,N_23247,N_23875);
xnor U24275 (N_24275,N_23149,N_23801);
nor U24276 (N_24276,N_23761,N_23200);
nor U24277 (N_24277,N_23303,N_23964);
xor U24278 (N_24278,N_23746,N_23836);
or U24279 (N_24279,N_23471,N_23585);
or U24280 (N_24280,N_23538,N_23711);
xnor U24281 (N_24281,N_23653,N_23715);
or U24282 (N_24282,N_23662,N_23298);
xnor U24283 (N_24283,N_23516,N_23556);
nand U24284 (N_24284,N_23452,N_23643);
and U24285 (N_24285,N_23705,N_23749);
nor U24286 (N_24286,N_23102,N_23696);
and U24287 (N_24287,N_23393,N_23287);
or U24288 (N_24288,N_23661,N_23501);
xnor U24289 (N_24289,N_23160,N_23377);
and U24290 (N_24290,N_23349,N_23884);
xnor U24291 (N_24291,N_23672,N_23180);
or U24292 (N_24292,N_23418,N_23508);
nor U24293 (N_24293,N_23685,N_23438);
xor U24294 (N_24294,N_23429,N_23536);
xnor U24295 (N_24295,N_23348,N_23044);
or U24296 (N_24296,N_23382,N_23052);
and U24297 (N_24297,N_23897,N_23985);
or U24298 (N_24298,N_23928,N_23598);
xnor U24299 (N_24299,N_23450,N_23514);
nor U24300 (N_24300,N_23273,N_23567);
and U24301 (N_24301,N_23954,N_23594);
nor U24302 (N_24302,N_23640,N_23970);
and U24303 (N_24303,N_23554,N_23109);
nand U24304 (N_24304,N_23307,N_23346);
nor U24305 (N_24305,N_23480,N_23802);
nand U24306 (N_24306,N_23903,N_23787);
and U24307 (N_24307,N_23331,N_23276);
or U24308 (N_24308,N_23732,N_23603);
nand U24309 (N_24309,N_23948,N_23214);
xnor U24310 (N_24310,N_23193,N_23159);
nor U24311 (N_24311,N_23462,N_23019);
or U24312 (N_24312,N_23612,N_23958);
nor U24313 (N_24313,N_23979,N_23517);
nor U24314 (N_24314,N_23336,N_23269);
and U24315 (N_24315,N_23482,N_23871);
nand U24316 (N_24316,N_23258,N_23651);
nor U24317 (N_24317,N_23259,N_23925);
xnor U24318 (N_24318,N_23391,N_23973);
and U24319 (N_24319,N_23427,N_23045);
xnor U24320 (N_24320,N_23457,N_23386);
nor U24321 (N_24321,N_23138,N_23571);
or U24322 (N_24322,N_23127,N_23957);
nor U24323 (N_24323,N_23494,N_23135);
or U24324 (N_24324,N_23345,N_23363);
or U24325 (N_24325,N_23778,N_23626);
and U24326 (N_24326,N_23455,N_23854);
nor U24327 (N_24327,N_23691,N_23996);
and U24328 (N_24328,N_23347,N_23392);
nand U24329 (N_24329,N_23332,N_23009);
and U24330 (N_24330,N_23428,N_23130);
xor U24331 (N_24331,N_23564,N_23541);
nor U24332 (N_24332,N_23489,N_23426);
xnor U24333 (N_24333,N_23818,N_23198);
xor U24334 (N_24334,N_23968,N_23415);
nand U24335 (N_24335,N_23325,N_23522);
nor U24336 (N_24336,N_23490,N_23865);
and U24337 (N_24337,N_23449,N_23184);
xor U24338 (N_24338,N_23375,N_23297);
or U24339 (N_24339,N_23069,N_23799);
or U24340 (N_24340,N_23789,N_23168);
or U24341 (N_24341,N_23931,N_23227);
and U24342 (N_24342,N_23488,N_23208);
and U24343 (N_24343,N_23704,N_23648);
nor U24344 (N_24344,N_23988,N_23820);
xor U24345 (N_24345,N_23240,N_23364);
xor U24346 (N_24346,N_23093,N_23081);
nor U24347 (N_24347,N_23669,N_23318);
nor U24348 (N_24348,N_23756,N_23539);
xnor U24349 (N_24349,N_23609,N_23296);
xor U24350 (N_24350,N_23366,N_23687);
xor U24351 (N_24351,N_23620,N_23962);
nand U24352 (N_24352,N_23233,N_23726);
or U24353 (N_24353,N_23262,N_23383);
nor U24354 (N_24354,N_23001,N_23832);
or U24355 (N_24355,N_23051,N_23217);
nand U24356 (N_24356,N_23408,N_23152);
and U24357 (N_24357,N_23454,N_23833);
nor U24358 (N_24358,N_23443,N_23413);
and U24359 (N_24359,N_23663,N_23493);
nor U24360 (N_24360,N_23717,N_23566);
or U24361 (N_24361,N_23739,N_23181);
nand U24362 (N_24362,N_23249,N_23000);
or U24363 (N_24363,N_23782,N_23112);
and U24364 (N_24364,N_23421,N_23646);
or U24365 (N_24365,N_23572,N_23196);
nor U24366 (N_24366,N_23272,N_23936);
nor U24367 (N_24367,N_23975,N_23673);
nor U24368 (N_24368,N_23192,N_23255);
and U24369 (N_24369,N_23024,N_23351);
nor U24370 (N_24370,N_23183,N_23859);
nor U24371 (N_24371,N_23808,N_23030);
nand U24372 (N_24372,N_23509,N_23681);
or U24373 (N_24373,N_23674,N_23683);
nand U24374 (N_24374,N_23729,N_23257);
nor U24375 (N_24375,N_23882,N_23074);
xnor U24376 (N_24376,N_23838,N_23707);
xor U24377 (N_24377,N_23479,N_23400);
or U24378 (N_24378,N_23100,N_23686);
nand U24379 (N_24379,N_23915,N_23178);
nand U24380 (N_24380,N_23254,N_23304);
and U24381 (N_24381,N_23466,N_23004);
or U24382 (N_24382,N_23280,N_23534);
nor U24383 (N_24383,N_23798,N_23943);
and U24384 (N_24384,N_23880,N_23284);
or U24385 (N_24385,N_23667,N_23803);
nand U24386 (N_24386,N_23360,N_23486);
xnor U24387 (N_24387,N_23498,N_23692);
or U24388 (N_24388,N_23121,N_23436);
nor U24389 (N_24389,N_23881,N_23315);
and U24390 (N_24390,N_23666,N_23026);
xor U24391 (N_24391,N_23664,N_23775);
xor U24392 (N_24392,N_23172,N_23146);
nand U24393 (N_24393,N_23913,N_23260);
xnor U24394 (N_24394,N_23440,N_23092);
nor U24395 (N_24395,N_23188,N_23752);
or U24396 (N_24396,N_23342,N_23147);
nand U24397 (N_24397,N_23374,N_23895);
xnor U24398 (N_24398,N_23048,N_23224);
or U24399 (N_24399,N_23533,N_23055);
nand U24400 (N_24400,N_23021,N_23675);
nand U24401 (N_24401,N_23916,N_23899);
nor U24402 (N_24402,N_23072,N_23606);
or U24403 (N_24403,N_23748,N_23837);
or U24404 (N_24404,N_23136,N_23821);
xnor U24405 (N_24405,N_23119,N_23892);
nand U24406 (N_24406,N_23507,N_23033);
xnor U24407 (N_24407,N_23984,N_23737);
nand U24408 (N_24408,N_23190,N_23898);
nand U24409 (N_24409,N_23226,N_23197);
and U24410 (N_24410,N_23921,N_23532);
xnor U24411 (N_24411,N_23978,N_23195);
or U24412 (N_24412,N_23236,N_23316);
xnor U24413 (N_24413,N_23199,N_23271);
nand U24414 (N_24414,N_23560,N_23698);
xor U24415 (N_24415,N_23054,N_23246);
nand U24416 (N_24416,N_23581,N_23568);
nor U24417 (N_24417,N_23524,N_23463);
and U24418 (N_24418,N_23474,N_23946);
nor U24419 (N_24419,N_23085,N_23788);
and U24420 (N_24420,N_23091,N_23483);
nand U24421 (N_24421,N_23905,N_23222);
nor U24422 (N_24422,N_23615,N_23814);
or U24423 (N_24423,N_23608,N_23173);
or U24424 (N_24424,N_23910,N_23792);
nor U24425 (N_24425,N_23942,N_23396);
xnor U24426 (N_24426,N_23813,N_23974);
xnor U24427 (N_24427,N_23106,N_23017);
and U24428 (N_24428,N_23735,N_23213);
nor U24429 (N_24429,N_23293,N_23103);
nand U24430 (N_24430,N_23831,N_23857);
nand U24431 (N_24431,N_23743,N_23595);
xnor U24432 (N_24432,N_23768,N_23065);
nand U24433 (N_24433,N_23376,N_23095);
or U24434 (N_24434,N_23448,N_23301);
nand U24435 (N_24435,N_23248,N_23642);
and U24436 (N_24436,N_23420,N_23281);
nand U24437 (N_24437,N_23866,N_23174);
nor U24438 (N_24438,N_23586,N_23652);
and U24439 (N_24439,N_23817,N_23029);
nor U24440 (N_24440,N_23223,N_23231);
or U24441 (N_24441,N_23999,N_23725);
and U24442 (N_24442,N_23295,N_23896);
and U24443 (N_24443,N_23302,N_23718);
xor U24444 (N_24444,N_23108,N_23868);
and U24445 (N_24445,N_23058,N_23830);
or U24446 (N_24446,N_23139,N_23028);
nor U24447 (N_24447,N_23447,N_23078);
or U24448 (N_24448,N_23758,N_23133);
nor U24449 (N_24449,N_23552,N_23800);
nand U24450 (N_24450,N_23841,N_23423);
xnor U24451 (N_24451,N_23621,N_23870);
nand U24452 (N_24452,N_23576,N_23343);
xnor U24453 (N_24453,N_23034,N_23724);
and U24454 (N_24454,N_23230,N_23333);
and U24455 (N_24455,N_23277,N_23624);
nor U24456 (N_24456,N_23242,N_23221);
or U24457 (N_24457,N_23485,N_23158);
nor U24458 (N_24458,N_23550,N_23006);
or U24459 (N_24459,N_23409,N_23967);
or U24460 (N_24460,N_23694,N_23419);
xor U24461 (N_24461,N_23202,N_23933);
or U24462 (N_24462,N_23056,N_23879);
and U24463 (N_24463,N_23794,N_23834);
and U24464 (N_24464,N_23850,N_23616);
xor U24465 (N_24465,N_23031,N_23371);
nor U24466 (N_24466,N_23232,N_23589);
nor U24467 (N_24467,N_23437,N_23110);
xnor U24468 (N_24468,N_23660,N_23920);
or U24469 (N_24469,N_23701,N_23012);
nand U24470 (N_24470,N_23317,N_23639);
nor U24471 (N_24471,N_23888,N_23453);
and U24472 (N_24472,N_23544,N_23311);
nand U24473 (N_24473,N_23215,N_23289);
xor U24474 (N_24474,N_23790,N_23755);
or U24475 (N_24475,N_23140,N_23125);
nand U24476 (N_24476,N_23991,N_23037);
and U24477 (N_24477,N_23329,N_23362);
and U24478 (N_24478,N_23460,N_23890);
or U24479 (N_24479,N_23549,N_23175);
or U24480 (N_24480,N_23060,N_23938);
nor U24481 (N_24481,N_23601,N_23959);
nor U24482 (N_24482,N_23166,N_23404);
nor U24483 (N_24483,N_23104,N_23395);
nor U24484 (N_24484,N_23132,N_23839);
and U24485 (N_24485,N_23068,N_23784);
nand U24486 (N_24486,N_23981,N_23877);
xor U24487 (N_24487,N_23123,N_23689);
and U24488 (N_24488,N_23398,N_23327);
nor U24489 (N_24489,N_23577,N_23238);
and U24490 (N_24490,N_23700,N_23275);
nand U24491 (N_24491,N_23397,N_23309);
or U24492 (N_24492,N_23658,N_23165);
or U24493 (N_24493,N_23753,N_23210);
nand U24494 (N_24494,N_23279,N_23394);
or U24495 (N_24495,N_23709,N_23212);
nor U24496 (N_24496,N_23270,N_23456);
or U24497 (N_24497,N_23811,N_23562);
xor U24498 (N_24498,N_23883,N_23976);
xnor U24499 (N_24499,N_23372,N_23380);
nor U24500 (N_24500,N_23097,N_23194);
nand U24501 (N_24501,N_23518,N_23464);
xnor U24502 (N_24502,N_23841,N_23125);
xor U24503 (N_24503,N_23559,N_23349);
and U24504 (N_24504,N_23962,N_23179);
xor U24505 (N_24505,N_23372,N_23887);
xnor U24506 (N_24506,N_23949,N_23130);
and U24507 (N_24507,N_23881,N_23552);
or U24508 (N_24508,N_23958,N_23914);
xnor U24509 (N_24509,N_23858,N_23510);
nor U24510 (N_24510,N_23371,N_23686);
or U24511 (N_24511,N_23393,N_23879);
and U24512 (N_24512,N_23519,N_23491);
and U24513 (N_24513,N_23214,N_23145);
or U24514 (N_24514,N_23860,N_23919);
and U24515 (N_24515,N_23197,N_23788);
xor U24516 (N_24516,N_23765,N_23081);
nand U24517 (N_24517,N_23584,N_23401);
or U24518 (N_24518,N_23200,N_23564);
or U24519 (N_24519,N_23463,N_23439);
nand U24520 (N_24520,N_23436,N_23134);
nand U24521 (N_24521,N_23706,N_23993);
nand U24522 (N_24522,N_23906,N_23199);
nand U24523 (N_24523,N_23334,N_23636);
nor U24524 (N_24524,N_23801,N_23107);
nand U24525 (N_24525,N_23525,N_23197);
xor U24526 (N_24526,N_23069,N_23235);
xnor U24527 (N_24527,N_23084,N_23949);
nand U24528 (N_24528,N_23164,N_23383);
xnor U24529 (N_24529,N_23479,N_23550);
nand U24530 (N_24530,N_23920,N_23544);
nand U24531 (N_24531,N_23743,N_23444);
or U24532 (N_24532,N_23486,N_23506);
or U24533 (N_24533,N_23087,N_23152);
nand U24534 (N_24534,N_23916,N_23355);
or U24535 (N_24535,N_23465,N_23981);
xnor U24536 (N_24536,N_23822,N_23227);
xor U24537 (N_24537,N_23303,N_23610);
xor U24538 (N_24538,N_23405,N_23350);
nand U24539 (N_24539,N_23721,N_23684);
or U24540 (N_24540,N_23082,N_23210);
nor U24541 (N_24541,N_23386,N_23388);
xnor U24542 (N_24542,N_23287,N_23431);
or U24543 (N_24543,N_23750,N_23011);
or U24544 (N_24544,N_23968,N_23793);
nor U24545 (N_24545,N_23837,N_23054);
or U24546 (N_24546,N_23111,N_23257);
and U24547 (N_24547,N_23560,N_23603);
or U24548 (N_24548,N_23666,N_23068);
or U24549 (N_24549,N_23668,N_23749);
nor U24550 (N_24550,N_23476,N_23248);
xnor U24551 (N_24551,N_23000,N_23680);
nor U24552 (N_24552,N_23264,N_23778);
and U24553 (N_24553,N_23118,N_23230);
and U24554 (N_24554,N_23099,N_23274);
nand U24555 (N_24555,N_23965,N_23096);
nor U24556 (N_24556,N_23322,N_23297);
and U24557 (N_24557,N_23563,N_23676);
nor U24558 (N_24558,N_23160,N_23652);
and U24559 (N_24559,N_23822,N_23751);
or U24560 (N_24560,N_23827,N_23226);
and U24561 (N_24561,N_23294,N_23390);
xnor U24562 (N_24562,N_23894,N_23088);
and U24563 (N_24563,N_23273,N_23260);
nor U24564 (N_24564,N_23066,N_23551);
and U24565 (N_24565,N_23099,N_23158);
or U24566 (N_24566,N_23395,N_23164);
or U24567 (N_24567,N_23680,N_23727);
nand U24568 (N_24568,N_23151,N_23291);
and U24569 (N_24569,N_23788,N_23641);
xor U24570 (N_24570,N_23344,N_23378);
nor U24571 (N_24571,N_23691,N_23352);
xor U24572 (N_24572,N_23920,N_23254);
nand U24573 (N_24573,N_23390,N_23990);
or U24574 (N_24574,N_23948,N_23099);
nand U24575 (N_24575,N_23331,N_23617);
or U24576 (N_24576,N_23358,N_23732);
and U24577 (N_24577,N_23150,N_23431);
nand U24578 (N_24578,N_23357,N_23813);
or U24579 (N_24579,N_23693,N_23505);
nor U24580 (N_24580,N_23661,N_23804);
or U24581 (N_24581,N_23856,N_23494);
nor U24582 (N_24582,N_23874,N_23453);
nor U24583 (N_24583,N_23663,N_23661);
nand U24584 (N_24584,N_23685,N_23919);
and U24585 (N_24585,N_23538,N_23263);
or U24586 (N_24586,N_23844,N_23700);
nor U24587 (N_24587,N_23259,N_23234);
nor U24588 (N_24588,N_23838,N_23748);
nor U24589 (N_24589,N_23108,N_23484);
or U24590 (N_24590,N_23121,N_23853);
nand U24591 (N_24591,N_23519,N_23239);
nand U24592 (N_24592,N_23113,N_23001);
xnor U24593 (N_24593,N_23627,N_23664);
xor U24594 (N_24594,N_23159,N_23938);
nand U24595 (N_24595,N_23154,N_23624);
nor U24596 (N_24596,N_23480,N_23133);
or U24597 (N_24597,N_23456,N_23466);
or U24598 (N_24598,N_23627,N_23447);
and U24599 (N_24599,N_23286,N_23190);
and U24600 (N_24600,N_23692,N_23950);
xor U24601 (N_24601,N_23485,N_23453);
nor U24602 (N_24602,N_23415,N_23261);
or U24603 (N_24603,N_23729,N_23233);
nor U24604 (N_24604,N_23220,N_23071);
nand U24605 (N_24605,N_23339,N_23421);
nor U24606 (N_24606,N_23314,N_23945);
or U24607 (N_24607,N_23509,N_23841);
xnor U24608 (N_24608,N_23697,N_23111);
or U24609 (N_24609,N_23243,N_23285);
nor U24610 (N_24610,N_23596,N_23651);
and U24611 (N_24611,N_23835,N_23282);
nor U24612 (N_24612,N_23023,N_23884);
nor U24613 (N_24613,N_23955,N_23154);
and U24614 (N_24614,N_23343,N_23942);
xor U24615 (N_24615,N_23151,N_23324);
nor U24616 (N_24616,N_23782,N_23170);
nor U24617 (N_24617,N_23221,N_23804);
or U24618 (N_24618,N_23482,N_23372);
xor U24619 (N_24619,N_23784,N_23912);
and U24620 (N_24620,N_23782,N_23943);
or U24621 (N_24621,N_23649,N_23964);
and U24622 (N_24622,N_23679,N_23726);
nand U24623 (N_24623,N_23949,N_23828);
and U24624 (N_24624,N_23805,N_23605);
and U24625 (N_24625,N_23369,N_23392);
or U24626 (N_24626,N_23123,N_23466);
and U24627 (N_24627,N_23218,N_23920);
nor U24628 (N_24628,N_23987,N_23768);
nor U24629 (N_24629,N_23705,N_23050);
and U24630 (N_24630,N_23013,N_23798);
xor U24631 (N_24631,N_23538,N_23697);
or U24632 (N_24632,N_23625,N_23144);
and U24633 (N_24633,N_23363,N_23452);
xor U24634 (N_24634,N_23740,N_23074);
nand U24635 (N_24635,N_23161,N_23786);
nand U24636 (N_24636,N_23375,N_23640);
or U24637 (N_24637,N_23483,N_23351);
and U24638 (N_24638,N_23119,N_23116);
nor U24639 (N_24639,N_23617,N_23293);
nand U24640 (N_24640,N_23720,N_23510);
nor U24641 (N_24641,N_23937,N_23993);
nand U24642 (N_24642,N_23852,N_23380);
nor U24643 (N_24643,N_23879,N_23422);
xnor U24644 (N_24644,N_23472,N_23453);
nand U24645 (N_24645,N_23683,N_23924);
or U24646 (N_24646,N_23595,N_23955);
or U24647 (N_24647,N_23332,N_23745);
nand U24648 (N_24648,N_23615,N_23076);
nand U24649 (N_24649,N_23187,N_23140);
xnor U24650 (N_24650,N_23825,N_23251);
or U24651 (N_24651,N_23870,N_23779);
or U24652 (N_24652,N_23641,N_23045);
nor U24653 (N_24653,N_23816,N_23668);
or U24654 (N_24654,N_23521,N_23399);
or U24655 (N_24655,N_23669,N_23493);
and U24656 (N_24656,N_23380,N_23036);
and U24657 (N_24657,N_23337,N_23888);
and U24658 (N_24658,N_23657,N_23562);
xnor U24659 (N_24659,N_23274,N_23460);
nor U24660 (N_24660,N_23761,N_23285);
xnor U24661 (N_24661,N_23303,N_23089);
and U24662 (N_24662,N_23733,N_23245);
nand U24663 (N_24663,N_23652,N_23770);
nor U24664 (N_24664,N_23493,N_23320);
nand U24665 (N_24665,N_23367,N_23181);
xor U24666 (N_24666,N_23408,N_23470);
xnor U24667 (N_24667,N_23787,N_23428);
nor U24668 (N_24668,N_23976,N_23236);
and U24669 (N_24669,N_23245,N_23116);
xnor U24670 (N_24670,N_23363,N_23811);
and U24671 (N_24671,N_23110,N_23802);
nor U24672 (N_24672,N_23660,N_23324);
nand U24673 (N_24673,N_23497,N_23457);
and U24674 (N_24674,N_23685,N_23369);
nor U24675 (N_24675,N_23581,N_23883);
or U24676 (N_24676,N_23302,N_23488);
or U24677 (N_24677,N_23618,N_23499);
and U24678 (N_24678,N_23450,N_23598);
nor U24679 (N_24679,N_23990,N_23116);
xor U24680 (N_24680,N_23720,N_23060);
and U24681 (N_24681,N_23620,N_23930);
or U24682 (N_24682,N_23657,N_23108);
nor U24683 (N_24683,N_23700,N_23129);
nor U24684 (N_24684,N_23086,N_23921);
nand U24685 (N_24685,N_23851,N_23990);
and U24686 (N_24686,N_23008,N_23532);
xnor U24687 (N_24687,N_23340,N_23530);
and U24688 (N_24688,N_23501,N_23370);
xnor U24689 (N_24689,N_23429,N_23796);
xor U24690 (N_24690,N_23845,N_23988);
nor U24691 (N_24691,N_23644,N_23307);
xor U24692 (N_24692,N_23539,N_23714);
nor U24693 (N_24693,N_23626,N_23892);
and U24694 (N_24694,N_23372,N_23833);
and U24695 (N_24695,N_23292,N_23345);
nor U24696 (N_24696,N_23414,N_23195);
or U24697 (N_24697,N_23415,N_23204);
nand U24698 (N_24698,N_23739,N_23761);
or U24699 (N_24699,N_23454,N_23873);
xnor U24700 (N_24700,N_23612,N_23036);
or U24701 (N_24701,N_23310,N_23958);
nor U24702 (N_24702,N_23479,N_23317);
or U24703 (N_24703,N_23517,N_23938);
or U24704 (N_24704,N_23529,N_23298);
or U24705 (N_24705,N_23697,N_23557);
nand U24706 (N_24706,N_23622,N_23472);
or U24707 (N_24707,N_23563,N_23658);
or U24708 (N_24708,N_23678,N_23080);
nor U24709 (N_24709,N_23219,N_23714);
and U24710 (N_24710,N_23789,N_23045);
nand U24711 (N_24711,N_23677,N_23464);
xnor U24712 (N_24712,N_23646,N_23204);
xor U24713 (N_24713,N_23700,N_23584);
nand U24714 (N_24714,N_23616,N_23184);
or U24715 (N_24715,N_23103,N_23954);
and U24716 (N_24716,N_23720,N_23947);
xnor U24717 (N_24717,N_23745,N_23398);
or U24718 (N_24718,N_23995,N_23017);
and U24719 (N_24719,N_23104,N_23743);
or U24720 (N_24720,N_23943,N_23461);
nor U24721 (N_24721,N_23060,N_23173);
xor U24722 (N_24722,N_23804,N_23045);
nand U24723 (N_24723,N_23670,N_23583);
xor U24724 (N_24724,N_23598,N_23334);
and U24725 (N_24725,N_23730,N_23550);
nand U24726 (N_24726,N_23965,N_23167);
or U24727 (N_24727,N_23701,N_23264);
nor U24728 (N_24728,N_23194,N_23390);
and U24729 (N_24729,N_23505,N_23798);
nor U24730 (N_24730,N_23264,N_23149);
or U24731 (N_24731,N_23167,N_23689);
nor U24732 (N_24732,N_23192,N_23195);
and U24733 (N_24733,N_23353,N_23108);
and U24734 (N_24734,N_23893,N_23171);
nor U24735 (N_24735,N_23367,N_23372);
xor U24736 (N_24736,N_23412,N_23496);
and U24737 (N_24737,N_23411,N_23084);
xnor U24738 (N_24738,N_23731,N_23222);
xor U24739 (N_24739,N_23793,N_23468);
or U24740 (N_24740,N_23760,N_23239);
nand U24741 (N_24741,N_23292,N_23885);
and U24742 (N_24742,N_23370,N_23968);
xnor U24743 (N_24743,N_23030,N_23899);
and U24744 (N_24744,N_23972,N_23940);
nor U24745 (N_24745,N_23808,N_23168);
xnor U24746 (N_24746,N_23678,N_23560);
nand U24747 (N_24747,N_23537,N_23918);
nor U24748 (N_24748,N_23198,N_23567);
and U24749 (N_24749,N_23820,N_23870);
xnor U24750 (N_24750,N_23383,N_23569);
xor U24751 (N_24751,N_23350,N_23931);
and U24752 (N_24752,N_23817,N_23735);
nor U24753 (N_24753,N_23579,N_23875);
nand U24754 (N_24754,N_23207,N_23700);
and U24755 (N_24755,N_23675,N_23595);
xnor U24756 (N_24756,N_23856,N_23960);
nor U24757 (N_24757,N_23953,N_23877);
xor U24758 (N_24758,N_23155,N_23467);
nand U24759 (N_24759,N_23706,N_23201);
nand U24760 (N_24760,N_23043,N_23698);
xnor U24761 (N_24761,N_23295,N_23550);
nor U24762 (N_24762,N_23530,N_23390);
or U24763 (N_24763,N_23098,N_23781);
and U24764 (N_24764,N_23224,N_23223);
nand U24765 (N_24765,N_23225,N_23977);
and U24766 (N_24766,N_23062,N_23778);
nor U24767 (N_24767,N_23426,N_23171);
nor U24768 (N_24768,N_23192,N_23021);
nand U24769 (N_24769,N_23891,N_23090);
or U24770 (N_24770,N_23369,N_23695);
and U24771 (N_24771,N_23033,N_23458);
nand U24772 (N_24772,N_23780,N_23207);
or U24773 (N_24773,N_23554,N_23608);
nand U24774 (N_24774,N_23087,N_23562);
and U24775 (N_24775,N_23292,N_23861);
and U24776 (N_24776,N_23820,N_23035);
or U24777 (N_24777,N_23338,N_23538);
nand U24778 (N_24778,N_23604,N_23988);
or U24779 (N_24779,N_23258,N_23901);
and U24780 (N_24780,N_23998,N_23268);
nor U24781 (N_24781,N_23691,N_23651);
nand U24782 (N_24782,N_23640,N_23462);
xor U24783 (N_24783,N_23736,N_23285);
xor U24784 (N_24784,N_23180,N_23927);
and U24785 (N_24785,N_23216,N_23911);
and U24786 (N_24786,N_23050,N_23381);
or U24787 (N_24787,N_23193,N_23435);
xor U24788 (N_24788,N_23106,N_23204);
or U24789 (N_24789,N_23087,N_23823);
or U24790 (N_24790,N_23755,N_23051);
or U24791 (N_24791,N_23921,N_23620);
xor U24792 (N_24792,N_23518,N_23532);
or U24793 (N_24793,N_23405,N_23602);
xor U24794 (N_24794,N_23944,N_23567);
nor U24795 (N_24795,N_23417,N_23869);
and U24796 (N_24796,N_23861,N_23755);
and U24797 (N_24797,N_23691,N_23400);
xnor U24798 (N_24798,N_23312,N_23272);
or U24799 (N_24799,N_23642,N_23913);
or U24800 (N_24800,N_23875,N_23925);
nor U24801 (N_24801,N_23012,N_23598);
nand U24802 (N_24802,N_23431,N_23690);
nor U24803 (N_24803,N_23494,N_23541);
and U24804 (N_24804,N_23773,N_23381);
nor U24805 (N_24805,N_23207,N_23139);
xnor U24806 (N_24806,N_23522,N_23887);
xnor U24807 (N_24807,N_23986,N_23376);
nor U24808 (N_24808,N_23666,N_23744);
xor U24809 (N_24809,N_23224,N_23469);
nor U24810 (N_24810,N_23568,N_23065);
nor U24811 (N_24811,N_23662,N_23592);
nand U24812 (N_24812,N_23677,N_23029);
or U24813 (N_24813,N_23340,N_23219);
and U24814 (N_24814,N_23270,N_23512);
or U24815 (N_24815,N_23956,N_23603);
xor U24816 (N_24816,N_23465,N_23311);
xor U24817 (N_24817,N_23532,N_23013);
nor U24818 (N_24818,N_23660,N_23014);
or U24819 (N_24819,N_23774,N_23603);
and U24820 (N_24820,N_23492,N_23858);
or U24821 (N_24821,N_23920,N_23418);
xor U24822 (N_24822,N_23844,N_23957);
xor U24823 (N_24823,N_23817,N_23602);
nor U24824 (N_24824,N_23547,N_23595);
nand U24825 (N_24825,N_23361,N_23513);
nor U24826 (N_24826,N_23292,N_23554);
and U24827 (N_24827,N_23077,N_23161);
nand U24828 (N_24828,N_23048,N_23981);
xnor U24829 (N_24829,N_23830,N_23121);
xor U24830 (N_24830,N_23177,N_23696);
and U24831 (N_24831,N_23981,N_23697);
nor U24832 (N_24832,N_23015,N_23433);
nor U24833 (N_24833,N_23569,N_23875);
nor U24834 (N_24834,N_23671,N_23860);
or U24835 (N_24835,N_23758,N_23435);
and U24836 (N_24836,N_23341,N_23326);
nor U24837 (N_24837,N_23914,N_23600);
nand U24838 (N_24838,N_23568,N_23730);
nor U24839 (N_24839,N_23254,N_23122);
nor U24840 (N_24840,N_23488,N_23707);
and U24841 (N_24841,N_23606,N_23642);
nor U24842 (N_24842,N_23312,N_23331);
xor U24843 (N_24843,N_23215,N_23722);
nor U24844 (N_24844,N_23923,N_23681);
or U24845 (N_24845,N_23581,N_23734);
xor U24846 (N_24846,N_23990,N_23960);
nor U24847 (N_24847,N_23662,N_23755);
nand U24848 (N_24848,N_23679,N_23132);
nor U24849 (N_24849,N_23901,N_23969);
xor U24850 (N_24850,N_23716,N_23202);
and U24851 (N_24851,N_23858,N_23790);
and U24852 (N_24852,N_23732,N_23084);
nand U24853 (N_24853,N_23380,N_23515);
nand U24854 (N_24854,N_23531,N_23451);
and U24855 (N_24855,N_23964,N_23209);
nor U24856 (N_24856,N_23061,N_23360);
and U24857 (N_24857,N_23191,N_23595);
nand U24858 (N_24858,N_23673,N_23749);
nand U24859 (N_24859,N_23339,N_23133);
or U24860 (N_24860,N_23354,N_23242);
or U24861 (N_24861,N_23219,N_23528);
and U24862 (N_24862,N_23021,N_23174);
xnor U24863 (N_24863,N_23754,N_23948);
and U24864 (N_24864,N_23801,N_23197);
nor U24865 (N_24865,N_23711,N_23378);
and U24866 (N_24866,N_23065,N_23822);
xor U24867 (N_24867,N_23540,N_23898);
or U24868 (N_24868,N_23395,N_23509);
nor U24869 (N_24869,N_23527,N_23174);
and U24870 (N_24870,N_23334,N_23005);
nor U24871 (N_24871,N_23616,N_23609);
and U24872 (N_24872,N_23129,N_23458);
xor U24873 (N_24873,N_23913,N_23382);
nand U24874 (N_24874,N_23137,N_23520);
and U24875 (N_24875,N_23226,N_23089);
and U24876 (N_24876,N_23525,N_23158);
nor U24877 (N_24877,N_23190,N_23416);
and U24878 (N_24878,N_23090,N_23726);
and U24879 (N_24879,N_23965,N_23944);
nor U24880 (N_24880,N_23205,N_23265);
and U24881 (N_24881,N_23361,N_23936);
or U24882 (N_24882,N_23699,N_23715);
nor U24883 (N_24883,N_23789,N_23648);
nor U24884 (N_24884,N_23116,N_23781);
nor U24885 (N_24885,N_23723,N_23775);
or U24886 (N_24886,N_23878,N_23415);
or U24887 (N_24887,N_23095,N_23101);
and U24888 (N_24888,N_23886,N_23766);
xnor U24889 (N_24889,N_23121,N_23164);
or U24890 (N_24890,N_23885,N_23776);
or U24891 (N_24891,N_23483,N_23551);
xor U24892 (N_24892,N_23563,N_23497);
and U24893 (N_24893,N_23938,N_23790);
nand U24894 (N_24894,N_23747,N_23061);
or U24895 (N_24895,N_23619,N_23801);
or U24896 (N_24896,N_23072,N_23671);
or U24897 (N_24897,N_23763,N_23642);
xnor U24898 (N_24898,N_23767,N_23308);
or U24899 (N_24899,N_23342,N_23072);
xnor U24900 (N_24900,N_23453,N_23612);
nor U24901 (N_24901,N_23051,N_23265);
nor U24902 (N_24902,N_23557,N_23206);
xor U24903 (N_24903,N_23761,N_23092);
or U24904 (N_24904,N_23528,N_23030);
nand U24905 (N_24905,N_23943,N_23600);
and U24906 (N_24906,N_23032,N_23846);
and U24907 (N_24907,N_23911,N_23726);
nand U24908 (N_24908,N_23382,N_23361);
xor U24909 (N_24909,N_23460,N_23008);
nor U24910 (N_24910,N_23174,N_23992);
and U24911 (N_24911,N_23387,N_23183);
and U24912 (N_24912,N_23280,N_23140);
nand U24913 (N_24913,N_23725,N_23973);
xor U24914 (N_24914,N_23510,N_23168);
nor U24915 (N_24915,N_23836,N_23173);
xor U24916 (N_24916,N_23287,N_23861);
or U24917 (N_24917,N_23100,N_23895);
xor U24918 (N_24918,N_23383,N_23520);
and U24919 (N_24919,N_23527,N_23676);
and U24920 (N_24920,N_23446,N_23765);
nand U24921 (N_24921,N_23349,N_23397);
nand U24922 (N_24922,N_23210,N_23002);
nor U24923 (N_24923,N_23319,N_23365);
and U24924 (N_24924,N_23369,N_23159);
xor U24925 (N_24925,N_23891,N_23952);
xor U24926 (N_24926,N_23593,N_23114);
and U24927 (N_24927,N_23170,N_23073);
nand U24928 (N_24928,N_23440,N_23355);
nand U24929 (N_24929,N_23960,N_23169);
or U24930 (N_24930,N_23286,N_23704);
nor U24931 (N_24931,N_23300,N_23622);
nor U24932 (N_24932,N_23497,N_23507);
and U24933 (N_24933,N_23114,N_23334);
and U24934 (N_24934,N_23854,N_23883);
or U24935 (N_24935,N_23329,N_23750);
nand U24936 (N_24936,N_23223,N_23051);
or U24937 (N_24937,N_23566,N_23218);
nor U24938 (N_24938,N_23147,N_23153);
and U24939 (N_24939,N_23498,N_23490);
and U24940 (N_24940,N_23558,N_23341);
nand U24941 (N_24941,N_23671,N_23244);
xor U24942 (N_24942,N_23511,N_23785);
or U24943 (N_24943,N_23503,N_23309);
nor U24944 (N_24944,N_23827,N_23648);
or U24945 (N_24945,N_23166,N_23416);
and U24946 (N_24946,N_23113,N_23106);
nor U24947 (N_24947,N_23147,N_23904);
or U24948 (N_24948,N_23919,N_23023);
nand U24949 (N_24949,N_23137,N_23846);
or U24950 (N_24950,N_23912,N_23457);
xor U24951 (N_24951,N_23768,N_23188);
nor U24952 (N_24952,N_23909,N_23911);
xor U24953 (N_24953,N_23702,N_23306);
and U24954 (N_24954,N_23906,N_23817);
and U24955 (N_24955,N_23261,N_23675);
and U24956 (N_24956,N_23487,N_23071);
nand U24957 (N_24957,N_23049,N_23628);
or U24958 (N_24958,N_23954,N_23685);
or U24959 (N_24959,N_23920,N_23558);
nor U24960 (N_24960,N_23784,N_23531);
or U24961 (N_24961,N_23091,N_23002);
nand U24962 (N_24962,N_23242,N_23325);
or U24963 (N_24963,N_23812,N_23746);
nand U24964 (N_24964,N_23644,N_23855);
xnor U24965 (N_24965,N_23781,N_23073);
or U24966 (N_24966,N_23617,N_23944);
nor U24967 (N_24967,N_23524,N_23648);
or U24968 (N_24968,N_23749,N_23820);
nand U24969 (N_24969,N_23189,N_23660);
xnor U24970 (N_24970,N_23963,N_23869);
or U24971 (N_24971,N_23288,N_23479);
nand U24972 (N_24972,N_23911,N_23013);
nor U24973 (N_24973,N_23298,N_23367);
nor U24974 (N_24974,N_23613,N_23088);
nand U24975 (N_24975,N_23661,N_23685);
and U24976 (N_24976,N_23624,N_23740);
xor U24977 (N_24977,N_23150,N_23689);
nor U24978 (N_24978,N_23637,N_23366);
and U24979 (N_24979,N_23164,N_23286);
and U24980 (N_24980,N_23916,N_23156);
xor U24981 (N_24981,N_23854,N_23715);
or U24982 (N_24982,N_23655,N_23293);
and U24983 (N_24983,N_23640,N_23260);
nand U24984 (N_24984,N_23978,N_23618);
nor U24985 (N_24985,N_23737,N_23073);
nand U24986 (N_24986,N_23320,N_23301);
nor U24987 (N_24987,N_23034,N_23733);
xor U24988 (N_24988,N_23407,N_23349);
and U24989 (N_24989,N_23901,N_23398);
nand U24990 (N_24990,N_23849,N_23121);
xnor U24991 (N_24991,N_23366,N_23535);
or U24992 (N_24992,N_23072,N_23447);
xnor U24993 (N_24993,N_23491,N_23209);
or U24994 (N_24994,N_23726,N_23897);
and U24995 (N_24995,N_23713,N_23012);
nor U24996 (N_24996,N_23822,N_23792);
nor U24997 (N_24997,N_23948,N_23265);
xor U24998 (N_24998,N_23316,N_23023);
nand U24999 (N_24999,N_23890,N_23341);
xnor UO_0 (O_0,N_24466,N_24614);
and UO_1 (O_1,N_24662,N_24866);
or UO_2 (O_2,N_24914,N_24457);
or UO_3 (O_3,N_24709,N_24968);
nor UO_4 (O_4,N_24188,N_24855);
nand UO_5 (O_5,N_24006,N_24375);
xor UO_6 (O_6,N_24035,N_24779);
nor UO_7 (O_7,N_24985,N_24969);
nand UO_8 (O_8,N_24094,N_24763);
or UO_9 (O_9,N_24178,N_24025);
xnor UO_10 (O_10,N_24912,N_24499);
nor UO_11 (O_11,N_24850,N_24449);
xnor UO_12 (O_12,N_24257,N_24999);
nor UO_13 (O_13,N_24562,N_24910);
and UO_14 (O_14,N_24019,N_24388);
and UO_15 (O_15,N_24377,N_24345);
nor UO_16 (O_16,N_24984,N_24471);
and UO_17 (O_17,N_24795,N_24229);
xnor UO_18 (O_18,N_24085,N_24817);
and UO_19 (O_19,N_24517,N_24897);
nand UO_20 (O_20,N_24186,N_24874);
nor UO_21 (O_21,N_24551,N_24120);
or UO_22 (O_22,N_24991,N_24421);
xor UO_23 (O_23,N_24931,N_24550);
xor UO_24 (O_24,N_24729,N_24980);
nor UO_25 (O_25,N_24141,N_24465);
nand UO_26 (O_26,N_24223,N_24370);
or UO_27 (O_27,N_24190,N_24732);
and UO_28 (O_28,N_24868,N_24800);
nor UO_29 (O_29,N_24137,N_24804);
xnor UO_30 (O_30,N_24444,N_24445);
nand UO_31 (O_31,N_24052,N_24327);
nand UO_32 (O_32,N_24539,N_24424);
xnor UO_33 (O_33,N_24121,N_24862);
or UO_34 (O_34,N_24658,N_24209);
or UO_35 (O_35,N_24703,N_24612);
nand UO_36 (O_36,N_24669,N_24100);
or UO_37 (O_37,N_24840,N_24216);
and UO_38 (O_38,N_24607,N_24900);
nor UO_39 (O_39,N_24005,N_24988);
or UO_40 (O_40,N_24233,N_24839);
nor UO_41 (O_41,N_24435,N_24953);
or UO_42 (O_42,N_24611,N_24632);
nand UO_43 (O_43,N_24749,N_24210);
or UO_44 (O_44,N_24407,N_24125);
nor UO_45 (O_45,N_24686,N_24700);
or UO_46 (O_46,N_24187,N_24847);
xnor UO_47 (O_47,N_24313,N_24751);
xnor UO_48 (O_48,N_24123,N_24308);
nand UO_49 (O_49,N_24107,N_24018);
nand UO_50 (O_50,N_24485,N_24571);
or UO_51 (O_51,N_24264,N_24320);
nand UO_52 (O_52,N_24856,N_24629);
or UO_53 (O_53,N_24057,N_24108);
and UO_54 (O_54,N_24939,N_24387);
or UO_55 (O_55,N_24343,N_24650);
xnor UO_56 (O_56,N_24268,N_24563);
xor UO_57 (O_57,N_24532,N_24604);
nand UO_58 (O_58,N_24110,N_24322);
and UO_59 (O_59,N_24506,N_24519);
or UO_60 (O_60,N_24000,N_24641);
xnor UO_61 (O_61,N_24762,N_24739);
nor UO_62 (O_62,N_24545,N_24974);
nand UO_63 (O_63,N_24194,N_24525);
nand UO_64 (O_64,N_24310,N_24920);
nand UO_65 (O_65,N_24728,N_24538);
nor UO_66 (O_66,N_24116,N_24936);
or UO_67 (O_67,N_24603,N_24023);
xor UO_68 (O_68,N_24064,N_24542);
nor UO_69 (O_69,N_24970,N_24761);
and UO_70 (O_70,N_24301,N_24513);
xnor UO_71 (O_71,N_24128,N_24886);
or UO_72 (O_72,N_24371,N_24047);
nand UO_73 (O_73,N_24083,N_24438);
xor UO_74 (O_74,N_24828,N_24176);
or UO_75 (O_75,N_24724,N_24189);
or UO_76 (O_76,N_24976,N_24099);
and UO_77 (O_77,N_24164,N_24262);
nor UO_78 (O_78,N_24369,N_24258);
nand UO_79 (O_79,N_24479,N_24699);
nand UO_80 (O_80,N_24736,N_24593);
nor UO_81 (O_81,N_24385,N_24959);
and UO_82 (O_82,N_24281,N_24381);
and UO_83 (O_83,N_24256,N_24587);
nor UO_84 (O_84,N_24860,N_24994);
or UO_85 (O_85,N_24655,N_24030);
nor UO_86 (O_86,N_24211,N_24267);
or UO_87 (O_87,N_24716,N_24225);
xor UO_88 (O_88,N_24311,N_24677);
and UO_89 (O_89,N_24086,N_24789);
nand UO_90 (O_90,N_24417,N_24754);
xnor UO_91 (O_91,N_24637,N_24857);
or UO_92 (O_92,N_24785,N_24863);
xor UO_93 (O_93,N_24460,N_24576);
and UO_94 (O_94,N_24536,N_24140);
xor UO_95 (O_95,N_24772,N_24364);
or UO_96 (O_96,N_24544,N_24305);
and UO_97 (O_97,N_24118,N_24302);
nor UO_98 (O_98,N_24306,N_24119);
and UO_99 (O_99,N_24454,N_24774);
nand UO_100 (O_100,N_24228,N_24938);
nand UO_101 (O_101,N_24656,N_24742);
or UO_102 (O_102,N_24244,N_24704);
nor UO_103 (O_103,N_24312,N_24437);
and UO_104 (O_104,N_24596,N_24134);
nand UO_105 (O_105,N_24464,N_24303);
nor UO_106 (O_106,N_24197,N_24824);
xnor UO_107 (O_107,N_24977,N_24284);
xor UO_108 (O_108,N_24516,N_24933);
xnor UO_109 (O_109,N_24923,N_24271);
or UO_110 (O_110,N_24055,N_24446);
nor UO_111 (O_111,N_24250,N_24565);
xnor UO_112 (O_112,N_24149,N_24033);
nor UO_113 (O_113,N_24770,N_24652);
or UO_114 (O_114,N_24916,N_24937);
nor UO_115 (O_115,N_24196,N_24971);
and UO_116 (O_116,N_24721,N_24461);
and UO_117 (O_117,N_24515,N_24872);
and UO_118 (O_118,N_24534,N_24053);
or UO_119 (O_119,N_24017,N_24351);
and UO_120 (O_120,N_24812,N_24034);
nand UO_121 (O_121,N_24255,N_24661);
or UO_122 (O_122,N_24090,N_24031);
nand UO_123 (O_123,N_24245,N_24152);
and UO_124 (O_124,N_24335,N_24326);
and UO_125 (O_125,N_24952,N_24111);
nor UO_126 (O_126,N_24476,N_24217);
nor UO_127 (O_127,N_24822,N_24929);
and UO_128 (O_128,N_24963,N_24958);
or UO_129 (O_129,N_24675,N_24441);
nor UO_130 (O_130,N_24877,N_24676);
and UO_131 (O_131,N_24115,N_24610);
xnor UO_132 (O_132,N_24051,N_24882);
nor UO_133 (O_133,N_24003,N_24391);
and UO_134 (O_134,N_24702,N_24630);
nor UO_135 (O_135,N_24296,N_24657);
xnor UO_136 (O_136,N_24674,N_24269);
or UO_137 (O_137,N_24741,N_24807);
xnor UO_138 (O_138,N_24531,N_24265);
and UO_139 (O_139,N_24957,N_24636);
or UO_140 (O_140,N_24172,N_24904);
and UO_141 (O_141,N_24291,N_24040);
xnor UO_142 (O_142,N_24433,N_24073);
nand UO_143 (O_143,N_24726,N_24713);
xor UO_144 (O_144,N_24214,N_24734);
nor UO_145 (O_145,N_24484,N_24103);
or UO_146 (O_146,N_24917,N_24841);
xor UO_147 (O_147,N_24443,N_24638);
and UO_148 (O_148,N_24913,N_24801);
and UO_149 (O_149,N_24678,N_24300);
and UO_150 (O_150,N_24207,N_24792);
and UO_151 (O_151,N_24832,N_24406);
or UO_152 (O_152,N_24242,N_24474);
nor UO_153 (O_153,N_24777,N_24237);
nand UO_154 (O_154,N_24069,N_24592);
xnor UO_155 (O_155,N_24878,N_24340);
nand UO_156 (O_156,N_24520,N_24213);
nor UO_157 (O_157,N_24028,N_24379);
and UO_158 (O_158,N_24292,N_24234);
xor UO_159 (O_159,N_24136,N_24114);
or UO_160 (O_160,N_24583,N_24773);
nand UO_161 (O_161,N_24378,N_24428);
xnor UO_162 (O_162,N_24497,N_24620);
nand UO_163 (O_163,N_24588,N_24329);
or UO_164 (O_164,N_24835,N_24180);
or UO_165 (O_165,N_24087,N_24082);
or UO_166 (O_166,N_24135,N_24272);
and UO_167 (O_167,N_24715,N_24434);
or UO_168 (O_168,N_24270,N_24227);
and UO_169 (O_169,N_24317,N_24293);
or UO_170 (O_170,N_24618,N_24448);
xor UO_171 (O_171,N_24405,N_24394);
nand UO_172 (O_172,N_24191,N_24429);
and UO_173 (O_173,N_24978,N_24092);
xnor UO_174 (O_174,N_24404,N_24949);
nand UO_175 (O_175,N_24459,N_24376);
and UO_176 (O_176,N_24767,N_24831);
or UO_177 (O_177,N_24590,N_24950);
and UO_178 (O_178,N_24667,N_24275);
nor UO_179 (O_179,N_24122,N_24791);
xnor UO_180 (O_180,N_24842,N_24456);
or UO_181 (O_181,N_24145,N_24560);
xnor UO_182 (O_182,N_24261,N_24737);
and UO_183 (O_183,N_24809,N_24338);
nor UO_184 (O_184,N_24646,N_24557);
and UO_185 (O_185,N_24947,N_24089);
or UO_186 (O_186,N_24887,N_24481);
and UO_187 (O_187,N_24347,N_24797);
nand UO_188 (O_188,N_24491,N_24352);
nor UO_189 (O_189,N_24436,N_24598);
xnor UO_190 (O_190,N_24230,N_24625);
nor UO_191 (O_191,N_24450,N_24836);
nand UO_192 (O_192,N_24594,N_24130);
or UO_193 (O_193,N_24526,N_24399);
xor UO_194 (O_194,N_24711,N_24823);
nand UO_195 (O_195,N_24483,N_24908);
nor UO_196 (O_196,N_24541,N_24597);
xor UO_197 (O_197,N_24537,N_24825);
xnor UO_198 (O_198,N_24496,N_24624);
xor UO_199 (O_199,N_24595,N_24467);
xor UO_200 (O_200,N_24009,N_24163);
nand UO_201 (O_201,N_24339,N_24723);
nor UO_202 (O_202,N_24026,N_24374);
and UO_203 (O_203,N_24362,N_24021);
xor UO_204 (O_204,N_24813,N_24166);
nand UO_205 (O_205,N_24993,N_24631);
xnor UO_206 (O_206,N_24333,N_24966);
nand UO_207 (O_207,N_24902,N_24852);
nor UO_208 (O_208,N_24577,N_24747);
nand UO_209 (O_209,N_24038,N_24698);
xnor UO_210 (O_210,N_24654,N_24368);
and UO_211 (O_211,N_24162,N_24580);
nand UO_212 (O_212,N_24240,N_24494);
nor UO_213 (O_213,N_24668,N_24046);
and UO_214 (O_214,N_24919,N_24752);
or UO_215 (O_215,N_24024,N_24748);
or UO_216 (O_216,N_24547,N_24851);
or UO_217 (O_217,N_24648,N_24815);
nand UO_218 (O_218,N_24037,N_24181);
and UO_219 (O_219,N_24442,N_24175);
xor UO_220 (O_220,N_24644,N_24556);
xor UO_221 (O_221,N_24403,N_24361);
xor UO_222 (O_222,N_24572,N_24451);
nor UO_223 (O_223,N_24357,N_24972);
nor UO_224 (O_224,N_24044,N_24853);
nand UO_225 (O_225,N_24011,N_24170);
nand UO_226 (O_226,N_24820,N_24384);
and UO_227 (O_227,N_24543,N_24503);
and UO_228 (O_228,N_24858,N_24778);
or UO_229 (O_229,N_24062,N_24869);
xor UO_230 (O_230,N_24876,N_24643);
and UO_231 (O_231,N_24712,N_24029);
nand UO_232 (O_232,N_24983,N_24918);
nor UO_233 (O_233,N_24290,N_24621);
xor UO_234 (O_234,N_24282,N_24490);
nor UO_235 (O_235,N_24295,N_24478);
or UO_236 (O_236,N_24027,N_24498);
nand UO_237 (O_237,N_24833,N_24967);
xor UO_238 (O_238,N_24492,N_24117);
or UO_239 (O_239,N_24389,N_24336);
nor UO_240 (O_240,N_24780,N_24154);
or UO_241 (O_241,N_24873,N_24248);
or UO_242 (O_242,N_24907,N_24951);
and UO_243 (O_243,N_24273,N_24973);
or UO_244 (O_244,N_24619,N_24666);
xor UO_245 (O_245,N_24294,N_24309);
xnor UO_246 (O_246,N_24808,N_24719);
xnor UO_247 (O_247,N_24330,N_24743);
xor UO_248 (O_248,N_24722,N_24109);
or UO_249 (O_249,N_24796,N_24591);
nand UO_250 (O_250,N_24226,N_24731);
and UO_251 (O_251,N_24144,N_24806);
nand UO_252 (O_252,N_24059,N_24221);
or UO_253 (O_253,N_24799,N_24096);
xnor UO_254 (O_254,N_24906,N_24725);
nor UO_255 (O_255,N_24150,N_24093);
and UO_256 (O_256,N_24696,N_24393);
xnor UO_257 (O_257,N_24156,N_24418);
and UO_258 (O_258,N_24627,N_24605);
or UO_259 (O_259,N_24208,N_24049);
nand UO_260 (O_260,N_24063,N_24198);
nand UO_261 (O_261,N_24319,N_24318);
nor UO_262 (O_262,N_24527,N_24710);
or UO_263 (O_263,N_24680,N_24472);
and UO_264 (O_264,N_24167,N_24133);
and UO_265 (O_265,N_24241,N_24871);
nor UO_266 (O_266,N_24996,N_24690);
and UO_267 (O_267,N_24578,N_24932);
and UO_268 (O_268,N_24380,N_24341);
nand UO_269 (O_269,N_24243,N_24246);
and UO_270 (O_270,N_24112,N_24689);
xor UO_271 (O_271,N_24819,N_24095);
nand UO_272 (O_272,N_24896,N_24990);
nor UO_273 (O_273,N_24054,N_24505);
nand UO_274 (O_274,N_24222,N_24299);
nor UO_275 (O_275,N_24081,N_24402);
xor UO_276 (O_276,N_24665,N_24899);
or UO_277 (O_277,N_24567,N_24487);
nor UO_278 (O_278,N_24158,N_24755);
and UO_279 (O_279,N_24925,N_24323);
xnor UO_280 (O_280,N_24200,N_24409);
and UO_281 (O_281,N_24279,N_24660);
nand UO_282 (O_282,N_24165,N_24821);
or UO_283 (O_283,N_24615,N_24373);
and UO_284 (O_284,N_24132,N_24427);
or UO_285 (O_285,N_24717,N_24139);
xnor UO_286 (O_286,N_24043,N_24500);
nor UO_287 (O_287,N_24431,N_24013);
and UO_288 (O_288,N_24192,N_24798);
nand UO_289 (O_289,N_24834,N_24760);
xnor UO_290 (O_290,N_24365,N_24639);
xnor UO_291 (O_291,N_24982,N_24775);
or UO_292 (O_292,N_24559,N_24253);
and UO_293 (O_293,N_24344,N_24909);
nor UO_294 (O_294,N_24286,N_24837);
nand UO_295 (O_295,N_24452,N_24287);
or UO_296 (O_296,N_24259,N_24201);
nand UO_297 (O_297,N_24477,N_24626);
and UO_298 (O_298,N_24420,N_24695);
nand UO_299 (O_299,N_24101,N_24782);
xnor UO_300 (O_300,N_24354,N_24470);
or UO_301 (O_301,N_24415,N_24768);
nand UO_302 (O_302,N_24535,N_24432);
or UO_303 (O_303,N_24533,N_24398);
or UO_304 (O_304,N_24382,N_24784);
or UO_305 (O_305,N_24826,N_24185);
xor UO_306 (O_306,N_24681,N_24169);
nand UO_307 (O_307,N_24179,N_24072);
nand UO_308 (O_308,N_24769,N_24964);
and UO_309 (O_309,N_24956,N_24151);
or UO_310 (O_310,N_24783,N_24579);
and UO_311 (O_311,N_24050,N_24501);
nand UO_312 (O_312,N_24905,N_24671);
and UO_313 (O_313,N_24707,N_24705);
nand UO_314 (O_314,N_24014,N_24986);
or UO_315 (O_315,N_24419,N_24584);
or UO_316 (O_316,N_24663,N_24235);
nor UO_317 (O_317,N_24602,N_24414);
and UO_318 (O_318,N_24898,N_24220);
nand UO_319 (O_319,N_24864,N_24056);
xnor UO_320 (O_320,N_24146,N_24942);
nor UO_321 (O_321,N_24193,N_24488);
or UO_322 (O_322,N_24001,N_24880);
nand UO_323 (O_323,N_24041,N_24744);
xor UO_324 (O_324,N_24586,N_24098);
nor UO_325 (O_325,N_24530,N_24890);
xnor UO_326 (O_326,N_24411,N_24915);
nand UO_327 (O_327,N_24350,N_24575);
nor UO_328 (O_328,N_24975,N_24482);
nor UO_329 (O_329,N_24195,N_24844);
and UO_330 (O_330,N_24480,N_24153);
nand UO_331 (O_331,N_24079,N_24355);
nor UO_332 (O_332,N_24574,N_24827);
or UO_333 (O_333,N_24386,N_24911);
and UO_334 (O_334,N_24439,N_24753);
and UO_335 (O_335,N_24314,N_24032);
nand UO_336 (O_336,N_24582,N_24892);
nand UO_337 (O_337,N_24570,N_24616);
nand UO_338 (O_338,N_24838,N_24203);
nor UO_339 (O_339,N_24458,N_24928);
xor UO_340 (O_340,N_24440,N_24647);
and UO_341 (O_341,N_24015,N_24004);
and UO_342 (O_342,N_24701,N_24202);
nor UO_343 (O_343,N_24113,N_24771);
nand UO_344 (O_344,N_24468,N_24413);
nand UO_345 (O_345,N_24549,N_24348);
or UO_346 (O_346,N_24462,N_24342);
or UO_347 (O_347,N_24182,N_24664);
or UO_348 (O_348,N_24634,N_24159);
nor UO_349 (O_349,N_24889,N_24080);
and UO_350 (O_350,N_24346,N_24510);
nand UO_351 (O_351,N_24585,N_24410);
and UO_352 (O_352,N_24622,N_24683);
nand UO_353 (O_353,N_24830,N_24861);
or UO_354 (O_354,N_24097,N_24447);
or UO_355 (O_355,N_24084,N_24071);
nand UO_356 (O_356,N_24816,N_24074);
and UO_357 (O_357,N_24065,N_24328);
nor UO_358 (O_358,N_24020,N_24766);
or UO_359 (O_359,N_24759,N_24514);
xnor UO_360 (O_360,N_24315,N_24802);
and UO_361 (O_361,N_24962,N_24921);
or UO_362 (O_362,N_24254,N_24218);
xor UO_363 (O_363,N_24989,N_24757);
or UO_364 (O_364,N_24843,N_24756);
and UO_365 (O_365,N_24885,N_24367);
and UO_366 (O_366,N_24568,N_24697);
and UO_367 (O_367,N_24174,N_24408);
or UO_368 (O_368,N_24787,N_24883);
and UO_369 (O_369,N_24845,N_24102);
nor UO_370 (O_370,N_24922,N_24016);
and UO_371 (O_371,N_24682,N_24160);
nand UO_372 (O_372,N_24940,N_24651);
nor UO_373 (O_373,N_24891,N_24276);
nand UO_374 (O_374,N_24998,N_24173);
nand UO_375 (O_375,N_24392,N_24495);
and UO_376 (O_376,N_24231,N_24171);
xor UO_377 (O_377,N_24215,N_24727);
nor UO_378 (O_378,N_24829,N_24334);
nand UO_379 (O_379,N_24316,N_24692);
nand UO_380 (O_380,N_24012,N_24008);
nand UO_381 (O_381,N_24718,N_24337);
or UO_382 (O_382,N_24613,N_24529);
and UO_383 (O_383,N_24358,N_24961);
and UO_384 (O_384,N_24486,N_24521);
or UO_385 (O_385,N_24635,N_24848);
nor UO_386 (O_386,N_24060,N_24219);
and UO_387 (O_387,N_24426,N_24688);
or UO_388 (O_388,N_24548,N_24781);
nor UO_389 (O_389,N_24623,N_24204);
and UO_390 (O_390,N_24157,N_24475);
and UO_391 (O_391,N_24205,N_24042);
or UO_392 (O_392,N_24168,N_24554);
xnor UO_393 (O_393,N_24992,N_24493);
and UO_394 (O_394,N_24672,N_24522);
or UO_395 (O_395,N_24423,N_24706);
nor UO_396 (O_396,N_24566,N_24184);
nand UO_397 (O_397,N_24670,N_24036);
nand UO_398 (O_398,N_24687,N_24552);
xnor UO_399 (O_399,N_24555,N_24924);
xnor UO_400 (O_400,N_24070,N_24078);
and UO_401 (O_401,N_24104,N_24776);
nor UO_402 (O_402,N_24504,N_24236);
or UO_403 (O_403,N_24608,N_24177);
nor UO_404 (O_404,N_24894,N_24277);
or UO_405 (O_405,N_24359,N_24564);
nor UO_406 (O_406,N_24524,N_24875);
nand UO_407 (O_407,N_24927,N_24366);
or UO_408 (O_408,N_24943,N_24091);
nor UO_409 (O_409,N_24068,N_24846);
nand UO_410 (O_410,N_24573,N_24758);
xor UO_411 (O_411,N_24263,N_24659);
xnor UO_412 (O_412,N_24685,N_24965);
xor UO_413 (O_413,N_24331,N_24280);
or UO_414 (O_414,N_24765,N_24561);
and UO_415 (O_415,N_24260,N_24395);
and UO_416 (O_416,N_24730,N_24239);
and UO_417 (O_417,N_24455,N_24383);
or UO_418 (O_418,N_24304,N_24649);
or UO_419 (O_419,N_24285,N_24349);
and UO_420 (O_420,N_24708,N_24142);
or UO_421 (O_421,N_24131,N_24935);
xor UO_422 (O_422,N_24396,N_24401);
nand UO_423 (O_423,N_24143,N_24199);
nand UO_424 (O_424,N_24283,N_24356);
nand UO_425 (O_425,N_24987,N_24212);
and UO_426 (O_426,N_24589,N_24129);
nand UO_427 (O_427,N_24224,N_24289);
nand UO_428 (O_428,N_24810,N_24425);
xnor UO_429 (O_429,N_24979,N_24581);
xnor UO_430 (O_430,N_24870,N_24934);
nand UO_431 (O_431,N_24617,N_24679);
nand UO_432 (O_432,N_24764,N_24297);
or UO_433 (O_433,N_24048,N_24512);
xnor UO_434 (O_434,N_24944,N_24463);
nor UO_435 (O_435,N_24879,N_24509);
or UO_436 (O_436,N_24805,N_24148);
nand UO_437 (O_437,N_24105,N_24266);
or UO_438 (O_438,N_24416,N_24794);
or UO_439 (O_439,N_24278,N_24948);
xor UO_440 (O_440,N_24945,N_24489);
nor UO_441 (O_441,N_24360,N_24955);
nor UO_442 (O_442,N_24232,N_24075);
and UO_443 (O_443,N_24738,N_24553);
xnor UO_444 (O_444,N_24884,N_24127);
nor UO_445 (O_445,N_24077,N_24997);
nand UO_446 (O_446,N_24453,N_24390);
xnor UO_447 (O_447,N_24247,N_24600);
nor UO_448 (O_448,N_24251,N_24628);
nor UO_449 (O_449,N_24067,N_24002);
xor UO_450 (O_450,N_24941,N_24606);
xnor UO_451 (O_451,N_24930,N_24558);
nor UO_452 (O_452,N_24865,N_24811);
nor UO_453 (O_453,N_24714,N_24502);
nor UO_454 (O_454,N_24693,N_24981);
nor UO_455 (O_455,N_24206,N_24058);
xor UO_456 (O_456,N_24735,N_24161);
nand UO_457 (O_457,N_24353,N_24745);
or UO_458 (O_458,N_24088,N_24147);
nor UO_459 (O_459,N_24903,N_24788);
and UO_460 (O_460,N_24733,N_24691);
xor UO_461 (O_461,N_24400,N_24960);
nor UO_462 (O_462,N_24633,N_24803);
nand UO_463 (O_463,N_24298,N_24645);
nand UO_464 (O_464,N_24332,N_24546);
nand UO_465 (O_465,N_24412,N_24893);
and UO_466 (O_466,N_24793,N_24750);
nor UO_467 (O_467,N_24039,N_24010);
nand UO_468 (O_468,N_24995,N_24249);
or UO_469 (O_469,N_24849,N_24307);
xnor UO_470 (O_470,N_24881,N_24473);
or UO_471 (O_471,N_24601,N_24507);
nand UO_472 (O_472,N_24126,N_24518);
xor UO_473 (O_473,N_24397,N_24640);
nor UO_474 (O_474,N_24183,N_24609);
or UO_475 (O_475,N_24325,N_24076);
nor UO_476 (O_476,N_24814,N_24854);
xnor UO_477 (O_477,N_24430,N_24106);
nor UO_478 (O_478,N_24022,N_24867);
nor UO_479 (O_479,N_24511,N_24859);
and UO_480 (O_480,N_24523,N_24469);
nand UO_481 (O_481,N_24422,N_24274);
nor UO_482 (O_482,N_24288,N_24954);
and UO_483 (O_483,N_24508,N_24926);
xor UO_484 (O_484,N_24720,N_24238);
and UO_485 (O_485,N_24061,N_24569);
or UO_486 (O_486,N_24642,N_24066);
nor UO_487 (O_487,N_24155,N_24790);
and UO_488 (O_488,N_24372,N_24694);
xnor UO_489 (O_489,N_24252,N_24746);
nand UO_490 (O_490,N_24740,N_24007);
and UO_491 (O_491,N_24673,N_24818);
or UO_492 (O_492,N_24528,N_24124);
xnor UO_493 (O_493,N_24946,N_24540);
nor UO_494 (O_494,N_24653,N_24363);
nor UO_495 (O_495,N_24321,N_24901);
and UO_496 (O_496,N_24888,N_24895);
xor UO_497 (O_497,N_24324,N_24138);
or UO_498 (O_498,N_24599,N_24045);
and UO_499 (O_499,N_24684,N_24786);
and UO_500 (O_500,N_24419,N_24922);
and UO_501 (O_501,N_24443,N_24282);
nand UO_502 (O_502,N_24966,N_24709);
nor UO_503 (O_503,N_24830,N_24493);
and UO_504 (O_504,N_24929,N_24631);
and UO_505 (O_505,N_24865,N_24201);
xnor UO_506 (O_506,N_24073,N_24950);
nor UO_507 (O_507,N_24662,N_24006);
xor UO_508 (O_508,N_24320,N_24495);
or UO_509 (O_509,N_24978,N_24279);
nor UO_510 (O_510,N_24789,N_24574);
xnor UO_511 (O_511,N_24218,N_24847);
and UO_512 (O_512,N_24215,N_24427);
and UO_513 (O_513,N_24275,N_24987);
and UO_514 (O_514,N_24833,N_24723);
xnor UO_515 (O_515,N_24267,N_24345);
nand UO_516 (O_516,N_24417,N_24527);
or UO_517 (O_517,N_24063,N_24446);
or UO_518 (O_518,N_24246,N_24722);
and UO_519 (O_519,N_24664,N_24217);
nand UO_520 (O_520,N_24275,N_24984);
and UO_521 (O_521,N_24598,N_24474);
or UO_522 (O_522,N_24547,N_24368);
nor UO_523 (O_523,N_24825,N_24334);
nand UO_524 (O_524,N_24350,N_24854);
nand UO_525 (O_525,N_24367,N_24156);
and UO_526 (O_526,N_24610,N_24810);
or UO_527 (O_527,N_24502,N_24020);
and UO_528 (O_528,N_24802,N_24930);
or UO_529 (O_529,N_24761,N_24363);
nand UO_530 (O_530,N_24733,N_24343);
xnor UO_531 (O_531,N_24453,N_24130);
or UO_532 (O_532,N_24680,N_24033);
xnor UO_533 (O_533,N_24906,N_24998);
nand UO_534 (O_534,N_24905,N_24360);
nand UO_535 (O_535,N_24435,N_24918);
and UO_536 (O_536,N_24308,N_24054);
and UO_537 (O_537,N_24674,N_24089);
and UO_538 (O_538,N_24397,N_24872);
nor UO_539 (O_539,N_24440,N_24524);
or UO_540 (O_540,N_24151,N_24449);
nor UO_541 (O_541,N_24165,N_24900);
and UO_542 (O_542,N_24974,N_24446);
nand UO_543 (O_543,N_24027,N_24362);
or UO_544 (O_544,N_24572,N_24767);
or UO_545 (O_545,N_24239,N_24218);
and UO_546 (O_546,N_24833,N_24298);
and UO_547 (O_547,N_24946,N_24306);
nand UO_548 (O_548,N_24146,N_24314);
nand UO_549 (O_549,N_24332,N_24770);
xnor UO_550 (O_550,N_24631,N_24500);
or UO_551 (O_551,N_24402,N_24288);
xor UO_552 (O_552,N_24946,N_24896);
or UO_553 (O_553,N_24733,N_24014);
nor UO_554 (O_554,N_24293,N_24471);
and UO_555 (O_555,N_24384,N_24755);
and UO_556 (O_556,N_24633,N_24167);
xor UO_557 (O_557,N_24446,N_24278);
nor UO_558 (O_558,N_24474,N_24789);
xnor UO_559 (O_559,N_24850,N_24082);
nand UO_560 (O_560,N_24044,N_24961);
nand UO_561 (O_561,N_24381,N_24410);
and UO_562 (O_562,N_24528,N_24853);
nand UO_563 (O_563,N_24756,N_24974);
xnor UO_564 (O_564,N_24210,N_24052);
or UO_565 (O_565,N_24392,N_24325);
xnor UO_566 (O_566,N_24077,N_24665);
or UO_567 (O_567,N_24576,N_24950);
nor UO_568 (O_568,N_24916,N_24912);
xnor UO_569 (O_569,N_24720,N_24607);
nor UO_570 (O_570,N_24114,N_24308);
nand UO_571 (O_571,N_24664,N_24219);
nand UO_572 (O_572,N_24325,N_24008);
nand UO_573 (O_573,N_24811,N_24109);
nand UO_574 (O_574,N_24545,N_24358);
nor UO_575 (O_575,N_24531,N_24954);
or UO_576 (O_576,N_24246,N_24669);
or UO_577 (O_577,N_24796,N_24376);
nor UO_578 (O_578,N_24296,N_24060);
and UO_579 (O_579,N_24967,N_24845);
or UO_580 (O_580,N_24015,N_24166);
xor UO_581 (O_581,N_24843,N_24288);
nand UO_582 (O_582,N_24509,N_24597);
or UO_583 (O_583,N_24093,N_24599);
nor UO_584 (O_584,N_24972,N_24463);
nand UO_585 (O_585,N_24358,N_24863);
nand UO_586 (O_586,N_24614,N_24476);
nand UO_587 (O_587,N_24730,N_24202);
and UO_588 (O_588,N_24453,N_24127);
and UO_589 (O_589,N_24952,N_24147);
or UO_590 (O_590,N_24648,N_24632);
xor UO_591 (O_591,N_24590,N_24969);
and UO_592 (O_592,N_24721,N_24345);
and UO_593 (O_593,N_24369,N_24609);
nand UO_594 (O_594,N_24033,N_24931);
xnor UO_595 (O_595,N_24600,N_24768);
and UO_596 (O_596,N_24157,N_24733);
nand UO_597 (O_597,N_24921,N_24965);
nor UO_598 (O_598,N_24047,N_24363);
and UO_599 (O_599,N_24706,N_24245);
or UO_600 (O_600,N_24500,N_24908);
xor UO_601 (O_601,N_24408,N_24478);
or UO_602 (O_602,N_24028,N_24340);
nand UO_603 (O_603,N_24059,N_24145);
or UO_604 (O_604,N_24611,N_24693);
nand UO_605 (O_605,N_24525,N_24248);
or UO_606 (O_606,N_24664,N_24737);
nor UO_607 (O_607,N_24397,N_24570);
and UO_608 (O_608,N_24940,N_24138);
xnor UO_609 (O_609,N_24888,N_24452);
nand UO_610 (O_610,N_24994,N_24779);
nand UO_611 (O_611,N_24395,N_24068);
nor UO_612 (O_612,N_24141,N_24366);
or UO_613 (O_613,N_24973,N_24823);
or UO_614 (O_614,N_24613,N_24676);
nand UO_615 (O_615,N_24989,N_24635);
xor UO_616 (O_616,N_24293,N_24356);
or UO_617 (O_617,N_24860,N_24509);
nor UO_618 (O_618,N_24371,N_24324);
and UO_619 (O_619,N_24338,N_24517);
nor UO_620 (O_620,N_24413,N_24540);
and UO_621 (O_621,N_24893,N_24876);
nand UO_622 (O_622,N_24736,N_24204);
nor UO_623 (O_623,N_24051,N_24501);
and UO_624 (O_624,N_24611,N_24472);
xnor UO_625 (O_625,N_24993,N_24999);
or UO_626 (O_626,N_24867,N_24530);
and UO_627 (O_627,N_24693,N_24431);
xor UO_628 (O_628,N_24191,N_24744);
nand UO_629 (O_629,N_24864,N_24896);
nor UO_630 (O_630,N_24480,N_24303);
xor UO_631 (O_631,N_24434,N_24504);
xnor UO_632 (O_632,N_24682,N_24158);
nor UO_633 (O_633,N_24636,N_24133);
and UO_634 (O_634,N_24875,N_24225);
and UO_635 (O_635,N_24016,N_24490);
nand UO_636 (O_636,N_24842,N_24535);
nor UO_637 (O_637,N_24643,N_24833);
nand UO_638 (O_638,N_24555,N_24326);
nand UO_639 (O_639,N_24784,N_24721);
or UO_640 (O_640,N_24572,N_24712);
nand UO_641 (O_641,N_24377,N_24998);
or UO_642 (O_642,N_24983,N_24761);
nor UO_643 (O_643,N_24525,N_24988);
xnor UO_644 (O_644,N_24210,N_24941);
nand UO_645 (O_645,N_24121,N_24397);
nor UO_646 (O_646,N_24139,N_24101);
nand UO_647 (O_647,N_24018,N_24879);
nor UO_648 (O_648,N_24016,N_24316);
xor UO_649 (O_649,N_24090,N_24634);
or UO_650 (O_650,N_24187,N_24290);
xnor UO_651 (O_651,N_24118,N_24665);
or UO_652 (O_652,N_24418,N_24461);
nand UO_653 (O_653,N_24765,N_24679);
xor UO_654 (O_654,N_24368,N_24178);
or UO_655 (O_655,N_24212,N_24037);
and UO_656 (O_656,N_24762,N_24934);
nand UO_657 (O_657,N_24990,N_24410);
nor UO_658 (O_658,N_24100,N_24665);
or UO_659 (O_659,N_24566,N_24717);
or UO_660 (O_660,N_24477,N_24898);
nor UO_661 (O_661,N_24286,N_24359);
nor UO_662 (O_662,N_24566,N_24907);
nand UO_663 (O_663,N_24339,N_24170);
nand UO_664 (O_664,N_24595,N_24817);
nand UO_665 (O_665,N_24897,N_24804);
nand UO_666 (O_666,N_24554,N_24178);
nand UO_667 (O_667,N_24247,N_24408);
or UO_668 (O_668,N_24421,N_24720);
xor UO_669 (O_669,N_24244,N_24554);
nand UO_670 (O_670,N_24742,N_24227);
xor UO_671 (O_671,N_24140,N_24420);
nor UO_672 (O_672,N_24502,N_24268);
or UO_673 (O_673,N_24624,N_24671);
nor UO_674 (O_674,N_24439,N_24783);
nor UO_675 (O_675,N_24291,N_24827);
nand UO_676 (O_676,N_24951,N_24163);
nor UO_677 (O_677,N_24218,N_24838);
and UO_678 (O_678,N_24268,N_24524);
or UO_679 (O_679,N_24960,N_24636);
or UO_680 (O_680,N_24408,N_24363);
or UO_681 (O_681,N_24742,N_24792);
nand UO_682 (O_682,N_24931,N_24633);
nand UO_683 (O_683,N_24112,N_24651);
and UO_684 (O_684,N_24103,N_24224);
nor UO_685 (O_685,N_24124,N_24216);
nor UO_686 (O_686,N_24549,N_24053);
or UO_687 (O_687,N_24374,N_24408);
nor UO_688 (O_688,N_24711,N_24729);
and UO_689 (O_689,N_24197,N_24708);
nor UO_690 (O_690,N_24789,N_24248);
or UO_691 (O_691,N_24706,N_24049);
xor UO_692 (O_692,N_24586,N_24198);
and UO_693 (O_693,N_24293,N_24641);
nand UO_694 (O_694,N_24267,N_24694);
and UO_695 (O_695,N_24048,N_24273);
nand UO_696 (O_696,N_24116,N_24133);
and UO_697 (O_697,N_24968,N_24041);
nor UO_698 (O_698,N_24644,N_24495);
nand UO_699 (O_699,N_24841,N_24299);
xnor UO_700 (O_700,N_24564,N_24790);
xor UO_701 (O_701,N_24348,N_24441);
nand UO_702 (O_702,N_24900,N_24100);
xnor UO_703 (O_703,N_24107,N_24048);
and UO_704 (O_704,N_24546,N_24539);
xor UO_705 (O_705,N_24577,N_24850);
or UO_706 (O_706,N_24734,N_24764);
or UO_707 (O_707,N_24609,N_24113);
nand UO_708 (O_708,N_24212,N_24879);
nor UO_709 (O_709,N_24803,N_24269);
xnor UO_710 (O_710,N_24631,N_24411);
or UO_711 (O_711,N_24046,N_24797);
or UO_712 (O_712,N_24019,N_24177);
xor UO_713 (O_713,N_24756,N_24583);
nand UO_714 (O_714,N_24341,N_24915);
nor UO_715 (O_715,N_24091,N_24570);
nor UO_716 (O_716,N_24838,N_24137);
xnor UO_717 (O_717,N_24616,N_24890);
and UO_718 (O_718,N_24140,N_24199);
nor UO_719 (O_719,N_24780,N_24525);
nand UO_720 (O_720,N_24225,N_24131);
nand UO_721 (O_721,N_24012,N_24841);
nor UO_722 (O_722,N_24426,N_24570);
nor UO_723 (O_723,N_24369,N_24292);
nor UO_724 (O_724,N_24809,N_24428);
nor UO_725 (O_725,N_24621,N_24204);
xnor UO_726 (O_726,N_24778,N_24809);
and UO_727 (O_727,N_24709,N_24184);
xor UO_728 (O_728,N_24666,N_24958);
or UO_729 (O_729,N_24407,N_24727);
or UO_730 (O_730,N_24945,N_24823);
and UO_731 (O_731,N_24580,N_24852);
and UO_732 (O_732,N_24547,N_24231);
nor UO_733 (O_733,N_24856,N_24306);
xor UO_734 (O_734,N_24815,N_24919);
xor UO_735 (O_735,N_24800,N_24460);
nand UO_736 (O_736,N_24024,N_24424);
and UO_737 (O_737,N_24302,N_24133);
nand UO_738 (O_738,N_24214,N_24327);
or UO_739 (O_739,N_24673,N_24150);
nor UO_740 (O_740,N_24490,N_24345);
nor UO_741 (O_741,N_24031,N_24649);
nor UO_742 (O_742,N_24614,N_24917);
nand UO_743 (O_743,N_24602,N_24572);
and UO_744 (O_744,N_24238,N_24370);
or UO_745 (O_745,N_24406,N_24963);
xor UO_746 (O_746,N_24890,N_24087);
and UO_747 (O_747,N_24151,N_24963);
or UO_748 (O_748,N_24369,N_24298);
nand UO_749 (O_749,N_24584,N_24179);
nor UO_750 (O_750,N_24219,N_24683);
or UO_751 (O_751,N_24977,N_24862);
or UO_752 (O_752,N_24097,N_24762);
or UO_753 (O_753,N_24294,N_24576);
nand UO_754 (O_754,N_24148,N_24339);
and UO_755 (O_755,N_24926,N_24229);
or UO_756 (O_756,N_24080,N_24558);
xor UO_757 (O_757,N_24103,N_24888);
nand UO_758 (O_758,N_24656,N_24197);
xnor UO_759 (O_759,N_24411,N_24421);
and UO_760 (O_760,N_24728,N_24122);
or UO_761 (O_761,N_24743,N_24398);
or UO_762 (O_762,N_24734,N_24808);
or UO_763 (O_763,N_24009,N_24115);
or UO_764 (O_764,N_24590,N_24462);
nand UO_765 (O_765,N_24604,N_24829);
and UO_766 (O_766,N_24894,N_24484);
and UO_767 (O_767,N_24546,N_24105);
and UO_768 (O_768,N_24671,N_24987);
and UO_769 (O_769,N_24602,N_24574);
nor UO_770 (O_770,N_24505,N_24567);
nand UO_771 (O_771,N_24896,N_24367);
nand UO_772 (O_772,N_24053,N_24398);
nand UO_773 (O_773,N_24587,N_24260);
and UO_774 (O_774,N_24883,N_24414);
nand UO_775 (O_775,N_24570,N_24448);
nand UO_776 (O_776,N_24245,N_24266);
xor UO_777 (O_777,N_24212,N_24986);
xnor UO_778 (O_778,N_24726,N_24146);
nand UO_779 (O_779,N_24562,N_24173);
nand UO_780 (O_780,N_24890,N_24157);
nor UO_781 (O_781,N_24690,N_24085);
nand UO_782 (O_782,N_24667,N_24870);
nor UO_783 (O_783,N_24474,N_24824);
xor UO_784 (O_784,N_24639,N_24235);
xor UO_785 (O_785,N_24813,N_24657);
or UO_786 (O_786,N_24012,N_24242);
xnor UO_787 (O_787,N_24208,N_24148);
xnor UO_788 (O_788,N_24891,N_24375);
nor UO_789 (O_789,N_24712,N_24448);
nor UO_790 (O_790,N_24334,N_24221);
and UO_791 (O_791,N_24899,N_24621);
and UO_792 (O_792,N_24774,N_24389);
nor UO_793 (O_793,N_24385,N_24298);
xnor UO_794 (O_794,N_24780,N_24060);
nor UO_795 (O_795,N_24181,N_24924);
nor UO_796 (O_796,N_24985,N_24108);
xor UO_797 (O_797,N_24808,N_24379);
xnor UO_798 (O_798,N_24321,N_24091);
nand UO_799 (O_799,N_24099,N_24379);
nor UO_800 (O_800,N_24111,N_24199);
and UO_801 (O_801,N_24704,N_24675);
xor UO_802 (O_802,N_24568,N_24998);
or UO_803 (O_803,N_24651,N_24352);
nand UO_804 (O_804,N_24052,N_24414);
or UO_805 (O_805,N_24300,N_24192);
nor UO_806 (O_806,N_24301,N_24052);
nor UO_807 (O_807,N_24353,N_24868);
or UO_808 (O_808,N_24218,N_24896);
xnor UO_809 (O_809,N_24598,N_24078);
and UO_810 (O_810,N_24795,N_24331);
and UO_811 (O_811,N_24051,N_24331);
nor UO_812 (O_812,N_24865,N_24113);
and UO_813 (O_813,N_24389,N_24901);
nor UO_814 (O_814,N_24117,N_24504);
or UO_815 (O_815,N_24993,N_24701);
or UO_816 (O_816,N_24770,N_24326);
and UO_817 (O_817,N_24941,N_24398);
nor UO_818 (O_818,N_24725,N_24629);
nor UO_819 (O_819,N_24905,N_24744);
and UO_820 (O_820,N_24806,N_24261);
and UO_821 (O_821,N_24105,N_24558);
and UO_822 (O_822,N_24449,N_24093);
and UO_823 (O_823,N_24069,N_24943);
or UO_824 (O_824,N_24230,N_24839);
and UO_825 (O_825,N_24142,N_24613);
nand UO_826 (O_826,N_24458,N_24010);
or UO_827 (O_827,N_24105,N_24901);
nor UO_828 (O_828,N_24182,N_24045);
nand UO_829 (O_829,N_24441,N_24869);
or UO_830 (O_830,N_24905,N_24030);
nor UO_831 (O_831,N_24554,N_24283);
nor UO_832 (O_832,N_24609,N_24005);
and UO_833 (O_833,N_24416,N_24274);
and UO_834 (O_834,N_24066,N_24605);
nand UO_835 (O_835,N_24613,N_24325);
nand UO_836 (O_836,N_24697,N_24109);
and UO_837 (O_837,N_24419,N_24964);
or UO_838 (O_838,N_24145,N_24931);
nand UO_839 (O_839,N_24991,N_24543);
nand UO_840 (O_840,N_24888,N_24367);
and UO_841 (O_841,N_24998,N_24113);
nand UO_842 (O_842,N_24315,N_24033);
or UO_843 (O_843,N_24982,N_24930);
or UO_844 (O_844,N_24024,N_24081);
nor UO_845 (O_845,N_24904,N_24749);
or UO_846 (O_846,N_24457,N_24678);
and UO_847 (O_847,N_24947,N_24341);
nor UO_848 (O_848,N_24098,N_24377);
and UO_849 (O_849,N_24085,N_24040);
nand UO_850 (O_850,N_24052,N_24905);
or UO_851 (O_851,N_24418,N_24232);
xor UO_852 (O_852,N_24901,N_24341);
nand UO_853 (O_853,N_24588,N_24163);
or UO_854 (O_854,N_24789,N_24293);
xnor UO_855 (O_855,N_24520,N_24872);
xnor UO_856 (O_856,N_24833,N_24544);
nand UO_857 (O_857,N_24323,N_24264);
nand UO_858 (O_858,N_24951,N_24511);
nand UO_859 (O_859,N_24186,N_24505);
nand UO_860 (O_860,N_24522,N_24693);
and UO_861 (O_861,N_24743,N_24445);
and UO_862 (O_862,N_24674,N_24162);
or UO_863 (O_863,N_24143,N_24434);
nand UO_864 (O_864,N_24309,N_24410);
or UO_865 (O_865,N_24467,N_24141);
xor UO_866 (O_866,N_24422,N_24095);
and UO_867 (O_867,N_24958,N_24063);
nor UO_868 (O_868,N_24989,N_24588);
and UO_869 (O_869,N_24403,N_24219);
xor UO_870 (O_870,N_24163,N_24748);
nor UO_871 (O_871,N_24663,N_24317);
nor UO_872 (O_872,N_24356,N_24671);
and UO_873 (O_873,N_24792,N_24981);
and UO_874 (O_874,N_24373,N_24056);
or UO_875 (O_875,N_24540,N_24606);
or UO_876 (O_876,N_24593,N_24862);
or UO_877 (O_877,N_24712,N_24080);
or UO_878 (O_878,N_24455,N_24353);
xnor UO_879 (O_879,N_24821,N_24076);
or UO_880 (O_880,N_24788,N_24492);
or UO_881 (O_881,N_24835,N_24377);
nor UO_882 (O_882,N_24082,N_24553);
nand UO_883 (O_883,N_24013,N_24899);
nand UO_884 (O_884,N_24574,N_24353);
nor UO_885 (O_885,N_24289,N_24418);
nor UO_886 (O_886,N_24534,N_24327);
or UO_887 (O_887,N_24351,N_24921);
and UO_888 (O_888,N_24835,N_24218);
and UO_889 (O_889,N_24332,N_24148);
and UO_890 (O_890,N_24328,N_24359);
or UO_891 (O_891,N_24197,N_24463);
nand UO_892 (O_892,N_24798,N_24871);
and UO_893 (O_893,N_24280,N_24340);
and UO_894 (O_894,N_24658,N_24476);
xor UO_895 (O_895,N_24881,N_24660);
and UO_896 (O_896,N_24386,N_24405);
and UO_897 (O_897,N_24824,N_24796);
xor UO_898 (O_898,N_24958,N_24827);
nand UO_899 (O_899,N_24169,N_24621);
xor UO_900 (O_900,N_24000,N_24842);
nand UO_901 (O_901,N_24099,N_24572);
nor UO_902 (O_902,N_24751,N_24599);
xor UO_903 (O_903,N_24387,N_24256);
xor UO_904 (O_904,N_24284,N_24586);
or UO_905 (O_905,N_24171,N_24856);
or UO_906 (O_906,N_24105,N_24179);
or UO_907 (O_907,N_24904,N_24511);
or UO_908 (O_908,N_24774,N_24799);
or UO_909 (O_909,N_24322,N_24288);
nor UO_910 (O_910,N_24128,N_24759);
or UO_911 (O_911,N_24023,N_24793);
and UO_912 (O_912,N_24680,N_24121);
nor UO_913 (O_913,N_24989,N_24036);
nor UO_914 (O_914,N_24134,N_24890);
nand UO_915 (O_915,N_24031,N_24844);
nand UO_916 (O_916,N_24659,N_24104);
and UO_917 (O_917,N_24819,N_24065);
or UO_918 (O_918,N_24550,N_24492);
or UO_919 (O_919,N_24269,N_24454);
nor UO_920 (O_920,N_24188,N_24401);
xor UO_921 (O_921,N_24066,N_24874);
or UO_922 (O_922,N_24979,N_24984);
and UO_923 (O_923,N_24048,N_24658);
or UO_924 (O_924,N_24389,N_24087);
nand UO_925 (O_925,N_24257,N_24501);
nand UO_926 (O_926,N_24797,N_24673);
and UO_927 (O_927,N_24806,N_24786);
xor UO_928 (O_928,N_24814,N_24828);
nor UO_929 (O_929,N_24187,N_24759);
xnor UO_930 (O_930,N_24998,N_24491);
or UO_931 (O_931,N_24916,N_24783);
xor UO_932 (O_932,N_24817,N_24823);
xnor UO_933 (O_933,N_24315,N_24433);
and UO_934 (O_934,N_24382,N_24028);
and UO_935 (O_935,N_24688,N_24653);
xnor UO_936 (O_936,N_24685,N_24754);
nor UO_937 (O_937,N_24153,N_24975);
and UO_938 (O_938,N_24853,N_24333);
and UO_939 (O_939,N_24184,N_24635);
xor UO_940 (O_940,N_24555,N_24268);
nand UO_941 (O_941,N_24574,N_24228);
or UO_942 (O_942,N_24008,N_24602);
nor UO_943 (O_943,N_24419,N_24043);
or UO_944 (O_944,N_24551,N_24039);
or UO_945 (O_945,N_24051,N_24597);
or UO_946 (O_946,N_24566,N_24434);
or UO_947 (O_947,N_24948,N_24244);
nor UO_948 (O_948,N_24649,N_24035);
and UO_949 (O_949,N_24794,N_24822);
and UO_950 (O_950,N_24643,N_24574);
and UO_951 (O_951,N_24298,N_24121);
or UO_952 (O_952,N_24911,N_24877);
xnor UO_953 (O_953,N_24641,N_24060);
nand UO_954 (O_954,N_24819,N_24661);
xnor UO_955 (O_955,N_24682,N_24679);
and UO_956 (O_956,N_24653,N_24974);
nand UO_957 (O_957,N_24999,N_24673);
nand UO_958 (O_958,N_24078,N_24348);
xor UO_959 (O_959,N_24256,N_24042);
xnor UO_960 (O_960,N_24395,N_24201);
xnor UO_961 (O_961,N_24348,N_24621);
nand UO_962 (O_962,N_24170,N_24654);
nand UO_963 (O_963,N_24339,N_24052);
nand UO_964 (O_964,N_24447,N_24782);
or UO_965 (O_965,N_24301,N_24265);
nor UO_966 (O_966,N_24311,N_24034);
nand UO_967 (O_967,N_24897,N_24493);
and UO_968 (O_968,N_24809,N_24993);
or UO_969 (O_969,N_24818,N_24459);
xnor UO_970 (O_970,N_24891,N_24372);
nand UO_971 (O_971,N_24909,N_24845);
nand UO_972 (O_972,N_24182,N_24106);
and UO_973 (O_973,N_24323,N_24318);
and UO_974 (O_974,N_24995,N_24402);
or UO_975 (O_975,N_24818,N_24781);
nor UO_976 (O_976,N_24781,N_24843);
xor UO_977 (O_977,N_24196,N_24968);
nor UO_978 (O_978,N_24804,N_24926);
and UO_979 (O_979,N_24584,N_24214);
and UO_980 (O_980,N_24398,N_24545);
or UO_981 (O_981,N_24181,N_24199);
xnor UO_982 (O_982,N_24793,N_24382);
or UO_983 (O_983,N_24744,N_24461);
or UO_984 (O_984,N_24493,N_24676);
xnor UO_985 (O_985,N_24719,N_24478);
and UO_986 (O_986,N_24773,N_24315);
nand UO_987 (O_987,N_24005,N_24986);
or UO_988 (O_988,N_24952,N_24155);
and UO_989 (O_989,N_24270,N_24956);
and UO_990 (O_990,N_24320,N_24786);
and UO_991 (O_991,N_24274,N_24982);
or UO_992 (O_992,N_24351,N_24211);
nand UO_993 (O_993,N_24818,N_24926);
xor UO_994 (O_994,N_24949,N_24683);
nor UO_995 (O_995,N_24436,N_24636);
nor UO_996 (O_996,N_24667,N_24441);
nand UO_997 (O_997,N_24940,N_24315);
nand UO_998 (O_998,N_24763,N_24888);
or UO_999 (O_999,N_24385,N_24427);
nand UO_1000 (O_1000,N_24971,N_24410);
and UO_1001 (O_1001,N_24512,N_24406);
xnor UO_1002 (O_1002,N_24831,N_24285);
nand UO_1003 (O_1003,N_24585,N_24554);
and UO_1004 (O_1004,N_24884,N_24160);
xnor UO_1005 (O_1005,N_24879,N_24776);
and UO_1006 (O_1006,N_24949,N_24294);
and UO_1007 (O_1007,N_24345,N_24086);
nand UO_1008 (O_1008,N_24753,N_24918);
nor UO_1009 (O_1009,N_24632,N_24763);
nand UO_1010 (O_1010,N_24608,N_24431);
and UO_1011 (O_1011,N_24148,N_24405);
xor UO_1012 (O_1012,N_24957,N_24934);
and UO_1013 (O_1013,N_24645,N_24101);
nor UO_1014 (O_1014,N_24877,N_24424);
xnor UO_1015 (O_1015,N_24024,N_24705);
xor UO_1016 (O_1016,N_24521,N_24232);
nand UO_1017 (O_1017,N_24636,N_24244);
and UO_1018 (O_1018,N_24709,N_24620);
and UO_1019 (O_1019,N_24562,N_24346);
nor UO_1020 (O_1020,N_24366,N_24610);
and UO_1021 (O_1021,N_24987,N_24760);
xnor UO_1022 (O_1022,N_24472,N_24479);
or UO_1023 (O_1023,N_24628,N_24154);
nand UO_1024 (O_1024,N_24644,N_24930);
or UO_1025 (O_1025,N_24287,N_24121);
nand UO_1026 (O_1026,N_24607,N_24760);
or UO_1027 (O_1027,N_24035,N_24302);
or UO_1028 (O_1028,N_24942,N_24021);
nand UO_1029 (O_1029,N_24005,N_24599);
xor UO_1030 (O_1030,N_24044,N_24019);
nand UO_1031 (O_1031,N_24259,N_24105);
xnor UO_1032 (O_1032,N_24922,N_24426);
or UO_1033 (O_1033,N_24842,N_24767);
xor UO_1034 (O_1034,N_24948,N_24693);
or UO_1035 (O_1035,N_24819,N_24300);
nor UO_1036 (O_1036,N_24976,N_24361);
or UO_1037 (O_1037,N_24072,N_24573);
or UO_1038 (O_1038,N_24412,N_24254);
nand UO_1039 (O_1039,N_24650,N_24536);
xnor UO_1040 (O_1040,N_24927,N_24420);
nand UO_1041 (O_1041,N_24369,N_24704);
nand UO_1042 (O_1042,N_24909,N_24459);
nor UO_1043 (O_1043,N_24771,N_24571);
or UO_1044 (O_1044,N_24633,N_24307);
nor UO_1045 (O_1045,N_24057,N_24116);
or UO_1046 (O_1046,N_24300,N_24608);
and UO_1047 (O_1047,N_24816,N_24411);
or UO_1048 (O_1048,N_24068,N_24822);
or UO_1049 (O_1049,N_24865,N_24164);
xnor UO_1050 (O_1050,N_24578,N_24594);
nor UO_1051 (O_1051,N_24135,N_24281);
nor UO_1052 (O_1052,N_24636,N_24717);
nor UO_1053 (O_1053,N_24663,N_24151);
nor UO_1054 (O_1054,N_24250,N_24416);
nand UO_1055 (O_1055,N_24065,N_24679);
or UO_1056 (O_1056,N_24694,N_24730);
nand UO_1057 (O_1057,N_24687,N_24932);
nor UO_1058 (O_1058,N_24032,N_24909);
nand UO_1059 (O_1059,N_24190,N_24996);
nand UO_1060 (O_1060,N_24634,N_24551);
nand UO_1061 (O_1061,N_24121,N_24575);
xor UO_1062 (O_1062,N_24464,N_24519);
nand UO_1063 (O_1063,N_24262,N_24310);
nand UO_1064 (O_1064,N_24357,N_24373);
nand UO_1065 (O_1065,N_24249,N_24756);
and UO_1066 (O_1066,N_24223,N_24848);
xor UO_1067 (O_1067,N_24817,N_24701);
nor UO_1068 (O_1068,N_24069,N_24042);
nand UO_1069 (O_1069,N_24848,N_24266);
and UO_1070 (O_1070,N_24002,N_24297);
nor UO_1071 (O_1071,N_24985,N_24081);
nor UO_1072 (O_1072,N_24788,N_24490);
xnor UO_1073 (O_1073,N_24311,N_24465);
and UO_1074 (O_1074,N_24843,N_24493);
xnor UO_1075 (O_1075,N_24968,N_24909);
and UO_1076 (O_1076,N_24886,N_24971);
or UO_1077 (O_1077,N_24849,N_24457);
xnor UO_1078 (O_1078,N_24872,N_24075);
nor UO_1079 (O_1079,N_24748,N_24448);
xnor UO_1080 (O_1080,N_24727,N_24840);
and UO_1081 (O_1081,N_24795,N_24085);
xnor UO_1082 (O_1082,N_24557,N_24999);
nor UO_1083 (O_1083,N_24532,N_24962);
and UO_1084 (O_1084,N_24606,N_24932);
xor UO_1085 (O_1085,N_24671,N_24174);
nor UO_1086 (O_1086,N_24777,N_24215);
nand UO_1087 (O_1087,N_24133,N_24776);
nand UO_1088 (O_1088,N_24186,N_24197);
xor UO_1089 (O_1089,N_24267,N_24965);
and UO_1090 (O_1090,N_24402,N_24429);
nand UO_1091 (O_1091,N_24887,N_24106);
and UO_1092 (O_1092,N_24646,N_24510);
or UO_1093 (O_1093,N_24482,N_24591);
nor UO_1094 (O_1094,N_24737,N_24498);
xnor UO_1095 (O_1095,N_24630,N_24094);
xnor UO_1096 (O_1096,N_24544,N_24348);
nand UO_1097 (O_1097,N_24347,N_24573);
xor UO_1098 (O_1098,N_24750,N_24115);
and UO_1099 (O_1099,N_24320,N_24010);
xor UO_1100 (O_1100,N_24277,N_24457);
or UO_1101 (O_1101,N_24787,N_24596);
nor UO_1102 (O_1102,N_24526,N_24799);
nor UO_1103 (O_1103,N_24448,N_24780);
nor UO_1104 (O_1104,N_24534,N_24462);
nor UO_1105 (O_1105,N_24746,N_24178);
nor UO_1106 (O_1106,N_24106,N_24935);
or UO_1107 (O_1107,N_24265,N_24644);
nand UO_1108 (O_1108,N_24565,N_24201);
and UO_1109 (O_1109,N_24237,N_24505);
xor UO_1110 (O_1110,N_24993,N_24587);
nor UO_1111 (O_1111,N_24434,N_24580);
nor UO_1112 (O_1112,N_24533,N_24482);
nand UO_1113 (O_1113,N_24735,N_24364);
and UO_1114 (O_1114,N_24626,N_24609);
xor UO_1115 (O_1115,N_24481,N_24182);
xnor UO_1116 (O_1116,N_24811,N_24156);
xor UO_1117 (O_1117,N_24112,N_24195);
nand UO_1118 (O_1118,N_24648,N_24998);
nor UO_1119 (O_1119,N_24071,N_24515);
and UO_1120 (O_1120,N_24627,N_24428);
nand UO_1121 (O_1121,N_24057,N_24014);
nor UO_1122 (O_1122,N_24950,N_24510);
xor UO_1123 (O_1123,N_24021,N_24853);
nand UO_1124 (O_1124,N_24057,N_24679);
nor UO_1125 (O_1125,N_24181,N_24881);
or UO_1126 (O_1126,N_24407,N_24527);
nand UO_1127 (O_1127,N_24312,N_24799);
nand UO_1128 (O_1128,N_24390,N_24303);
nand UO_1129 (O_1129,N_24508,N_24784);
nand UO_1130 (O_1130,N_24961,N_24416);
nor UO_1131 (O_1131,N_24439,N_24450);
nor UO_1132 (O_1132,N_24304,N_24356);
xor UO_1133 (O_1133,N_24993,N_24225);
or UO_1134 (O_1134,N_24277,N_24350);
nand UO_1135 (O_1135,N_24919,N_24871);
xor UO_1136 (O_1136,N_24718,N_24825);
nand UO_1137 (O_1137,N_24615,N_24381);
and UO_1138 (O_1138,N_24003,N_24594);
or UO_1139 (O_1139,N_24148,N_24432);
and UO_1140 (O_1140,N_24993,N_24794);
or UO_1141 (O_1141,N_24425,N_24154);
or UO_1142 (O_1142,N_24752,N_24421);
or UO_1143 (O_1143,N_24652,N_24653);
or UO_1144 (O_1144,N_24724,N_24677);
nor UO_1145 (O_1145,N_24680,N_24001);
and UO_1146 (O_1146,N_24324,N_24774);
xnor UO_1147 (O_1147,N_24074,N_24766);
xnor UO_1148 (O_1148,N_24376,N_24094);
nand UO_1149 (O_1149,N_24682,N_24876);
xnor UO_1150 (O_1150,N_24872,N_24863);
nor UO_1151 (O_1151,N_24145,N_24710);
nor UO_1152 (O_1152,N_24583,N_24656);
nand UO_1153 (O_1153,N_24117,N_24295);
nor UO_1154 (O_1154,N_24401,N_24255);
or UO_1155 (O_1155,N_24509,N_24267);
and UO_1156 (O_1156,N_24140,N_24681);
or UO_1157 (O_1157,N_24537,N_24478);
and UO_1158 (O_1158,N_24596,N_24739);
nor UO_1159 (O_1159,N_24422,N_24402);
nor UO_1160 (O_1160,N_24942,N_24656);
and UO_1161 (O_1161,N_24727,N_24739);
nor UO_1162 (O_1162,N_24184,N_24457);
nor UO_1163 (O_1163,N_24922,N_24905);
or UO_1164 (O_1164,N_24329,N_24354);
or UO_1165 (O_1165,N_24538,N_24269);
nor UO_1166 (O_1166,N_24157,N_24726);
xnor UO_1167 (O_1167,N_24138,N_24078);
nand UO_1168 (O_1168,N_24090,N_24599);
or UO_1169 (O_1169,N_24294,N_24276);
nor UO_1170 (O_1170,N_24969,N_24020);
nand UO_1171 (O_1171,N_24930,N_24684);
and UO_1172 (O_1172,N_24556,N_24965);
or UO_1173 (O_1173,N_24888,N_24080);
xor UO_1174 (O_1174,N_24977,N_24055);
or UO_1175 (O_1175,N_24494,N_24485);
nand UO_1176 (O_1176,N_24856,N_24646);
and UO_1177 (O_1177,N_24321,N_24302);
xnor UO_1178 (O_1178,N_24689,N_24674);
nand UO_1179 (O_1179,N_24510,N_24871);
and UO_1180 (O_1180,N_24680,N_24661);
nor UO_1181 (O_1181,N_24444,N_24386);
and UO_1182 (O_1182,N_24077,N_24917);
xnor UO_1183 (O_1183,N_24506,N_24438);
nor UO_1184 (O_1184,N_24387,N_24499);
and UO_1185 (O_1185,N_24149,N_24562);
nand UO_1186 (O_1186,N_24737,N_24340);
and UO_1187 (O_1187,N_24746,N_24314);
xor UO_1188 (O_1188,N_24259,N_24742);
or UO_1189 (O_1189,N_24591,N_24029);
nand UO_1190 (O_1190,N_24916,N_24496);
nand UO_1191 (O_1191,N_24421,N_24229);
and UO_1192 (O_1192,N_24616,N_24831);
and UO_1193 (O_1193,N_24755,N_24663);
and UO_1194 (O_1194,N_24811,N_24495);
or UO_1195 (O_1195,N_24202,N_24879);
xnor UO_1196 (O_1196,N_24122,N_24850);
and UO_1197 (O_1197,N_24540,N_24798);
or UO_1198 (O_1198,N_24487,N_24013);
xnor UO_1199 (O_1199,N_24382,N_24159);
xor UO_1200 (O_1200,N_24020,N_24817);
and UO_1201 (O_1201,N_24898,N_24356);
xor UO_1202 (O_1202,N_24853,N_24226);
and UO_1203 (O_1203,N_24193,N_24565);
nand UO_1204 (O_1204,N_24293,N_24400);
nand UO_1205 (O_1205,N_24442,N_24079);
xnor UO_1206 (O_1206,N_24765,N_24354);
nor UO_1207 (O_1207,N_24209,N_24793);
nor UO_1208 (O_1208,N_24642,N_24576);
nor UO_1209 (O_1209,N_24219,N_24956);
nor UO_1210 (O_1210,N_24976,N_24852);
xor UO_1211 (O_1211,N_24552,N_24378);
nand UO_1212 (O_1212,N_24279,N_24771);
nor UO_1213 (O_1213,N_24955,N_24203);
and UO_1214 (O_1214,N_24233,N_24488);
nand UO_1215 (O_1215,N_24847,N_24575);
nor UO_1216 (O_1216,N_24783,N_24032);
and UO_1217 (O_1217,N_24050,N_24558);
nor UO_1218 (O_1218,N_24285,N_24578);
or UO_1219 (O_1219,N_24406,N_24147);
or UO_1220 (O_1220,N_24515,N_24979);
xnor UO_1221 (O_1221,N_24242,N_24829);
nand UO_1222 (O_1222,N_24833,N_24864);
nor UO_1223 (O_1223,N_24006,N_24206);
nor UO_1224 (O_1224,N_24249,N_24366);
or UO_1225 (O_1225,N_24188,N_24159);
xor UO_1226 (O_1226,N_24962,N_24148);
or UO_1227 (O_1227,N_24664,N_24139);
and UO_1228 (O_1228,N_24408,N_24604);
and UO_1229 (O_1229,N_24572,N_24862);
nand UO_1230 (O_1230,N_24274,N_24408);
or UO_1231 (O_1231,N_24140,N_24224);
nor UO_1232 (O_1232,N_24234,N_24049);
xnor UO_1233 (O_1233,N_24298,N_24449);
or UO_1234 (O_1234,N_24497,N_24674);
or UO_1235 (O_1235,N_24708,N_24150);
nand UO_1236 (O_1236,N_24936,N_24726);
nor UO_1237 (O_1237,N_24033,N_24800);
nand UO_1238 (O_1238,N_24286,N_24584);
or UO_1239 (O_1239,N_24037,N_24922);
or UO_1240 (O_1240,N_24134,N_24834);
and UO_1241 (O_1241,N_24954,N_24461);
nor UO_1242 (O_1242,N_24420,N_24966);
and UO_1243 (O_1243,N_24559,N_24104);
nand UO_1244 (O_1244,N_24481,N_24021);
xnor UO_1245 (O_1245,N_24539,N_24487);
xnor UO_1246 (O_1246,N_24801,N_24061);
nand UO_1247 (O_1247,N_24258,N_24442);
nor UO_1248 (O_1248,N_24528,N_24706);
nand UO_1249 (O_1249,N_24295,N_24394);
nor UO_1250 (O_1250,N_24135,N_24543);
nand UO_1251 (O_1251,N_24219,N_24107);
xor UO_1252 (O_1252,N_24632,N_24200);
xnor UO_1253 (O_1253,N_24367,N_24524);
xor UO_1254 (O_1254,N_24031,N_24834);
and UO_1255 (O_1255,N_24288,N_24581);
or UO_1256 (O_1256,N_24718,N_24023);
and UO_1257 (O_1257,N_24277,N_24871);
xor UO_1258 (O_1258,N_24532,N_24127);
nor UO_1259 (O_1259,N_24720,N_24179);
nand UO_1260 (O_1260,N_24923,N_24451);
and UO_1261 (O_1261,N_24533,N_24917);
nand UO_1262 (O_1262,N_24793,N_24356);
nor UO_1263 (O_1263,N_24695,N_24203);
nor UO_1264 (O_1264,N_24651,N_24336);
nand UO_1265 (O_1265,N_24079,N_24335);
or UO_1266 (O_1266,N_24472,N_24184);
or UO_1267 (O_1267,N_24736,N_24650);
and UO_1268 (O_1268,N_24808,N_24877);
nand UO_1269 (O_1269,N_24532,N_24055);
or UO_1270 (O_1270,N_24714,N_24027);
or UO_1271 (O_1271,N_24867,N_24291);
nor UO_1272 (O_1272,N_24467,N_24192);
nor UO_1273 (O_1273,N_24908,N_24525);
nor UO_1274 (O_1274,N_24382,N_24349);
nand UO_1275 (O_1275,N_24164,N_24796);
nand UO_1276 (O_1276,N_24574,N_24227);
nand UO_1277 (O_1277,N_24011,N_24609);
nand UO_1278 (O_1278,N_24002,N_24470);
nor UO_1279 (O_1279,N_24159,N_24344);
and UO_1280 (O_1280,N_24380,N_24815);
or UO_1281 (O_1281,N_24151,N_24744);
or UO_1282 (O_1282,N_24645,N_24928);
nand UO_1283 (O_1283,N_24428,N_24493);
or UO_1284 (O_1284,N_24648,N_24439);
nand UO_1285 (O_1285,N_24449,N_24579);
nand UO_1286 (O_1286,N_24256,N_24317);
nor UO_1287 (O_1287,N_24326,N_24861);
xor UO_1288 (O_1288,N_24607,N_24853);
or UO_1289 (O_1289,N_24999,N_24526);
or UO_1290 (O_1290,N_24665,N_24750);
and UO_1291 (O_1291,N_24921,N_24280);
or UO_1292 (O_1292,N_24550,N_24399);
nor UO_1293 (O_1293,N_24146,N_24101);
or UO_1294 (O_1294,N_24156,N_24767);
and UO_1295 (O_1295,N_24089,N_24566);
nor UO_1296 (O_1296,N_24944,N_24917);
or UO_1297 (O_1297,N_24500,N_24840);
and UO_1298 (O_1298,N_24484,N_24815);
nor UO_1299 (O_1299,N_24656,N_24680);
or UO_1300 (O_1300,N_24404,N_24885);
nand UO_1301 (O_1301,N_24830,N_24792);
xnor UO_1302 (O_1302,N_24041,N_24165);
xnor UO_1303 (O_1303,N_24638,N_24829);
nand UO_1304 (O_1304,N_24794,N_24475);
and UO_1305 (O_1305,N_24491,N_24371);
and UO_1306 (O_1306,N_24097,N_24159);
and UO_1307 (O_1307,N_24459,N_24550);
xnor UO_1308 (O_1308,N_24236,N_24496);
nand UO_1309 (O_1309,N_24870,N_24892);
and UO_1310 (O_1310,N_24697,N_24202);
xnor UO_1311 (O_1311,N_24545,N_24875);
nand UO_1312 (O_1312,N_24174,N_24858);
xor UO_1313 (O_1313,N_24772,N_24986);
or UO_1314 (O_1314,N_24595,N_24533);
and UO_1315 (O_1315,N_24926,N_24929);
nor UO_1316 (O_1316,N_24339,N_24561);
xnor UO_1317 (O_1317,N_24628,N_24494);
and UO_1318 (O_1318,N_24627,N_24957);
or UO_1319 (O_1319,N_24046,N_24729);
nand UO_1320 (O_1320,N_24371,N_24041);
nor UO_1321 (O_1321,N_24787,N_24908);
xnor UO_1322 (O_1322,N_24449,N_24849);
nand UO_1323 (O_1323,N_24966,N_24849);
nand UO_1324 (O_1324,N_24725,N_24803);
or UO_1325 (O_1325,N_24985,N_24314);
nor UO_1326 (O_1326,N_24037,N_24705);
nand UO_1327 (O_1327,N_24703,N_24990);
and UO_1328 (O_1328,N_24634,N_24613);
xnor UO_1329 (O_1329,N_24707,N_24809);
or UO_1330 (O_1330,N_24881,N_24960);
nand UO_1331 (O_1331,N_24284,N_24326);
and UO_1332 (O_1332,N_24736,N_24626);
xor UO_1333 (O_1333,N_24693,N_24985);
nor UO_1334 (O_1334,N_24692,N_24928);
xor UO_1335 (O_1335,N_24782,N_24509);
and UO_1336 (O_1336,N_24731,N_24574);
nand UO_1337 (O_1337,N_24950,N_24496);
and UO_1338 (O_1338,N_24965,N_24127);
nor UO_1339 (O_1339,N_24768,N_24516);
nor UO_1340 (O_1340,N_24664,N_24441);
xnor UO_1341 (O_1341,N_24894,N_24579);
nand UO_1342 (O_1342,N_24737,N_24960);
xnor UO_1343 (O_1343,N_24389,N_24822);
nand UO_1344 (O_1344,N_24013,N_24938);
nor UO_1345 (O_1345,N_24778,N_24670);
xnor UO_1346 (O_1346,N_24986,N_24111);
or UO_1347 (O_1347,N_24550,N_24907);
nor UO_1348 (O_1348,N_24891,N_24371);
or UO_1349 (O_1349,N_24947,N_24390);
and UO_1350 (O_1350,N_24938,N_24894);
or UO_1351 (O_1351,N_24999,N_24524);
and UO_1352 (O_1352,N_24076,N_24523);
nand UO_1353 (O_1353,N_24354,N_24250);
nor UO_1354 (O_1354,N_24021,N_24360);
xnor UO_1355 (O_1355,N_24335,N_24676);
nand UO_1356 (O_1356,N_24082,N_24807);
nor UO_1357 (O_1357,N_24867,N_24059);
xnor UO_1358 (O_1358,N_24508,N_24008);
and UO_1359 (O_1359,N_24325,N_24028);
or UO_1360 (O_1360,N_24131,N_24946);
nor UO_1361 (O_1361,N_24712,N_24320);
and UO_1362 (O_1362,N_24479,N_24508);
or UO_1363 (O_1363,N_24165,N_24096);
xor UO_1364 (O_1364,N_24284,N_24334);
or UO_1365 (O_1365,N_24368,N_24765);
nand UO_1366 (O_1366,N_24708,N_24888);
xor UO_1367 (O_1367,N_24971,N_24255);
nor UO_1368 (O_1368,N_24827,N_24480);
xnor UO_1369 (O_1369,N_24830,N_24700);
nor UO_1370 (O_1370,N_24083,N_24885);
and UO_1371 (O_1371,N_24052,N_24740);
and UO_1372 (O_1372,N_24283,N_24311);
nor UO_1373 (O_1373,N_24470,N_24790);
and UO_1374 (O_1374,N_24634,N_24329);
and UO_1375 (O_1375,N_24993,N_24382);
or UO_1376 (O_1376,N_24554,N_24813);
or UO_1377 (O_1377,N_24432,N_24746);
nand UO_1378 (O_1378,N_24796,N_24401);
xnor UO_1379 (O_1379,N_24493,N_24834);
or UO_1380 (O_1380,N_24960,N_24752);
nand UO_1381 (O_1381,N_24867,N_24287);
or UO_1382 (O_1382,N_24777,N_24001);
xnor UO_1383 (O_1383,N_24273,N_24165);
xnor UO_1384 (O_1384,N_24543,N_24335);
nor UO_1385 (O_1385,N_24599,N_24394);
xnor UO_1386 (O_1386,N_24987,N_24416);
nand UO_1387 (O_1387,N_24362,N_24137);
and UO_1388 (O_1388,N_24832,N_24811);
nor UO_1389 (O_1389,N_24393,N_24004);
nor UO_1390 (O_1390,N_24647,N_24218);
and UO_1391 (O_1391,N_24071,N_24883);
nor UO_1392 (O_1392,N_24936,N_24595);
xor UO_1393 (O_1393,N_24226,N_24374);
or UO_1394 (O_1394,N_24685,N_24790);
and UO_1395 (O_1395,N_24289,N_24260);
nand UO_1396 (O_1396,N_24340,N_24945);
and UO_1397 (O_1397,N_24905,N_24383);
nor UO_1398 (O_1398,N_24044,N_24074);
or UO_1399 (O_1399,N_24979,N_24813);
or UO_1400 (O_1400,N_24988,N_24449);
nor UO_1401 (O_1401,N_24388,N_24292);
and UO_1402 (O_1402,N_24761,N_24361);
xor UO_1403 (O_1403,N_24530,N_24923);
nand UO_1404 (O_1404,N_24107,N_24992);
nand UO_1405 (O_1405,N_24909,N_24220);
nand UO_1406 (O_1406,N_24676,N_24780);
nand UO_1407 (O_1407,N_24931,N_24777);
nor UO_1408 (O_1408,N_24808,N_24214);
or UO_1409 (O_1409,N_24279,N_24925);
xor UO_1410 (O_1410,N_24866,N_24207);
and UO_1411 (O_1411,N_24073,N_24191);
nand UO_1412 (O_1412,N_24106,N_24436);
nand UO_1413 (O_1413,N_24546,N_24774);
nor UO_1414 (O_1414,N_24202,N_24682);
xnor UO_1415 (O_1415,N_24505,N_24811);
or UO_1416 (O_1416,N_24251,N_24049);
nor UO_1417 (O_1417,N_24461,N_24077);
nand UO_1418 (O_1418,N_24273,N_24946);
nand UO_1419 (O_1419,N_24815,N_24822);
and UO_1420 (O_1420,N_24138,N_24056);
xnor UO_1421 (O_1421,N_24339,N_24189);
and UO_1422 (O_1422,N_24854,N_24693);
and UO_1423 (O_1423,N_24416,N_24535);
or UO_1424 (O_1424,N_24303,N_24818);
or UO_1425 (O_1425,N_24821,N_24363);
nor UO_1426 (O_1426,N_24613,N_24754);
and UO_1427 (O_1427,N_24496,N_24318);
nor UO_1428 (O_1428,N_24474,N_24823);
nor UO_1429 (O_1429,N_24544,N_24567);
nand UO_1430 (O_1430,N_24823,N_24693);
nor UO_1431 (O_1431,N_24524,N_24038);
xor UO_1432 (O_1432,N_24191,N_24389);
and UO_1433 (O_1433,N_24687,N_24477);
nor UO_1434 (O_1434,N_24005,N_24069);
and UO_1435 (O_1435,N_24484,N_24757);
xnor UO_1436 (O_1436,N_24934,N_24088);
xor UO_1437 (O_1437,N_24987,N_24532);
or UO_1438 (O_1438,N_24406,N_24975);
nand UO_1439 (O_1439,N_24384,N_24597);
or UO_1440 (O_1440,N_24470,N_24555);
nor UO_1441 (O_1441,N_24333,N_24265);
or UO_1442 (O_1442,N_24308,N_24539);
or UO_1443 (O_1443,N_24374,N_24106);
nand UO_1444 (O_1444,N_24135,N_24965);
or UO_1445 (O_1445,N_24274,N_24517);
nor UO_1446 (O_1446,N_24295,N_24234);
or UO_1447 (O_1447,N_24442,N_24456);
or UO_1448 (O_1448,N_24757,N_24882);
and UO_1449 (O_1449,N_24852,N_24813);
nand UO_1450 (O_1450,N_24105,N_24025);
nor UO_1451 (O_1451,N_24022,N_24877);
and UO_1452 (O_1452,N_24458,N_24033);
or UO_1453 (O_1453,N_24572,N_24297);
nand UO_1454 (O_1454,N_24588,N_24270);
or UO_1455 (O_1455,N_24778,N_24056);
or UO_1456 (O_1456,N_24894,N_24263);
nor UO_1457 (O_1457,N_24392,N_24983);
or UO_1458 (O_1458,N_24104,N_24371);
xor UO_1459 (O_1459,N_24379,N_24317);
nand UO_1460 (O_1460,N_24493,N_24999);
xor UO_1461 (O_1461,N_24355,N_24837);
xor UO_1462 (O_1462,N_24248,N_24395);
or UO_1463 (O_1463,N_24652,N_24803);
nor UO_1464 (O_1464,N_24628,N_24298);
or UO_1465 (O_1465,N_24022,N_24497);
nor UO_1466 (O_1466,N_24699,N_24126);
and UO_1467 (O_1467,N_24245,N_24808);
or UO_1468 (O_1468,N_24332,N_24786);
and UO_1469 (O_1469,N_24545,N_24893);
nand UO_1470 (O_1470,N_24622,N_24057);
or UO_1471 (O_1471,N_24366,N_24975);
and UO_1472 (O_1472,N_24958,N_24834);
xnor UO_1473 (O_1473,N_24277,N_24361);
and UO_1474 (O_1474,N_24161,N_24676);
xnor UO_1475 (O_1475,N_24496,N_24146);
or UO_1476 (O_1476,N_24638,N_24555);
nor UO_1477 (O_1477,N_24662,N_24023);
nor UO_1478 (O_1478,N_24189,N_24678);
and UO_1479 (O_1479,N_24726,N_24199);
nor UO_1480 (O_1480,N_24585,N_24873);
and UO_1481 (O_1481,N_24860,N_24749);
xor UO_1482 (O_1482,N_24052,N_24551);
and UO_1483 (O_1483,N_24754,N_24743);
and UO_1484 (O_1484,N_24587,N_24924);
and UO_1485 (O_1485,N_24700,N_24638);
xor UO_1486 (O_1486,N_24996,N_24104);
xor UO_1487 (O_1487,N_24724,N_24583);
and UO_1488 (O_1488,N_24633,N_24222);
nor UO_1489 (O_1489,N_24084,N_24397);
nor UO_1490 (O_1490,N_24919,N_24056);
or UO_1491 (O_1491,N_24645,N_24315);
nor UO_1492 (O_1492,N_24605,N_24902);
or UO_1493 (O_1493,N_24533,N_24701);
xnor UO_1494 (O_1494,N_24197,N_24532);
or UO_1495 (O_1495,N_24362,N_24781);
nand UO_1496 (O_1496,N_24111,N_24663);
or UO_1497 (O_1497,N_24199,N_24441);
nand UO_1498 (O_1498,N_24588,N_24168);
or UO_1499 (O_1499,N_24004,N_24659);
and UO_1500 (O_1500,N_24433,N_24174);
nand UO_1501 (O_1501,N_24153,N_24457);
and UO_1502 (O_1502,N_24196,N_24147);
or UO_1503 (O_1503,N_24832,N_24339);
and UO_1504 (O_1504,N_24667,N_24960);
or UO_1505 (O_1505,N_24084,N_24292);
nand UO_1506 (O_1506,N_24977,N_24885);
xnor UO_1507 (O_1507,N_24997,N_24688);
xor UO_1508 (O_1508,N_24291,N_24007);
nand UO_1509 (O_1509,N_24320,N_24883);
xor UO_1510 (O_1510,N_24411,N_24578);
and UO_1511 (O_1511,N_24037,N_24222);
or UO_1512 (O_1512,N_24359,N_24569);
or UO_1513 (O_1513,N_24128,N_24954);
or UO_1514 (O_1514,N_24982,N_24582);
nand UO_1515 (O_1515,N_24015,N_24259);
and UO_1516 (O_1516,N_24972,N_24022);
and UO_1517 (O_1517,N_24742,N_24073);
xor UO_1518 (O_1518,N_24751,N_24892);
xnor UO_1519 (O_1519,N_24387,N_24366);
xnor UO_1520 (O_1520,N_24648,N_24891);
xnor UO_1521 (O_1521,N_24501,N_24965);
xor UO_1522 (O_1522,N_24470,N_24468);
nand UO_1523 (O_1523,N_24655,N_24657);
xor UO_1524 (O_1524,N_24743,N_24048);
nor UO_1525 (O_1525,N_24685,N_24541);
nor UO_1526 (O_1526,N_24250,N_24421);
nand UO_1527 (O_1527,N_24205,N_24655);
or UO_1528 (O_1528,N_24191,N_24747);
nand UO_1529 (O_1529,N_24750,N_24554);
or UO_1530 (O_1530,N_24526,N_24805);
and UO_1531 (O_1531,N_24096,N_24972);
xnor UO_1532 (O_1532,N_24273,N_24628);
nor UO_1533 (O_1533,N_24374,N_24979);
nor UO_1534 (O_1534,N_24417,N_24114);
and UO_1535 (O_1535,N_24054,N_24963);
nand UO_1536 (O_1536,N_24348,N_24813);
and UO_1537 (O_1537,N_24072,N_24252);
or UO_1538 (O_1538,N_24136,N_24837);
nor UO_1539 (O_1539,N_24509,N_24866);
or UO_1540 (O_1540,N_24230,N_24107);
nor UO_1541 (O_1541,N_24297,N_24212);
or UO_1542 (O_1542,N_24270,N_24737);
nor UO_1543 (O_1543,N_24783,N_24893);
nor UO_1544 (O_1544,N_24287,N_24472);
nand UO_1545 (O_1545,N_24314,N_24408);
xnor UO_1546 (O_1546,N_24726,N_24817);
and UO_1547 (O_1547,N_24294,N_24993);
or UO_1548 (O_1548,N_24499,N_24502);
nor UO_1549 (O_1549,N_24561,N_24176);
nand UO_1550 (O_1550,N_24584,N_24538);
and UO_1551 (O_1551,N_24071,N_24614);
nand UO_1552 (O_1552,N_24415,N_24674);
and UO_1553 (O_1553,N_24743,N_24147);
xor UO_1554 (O_1554,N_24141,N_24550);
nor UO_1555 (O_1555,N_24244,N_24462);
xor UO_1556 (O_1556,N_24566,N_24913);
nand UO_1557 (O_1557,N_24942,N_24197);
and UO_1558 (O_1558,N_24328,N_24509);
and UO_1559 (O_1559,N_24005,N_24220);
nor UO_1560 (O_1560,N_24383,N_24812);
nand UO_1561 (O_1561,N_24734,N_24327);
or UO_1562 (O_1562,N_24853,N_24680);
or UO_1563 (O_1563,N_24424,N_24795);
or UO_1564 (O_1564,N_24336,N_24696);
and UO_1565 (O_1565,N_24040,N_24232);
or UO_1566 (O_1566,N_24854,N_24273);
xnor UO_1567 (O_1567,N_24665,N_24924);
nand UO_1568 (O_1568,N_24241,N_24921);
nand UO_1569 (O_1569,N_24657,N_24960);
and UO_1570 (O_1570,N_24557,N_24932);
nand UO_1571 (O_1571,N_24149,N_24573);
nand UO_1572 (O_1572,N_24152,N_24846);
and UO_1573 (O_1573,N_24810,N_24008);
xor UO_1574 (O_1574,N_24975,N_24017);
or UO_1575 (O_1575,N_24311,N_24761);
xor UO_1576 (O_1576,N_24994,N_24345);
nand UO_1577 (O_1577,N_24023,N_24281);
nor UO_1578 (O_1578,N_24875,N_24048);
and UO_1579 (O_1579,N_24332,N_24771);
nand UO_1580 (O_1580,N_24251,N_24691);
nor UO_1581 (O_1581,N_24357,N_24362);
nand UO_1582 (O_1582,N_24681,N_24014);
nor UO_1583 (O_1583,N_24281,N_24976);
nor UO_1584 (O_1584,N_24157,N_24660);
xor UO_1585 (O_1585,N_24824,N_24469);
and UO_1586 (O_1586,N_24060,N_24647);
xor UO_1587 (O_1587,N_24710,N_24139);
nor UO_1588 (O_1588,N_24181,N_24180);
nor UO_1589 (O_1589,N_24640,N_24194);
xnor UO_1590 (O_1590,N_24279,N_24670);
nor UO_1591 (O_1591,N_24013,N_24159);
xor UO_1592 (O_1592,N_24410,N_24789);
or UO_1593 (O_1593,N_24560,N_24538);
nor UO_1594 (O_1594,N_24531,N_24715);
and UO_1595 (O_1595,N_24955,N_24790);
and UO_1596 (O_1596,N_24744,N_24955);
xnor UO_1597 (O_1597,N_24192,N_24019);
nor UO_1598 (O_1598,N_24407,N_24130);
nor UO_1599 (O_1599,N_24618,N_24204);
or UO_1600 (O_1600,N_24671,N_24813);
and UO_1601 (O_1601,N_24743,N_24165);
nand UO_1602 (O_1602,N_24448,N_24703);
nand UO_1603 (O_1603,N_24207,N_24668);
xnor UO_1604 (O_1604,N_24287,N_24881);
or UO_1605 (O_1605,N_24190,N_24920);
nand UO_1606 (O_1606,N_24088,N_24713);
or UO_1607 (O_1607,N_24255,N_24348);
nor UO_1608 (O_1608,N_24452,N_24025);
nand UO_1609 (O_1609,N_24982,N_24063);
and UO_1610 (O_1610,N_24894,N_24104);
or UO_1611 (O_1611,N_24863,N_24074);
xnor UO_1612 (O_1612,N_24151,N_24592);
xnor UO_1613 (O_1613,N_24728,N_24606);
and UO_1614 (O_1614,N_24681,N_24913);
nand UO_1615 (O_1615,N_24780,N_24673);
and UO_1616 (O_1616,N_24251,N_24035);
or UO_1617 (O_1617,N_24989,N_24983);
nor UO_1618 (O_1618,N_24014,N_24773);
nor UO_1619 (O_1619,N_24189,N_24593);
nor UO_1620 (O_1620,N_24704,N_24812);
nor UO_1621 (O_1621,N_24565,N_24008);
nand UO_1622 (O_1622,N_24431,N_24173);
nor UO_1623 (O_1623,N_24569,N_24341);
or UO_1624 (O_1624,N_24745,N_24533);
nor UO_1625 (O_1625,N_24520,N_24700);
nor UO_1626 (O_1626,N_24319,N_24722);
nand UO_1627 (O_1627,N_24545,N_24380);
nand UO_1628 (O_1628,N_24626,N_24284);
nand UO_1629 (O_1629,N_24566,N_24725);
and UO_1630 (O_1630,N_24532,N_24187);
xnor UO_1631 (O_1631,N_24245,N_24162);
nand UO_1632 (O_1632,N_24417,N_24707);
nand UO_1633 (O_1633,N_24493,N_24586);
nor UO_1634 (O_1634,N_24763,N_24686);
or UO_1635 (O_1635,N_24172,N_24780);
and UO_1636 (O_1636,N_24702,N_24054);
or UO_1637 (O_1637,N_24501,N_24728);
nor UO_1638 (O_1638,N_24308,N_24087);
xor UO_1639 (O_1639,N_24673,N_24820);
xnor UO_1640 (O_1640,N_24252,N_24904);
nand UO_1641 (O_1641,N_24084,N_24227);
and UO_1642 (O_1642,N_24356,N_24625);
and UO_1643 (O_1643,N_24314,N_24171);
xnor UO_1644 (O_1644,N_24536,N_24724);
nand UO_1645 (O_1645,N_24678,N_24210);
nand UO_1646 (O_1646,N_24624,N_24910);
xnor UO_1647 (O_1647,N_24750,N_24365);
nor UO_1648 (O_1648,N_24971,N_24536);
nand UO_1649 (O_1649,N_24729,N_24877);
or UO_1650 (O_1650,N_24871,N_24832);
or UO_1651 (O_1651,N_24145,N_24073);
and UO_1652 (O_1652,N_24675,N_24801);
xor UO_1653 (O_1653,N_24891,N_24508);
and UO_1654 (O_1654,N_24643,N_24008);
xnor UO_1655 (O_1655,N_24591,N_24380);
or UO_1656 (O_1656,N_24783,N_24289);
or UO_1657 (O_1657,N_24967,N_24525);
nor UO_1658 (O_1658,N_24903,N_24787);
xnor UO_1659 (O_1659,N_24170,N_24277);
and UO_1660 (O_1660,N_24823,N_24220);
nand UO_1661 (O_1661,N_24834,N_24931);
nor UO_1662 (O_1662,N_24689,N_24848);
xnor UO_1663 (O_1663,N_24963,N_24643);
xor UO_1664 (O_1664,N_24913,N_24810);
nor UO_1665 (O_1665,N_24028,N_24220);
or UO_1666 (O_1666,N_24627,N_24334);
nor UO_1667 (O_1667,N_24069,N_24552);
nand UO_1668 (O_1668,N_24906,N_24113);
and UO_1669 (O_1669,N_24423,N_24345);
nand UO_1670 (O_1670,N_24039,N_24040);
nand UO_1671 (O_1671,N_24466,N_24403);
nand UO_1672 (O_1672,N_24875,N_24285);
and UO_1673 (O_1673,N_24280,N_24527);
xnor UO_1674 (O_1674,N_24015,N_24145);
and UO_1675 (O_1675,N_24407,N_24084);
or UO_1676 (O_1676,N_24625,N_24503);
or UO_1677 (O_1677,N_24105,N_24085);
nor UO_1678 (O_1678,N_24802,N_24154);
xor UO_1679 (O_1679,N_24931,N_24139);
xnor UO_1680 (O_1680,N_24543,N_24188);
or UO_1681 (O_1681,N_24562,N_24959);
nor UO_1682 (O_1682,N_24080,N_24372);
xnor UO_1683 (O_1683,N_24779,N_24094);
or UO_1684 (O_1684,N_24061,N_24390);
nand UO_1685 (O_1685,N_24573,N_24235);
xor UO_1686 (O_1686,N_24750,N_24293);
or UO_1687 (O_1687,N_24034,N_24168);
nand UO_1688 (O_1688,N_24553,N_24732);
xnor UO_1689 (O_1689,N_24740,N_24940);
nor UO_1690 (O_1690,N_24430,N_24606);
and UO_1691 (O_1691,N_24214,N_24054);
and UO_1692 (O_1692,N_24780,N_24217);
and UO_1693 (O_1693,N_24955,N_24926);
and UO_1694 (O_1694,N_24748,N_24485);
nor UO_1695 (O_1695,N_24368,N_24002);
and UO_1696 (O_1696,N_24650,N_24364);
nand UO_1697 (O_1697,N_24840,N_24993);
nor UO_1698 (O_1698,N_24696,N_24574);
xnor UO_1699 (O_1699,N_24279,N_24128);
nand UO_1700 (O_1700,N_24325,N_24707);
nand UO_1701 (O_1701,N_24017,N_24912);
nand UO_1702 (O_1702,N_24537,N_24419);
or UO_1703 (O_1703,N_24157,N_24255);
or UO_1704 (O_1704,N_24302,N_24634);
xor UO_1705 (O_1705,N_24855,N_24598);
xnor UO_1706 (O_1706,N_24466,N_24994);
nand UO_1707 (O_1707,N_24997,N_24274);
nand UO_1708 (O_1708,N_24197,N_24466);
or UO_1709 (O_1709,N_24740,N_24000);
nor UO_1710 (O_1710,N_24795,N_24326);
xor UO_1711 (O_1711,N_24241,N_24392);
xor UO_1712 (O_1712,N_24942,N_24423);
nor UO_1713 (O_1713,N_24815,N_24549);
nor UO_1714 (O_1714,N_24274,N_24509);
and UO_1715 (O_1715,N_24462,N_24184);
and UO_1716 (O_1716,N_24508,N_24351);
nand UO_1717 (O_1717,N_24876,N_24814);
or UO_1718 (O_1718,N_24017,N_24388);
nand UO_1719 (O_1719,N_24712,N_24156);
xor UO_1720 (O_1720,N_24735,N_24063);
nor UO_1721 (O_1721,N_24144,N_24932);
nor UO_1722 (O_1722,N_24908,N_24233);
xor UO_1723 (O_1723,N_24674,N_24828);
or UO_1724 (O_1724,N_24945,N_24937);
or UO_1725 (O_1725,N_24475,N_24252);
and UO_1726 (O_1726,N_24472,N_24579);
nor UO_1727 (O_1727,N_24456,N_24277);
nor UO_1728 (O_1728,N_24739,N_24480);
nor UO_1729 (O_1729,N_24203,N_24716);
nor UO_1730 (O_1730,N_24454,N_24848);
xnor UO_1731 (O_1731,N_24657,N_24656);
and UO_1732 (O_1732,N_24358,N_24605);
nor UO_1733 (O_1733,N_24833,N_24524);
xor UO_1734 (O_1734,N_24494,N_24741);
nand UO_1735 (O_1735,N_24745,N_24930);
nor UO_1736 (O_1736,N_24943,N_24169);
or UO_1737 (O_1737,N_24351,N_24072);
nor UO_1738 (O_1738,N_24497,N_24640);
nand UO_1739 (O_1739,N_24540,N_24970);
or UO_1740 (O_1740,N_24923,N_24726);
or UO_1741 (O_1741,N_24183,N_24318);
nand UO_1742 (O_1742,N_24692,N_24085);
nand UO_1743 (O_1743,N_24906,N_24623);
nor UO_1744 (O_1744,N_24338,N_24742);
nor UO_1745 (O_1745,N_24921,N_24101);
and UO_1746 (O_1746,N_24111,N_24424);
and UO_1747 (O_1747,N_24080,N_24352);
nor UO_1748 (O_1748,N_24511,N_24219);
or UO_1749 (O_1749,N_24950,N_24023);
and UO_1750 (O_1750,N_24289,N_24920);
and UO_1751 (O_1751,N_24814,N_24808);
xnor UO_1752 (O_1752,N_24326,N_24891);
and UO_1753 (O_1753,N_24390,N_24440);
or UO_1754 (O_1754,N_24520,N_24047);
nor UO_1755 (O_1755,N_24419,N_24767);
nor UO_1756 (O_1756,N_24195,N_24215);
and UO_1757 (O_1757,N_24474,N_24553);
nand UO_1758 (O_1758,N_24812,N_24178);
and UO_1759 (O_1759,N_24023,N_24306);
xnor UO_1760 (O_1760,N_24902,N_24614);
nand UO_1761 (O_1761,N_24994,N_24082);
nand UO_1762 (O_1762,N_24968,N_24694);
or UO_1763 (O_1763,N_24512,N_24132);
nor UO_1764 (O_1764,N_24204,N_24461);
nand UO_1765 (O_1765,N_24149,N_24758);
xor UO_1766 (O_1766,N_24358,N_24355);
nand UO_1767 (O_1767,N_24459,N_24730);
xnor UO_1768 (O_1768,N_24780,N_24945);
nand UO_1769 (O_1769,N_24051,N_24373);
nor UO_1770 (O_1770,N_24390,N_24362);
nor UO_1771 (O_1771,N_24692,N_24296);
nand UO_1772 (O_1772,N_24569,N_24587);
nand UO_1773 (O_1773,N_24995,N_24073);
xor UO_1774 (O_1774,N_24678,N_24859);
xor UO_1775 (O_1775,N_24755,N_24864);
and UO_1776 (O_1776,N_24337,N_24425);
nor UO_1777 (O_1777,N_24507,N_24804);
xnor UO_1778 (O_1778,N_24257,N_24134);
or UO_1779 (O_1779,N_24710,N_24407);
nand UO_1780 (O_1780,N_24363,N_24507);
and UO_1781 (O_1781,N_24928,N_24434);
nor UO_1782 (O_1782,N_24851,N_24977);
xor UO_1783 (O_1783,N_24409,N_24906);
nand UO_1784 (O_1784,N_24458,N_24264);
and UO_1785 (O_1785,N_24605,N_24154);
or UO_1786 (O_1786,N_24370,N_24031);
and UO_1787 (O_1787,N_24507,N_24819);
nand UO_1788 (O_1788,N_24351,N_24303);
nor UO_1789 (O_1789,N_24293,N_24916);
nor UO_1790 (O_1790,N_24768,N_24748);
and UO_1791 (O_1791,N_24045,N_24351);
nand UO_1792 (O_1792,N_24474,N_24482);
and UO_1793 (O_1793,N_24484,N_24936);
and UO_1794 (O_1794,N_24025,N_24865);
nand UO_1795 (O_1795,N_24912,N_24582);
and UO_1796 (O_1796,N_24687,N_24164);
nor UO_1797 (O_1797,N_24795,N_24891);
xnor UO_1798 (O_1798,N_24396,N_24558);
nand UO_1799 (O_1799,N_24881,N_24716);
and UO_1800 (O_1800,N_24910,N_24996);
nand UO_1801 (O_1801,N_24676,N_24477);
nand UO_1802 (O_1802,N_24977,N_24353);
xor UO_1803 (O_1803,N_24715,N_24142);
and UO_1804 (O_1804,N_24168,N_24340);
and UO_1805 (O_1805,N_24796,N_24787);
or UO_1806 (O_1806,N_24214,N_24850);
nand UO_1807 (O_1807,N_24519,N_24060);
or UO_1808 (O_1808,N_24314,N_24178);
and UO_1809 (O_1809,N_24018,N_24633);
nor UO_1810 (O_1810,N_24662,N_24490);
or UO_1811 (O_1811,N_24652,N_24206);
xnor UO_1812 (O_1812,N_24519,N_24036);
nor UO_1813 (O_1813,N_24448,N_24900);
or UO_1814 (O_1814,N_24723,N_24570);
or UO_1815 (O_1815,N_24543,N_24923);
nor UO_1816 (O_1816,N_24540,N_24164);
nand UO_1817 (O_1817,N_24824,N_24026);
nor UO_1818 (O_1818,N_24490,N_24829);
nor UO_1819 (O_1819,N_24581,N_24512);
nor UO_1820 (O_1820,N_24585,N_24981);
nor UO_1821 (O_1821,N_24757,N_24815);
and UO_1822 (O_1822,N_24188,N_24482);
nand UO_1823 (O_1823,N_24161,N_24125);
or UO_1824 (O_1824,N_24058,N_24103);
xnor UO_1825 (O_1825,N_24505,N_24168);
or UO_1826 (O_1826,N_24546,N_24339);
nor UO_1827 (O_1827,N_24836,N_24246);
or UO_1828 (O_1828,N_24925,N_24457);
xor UO_1829 (O_1829,N_24611,N_24954);
nand UO_1830 (O_1830,N_24283,N_24527);
nor UO_1831 (O_1831,N_24524,N_24083);
nand UO_1832 (O_1832,N_24089,N_24176);
nor UO_1833 (O_1833,N_24637,N_24519);
nor UO_1834 (O_1834,N_24731,N_24750);
xnor UO_1835 (O_1835,N_24078,N_24820);
or UO_1836 (O_1836,N_24349,N_24827);
nor UO_1837 (O_1837,N_24734,N_24436);
nor UO_1838 (O_1838,N_24631,N_24151);
nor UO_1839 (O_1839,N_24462,N_24772);
or UO_1840 (O_1840,N_24533,N_24381);
nand UO_1841 (O_1841,N_24858,N_24253);
or UO_1842 (O_1842,N_24210,N_24902);
nand UO_1843 (O_1843,N_24756,N_24639);
nor UO_1844 (O_1844,N_24529,N_24188);
xnor UO_1845 (O_1845,N_24130,N_24383);
or UO_1846 (O_1846,N_24202,N_24364);
or UO_1847 (O_1847,N_24011,N_24291);
nand UO_1848 (O_1848,N_24355,N_24523);
nand UO_1849 (O_1849,N_24856,N_24283);
nor UO_1850 (O_1850,N_24972,N_24397);
and UO_1851 (O_1851,N_24791,N_24197);
nor UO_1852 (O_1852,N_24914,N_24133);
nor UO_1853 (O_1853,N_24986,N_24991);
nor UO_1854 (O_1854,N_24299,N_24696);
nor UO_1855 (O_1855,N_24888,N_24005);
and UO_1856 (O_1856,N_24254,N_24955);
xor UO_1857 (O_1857,N_24557,N_24034);
nor UO_1858 (O_1858,N_24005,N_24798);
and UO_1859 (O_1859,N_24716,N_24174);
or UO_1860 (O_1860,N_24343,N_24080);
or UO_1861 (O_1861,N_24000,N_24033);
and UO_1862 (O_1862,N_24526,N_24032);
or UO_1863 (O_1863,N_24940,N_24437);
xnor UO_1864 (O_1864,N_24604,N_24457);
and UO_1865 (O_1865,N_24929,N_24861);
or UO_1866 (O_1866,N_24987,N_24044);
nor UO_1867 (O_1867,N_24443,N_24174);
and UO_1868 (O_1868,N_24743,N_24266);
xor UO_1869 (O_1869,N_24202,N_24557);
nor UO_1870 (O_1870,N_24593,N_24376);
xor UO_1871 (O_1871,N_24967,N_24364);
or UO_1872 (O_1872,N_24616,N_24825);
and UO_1873 (O_1873,N_24182,N_24046);
or UO_1874 (O_1874,N_24347,N_24979);
xnor UO_1875 (O_1875,N_24932,N_24136);
and UO_1876 (O_1876,N_24439,N_24679);
nand UO_1877 (O_1877,N_24853,N_24388);
nor UO_1878 (O_1878,N_24248,N_24876);
or UO_1879 (O_1879,N_24220,N_24889);
xor UO_1880 (O_1880,N_24341,N_24632);
nor UO_1881 (O_1881,N_24541,N_24816);
xnor UO_1882 (O_1882,N_24251,N_24361);
nand UO_1883 (O_1883,N_24084,N_24480);
nor UO_1884 (O_1884,N_24817,N_24129);
and UO_1885 (O_1885,N_24287,N_24534);
nand UO_1886 (O_1886,N_24456,N_24139);
xnor UO_1887 (O_1887,N_24325,N_24344);
xnor UO_1888 (O_1888,N_24827,N_24390);
and UO_1889 (O_1889,N_24402,N_24658);
or UO_1890 (O_1890,N_24383,N_24685);
nor UO_1891 (O_1891,N_24008,N_24879);
nand UO_1892 (O_1892,N_24416,N_24662);
xnor UO_1893 (O_1893,N_24668,N_24596);
nand UO_1894 (O_1894,N_24743,N_24357);
and UO_1895 (O_1895,N_24782,N_24254);
and UO_1896 (O_1896,N_24752,N_24810);
nor UO_1897 (O_1897,N_24172,N_24669);
or UO_1898 (O_1898,N_24112,N_24446);
nand UO_1899 (O_1899,N_24731,N_24259);
nand UO_1900 (O_1900,N_24290,N_24176);
nor UO_1901 (O_1901,N_24824,N_24718);
nor UO_1902 (O_1902,N_24200,N_24691);
nand UO_1903 (O_1903,N_24986,N_24617);
xnor UO_1904 (O_1904,N_24566,N_24721);
and UO_1905 (O_1905,N_24957,N_24376);
or UO_1906 (O_1906,N_24202,N_24733);
or UO_1907 (O_1907,N_24438,N_24661);
or UO_1908 (O_1908,N_24308,N_24595);
nor UO_1909 (O_1909,N_24097,N_24144);
nand UO_1910 (O_1910,N_24425,N_24398);
nand UO_1911 (O_1911,N_24920,N_24156);
nand UO_1912 (O_1912,N_24069,N_24047);
nand UO_1913 (O_1913,N_24318,N_24287);
nor UO_1914 (O_1914,N_24884,N_24379);
nand UO_1915 (O_1915,N_24096,N_24624);
or UO_1916 (O_1916,N_24010,N_24705);
xor UO_1917 (O_1917,N_24725,N_24412);
xnor UO_1918 (O_1918,N_24783,N_24380);
nand UO_1919 (O_1919,N_24115,N_24218);
xor UO_1920 (O_1920,N_24129,N_24779);
and UO_1921 (O_1921,N_24805,N_24284);
and UO_1922 (O_1922,N_24468,N_24376);
and UO_1923 (O_1923,N_24130,N_24555);
or UO_1924 (O_1924,N_24017,N_24802);
and UO_1925 (O_1925,N_24328,N_24166);
and UO_1926 (O_1926,N_24472,N_24686);
or UO_1927 (O_1927,N_24036,N_24385);
xnor UO_1928 (O_1928,N_24126,N_24059);
or UO_1929 (O_1929,N_24920,N_24484);
nand UO_1930 (O_1930,N_24955,N_24302);
and UO_1931 (O_1931,N_24072,N_24190);
or UO_1932 (O_1932,N_24996,N_24791);
nor UO_1933 (O_1933,N_24706,N_24867);
or UO_1934 (O_1934,N_24897,N_24583);
xnor UO_1935 (O_1935,N_24235,N_24695);
xnor UO_1936 (O_1936,N_24828,N_24410);
nand UO_1937 (O_1937,N_24786,N_24571);
nor UO_1938 (O_1938,N_24418,N_24800);
nand UO_1939 (O_1939,N_24220,N_24476);
nand UO_1940 (O_1940,N_24394,N_24799);
xnor UO_1941 (O_1941,N_24128,N_24982);
xor UO_1942 (O_1942,N_24287,N_24139);
nor UO_1943 (O_1943,N_24432,N_24527);
xor UO_1944 (O_1944,N_24292,N_24766);
nor UO_1945 (O_1945,N_24718,N_24114);
nor UO_1946 (O_1946,N_24705,N_24616);
and UO_1947 (O_1947,N_24611,N_24041);
nor UO_1948 (O_1948,N_24580,N_24568);
xnor UO_1949 (O_1949,N_24472,N_24283);
or UO_1950 (O_1950,N_24598,N_24620);
nand UO_1951 (O_1951,N_24097,N_24826);
and UO_1952 (O_1952,N_24441,N_24282);
nand UO_1953 (O_1953,N_24522,N_24866);
and UO_1954 (O_1954,N_24647,N_24239);
nor UO_1955 (O_1955,N_24827,N_24417);
and UO_1956 (O_1956,N_24529,N_24031);
or UO_1957 (O_1957,N_24246,N_24717);
or UO_1958 (O_1958,N_24812,N_24321);
nand UO_1959 (O_1959,N_24178,N_24821);
xnor UO_1960 (O_1960,N_24419,N_24106);
and UO_1961 (O_1961,N_24419,N_24975);
xnor UO_1962 (O_1962,N_24844,N_24853);
nor UO_1963 (O_1963,N_24890,N_24056);
or UO_1964 (O_1964,N_24356,N_24359);
nor UO_1965 (O_1965,N_24352,N_24814);
nor UO_1966 (O_1966,N_24713,N_24114);
nand UO_1967 (O_1967,N_24958,N_24693);
xnor UO_1968 (O_1968,N_24358,N_24286);
or UO_1969 (O_1969,N_24937,N_24395);
and UO_1970 (O_1970,N_24004,N_24471);
and UO_1971 (O_1971,N_24202,N_24605);
nor UO_1972 (O_1972,N_24246,N_24137);
or UO_1973 (O_1973,N_24369,N_24263);
or UO_1974 (O_1974,N_24416,N_24264);
and UO_1975 (O_1975,N_24962,N_24239);
and UO_1976 (O_1976,N_24886,N_24611);
and UO_1977 (O_1977,N_24149,N_24985);
xnor UO_1978 (O_1978,N_24050,N_24425);
nand UO_1979 (O_1979,N_24653,N_24282);
nor UO_1980 (O_1980,N_24894,N_24776);
nor UO_1981 (O_1981,N_24164,N_24318);
nand UO_1982 (O_1982,N_24404,N_24203);
and UO_1983 (O_1983,N_24301,N_24982);
nand UO_1984 (O_1984,N_24184,N_24032);
nand UO_1985 (O_1985,N_24101,N_24478);
and UO_1986 (O_1986,N_24569,N_24147);
nor UO_1987 (O_1987,N_24764,N_24439);
and UO_1988 (O_1988,N_24899,N_24634);
nand UO_1989 (O_1989,N_24805,N_24214);
nand UO_1990 (O_1990,N_24667,N_24385);
or UO_1991 (O_1991,N_24193,N_24944);
and UO_1992 (O_1992,N_24330,N_24533);
xor UO_1993 (O_1993,N_24715,N_24726);
nor UO_1994 (O_1994,N_24933,N_24333);
and UO_1995 (O_1995,N_24959,N_24724);
or UO_1996 (O_1996,N_24683,N_24416);
xnor UO_1997 (O_1997,N_24578,N_24458);
xor UO_1998 (O_1998,N_24227,N_24508);
xnor UO_1999 (O_1999,N_24050,N_24150);
or UO_2000 (O_2000,N_24324,N_24483);
and UO_2001 (O_2001,N_24581,N_24081);
and UO_2002 (O_2002,N_24117,N_24551);
xnor UO_2003 (O_2003,N_24280,N_24719);
nor UO_2004 (O_2004,N_24878,N_24770);
nor UO_2005 (O_2005,N_24918,N_24441);
xor UO_2006 (O_2006,N_24993,N_24186);
xnor UO_2007 (O_2007,N_24218,N_24926);
nor UO_2008 (O_2008,N_24170,N_24503);
nor UO_2009 (O_2009,N_24670,N_24828);
nand UO_2010 (O_2010,N_24596,N_24789);
or UO_2011 (O_2011,N_24989,N_24005);
nand UO_2012 (O_2012,N_24511,N_24214);
xor UO_2013 (O_2013,N_24118,N_24746);
xnor UO_2014 (O_2014,N_24846,N_24535);
nor UO_2015 (O_2015,N_24721,N_24405);
xnor UO_2016 (O_2016,N_24524,N_24821);
nor UO_2017 (O_2017,N_24188,N_24412);
nand UO_2018 (O_2018,N_24794,N_24231);
and UO_2019 (O_2019,N_24718,N_24308);
and UO_2020 (O_2020,N_24983,N_24573);
nor UO_2021 (O_2021,N_24889,N_24112);
and UO_2022 (O_2022,N_24727,N_24384);
xor UO_2023 (O_2023,N_24166,N_24421);
nor UO_2024 (O_2024,N_24572,N_24823);
or UO_2025 (O_2025,N_24665,N_24648);
xnor UO_2026 (O_2026,N_24900,N_24007);
xnor UO_2027 (O_2027,N_24564,N_24505);
nand UO_2028 (O_2028,N_24530,N_24074);
nand UO_2029 (O_2029,N_24335,N_24838);
xnor UO_2030 (O_2030,N_24048,N_24312);
nor UO_2031 (O_2031,N_24801,N_24625);
and UO_2032 (O_2032,N_24599,N_24300);
nand UO_2033 (O_2033,N_24675,N_24479);
nor UO_2034 (O_2034,N_24629,N_24079);
and UO_2035 (O_2035,N_24093,N_24171);
or UO_2036 (O_2036,N_24900,N_24979);
nor UO_2037 (O_2037,N_24285,N_24909);
nor UO_2038 (O_2038,N_24157,N_24514);
nand UO_2039 (O_2039,N_24502,N_24799);
xnor UO_2040 (O_2040,N_24688,N_24042);
nand UO_2041 (O_2041,N_24653,N_24828);
and UO_2042 (O_2042,N_24326,N_24320);
xnor UO_2043 (O_2043,N_24379,N_24080);
or UO_2044 (O_2044,N_24232,N_24096);
and UO_2045 (O_2045,N_24586,N_24050);
xor UO_2046 (O_2046,N_24051,N_24594);
nand UO_2047 (O_2047,N_24710,N_24982);
nand UO_2048 (O_2048,N_24637,N_24423);
xor UO_2049 (O_2049,N_24271,N_24671);
xor UO_2050 (O_2050,N_24449,N_24173);
nor UO_2051 (O_2051,N_24268,N_24471);
and UO_2052 (O_2052,N_24136,N_24390);
xnor UO_2053 (O_2053,N_24486,N_24403);
nor UO_2054 (O_2054,N_24949,N_24805);
nand UO_2055 (O_2055,N_24824,N_24939);
nand UO_2056 (O_2056,N_24753,N_24407);
or UO_2057 (O_2057,N_24086,N_24781);
xnor UO_2058 (O_2058,N_24232,N_24015);
and UO_2059 (O_2059,N_24054,N_24020);
and UO_2060 (O_2060,N_24933,N_24569);
and UO_2061 (O_2061,N_24541,N_24095);
xor UO_2062 (O_2062,N_24461,N_24208);
or UO_2063 (O_2063,N_24558,N_24487);
nor UO_2064 (O_2064,N_24265,N_24272);
xnor UO_2065 (O_2065,N_24440,N_24623);
nand UO_2066 (O_2066,N_24035,N_24263);
and UO_2067 (O_2067,N_24778,N_24234);
and UO_2068 (O_2068,N_24924,N_24460);
and UO_2069 (O_2069,N_24403,N_24722);
or UO_2070 (O_2070,N_24498,N_24593);
nand UO_2071 (O_2071,N_24023,N_24787);
or UO_2072 (O_2072,N_24726,N_24617);
xnor UO_2073 (O_2073,N_24633,N_24841);
xnor UO_2074 (O_2074,N_24501,N_24969);
and UO_2075 (O_2075,N_24723,N_24149);
and UO_2076 (O_2076,N_24069,N_24300);
or UO_2077 (O_2077,N_24512,N_24166);
nand UO_2078 (O_2078,N_24347,N_24580);
nand UO_2079 (O_2079,N_24414,N_24523);
nor UO_2080 (O_2080,N_24522,N_24225);
nor UO_2081 (O_2081,N_24907,N_24377);
and UO_2082 (O_2082,N_24537,N_24446);
nand UO_2083 (O_2083,N_24552,N_24520);
nor UO_2084 (O_2084,N_24483,N_24808);
and UO_2085 (O_2085,N_24734,N_24075);
nand UO_2086 (O_2086,N_24337,N_24379);
nor UO_2087 (O_2087,N_24189,N_24008);
and UO_2088 (O_2088,N_24876,N_24667);
nor UO_2089 (O_2089,N_24410,N_24728);
nand UO_2090 (O_2090,N_24403,N_24111);
xnor UO_2091 (O_2091,N_24355,N_24841);
or UO_2092 (O_2092,N_24256,N_24987);
and UO_2093 (O_2093,N_24323,N_24241);
xnor UO_2094 (O_2094,N_24262,N_24298);
nand UO_2095 (O_2095,N_24722,N_24549);
nor UO_2096 (O_2096,N_24165,N_24493);
nand UO_2097 (O_2097,N_24328,N_24475);
and UO_2098 (O_2098,N_24923,N_24365);
nor UO_2099 (O_2099,N_24401,N_24808);
nand UO_2100 (O_2100,N_24775,N_24215);
and UO_2101 (O_2101,N_24666,N_24192);
nand UO_2102 (O_2102,N_24388,N_24538);
nor UO_2103 (O_2103,N_24596,N_24621);
nor UO_2104 (O_2104,N_24386,N_24580);
and UO_2105 (O_2105,N_24681,N_24634);
and UO_2106 (O_2106,N_24515,N_24505);
nand UO_2107 (O_2107,N_24875,N_24925);
and UO_2108 (O_2108,N_24882,N_24232);
and UO_2109 (O_2109,N_24286,N_24295);
and UO_2110 (O_2110,N_24267,N_24632);
nand UO_2111 (O_2111,N_24881,N_24321);
nor UO_2112 (O_2112,N_24023,N_24985);
or UO_2113 (O_2113,N_24610,N_24916);
xor UO_2114 (O_2114,N_24598,N_24060);
nor UO_2115 (O_2115,N_24406,N_24064);
and UO_2116 (O_2116,N_24886,N_24516);
nand UO_2117 (O_2117,N_24874,N_24042);
xor UO_2118 (O_2118,N_24927,N_24475);
or UO_2119 (O_2119,N_24916,N_24711);
nor UO_2120 (O_2120,N_24158,N_24878);
nor UO_2121 (O_2121,N_24241,N_24595);
nor UO_2122 (O_2122,N_24989,N_24948);
or UO_2123 (O_2123,N_24971,N_24980);
nor UO_2124 (O_2124,N_24616,N_24384);
and UO_2125 (O_2125,N_24310,N_24822);
xnor UO_2126 (O_2126,N_24862,N_24057);
nand UO_2127 (O_2127,N_24021,N_24919);
nand UO_2128 (O_2128,N_24109,N_24902);
nor UO_2129 (O_2129,N_24903,N_24930);
or UO_2130 (O_2130,N_24973,N_24935);
and UO_2131 (O_2131,N_24465,N_24561);
xor UO_2132 (O_2132,N_24405,N_24253);
xnor UO_2133 (O_2133,N_24042,N_24801);
or UO_2134 (O_2134,N_24975,N_24066);
nand UO_2135 (O_2135,N_24819,N_24624);
nor UO_2136 (O_2136,N_24658,N_24837);
nand UO_2137 (O_2137,N_24406,N_24704);
xnor UO_2138 (O_2138,N_24281,N_24382);
nor UO_2139 (O_2139,N_24654,N_24126);
nand UO_2140 (O_2140,N_24575,N_24235);
xor UO_2141 (O_2141,N_24812,N_24240);
and UO_2142 (O_2142,N_24012,N_24579);
nor UO_2143 (O_2143,N_24508,N_24320);
and UO_2144 (O_2144,N_24303,N_24638);
or UO_2145 (O_2145,N_24061,N_24827);
or UO_2146 (O_2146,N_24277,N_24919);
nor UO_2147 (O_2147,N_24080,N_24924);
nand UO_2148 (O_2148,N_24520,N_24609);
nor UO_2149 (O_2149,N_24763,N_24373);
nand UO_2150 (O_2150,N_24954,N_24894);
and UO_2151 (O_2151,N_24916,N_24206);
and UO_2152 (O_2152,N_24948,N_24357);
and UO_2153 (O_2153,N_24856,N_24402);
xor UO_2154 (O_2154,N_24593,N_24183);
or UO_2155 (O_2155,N_24666,N_24862);
xor UO_2156 (O_2156,N_24196,N_24256);
xnor UO_2157 (O_2157,N_24486,N_24917);
xnor UO_2158 (O_2158,N_24035,N_24192);
and UO_2159 (O_2159,N_24251,N_24842);
nor UO_2160 (O_2160,N_24735,N_24138);
nand UO_2161 (O_2161,N_24357,N_24111);
and UO_2162 (O_2162,N_24864,N_24365);
or UO_2163 (O_2163,N_24830,N_24866);
and UO_2164 (O_2164,N_24517,N_24625);
or UO_2165 (O_2165,N_24097,N_24391);
nand UO_2166 (O_2166,N_24763,N_24690);
nand UO_2167 (O_2167,N_24458,N_24752);
and UO_2168 (O_2168,N_24619,N_24931);
nand UO_2169 (O_2169,N_24278,N_24835);
nor UO_2170 (O_2170,N_24804,N_24644);
and UO_2171 (O_2171,N_24307,N_24078);
nand UO_2172 (O_2172,N_24032,N_24683);
nand UO_2173 (O_2173,N_24950,N_24746);
nor UO_2174 (O_2174,N_24339,N_24531);
nor UO_2175 (O_2175,N_24134,N_24872);
and UO_2176 (O_2176,N_24376,N_24859);
nor UO_2177 (O_2177,N_24024,N_24644);
or UO_2178 (O_2178,N_24923,N_24476);
nand UO_2179 (O_2179,N_24633,N_24183);
nand UO_2180 (O_2180,N_24161,N_24841);
and UO_2181 (O_2181,N_24759,N_24432);
nand UO_2182 (O_2182,N_24304,N_24231);
or UO_2183 (O_2183,N_24077,N_24227);
and UO_2184 (O_2184,N_24444,N_24955);
nor UO_2185 (O_2185,N_24435,N_24537);
nand UO_2186 (O_2186,N_24602,N_24713);
xor UO_2187 (O_2187,N_24718,N_24699);
nor UO_2188 (O_2188,N_24152,N_24243);
xor UO_2189 (O_2189,N_24393,N_24408);
or UO_2190 (O_2190,N_24185,N_24291);
nor UO_2191 (O_2191,N_24435,N_24719);
nor UO_2192 (O_2192,N_24913,N_24509);
nand UO_2193 (O_2193,N_24047,N_24134);
xor UO_2194 (O_2194,N_24055,N_24069);
nor UO_2195 (O_2195,N_24298,N_24005);
xnor UO_2196 (O_2196,N_24928,N_24250);
or UO_2197 (O_2197,N_24264,N_24188);
and UO_2198 (O_2198,N_24086,N_24620);
nor UO_2199 (O_2199,N_24511,N_24320);
or UO_2200 (O_2200,N_24800,N_24100);
nand UO_2201 (O_2201,N_24987,N_24861);
or UO_2202 (O_2202,N_24604,N_24549);
and UO_2203 (O_2203,N_24487,N_24613);
or UO_2204 (O_2204,N_24118,N_24014);
nand UO_2205 (O_2205,N_24742,N_24911);
or UO_2206 (O_2206,N_24333,N_24770);
nor UO_2207 (O_2207,N_24991,N_24854);
xnor UO_2208 (O_2208,N_24458,N_24842);
nor UO_2209 (O_2209,N_24202,N_24668);
nand UO_2210 (O_2210,N_24147,N_24895);
nand UO_2211 (O_2211,N_24301,N_24669);
nor UO_2212 (O_2212,N_24459,N_24167);
or UO_2213 (O_2213,N_24423,N_24994);
xnor UO_2214 (O_2214,N_24979,N_24852);
nor UO_2215 (O_2215,N_24349,N_24574);
nand UO_2216 (O_2216,N_24965,N_24987);
nand UO_2217 (O_2217,N_24405,N_24584);
xnor UO_2218 (O_2218,N_24039,N_24401);
and UO_2219 (O_2219,N_24218,N_24112);
or UO_2220 (O_2220,N_24138,N_24839);
nor UO_2221 (O_2221,N_24870,N_24189);
and UO_2222 (O_2222,N_24307,N_24606);
or UO_2223 (O_2223,N_24787,N_24220);
and UO_2224 (O_2224,N_24848,N_24326);
and UO_2225 (O_2225,N_24723,N_24502);
or UO_2226 (O_2226,N_24328,N_24120);
and UO_2227 (O_2227,N_24476,N_24305);
xor UO_2228 (O_2228,N_24991,N_24504);
nand UO_2229 (O_2229,N_24573,N_24671);
xor UO_2230 (O_2230,N_24775,N_24233);
and UO_2231 (O_2231,N_24407,N_24261);
xor UO_2232 (O_2232,N_24583,N_24911);
nand UO_2233 (O_2233,N_24851,N_24424);
xnor UO_2234 (O_2234,N_24285,N_24753);
nor UO_2235 (O_2235,N_24802,N_24152);
or UO_2236 (O_2236,N_24568,N_24015);
nand UO_2237 (O_2237,N_24266,N_24251);
nand UO_2238 (O_2238,N_24568,N_24275);
xor UO_2239 (O_2239,N_24862,N_24446);
nand UO_2240 (O_2240,N_24705,N_24524);
nor UO_2241 (O_2241,N_24316,N_24998);
or UO_2242 (O_2242,N_24936,N_24824);
nor UO_2243 (O_2243,N_24069,N_24168);
nor UO_2244 (O_2244,N_24302,N_24933);
or UO_2245 (O_2245,N_24952,N_24879);
nand UO_2246 (O_2246,N_24837,N_24132);
nand UO_2247 (O_2247,N_24065,N_24814);
nand UO_2248 (O_2248,N_24412,N_24043);
nor UO_2249 (O_2249,N_24805,N_24224);
nand UO_2250 (O_2250,N_24787,N_24901);
or UO_2251 (O_2251,N_24910,N_24651);
nor UO_2252 (O_2252,N_24467,N_24456);
and UO_2253 (O_2253,N_24050,N_24095);
nor UO_2254 (O_2254,N_24816,N_24473);
or UO_2255 (O_2255,N_24040,N_24575);
and UO_2256 (O_2256,N_24533,N_24504);
nand UO_2257 (O_2257,N_24122,N_24683);
xor UO_2258 (O_2258,N_24468,N_24418);
and UO_2259 (O_2259,N_24915,N_24646);
and UO_2260 (O_2260,N_24954,N_24866);
and UO_2261 (O_2261,N_24391,N_24867);
xor UO_2262 (O_2262,N_24703,N_24820);
nor UO_2263 (O_2263,N_24224,N_24225);
xor UO_2264 (O_2264,N_24960,N_24546);
nand UO_2265 (O_2265,N_24887,N_24132);
xnor UO_2266 (O_2266,N_24388,N_24929);
or UO_2267 (O_2267,N_24262,N_24765);
or UO_2268 (O_2268,N_24456,N_24288);
xnor UO_2269 (O_2269,N_24492,N_24481);
or UO_2270 (O_2270,N_24395,N_24823);
and UO_2271 (O_2271,N_24260,N_24490);
nand UO_2272 (O_2272,N_24449,N_24385);
xor UO_2273 (O_2273,N_24665,N_24804);
nor UO_2274 (O_2274,N_24057,N_24961);
nor UO_2275 (O_2275,N_24323,N_24136);
or UO_2276 (O_2276,N_24875,N_24176);
nor UO_2277 (O_2277,N_24168,N_24810);
and UO_2278 (O_2278,N_24799,N_24191);
nand UO_2279 (O_2279,N_24134,N_24516);
or UO_2280 (O_2280,N_24807,N_24682);
and UO_2281 (O_2281,N_24673,N_24020);
and UO_2282 (O_2282,N_24608,N_24703);
and UO_2283 (O_2283,N_24174,N_24350);
or UO_2284 (O_2284,N_24980,N_24754);
nor UO_2285 (O_2285,N_24960,N_24922);
nor UO_2286 (O_2286,N_24610,N_24249);
or UO_2287 (O_2287,N_24190,N_24630);
xnor UO_2288 (O_2288,N_24908,N_24573);
or UO_2289 (O_2289,N_24417,N_24684);
or UO_2290 (O_2290,N_24493,N_24971);
xor UO_2291 (O_2291,N_24563,N_24559);
or UO_2292 (O_2292,N_24020,N_24080);
and UO_2293 (O_2293,N_24260,N_24233);
xnor UO_2294 (O_2294,N_24198,N_24463);
xor UO_2295 (O_2295,N_24295,N_24819);
and UO_2296 (O_2296,N_24571,N_24860);
or UO_2297 (O_2297,N_24333,N_24149);
and UO_2298 (O_2298,N_24815,N_24112);
xor UO_2299 (O_2299,N_24312,N_24862);
nand UO_2300 (O_2300,N_24784,N_24301);
nand UO_2301 (O_2301,N_24984,N_24444);
or UO_2302 (O_2302,N_24410,N_24618);
nand UO_2303 (O_2303,N_24881,N_24942);
xor UO_2304 (O_2304,N_24321,N_24266);
and UO_2305 (O_2305,N_24116,N_24559);
xnor UO_2306 (O_2306,N_24700,N_24045);
or UO_2307 (O_2307,N_24468,N_24171);
nor UO_2308 (O_2308,N_24432,N_24512);
and UO_2309 (O_2309,N_24093,N_24404);
or UO_2310 (O_2310,N_24129,N_24108);
nor UO_2311 (O_2311,N_24173,N_24379);
nor UO_2312 (O_2312,N_24463,N_24265);
or UO_2313 (O_2313,N_24720,N_24438);
and UO_2314 (O_2314,N_24754,N_24942);
nor UO_2315 (O_2315,N_24351,N_24313);
or UO_2316 (O_2316,N_24416,N_24247);
or UO_2317 (O_2317,N_24649,N_24635);
nand UO_2318 (O_2318,N_24416,N_24760);
nor UO_2319 (O_2319,N_24462,N_24033);
and UO_2320 (O_2320,N_24939,N_24316);
nand UO_2321 (O_2321,N_24535,N_24276);
nor UO_2322 (O_2322,N_24884,N_24691);
or UO_2323 (O_2323,N_24553,N_24294);
nor UO_2324 (O_2324,N_24029,N_24306);
or UO_2325 (O_2325,N_24283,N_24726);
nor UO_2326 (O_2326,N_24508,N_24495);
xnor UO_2327 (O_2327,N_24223,N_24589);
nand UO_2328 (O_2328,N_24923,N_24979);
nor UO_2329 (O_2329,N_24887,N_24489);
nor UO_2330 (O_2330,N_24394,N_24847);
nor UO_2331 (O_2331,N_24487,N_24373);
nand UO_2332 (O_2332,N_24943,N_24160);
or UO_2333 (O_2333,N_24795,N_24159);
nand UO_2334 (O_2334,N_24685,N_24368);
nor UO_2335 (O_2335,N_24032,N_24121);
nor UO_2336 (O_2336,N_24131,N_24887);
xor UO_2337 (O_2337,N_24555,N_24116);
nand UO_2338 (O_2338,N_24384,N_24301);
nand UO_2339 (O_2339,N_24662,N_24392);
or UO_2340 (O_2340,N_24310,N_24509);
and UO_2341 (O_2341,N_24873,N_24250);
and UO_2342 (O_2342,N_24481,N_24098);
nand UO_2343 (O_2343,N_24019,N_24082);
xor UO_2344 (O_2344,N_24109,N_24447);
xnor UO_2345 (O_2345,N_24490,N_24161);
or UO_2346 (O_2346,N_24889,N_24862);
and UO_2347 (O_2347,N_24679,N_24622);
or UO_2348 (O_2348,N_24594,N_24298);
nand UO_2349 (O_2349,N_24877,N_24495);
nor UO_2350 (O_2350,N_24618,N_24095);
xor UO_2351 (O_2351,N_24742,N_24866);
and UO_2352 (O_2352,N_24395,N_24953);
xor UO_2353 (O_2353,N_24630,N_24316);
and UO_2354 (O_2354,N_24293,N_24780);
or UO_2355 (O_2355,N_24166,N_24119);
nor UO_2356 (O_2356,N_24491,N_24172);
nor UO_2357 (O_2357,N_24003,N_24359);
nor UO_2358 (O_2358,N_24947,N_24522);
or UO_2359 (O_2359,N_24859,N_24226);
nor UO_2360 (O_2360,N_24282,N_24969);
nand UO_2361 (O_2361,N_24465,N_24562);
nor UO_2362 (O_2362,N_24592,N_24710);
or UO_2363 (O_2363,N_24931,N_24447);
nand UO_2364 (O_2364,N_24045,N_24686);
nor UO_2365 (O_2365,N_24074,N_24462);
nand UO_2366 (O_2366,N_24687,N_24395);
nor UO_2367 (O_2367,N_24883,N_24158);
and UO_2368 (O_2368,N_24029,N_24656);
or UO_2369 (O_2369,N_24633,N_24819);
xor UO_2370 (O_2370,N_24827,N_24137);
and UO_2371 (O_2371,N_24061,N_24009);
nand UO_2372 (O_2372,N_24455,N_24529);
xor UO_2373 (O_2373,N_24699,N_24424);
nand UO_2374 (O_2374,N_24894,N_24069);
and UO_2375 (O_2375,N_24670,N_24743);
xor UO_2376 (O_2376,N_24456,N_24187);
and UO_2377 (O_2377,N_24343,N_24724);
xnor UO_2378 (O_2378,N_24319,N_24362);
xor UO_2379 (O_2379,N_24622,N_24813);
and UO_2380 (O_2380,N_24583,N_24381);
and UO_2381 (O_2381,N_24635,N_24276);
or UO_2382 (O_2382,N_24778,N_24105);
nand UO_2383 (O_2383,N_24868,N_24395);
nand UO_2384 (O_2384,N_24077,N_24538);
or UO_2385 (O_2385,N_24170,N_24784);
nor UO_2386 (O_2386,N_24819,N_24196);
xnor UO_2387 (O_2387,N_24974,N_24326);
nor UO_2388 (O_2388,N_24226,N_24155);
xor UO_2389 (O_2389,N_24617,N_24735);
xor UO_2390 (O_2390,N_24297,N_24252);
xor UO_2391 (O_2391,N_24688,N_24839);
and UO_2392 (O_2392,N_24409,N_24537);
nand UO_2393 (O_2393,N_24967,N_24342);
and UO_2394 (O_2394,N_24174,N_24291);
or UO_2395 (O_2395,N_24991,N_24142);
nor UO_2396 (O_2396,N_24574,N_24338);
and UO_2397 (O_2397,N_24906,N_24621);
xor UO_2398 (O_2398,N_24714,N_24899);
and UO_2399 (O_2399,N_24343,N_24354);
xnor UO_2400 (O_2400,N_24174,N_24954);
xnor UO_2401 (O_2401,N_24540,N_24410);
nand UO_2402 (O_2402,N_24517,N_24752);
or UO_2403 (O_2403,N_24630,N_24789);
and UO_2404 (O_2404,N_24769,N_24374);
and UO_2405 (O_2405,N_24854,N_24330);
and UO_2406 (O_2406,N_24031,N_24159);
nor UO_2407 (O_2407,N_24372,N_24194);
and UO_2408 (O_2408,N_24605,N_24150);
and UO_2409 (O_2409,N_24723,N_24172);
nor UO_2410 (O_2410,N_24319,N_24044);
nor UO_2411 (O_2411,N_24015,N_24053);
or UO_2412 (O_2412,N_24693,N_24844);
nor UO_2413 (O_2413,N_24038,N_24154);
nor UO_2414 (O_2414,N_24293,N_24990);
nor UO_2415 (O_2415,N_24001,N_24396);
xnor UO_2416 (O_2416,N_24166,N_24012);
xnor UO_2417 (O_2417,N_24862,N_24545);
or UO_2418 (O_2418,N_24461,N_24657);
or UO_2419 (O_2419,N_24879,N_24363);
or UO_2420 (O_2420,N_24927,N_24304);
or UO_2421 (O_2421,N_24576,N_24020);
xnor UO_2422 (O_2422,N_24177,N_24939);
or UO_2423 (O_2423,N_24763,N_24981);
and UO_2424 (O_2424,N_24725,N_24450);
and UO_2425 (O_2425,N_24828,N_24062);
xnor UO_2426 (O_2426,N_24117,N_24807);
and UO_2427 (O_2427,N_24201,N_24240);
or UO_2428 (O_2428,N_24897,N_24965);
and UO_2429 (O_2429,N_24318,N_24871);
nand UO_2430 (O_2430,N_24164,N_24485);
or UO_2431 (O_2431,N_24155,N_24802);
and UO_2432 (O_2432,N_24469,N_24043);
nand UO_2433 (O_2433,N_24473,N_24634);
and UO_2434 (O_2434,N_24274,N_24512);
nand UO_2435 (O_2435,N_24514,N_24530);
or UO_2436 (O_2436,N_24509,N_24653);
or UO_2437 (O_2437,N_24437,N_24352);
nor UO_2438 (O_2438,N_24566,N_24742);
and UO_2439 (O_2439,N_24845,N_24351);
xnor UO_2440 (O_2440,N_24406,N_24559);
and UO_2441 (O_2441,N_24040,N_24602);
nor UO_2442 (O_2442,N_24166,N_24710);
xor UO_2443 (O_2443,N_24526,N_24577);
nand UO_2444 (O_2444,N_24126,N_24683);
nand UO_2445 (O_2445,N_24987,N_24710);
and UO_2446 (O_2446,N_24932,N_24795);
and UO_2447 (O_2447,N_24031,N_24892);
and UO_2448 (O_2448,N_24751,N_24208);
nand UO_2449 (O_2449,N_24638,N_24180);
and UO_2450 (O_2450,N_24552,N_24477);
xor UO_2451 (O_2451,N_24549,N_24920);
nand UO_2452 (O_2452,N_24186,N_24809);
or UO_2453 (O_2453,N_24278,N_24687);
and UO_2454 (O_2454,N_24367,N_24607);
xor UO_2455 (O_2455,N_24279,N_24317);
nor UO_2456 (O_2456,N_24147,N_24866);
xnor UO_2457 (O_2457,N_24053,N_24983);
or UO_2458 (O_2458,N_24468,N_24604);
nand UO_2459 (O_2459,N_24373,N_24493);
xnor UO_2460 (O_2460,N_24502,N_24777);
or UO_2461 (O_2461,N_24559,N_24742);
xnor UO_2462 (O_2462,N_24838,N_24962);
nor UO_2463 (O_2463,N_24433,N_24027);
and UO_2464 (O_2464,N_24968,N_24797);
nor UO_2465 (O_2465,N_24182,N_24731);
xnor UO_2466 (O_2466,N_24766,N_24719);
and UO_2467 (O_2467,N_24327,N_24633);
xor UO_2468 (O_2468,N_24260,N_24713);
nor UO_2469 (O_2469,N_24951,N_24414);
nand UO_2470 (O_2470,N_24119,N_24525);
nor UO_2471 (O_2471,N_24775,N_24182);
and UO_2472 (O_2472,N_24179,N_24728);
and UO_2473 (O_2473,N_24050,N_24752);
nor UO_2474 (O_2474,N_24028,N_24015);
nand UO_2475 (O_2475,N_24545,N_24729);
nor UO_2476 (O_2476,N_24760,N_24559);
xnor UO_2477 (O_2477,N_24147,N_24664);
nand UO_2478 (O_2478,N_24031,N_24740);
or UO_2479 (O_2479,N_24652,N_24364);
nand UO_2480 (O_2480,N_24452,N_24511);
nand UO_2481 (O_2481,N_24109,N_24593);
nand UO_2482 (O_2482,N_24019,N_24383);
and UO_2483 (O_2483,N_24165,N_24476);
and UO_2484 (O_2484,N_24849,N_24961);
or UO_2485 (O_2485,N_24205,N_24387);
nand UO_2486 (O_2486,N_24559,N_24818);
nand UO_2487 (O_2487,N_24645,N_24312);
and UO_2488 (O_2488,N_24667,N_24166);
or UO_2489 (O_2489,N_24295,N_24001);
or UO_2490 (O_2490,N_24683,N_24094);
nand UO_2491 (O_2491,N_24003,N_24740);
and UO_2492 (O_2492,N_24363,N_24286);
or UO_2493 (O_2493,N_24892,N_24917);
xnor UO_2494 (O_2494,N_24353,N_24029);
nor UO_2495 (O_2495,N_24687,N_24631);
and UO_2496 (O_2496,N_24531,N_24329);
or UO_2497 (O_2497,N_24204,N_24009);
or UO_2498 (O_2498,N_24728,N_24083);
or UO_2499 (O_2499,N_24812,N_24431);
xnor UO_2500 (O_2500,N_24891,N_24881);
nand UO_2501 (O_2501,N_24461,N_24951);
nand UO_2502 (O_2502,N_24854,N_24861);
xor UO_2503 (O_2503,N_24545,N_24775);
or UO_2504 (O_2504,N_24839,N_24442);
nor UO_2505 (O_2505,N_24739,N_24011);
nor UO_2506 (O_2506,N_24992,N_24478);
nor UO_2507 (O_2507,N_24818,N_24480);
nor UO_2508 (O_2508,N_24697,N_24013);
or UO_2509 (O_2509,N_24097,N_24334);
xnor UO_2510 (O_2510,N_24228,N_24855);
and UO_2511 (O_2511,N_24217,N_24944);
nor UO_2512 (O_2512,N_24456,N_24073);
nor UO_2513 (O_2513,N_24280,N_24420);
or UO_2514 (O_2514,N_24535,N_24211);
nand UO_2515 (O_2515,N_24678,N_24724);
nor UO_2516 (O_2516,N_24146,N_24748);
or UO_2517 (O_2517,N_24786,N_24087);
xor UO_2518 (O_2518,N_24346,N_24038);
or UO_2519 (O_2519,N_24036,N_24880);
nor UO_2520 (O_2520,N_24416,N_24335);
or UO_2521 (O_2521,N_24501,N_24940);
nor UO_2522 (O_2522,N_24234,N_24078);
or UO_2523 (O_2523,N_24810,N_24238);
nand UO_2524 (O_2524,N_24129,N_24627);
nand UO_2525 (O_2525,N_24258,N_24893);
nand UO_2526 (O_2526,N_24754,N_24552);
nor UO_2527 (O_2527,N_24896,N_24287);
nor UO_2528 (O_2528,N_24123,N_24990);
xnor UO_2529 (O_2529,N_24249,N_24110);
nand UO_2530 (O_2530,N_24976,N_24497);
nand UO_2531 (O_2531,N_24312,N_24470);
xnor UO_2532 (O_2532,N_24708,N_24854);
nor UO_2533 (O_2533,N_24166,N_24995);
nand UO_2534 (O_2534,N_24423,N_24754);
xnor UO_2535 (O_2535,N_24599,N_24064);
and UO_2536 (O_2536,N_24140,N_24099);
xnor UO_2537 (O_2537,N_24176,N_24299);
nand UO_2538 (O_2538,N_24985,N_24494);
nand UO_2539 (O_2539,N_24476,N_24735);
nand UO_2540 (O_2540,N_24720,N_24328);
and UO_2541 (O_2541,N_24863,N_24587);
or UO_2542 (O_2542,N_24802,N_24690);
and UO_2543 (O_2543,N_24936,N_24883);
nand UO_2544 (O_2544,N_24547,N_24573);
and UO_2545 (O_2545,N_24550,N_24372);
xnor UO_2546 (O_2546,N_24522,N_24337);
or UO_2547 (O_2547,N_24551,N_24267);
xnor UO_2548 (O_2548,N_24545,N_24242);
and UO_2549 (O_2549,N_24077,N_24739);
nor UO_2550 (O_2550,N_24971,N_24297);
xnor UO_2551 (O_2551,N_24907,N_24964);
nor UO_2552 (O_2552,N_24029,N_24490);
nor UO_2553 (O_2553,N_24270,N_24546);
nor UO_2554 (O_2554,N_24106,N_24804);
or UO_2555 (O_2555,N_24582,N_24084);
or UO_2556 (O_2556,N_24393,N_24253);
or UO_2557 (O_2557,N_24218,N_24842);
xnor UO_2558 (O_2558,N_24630,N_24580);
or UO_2559 (O_2559,N_24843,N_24320);
nand UO_2560 (O_2560,N_24180,N_24078);
xnor UO_2561 (O_2561,N_24228,N_24150);
and UO_2562 (O_2562,N_24780,N_24092);
nand UO_2563 (O_2563,N_24727,N_24311);
nor UO_2564 (O_2564,N_24036,N_24199);
nand UO_2565 (O_2565,N_24595,N_24355);
xor UO_2566 (O_2566,N_24073,N_24020);
nor UO_2567 (O_2567,N_24847,N_24369);
nor UO_2568 (O_2568,N_24352,N_24020);
xor UO_2569 (O_2569,N_24914,N_24569);
and UO_2570 (O_2570,N_24990,N_24500);
and UO_2571 (O_2571,N_24503,N_24760);
and UO_2572 (O_2572,N_24616,N_24979);
or UO_2573 (O_2573,N_24934,N_24166);
xor UO_2574 (O_2574,N_24082,N_24625);
nand UO_2575 (O_2575,N_24260,N_24818);
xor UO_2576 (O_2576,N_24283,N_24575);
nor UO_2577 (O_2577,N_24491,N_24530);
nand UO_2578 (O_2578,N_24943,N_24076);
or UO_2579 (O_2579,N_24554,N_24172);
xnor UO_2580 (O_2580,N_24948,N_24621);
or UO_2581 (O_2581,N_24808,N_24368);
nand UO_2582 (O_2582,N_24013,N_24386);
nor UO_2583 (O_2583,N_24065,N_24208);
xor UO_2584 (O_2584,N_24572,N_24594);
or UO_2585 (O_2585,N_24124,N_24397);
nor UO_2586 (O_2586,N_24238,N_24384);
nand UO_2587 (O_2587,N_24517,N_24765);
or UO_2588 (O_2588,N_24576,N_24667);
nand UO_2589 (O_2589,N_24732,N_24631);
or UO_2590 (O_2590,N_24361,N_24924);
xnor UO_2591 (O_2591,N_24195,N_24129);
xor UO_2592 (O_2592,N_24547,N_24257);
xnor UO_2593 (O_2593,N_24259,N_24012);
or UO_2594 (O_2594,N_24449,N_24078);
or UO_2595 (O_2595,N_24309,N_24043);
or UO_2596 (O_2596,N_24041,N_24879);
nand UO_2597 (O_2597,N_24199,N_24229);
or UO_2598 (O_2598,N_24697,N_24267);
nand UO_2599 (O_2599,N_24701,N_24859);
nand UO_2600 (O_2600,N_24997,N_24052);
or UO_2601 (O_2601,N_24789,N_24479);
nand UO_2602 (O_2602,N_24970,N_24208);
nand UO_2603 (O_2603,N_24679,N_24223);
nor UO_2604 (O_2604,N_24981,N_24370);
or UO_2605 (O_2605,N_24394,N_24901);
nand UO_2606 (O_2606,N_24331,N_24358);
nand UO_2607 (O_2607,N_24041,N_24674);
nor UO_2608 (O_2608,N_24086,N_24511);
nor UO_2609 (O_2609,N_24045,N_24129);
xnor UO_2610 (O_2610,N_24950,N_24208);
or UO_2611 (O_2611,N_24950,N_24583);
xnor UO_2612 (O_2612,N_24427,N_24319);
nor UO_2613 (O_2613,N_24165,N_24149);
xnor UO_2614 (O_2614,N_24447,N_24647);
and UO_2615 (O_2615,N_24321,N_24428);
and UO_2616 (O_2616,N_24415,N_24803);
nor UO_2617 (O_2617,N_24382,N_24178);
nand UO_2618 (O_2618,N_24832,N_24014);
nand UO_2619 (O_2619,N_24649,N_24739);
and UO_2620 (O_2620,N_24279,N_24442);
nand UO_2621 (O_2621,N_24359,N_24835);
xnor UO_2622 (O_2622,N_24356,N_24938);
xnor UO_2623 (O_2623,N_24524,N_24087);
nor UO_2624 (O_2624,N_24011,N_24740);
or UO_2625 (O_2625,N_24755,N_24819);
nand UO_2626 (O_2626,N_24245,N_24950);
xor UO_2627 (O_2627,N_24369,N_24523);
and UO_2628 (O_2628,N_24324,N_24458);
nor UO_2629 (O_2629,N_24613,N_24280);
xor UO_2630 (O_2630,N_24461,N_24021);
nand UO_2631 (O_2631,N_24439,N_24732);
nor UO_2632 (O_2632,N_24714,N_24689);
nand UO_2633 (O_2633,N_24506,N_24214);
xnor UO_2634 (O_2634,N_24265,N_24562);
nor UO_2635 (O_2635,N_24874,N_24236);
nand UO_2636 (O_2636,N_24539,N_24658);
xnor UO_2637 (O_2637,N_24702,N_24041);
nand UO_2638 (O_2638,N_24448,N_24638);
nand UO_2639 (O_2639,N_24895,N_24002);
and UO_2640 (O_2640,N_24471,N_24315);
xnor UO_2641 (O_2641,N_24730,N_24532);
nand UO_2642 (O_2642,N_24712,N_24409);
and UO_2643 (O_2643,N_24285,N_24564);
and UO_2644 (O_2644,N_24149,N_24256);
xor UO_2645 (O_2645,N_24667,N_24079);
nor UO_2646 (O_2646,N_24622,N_24764);
nor UO_2647 (O_2647,N_24495,N_24446);
nand UO_2648 (O_2648,N_24151,N_24314);
and UO_2649 (O_2649,N_24753,N_24456);
or UO_2650 (O_2650,N_24237,N_24934);
nor UO_2651 (O_2651,N_24921,N_24475);
or UO_2652 (O_2652,N_24091,N_24874);
nand UO_2653 (O_2653,N_24697,N_24053);
or UO_2654 (O_2654,N_24990,N_24021);
nor UO_2655 (O_2655,N_24978,N_24824);
nand UO_2656 (O_2656,N_24238,N_24915);
xnor UO_2657 (O_2657,N_24271,N_24784);
or UO_2658 (O_2658,N_24014,N_24499);
and UO_2659 (O_2659,N_24415,N_24877);
nor UO_2660 (O_2660,N_24276,N_24326);
nor UO_2661 (O_2661,N_24744,N_24628);
or UO_2662 (O_2662,N_24187,N_24516);
nand UO_2663 (O_2663,N_24784,N_24951);
and UO_2664 (O_2664,N_24527,N_24022);
nand UO_2665 (O_2665,N_24817,N_24659);
xor UO_2666 (O_2666,N_24713,N_24775);
and UO_2667 (O_2667,N_24129,N_24642);
xnor UO_2668 (O_2668,N_24799,N_24880);
or UO_2669 (O_2669,N_24065,N_24941);
nand UO_2670 (O_2670,N_24795,N_24895);
and UO_2671 (O_2671,N_24177,N_24985);
xor UO_2672 (O_2672,N_24170,N_24731);
nor UO_2673 (O_2673,N_24357,N_24158);
nor UO_2674 (O_2674,N_24134,N_24962);
or UO_2675 (O_2675,N_24921,N_24276);
or UO_2676 (O_2676,N_24390,N_24406);
xnor UO_2677 (O_2677,N_24297,N_24927);
nor UO_2678 (O_2678,N_24775,N_24605);
or UO_2679 (O_2679,N_24809,N_24676);
nand UO_2680 (O_2680,N_24787,N_24225);
and UO_2681 (O_2681,N_24615,N_24892);
or UO_2682 (O_2682,N_24272,N_24540);
nor UO_2683 (O_2683,N_24451,N_24508);
nor UO_2684 (O_2684,N_24494,N_24387);
or UO_2685 (O_2685,N_24267,N_24826);
nor UO_2686 (O_2686,N_24161,N_24291);
xnor UO_2687 (O_2687,N_24155,N_24836);
nor UO_2688 (O_2688,N_24497,N_24987);
xor UO_2689 (O_2689,N_24906,N_24580);
nor UO_2690 (O_2690,N_24992,N_24878);
nand UO_2691 (O_2691,N_24462,N_24771);
or UO_2692 (O_2692,N_24465,N_24430);
and UO_2693 (O_2693,N_24128,N_24141);
nor UO_2694 (O_2694,N_24789,N_24206);
or UO_2695 (O_2695,N_24503,N_24629);
nor UO_2696 (O_2696,N_24092,N_24468);
and UO_2697 (O_2697,N_24121,N_24299);
or UO_2698 (O_2698,N_24674,N_24038);
and UO_2699 (O_2699,N_24858,N_24006);
or UO_2700 (O_2700,N_24242,N_24052);
and UO_2701 (O_2701,N_24728,N_24356);
xor UO_2702 (O_2702,N_24410,N_24128);
or UO_2703 (O_2703,N_24256,N_24436);
or UO_2704 (O_2704,N_24917,N_24192);
or UO_2705 (O_2705,N_24973,N_24624);
nand UO_2706 (O_2706,N_24575,N_24317);
nand UO_2707 (O_2707,N_24868,N_24335);
or UO_2708 (O_2708,N_24588,N_24640);
xor UO_2709 (O_2709,N_24554,N_24835);
nand UO_2710 (O_2710,N_24406,N_24980);
and UO_2711 (O_2711,N_24479,N_24868);
or UO_2712 (O_2712,N_24319,N_24929);
and UO_2713 (O_2713,N_24150,N_24766);
nand UO_2714 (O_2714,N_24487,N_24583);
and UO_2715 (O_2715,N_24666,N_24294);
nand UO_2716 (O_2716,N_24145,N_24420);
nor UO_2717 (O_2717,N_24914,N_24583);
nor UO_2718 (O_2718,N_24920,N_24443);
or UO_2719 (O_2719,N_24668,N_24376);
nand UO_2720 (O_2720,N_24980,N_24312);
or UO_2721 (O_2721,N_24882,N_24281);
and UO_2722 (O_2722,N_24109,N_24512);
nand UO_2723 (O_2723,N_24259,N_24570);
xor UO_2724 (O_2724,N_24902,N_24165);
nand UO_2725 (O_2725,N_24052,N_24187);
xor UO_2726 (O_2726,N_24500,N_24509);
xor UO_2727 (O_2727,N_24597,N_24043);
and UO_2728 (O_2728,N_24623,N_24106);
xor UO_2729 (O_2729,N_24607,N_24487);
or UO_2730 (O_2730,N_24552,N_24781);
and UO_2731 (O_2731,N_24903,N_24334);
or UO_2732 (O_2732,N_24489,N_24268);
nand UO_2733 (O_2733,N_24199,N_24012);
nor UO_2734 (O_2734,N_24960,N_24760);
nand UO_2735 (O_2735,N_24327,N_24168);
nor UO_2736 (O_2736,N_24312,N_24952);
nand UO_2737 (O_2737,N_24239,N_24434);
xor UO_2738 (O_2738,N_24242,N_24659);
xor UO_2739 (O_2739,N_24077,N_24272);
nand UO_2740 (O_2740,N_24637,N_24358);
nand UO_2741 (O_2741,N_24348,N_24391);
xnor UO_2742 (O_2742,N_24432,N_24341);
nand UO_2743 (O_2743,N_24405,N_24541);
and UO_2744 (O_2744,N_24491,N_24924);
nor UO_2745 (O_2745,N_24007,N_24456);
nand UO_2746 (O_2746,N_24138,N_24444);
xnor UO_2747 (O_2747,N_24942,N_24906);
or UO_2748 (O_2748,N_24498,N_24541);
nor UO_2749 (O_2749,N_24170,N_24809);
or UO_2750 (O_2750,N_24721,N_24757);
or UO_2751 (O_2751,N_24587,N_24648);
nor UO_2752 (O_2752,N_24937,N_24209);
xor UO_2753 (O_2753,N_24032,N_24240);
nor UO_2754 (O_2754,N_24080,N_24807);
nor UO_2755 (O_2755,N_24633,N_24690);
or UO_2756 (O_2756,N_24749,N_24306);
nand UO_2757 (O_2757,N_24661,N_24977);
nand UO_2758 (O_2758,N_24792,N_24722);
and UO_2759 (O_2759,N_24410,N_24082);
and UO_2760 (O_2760,N_24076,N_24297);
xor UO_2761 (O_2761,N_24013,N_24407);
nand UO_2762 (O_2762,N_24331,N_24844);
and UO_2763 (O_2763,N_24082,N_24873);
or UO_2764 (O_2764,N_24778,N_24213);
and UO_2765 (O_2765,N_24533,N_24802);
and UO_2766 (O_2766,N_24246,N_24268);
and UO_2767 (O_2767,N_24082,N_24357);
or UO_2768 (O_2768,N_24041,N_24196);
nor UO_2769 (O_2769,N_24857,N_24326);
or UO_2770 (O_2770,N_24252,N_24333);
xor UO_2771 (O_2771,N_24335,N_24433);
or UO_2772 (O_2772,N_24054,N_24010);
nand UO_2773 (O_2773,N_24179,N_24339);
xnor UO_2774 (O_2774,N_24668,N_24497);
xnor UO_2775 (O_2775,N_24234,N_24663);
xor UO_2776 (O_2776,N_24982,N_24762);
and UO_2777 (O_2777,N_24989,N_24062);
or UO_2778 (O_2778,N_24841,N_24953);
and UO_2779 (O_2779,N_24923,N_24038);
nor UO_2780 (O_2780,N_24904,N_24266);
xor UO_2781 (O_2781,N_24374,N_24775);
and UO_2782 (O_2782,N_24473,N_24483);
or UO_2783 (O_2783,N_24721,N_24755);
or UO_2784 (O_2784,N_24207,N_24892);
or UO_2785 (O_2785,N_24111,N_24733);
or UO_2786 (O_2786,N_24663,N_24835);
nand UO_2787 (O_2787,N_24452,N_24796);
nand UO_2788 (O_2788,N_24885,N_24080);
or UO_2789 (O_2789,N_24720,N_24368);
or UO_2790 (O_2790,N_24525,N_24326);
nand UO_2791 (O_2791,N_24769,N_24720);
nor UO_2792 (O_2792,N_24874,N_24544);
or UO_2793 (O_2793,N_24926,N_24814);
nand UO_2794 (O_2794,N_24417,N_24004);
nand UO_2795 (O_2795,N_24636,N_24095);
nand UO_2796 (O_2796,N_24026,N_24968);
nand UO_2797 (O_2797,N_24683,N_24051);
nor UO_2798 (O_2798,N_24627,N_24385);
nor UO_2799 (O_2799,N_24441,N_24991);
nor UO_2800 (O_2800,N_24818,N_24501);
nand UO_2801 (O_2801,N_24222,N_24899);
nor UO_2802 (O_2802,N_24411,N_24830);
nor UO_2803 (O_2803,N_24713,N_24995);
nand UO_2804 (O_2804,N_24320,N_24244);
nor UO_2805 (O_2805,N_24647,N_24772);
xnor UO_2806 (O_2806,N_24971,N_24902);
and UO_2807 (O_2807,N_24826,N_24215);
and UO_2808 (O_2808,N_24413,N_24137);
nor UO_2809 (O_2809,N_24951,N_24248);
nor UO_2810 (O_2810,N_24259,N_24755);
and UO_2811 (O_2811,N_24977,N_24739);
xnor UO_2812 (O_2812,N_24445,N_24211);
xnor UO_2813 (O_2813,N_24267,N_24543);
nand UO_2814 (O_2814,N_24932,N_24024);
or UO_2815 (O_2815,N_24553,N_24163);
nand UO_2816 (O_2816,N_24530,N_24941);
or UO_2817 (O_2817,N_24730,N_24317);
nand UO_2818 (O_2818,N_24548,N_24194);
nor UO_2819 (O_2819,N_24874,N_24900);
nor UO_2820 (O_2820,N_24547,N_24176);
and UO_2821 (O_2821,N_24483,N_24755);
nand UO_2822 (O_2822,N_24208,N_24875);
or UO_2823 (O_2823,N_24032,N_24164);
or UO_2824 (O_2824,N_24449,N_24675);
or UO_2825 (O_2825,N_24251,N_24136);
xnor UO_2826 (O_2826,N_24826,N_24989);
and UO_2827 (O_2827,N_24744,N_24507);
xor UO_2828 (O_2828,N_24983,N_24125);
xor UO_2829 (O_2829,N_24412,N_24017);
and UO_2830 (O_2830,N_24067,N_24707);
or UO_2831 (O_2831,N_24004,N_24622);
or UO_2832 (O_2832,N_24422,N_24716);
nand UO_2833 (O_2833,N_24365,N_24770);
and UO_2834 (O_2834,N_24372,N_24553);
nand UO_2835 (O_2835,N_24627,N_24965);
xor UO_2836 (O_2836,N_24915,N_24095);
nand UO_2837 (O_2837,N_24056,N_24758);
and UO_2838 (O_2838,N_24323,N_24812);
xor UO_2839 (O_2839,N_24017,N_24915);
nand UO_2840 (O_2840,N_24389,N_24999);
xnor UO_2841 (O_2841,N_24736,N_24401);
and UO_2842 (O_2842,N_24341,N_24895);
or UO_2843 (O_2843,N_24298,N_24982);
xnor UO_2844 (O_2844,N_24230,N_24730);
nor UO_2845 (O_2845,N_24402,N_24517);
xor UO_2846 (O_2846,N_24805,N_24201);
and UO_2847 (O_2847,N_24873,N_24311);
or UO_2848 (O_2848,N_24550,N_24308);
nor UO_2849 (O_2849,N_24322,N_24231);
xor UO_2850 (O_2850,N_24632,N_24551);
or UO_2851 (O_2851,N_24710,N_24339);
and UO_2852 (O_2852,N_24431,N_24636);
nor UO_2853 (O_2853,N_24588,N_24454);
xor UO_2854 (O_2854,N_24572,N_24942);
xnor UO_2855 (O_2855,N_24658,N_24780);
nand UO_2856 (O_2856,N_24022,N_24991);
and UO_2857 (O_2857,N_24198,N_24081);
or UO_2858 (O_2858,N_24154,N_24673);
xor UO_2859 (O_2859,N_24707,N_24072);
nand UO_2860 (O_2860,N_24197,N_24492);
and UO_2861 (O_2861,N_24389,N_24147);
nand UO_2862 (O_2862,N_24635,N_24392);
nor UO_2863 (O_2863,N_24829,N_24869);
or UO_2864 (O_2864,N_24339,N_24114);
xnor UO_2865 (O_2865,N_24918,N_24660);
nor UO_2866 (O_2866,N_24872,N_24159);
or UO_2867 (O_2867,N_24672,N_24001);
or UO_2868 (O_2868,N_24018,N_24552);
nand UO_2869 (O_2869,N_24244,N_24416);
and UO_2870 (O_2870,N_24972,N_24958);
xnor UO_2871 (O_2871,N_24173,N_24685);
xnor UO_2872 (O_2872,N_24628,N_24352);
and UO_2873 (O_2873,N_24616,N_24238);
xnor UO_2874 (O_2874,N_24907,N_24543);
nor UO_2875 (O_2875,N_24595,N_24217);
and UO_2876 (O_2876,N_24196,N_24716);
and UO_2877 (O_2877,N_24272,N_24047);
nand UO_2878 (O_2878,N_24162,N_24187);
nand UO_2879 (O_2879,N_24170,N_24860);
xnor UO_2880 (O_2880,N_24858,N_24777);
and UO_2881 (O_2881,N_24248,N_24553);
nand UO_2882 (O_2882,N_24034,N_24849);
xnor UO_2883 (O_2883,N_24719,N_24197);
nand UO_2884 (O_2884,N_24099,N_24941);
nor UO_2885 (O_2885,N_24333,N_24135);
and UO_2886 (O_2886,N_24507,N_24634);
nand UO_2887 (O_2887,N_24394,N_24556);
nor UO_2888 (O_2888,N_24854,N_24898);
and UO_2889 (O_2889,N_24790,N_24098);
nor UO_2890 (O_2890,N_24598,N_24320);
nand UO_2891 (O_2891,N_24058,N_24081);
xor UO_2892 (O_2892,N_24673,N_24125);
and UO_2893 (O_2893,N_24583,N_24746);
and UO_2894 (O_2894,N_24425,N_24115);
xnor UO_2895 (O_2895,N_24699,N_24190);
nand UO_2896 (O_2896,N_24761,N_24463);
xor UO_2897 (O_2897,N_24408,N_24458);
nor UO_2898 (O_2898,N_24076,N_24684);
nor UO_2899 (O_2899,N_24487,N_24404);
xnor UO_2900 (O_2900,N_24712,N_24887);
xnor UO_2901 (O_2901,N_24068,N_24965);
xnor UO_2902 (O_2902,N_24839,N_24605);
xor UO_2903 (O_2903,N_24655,N_24737);
and UO_2904 (O_2904,N_24609,N_24658);
and UO_2905 (O_2905,N_24691,N_24089);
or UO_2906 (O_2906,N_24586,N_24726);
xor UO_2907 (O_2907,N_24956,N_24284);
nand UO_2908 (O_2908,N_24063,N_24044);
nor UO_2909 (O_2909,N_24129,N_24365);
xor UO_2910 (O_2910,N_24064,N_24225);
nand UO_2911 (O_2911,N_24711,N_24872);
nand UO_2912 (O_2912,N_24680,N_24780);
nand UO_2913 (O_2913,N_24487,N_24739);
nor UO_2914 (O_2914,N_24757,N_24479);
nor UO_2915 (O_2915,N_24383,N_24933);
and UO_2916 (O_2916,N_24625,N_24399);
and UO_2917 (O_2917,N_24364,N_24585);
and UO_2918 (O_2918,N_24145,N_24084);
xor UO_2919 (O_2919,N_24004,N_24048);
nand UO_2920 (O_2920,N_24755,N_24143);
nand UO_2921 (O_2921,N_24811,N_24081);
nor UO_2922 (O_2922,N_24090,N_24924);
and UO_2923 (O_2923,N_24596,N_24648);
or UO_2924 (O_2924,N_24489,N_24590);
and UO_2925 (O_2925,N_24126,N_24913);
xnor UO_2926 (O_2926,N_24028,N_24662);
nor UO_2927 (O_2927,N_24002,N_24429);
nand UO_2928 (O_2928,N_24201,N_24111);
xnor UO_2929 (O_2929,N_24527,N_24964);
nor UO_2930 (O_2930,N_24805,N_24921);
and UO_2931 (O_2931,N_24918,N_24720);
or UO_2932 (O_2932,N_24483,N_24451);
nand UO_2933 (O_2933,N_24690,N_24626);
xor UO_2934 (O_2934,N_24412,N_24537);
or UO_2935 (O_2935,N_24748,N_24339);
nor UO_2936 (O_2936,N_24139,N_24993);
and UO_2937 (O_2937,N_24058,N_24259);
and UO_2938 (O_2938,N_24131,N_24687);
and UO_2939 (O_2939,N_24997,N_24331);
nand UO_2940 (O_2940,N_24185,N_24006);
nand UO_2941 (O_2941,N_24189,N_24847);
nor UO_2942 (O_2942,N_24121,N_24053);
or UO_2943 (O_2943,N_24415,N_24720);
or UO_2944 (O_2944,N_24179,N_24398);
or UO_2945 (O_2945,N_24890,N_24368);
nor UO_2946 (O_2946,N_24868,N_24433);
or UO_2947 (O_2947,N_24241,N_24902);
and UO_2948 (O_2948,N_24818,N_24297);
nor UO_2949 (O_2949,N_24962,N_24855);
nor UO_2950 (O_2950,N_24295,N_24284);
nand UO_2951 (O_2951,N_24054,N_24126);
nor UO_2952 (O_2952,N_24173,N_24138);
nand UO_2953 (O_2953,N_24176,N_24709);
nor UO_2954 (O_2954,N_24094,N_24637);
xor UO_2955 (O_2955,N_24633,N_24336);
nor UO_2956 (O_2956,N_24380,N_24969);
or UO_2957 (O_2957,N_24902,N_24104);
xnor UO_2958 (O_2958,N_24311,N_24077);
or UO_2959 (O_2959,N_24151,N_24905);
nand UO_2960 (O_2960,N_24213,N_24750);
nand UO_2961 (O_2961,N_24997,N_24157);
or UO_2962 (O_2962,N_24886,N_24643);
nor UO_2963 (O_2963,N_24181,N_24496);
nor UO_2964 (O_2964,N_24130,N_24178);
xor UO_2965 (O_2965,N_24621,N_24741);
and UO_2966 (O_2966,N_24918,N_24467);
nor UO_2967 (O_2967,N_24098,N_24265);
and UO_2968 (O_2968,N_24833,N_24417);
or UO_2969 (O_2969,N_24111,N_24931);
and UO_2970 (O_2970,N_24030,N_24489);
xnor UO_2971 (O_2971,N_24246,N_24025);
nand UO_2972 (O_2972,N_24614,N_24342);
nand UO_2973 (O_2973,N_24206,N_24619);
nor UO_2974 (O_2974,N_24089,N_24729);
and UO_2975 (O_2975,N_24074,N_24590);
or UO_2976 (O_2976,N_24274,N_24020);
nand UO_2977 (O_2977,N_24696,N_24905);
or UO_2978 (O_2978,N_24485,N_24258);
xor UO_2979 (O_2979,N_24772,N_24864);
and UO_2980 (O_2980,N_24062,N_24014);
nand UO_2981 (O_2981,N_24929,N_24879);
or UO_2982 (O_2982,N_24159,N_24939);
nor UO_2983 (O_2983,N_24031,N_24133);
and UO_2984 (O_2984,N_24470,N_24160);
xnor UO_2985 (O_2985,N_24309,N_24395);
or UO_2986 (O_2986,N_24146,N_24238);
nor UO_2987 (O_2987,N_24172,N_24313);
nor UO_2988 (O_2988,N_24834,N_24471);
and UO_2989 (O_2989,N_24300,N_24377);
nor UO_2990 (O_2990,N_24467,N_24947);
or UO_2991 (O_2991,N_24005,N_24192);
nor UO_2992 (O_2992,N_24140,N_24750);
or UO_2993 (O_2993,N_24616,N_24531);
or UO_2994 (O_2994,N_24967,N_24175);
and UO_2995 (O_2995,N_24438,N_24426);
nand UO_2996 (O_2996,N_24083,N_24410);
nor UO_2997 (O_2997,N_24772,N_24235);
or UO_2998 (O_2998,N_24057,N_24893);
xor UO_2999 (O_2999,N_24129,N_24789);
endmodule