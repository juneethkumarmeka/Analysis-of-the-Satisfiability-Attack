module basic_5000_50000_5000_20_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_27,In_388);
and U1 (N_1,In_4335,In_1422);
xor U2 (N_2,In_1694,In_4087);
or U3 (N_3,In_816,In_3507);
and U4 (N_4,In_3989,In_1120);
nor U5 (N_5,In_4590,In_3320);
xnor U6 (N_6,In_2266,In_2520);
nand U7 (N_7,In_2377,In_4659);
nor U8 (N_8,In_4854,In_213);
and U9 (N_9,In_2633,In_2616);
and U10 (N_10,In_2093,In_4143);
nand U11 (N_11,In_531,In_4060);
nand U12 (N_12,In_2521,In_3578);
or U13 (N_13,In_1272,In_2601);
or U14 (N_14,In_2823,In_4331);
and U15 (N_15,In_521,In_3251);
nor U16 (N_16,In_3565,In_1324);
xnor U17 (N_17,In_15,In_2358);
nand U18 (N_18,In_3272,In_4301);
or U19 (N_19,In_2865,In_4007);
xor U20 (N_20,In_3424,In_666);
and U21 (N_21,In_3038,In_580);
nor U22 (N_22,In_2537,In_1001);
nor U23 (N_23,In_2803,In_3802);
nand U24 (N_24,In_185,In_2594);
and U25 (N_25,In_4797,In_1091);
nor U26 (N_26,In_1160,In_786);
nor U27 (N_27,In_924,In_722);
xor U28 (N_28,In_2951,In_3872);
nand U29 (N_29,In_3267,In_1236);
nand U30 (N_30,In_3150,In_290);
and U31 (N_31,In_1306,In_1019);
nor U32 (N_32,In_4226,In_4651);
or U33 (N_33,In_276,In_3262);
xor U34 (N_34,In_3679,In_198);
nor U35 (N_35,In_2811,In_360);
xnor U36 (N_36,In_4295,In_1470);
nand U37 (N_37,In_2932,In_4555);
nor U38 (N_38,In_335,In_1279);
xnor U39 (N_39,In_2578,In_4862);
nand U40 (N_40,In_2718,In_2863);
or U41 (N_41,In_4100,In_1150);
or U42 (N_42,In_3081,In_240);
or U43 (N_43,In_4534,In_4210);
and U44 (N_44,In_4605,In_1217);
xor U45 (N_45,In_3454,In_1963);
nand U46 (N_46,In_1660,In_227);
nor U47 (N_47,In_927,In_1901);
nor U48 (N_48,In_1551,In_4182);
nor U49 (N_49,In_3514,In_4760);
or U50 (N_50,In_3299,In_2275);
or U51 (N_51,In_4003,In_43);
nor U52 (N_52,In_3619,In_624);
nor U53 (N_53,In_196,In_4468);
xnor U54 (N_54,In_919,In_3902);
and U55 (N_55,In_2693,In_3435);
nand U56 (N_56,In_432,In_1226);
or U57 (N_57,In_289,In_607);
xor U58 (N_58,In_4195,In_4307);
xor U59 (N_59,In_3254,In_3582);
xnor U60 (N_60,In_511,In_2373);
nor U61 (N_61,In_1305,In_1478);
or U62 (N_62,In_3512,In_433);
xnor U63 (N_63,In_2919,In_3371);
xnor U64 (N_64,In_2945,In_1555);
nor U65 (N_65,In_1987,In_2708);
or U66 (N_66,In_4937,In_4643);
nand U67 (N_67,In_2965,In_794);
or U68 (N_68,In_206,In_908);
xnor U69 (N_69,In_3640,In_2185);
nor U70 (N_70,In_1501,In_678);
and U71 (N_71,In_915,In_4022);
and U72 (N_72,In_3404,In_4571);
and U73 (N_73,In_125,In_324);
or U74 (N_74,In_1605,In_1618);
xor U75 (N_75,In_3645,In_4027);
nor U76 (N_76,In_1836,In_4709);
xor U77 (N_77,In_3309,In_3470);
and U78 (N_78,In_2286,In_2844);
nand U79 (N_79,In_771,In_4731);
nor U80 (N_80,In_3000,In_3303);
xor U81 (N_81,In_1566,In_749);
xor U82 (N_82,In_2488,In_824);
and U83 (N_83,In_68,In_54);
nor U84 (N_84,In_4650,In_3172);
or U85 (N_85,In_2943,In_3572);
or U86 (N_86,In_4313,In_172);
nand U87 (N_87,In_2478,In_1336);
or U88 (N_88,In_4603,In_3706);
nor U89 (N_89,In_3852,In_2716);
or U90 (N_90,In_3359,In_569);
nand U91 (N_91,In_4916,In_2273);
nor U92 (N_92,In_1585,In_4745);
xor U93 (N_93,In_1093,In_2098);
and U94 (N_94,In_1870,In_62);
or U95 (N_95,In_2729,In_67);
nor U96 (N_96,In_4469,In_4221);
nor U97 (N_97,In_4844,In_3346);
nor U98 (N_98,In_4722,In_3307);
xnor U99 (N_99,In_3928,In_3784);
nor U100 (N_100,In_2506,In_4621);
xor U101 (N_101,In_4547,In_4391);
and U102 (N_102,In_623,In_3310);
or U103 (N_103,In_1966,In_56);
and U104 (N_104,In_1500,In_4888);
nand U105 (N_105,In_3682,In_2356);
nand U106 (N_106,In_1223,In_469);
xor U107 (N_107,In_4193,In_1420);
nor U108 (N_108,In_1923,In_4244);
xor U109 (N_109,In_1925,In_853);
nand U110 (N_110,In_1601,In_1561);
nand U111 (N_111,In_1556,In_3164);
nand U112 (N_112,In_2649,In_262);
or U113 (N_113,In_2902,In_349);
and U114 (N_114,In_1543,In_4541);
or U115 (N_115,In_3003,In_4801);
nor U116 (N_116,In_1860,In_4302);
or U117 (N_117,In_2855,In_2330);
nand U118 (N_118,In_2542,In_2427);
or U119 (N_119,In_2894,In_4598);
nand U120 (N_120,In_3955,In_1774);
nand U121 (N_121,In_4150,In_800);
nand U122 (N_122,In_4356,In_4281);
nand U123 (N_123,In_2576,In_3407);
nor U124 (N_124,In_543,In_4405);
xnor U125 (N_125,In_2043,In_4373);
nand U126 (N_126,In_396,In_1434);
xnor U127 (N_127,In_4358,In_3510);
and U128 (N_128,In_2981,In_4719);
and U129 (N_129,In_4018,In_1675);
nand U130 (N_130,In_1303,In_2342);
nor U131 (N_131,In_1875,In_914);
and U132 (N_132,In_851,In_1291);
xor U133 (N_133,In_3838,In_2442);
nor U134 (N_134,In_3830,In_3213);
nor U135 (N_135,In_4668,In_3304);
and U136 (N_136,In_1273,In_4235);
xnor U137 (N_137,In_3867,In_3613);
nand U138 (N_138,In_1109,In_310);
and U139 (N_139,In_934,In_4699);
nor U140 (N_140,In_3035,In_353);
nand U141 (N_141,In_3440,In_719);
nor U142 (N_142,In_4248,In_2390);
or U143 (N_143,In_949,In_876);
xor U144 (N_144,In_402,In_418);
and U145 (N_145,In_3597,In_309);
or U146 (N_146,In_3399,In_242);
nor U147 (N_147,In_4136,In_3220);
nor U148 (N_148,In_2972,In_3764);
and U149 (N_149,In_1718,In_1611);
nand U150 (N_150,In_211,In_2928);
nand U151 (N_151,In_305,In_2210);
xnor U152 (N_152,In_319,In_2630);
and U153 (N_153,In_93,In_727);
and U154 (N_154,In_4480,In_3427);
or U155 (N_155,In_939,In_1803);
xnor U156 (N_156,In_3699,In_2942);
xnor U157 (N_157,In_2124,In_3810);
nor U158 (N_158,In_5,In_415);
and U159 (N_159,In_2704,In_4656);
or U160 (N_160,In_773,In_4697);
nor U161 (N_161,In_2446,In_891);
xnor U162 (N_162,In_1285,In_3455);
xor U163 (N_163,In_2084,In_2386);
nand U164 (N_164,In_2510,In_1945);
or U165 (N_165,In_3697,In_3244);
nor U166 (N_166,In_2949,In_1076);
or U167 (N_167,In_2264,In_401);
xor U168 (N_168,In_634,In_374);
or U169 (N_169,In_3696,In_1363);
or U170 (N_170,In_1587,In_3165);
nor U171 (N_171,In_3453,In_3538);
nand U172 (N_172,In_4247,In_1340);
nand U173 (N_173,In_1293,In_3231);
nand U174 (N_174,In_4735,In_2088);
xor U175 (N_175,In_1265,In_2192);
nand U176 (N_176,In_1145,In_435);
nor U177 (N_177,In_457,In_2870);
nand U178 (N_178,In_829,In_2899);
xor U179 (N_179,In_490,In_2156);
nor U180 (N_180,In_2692,In_3295);
nor U181 (N_181,In_1107,In_4300);
or U182 (N_182,In_2437,In_3936);
or U183 (N_183,In_4979,In_333);
or U184 (N_184,In_4073,In_2285);
nand U185 (N_185,In_1046,In_1616);
nand U186 (N_186,In_1043,In_3496);
or U187 (N_187,In_4428,In_2830);
nand U188 (N_188,In_3559,In_1827);
xnor U189 (N_189,In_651,In_3495);
nor U190 (N_190,In_2585,In_2355);
and U191 (N_191,In_3439,In_4496);
or U192 (N_192,In_3913,In_2208);
nand U193 (N_193,In_1231,In_444);
nand U194 (N_194,In_342,In_3414);
nand U195 (N_195,In_35,In_4524);
and U196 (N_196,In_2307,In_519);
or U197 (N_197,In_4520,In_4372);
or U198 (N_198,In_2690,In_843);
and U199 (N_199,In_4525,In_2831);
xnor U200 (N_200,In_2737,In_817);
and U201 (N_201,In_3073,In_2167);
or U202 (N_202,In_2219,In_1496);
nand U203 (N_203,In_2077,In_3327);
xnor U204 (N_204,In_4923,In_2021);
nand U205 (N_205,In_4947,In_1714);
nand U206 (N_206,In_1642,In_930);
xor U207 (N_207,In_4542,In_19);
or U208 (N_208,In_1845,In_4346);
nand U209 (N_209,In_4956,In_1036);
xnor U210 (N_210,In_4990,In_4453);
xnor U211 (N_211,In_462,In_164);
or U212 (N_212,In_759,In_1292);
or U213 (N_213,In_1890,In_2670);
nor U214 (N_214,In_1190,In_3798);
and U215 (N_215,In_2404,In_1450);
nor U216 (N_216,In_1189,In_2222);
or U217 (N_217,In_4974,In_2547);
or U218 (N_218,In_4749,In_3500);
nor U219 (N_219,In_2421,In_4583);
xnor U220 (N_220,In_1835,In_3467);
and U221 (N_221,In_3824,In_3876);
and U222 (N_222,In_2723,In_1258);
and U223 (N_223,In_796,In_1380);
xor U224 (N_224,In_793,In_3173);
or U225 (N_225,In_2051,In_3615);
and U226 (N_226,In_1307,In_479);
or U227 (N_227,In_3569,In_812);
nor U228 (N_228,In_294,In_1856);
nand U229 (N_229,In_4744,In_4807);
xnor U230 (N_230,In_1484,In_4532);
or U231 (N_231,In_4217,In_3808);
or U232 (N_232,In_254,In_471);
and U233 (N_233,In_2298,In_4781);
nor U234 (N_234,In_153,In_137);
or U235 (N_235,In_2560,In_2226);
or U236 (N_236,In_4811,In_74);
xor U237 (N_237,In_1913,In_1784);
nor U238 (N_238,In_1681,In_1800);
or U239 (N_239,In_3992,In_4283);
or U240 (N_240,In_1325,In_3016);
nand U241 (N_241,In_1719,In_328);
xor U242 (N_242,In_1425,In_3215);
nor U243 (N_243,In_2482,In_2497);
nand U244 (N_244,In_3058,In_752);
xnor U245 (N_245,In_1558,In_4051);
nand U246 (N_246,In_3873,In_1995);
nor U247 (N_247,In_3216,In_2995);
xnor U248 (N_248,In_3667,In_2502);
nand U249 (N_249,In_4602,In_4438);
nand U250 (N_250,In_4215,In_677);
nand U251 (N_251,In_4363,In_743);
xor U252 (N_252,In_3877,In_2287);
nor U253 (N_253,In_1244,In_4765);
and U254 (N_254,In_2522,In_725);
xnor U255 (N_255,In_1879,In_4871);
or U256 (N_256,In_2947,In_4834);
and U257 (N_257,In_3271,In_1703);
xnor U258 (N_258,In_3828,In_3647);
or U259 (N_259,In_3430,In_2667);
xor U260 (N_260,In_4086,In_2525);
nor U261 (N_261,In_1059,In_3140);
nand U262 (N_262,In_4312,In_4963);
nor U263 (N_263,In_2235,In_3214);
or U264 (N_264,In_3041,In_9);
or U265 (N_265,In_3446,In_4550);
or U266 (N_266,In_4543,In_1014);
nor U267 (N_267,In_1550,In_4848);
nor U268 (N_268,In_3780,In_2999);
and U269 (N_269,In_3546,In_3475);
xor U270 (N_270,In_2513,In_3920);
nand U271 (N_271,In_55,In_581);
and U272 (N_272,In_2706,In_1647);
and U273 (N_273,In_1485,In_158);
or U274 (N_274,In_3782,In_1338);
xor U275 (N_275,In_1376,In_4561);
and U276 (N_276,In_176,In_3580);
nand U277 (N_277,In_4667,In_512);
nand U278 (N_278,In_3366,In_3492);
nand U279 (N_279,In_2479,In_400);
xnor U280 (N_280,In_1950,In_3027);
and U281 (N_281,In_2184,In_2162);
nand U282 (N_282,In_1985,In_2982);
nor U283 (N_283,In_1175,In_4873);
nor U284 (N_284,In_865,In_981);
xnor U285 (N_285,In_3845,In_1104);
nand U286 (N_286,In_3627,In_233);
xnor U287 (N_287,In_3129,In_630);
or U288 (N_288,In_1546,In_3515);
xnor U289 (N_289,In_2925,In_4314);
or U290 (N_290,In_2895,In_509);
or U291 (N_291,In_3263,In_2860);
nand U292 (N_292,In_1115,In_3048);
nand U293 (N_293,In_3772,In_2799);
xor U294 (N_294,In_4914,In_1404);
nor U295 (N_295,In_4991,In_1176);
xnor U296 (N_296,In_4685,In_2114);
nand U297 (N_297,In_80,In_3266);
and U298 (N_298,In_3208,In_2662);
or U299 (N_299,In_3275,In_452);
or U300 (N_300,In_2372,In_2927);
nand U301 (N_301,In_1902,In_1168);
xor U302 (N_302,In_1643,In_4386);
and U303 (N_303,In_1531,In_1288);
nor U304 (N_304,In_3738,In_2890);
or U305 (N_305,In_4747,In_1955);
or U306 (N_306,In_4299,In_4806);
xnor U307 (N_307,In_1458,In_2282);
nor U308 (N_308,In_769,In_3278);
or U309 (N_309,In_138,In_1147);
nand U310 (N_310,In_3953,In_652);
xnor U311 (N_311,In_20,In_1362);
and U312 (N_312,In_627,In_3349);
nand U313 (N_313,In_825,In_4272);
xor U314 (N_314,In_2255,In_3516);
and U315 (N_315,In_3766,In_2239);
and U316 (N_316,In_341,In_460);
nand U317 (N_317,In_2906,In_405);
xnor U318 (N_318,In_177,In_3671);
nand U319 (N_319,In_1841,In_1783);
or U320 (N_320,In_1808,In_411);
xnor U321 (N_321,In_3526,In_4464);
nor U322 (N_322,In_3662,In_3408);
nor U323 (N_323,In_2936,In_1068);
nor U324 (N_324,In_3141,In_4995);
nor U325 (N_325,In_1944,In_1785);
or U326 (N_326,In_1529,In_3871);
nand U327 (N_327,In_3632,In_871);
xor U328 (N_328,In_3814,In_4306);
and U329 (N_329,In_36,In_139);
or U330 (N_330,In_4623,In_4946);
nor U331 (N_331,In_746,In_885);
nand U332 (N_332,In_1474,In_1028);
or U333 (N_333,In_2859,In_1655);
nor U334 (N_334,In_1113,In_1992);
or U335 (N_335,In_4098,In_268);
or U336 (N_336,In_4717,In_4596);
nand U337 (N_337,In_454,In_1121);
nor U338 (N_338,In_3380,In_505);
and U339 (N_339,In_4905,In_347);
or U340 (N_340,In_596,In_2258);
or U341 (N_341,In_53,In_1343);
nor U342 (N_342,In_2873,In_1462);
or U343 (N_343,In_2683,In_2935);
and U344 (N_344,In_2833,In_3945);
xnor U345 (N_345,In_665,In_2840);
nand U346 (N_346,In_2464,In_2841);
xor U347 (N_347,In_3923,In_4156);
nand U348 (N_348,In_763,In_712);
nand U349 (N_349,In_3544,In_1871);
or U350 (N_350,In_4752,In_155);
xor U351 (N_351,In_1917,In_2382);
nor U352 (N_352,In_2818,In_709);
and U353 (N_353,In_741,In_1699);
xor U354 (N_354,In_4929,In_3184);
nor U355 (N_355,In_4353,In_1998);
xnor U356 (N_356,In_803,In_942);
and U357 (N_357,In_2274,In_1154);
nand U358 (N_358,In_605,In_950);
and U359 (N_359,In_3833,In_3748);
nand U360 (N_360,In_4860,In_2637);
or U361 (N_361,In_3363,In_1665);
or U362 (N_362,In_4135,In_640);
or U363 (N_363,In_4218,In_3668);
nor U364 (N_364,In_1668,In_4279);
and U365 (N_365,In_1486,In_4230);
xor U366 (N_366,In_4506,In_3009);
xor U367 (N_367,In_3350,In_3686);
xnor U368 (N_368,In_474,In_2153);
or U369 (N_369,In_245,In_4336);
nor U370 (N_370,In_1878,In_3166);
or U371 (N_371,In_4113,In_210);
nand U372 (N_372,In_4096,In_2904);
xor U373 (N_373,In_2941,In_3223);
or U374 (N_374,In_2791,In_1040);
or U375 (N_375,In_1796,In_4388);
nand U376 (N_376,In_1858,In_4786);
nand U377 (N_377,In_4504,In_1097);
nand U378 (N_378,In_4519,In_445);
nand U379 (N_379,In_92,In_557);
nor U380 (N_380,In_2682,In_2804);
and U381 (N_381,In_4039,In_1911);
nor U382 (N_382,In_2106,In_3743);
nand U383 (N_383,In_3389,In_2284);
nand U384 (N_384,In_3752,In_3061);
nand U385 (N_385,In_810,In_2821);
xor U386 (N_386,In_1772,In_2086);
or U387 (N_387,In_3669,In_700);
xnor U388 (N_388,In_2487,In_1144);
nand U389 (N_389,In_2078,In_3617);
and U390 (N_390,In_3570,In_3202);
and U391 (N_391,In_1286,In_2558);
or U392 (N_392,In_3860,In_1063);
xnor U393 (N_393,In_1527,In_4433);
nor U394 (N_394,In_4494,In_2658);
xnor U395 (N_395,In_4907,In_3853);
nand U396 (N_396,In_248,In_1920);
xor U397 (N_397,In_2237,In_1523);
and U398 (N_398,In_3284,In_2292);
xnor U399 (N_399,In_4637,In_2322);
and U400 (N_400,In_3264,In_928);
nor U401 (N_401,In_4821,In_4687);
nand U402 (N_402,In_4791,In_2686);
nand U403 (N_403,In_4145,In_104);
xnor U404 (N_404,In_2620,In_3189);
nor U405 (N_405,In_2913,In_4622);
nor U406 (N_406,In_2344,In_1356);
or U407 (N_407,In_4800,In_1322);
or U408 (N_408,In_4138,In_3585);
nand U409 (N_409,In_2953,In_87);
xor U410 (N_410,In_869,In_2900);
xor U411 (N_411,In_2026,In_4264);
nand U412 (N_412,In_1249,In_3325);
or U413 (N_413,In_1415,In_893);
and U414 (N_414,In_4112,In_4951);
or U415 (N_415,In_458,In_1396);
nand U416 (N_416,In_2411,In_1666);
and U417 (N_417,In_762,In_3117);
or U418 (N_418,In_2606,In_260);
and U419 (N_419,In_4253,In_4944);
xor U420 (N_420,In_3300,In_2349);
xor U421 (N_421,In_1567,In_2592);
xnor U422 (N_422,In_4676,In_4323);
nand U423 (N_423,In_3967,In_4549);
nor U424 (N_424,In_597,In_767);
or U425 (N_425,In_2262,In_2265);
and U426 (N_426,In_170,In_3153);
xor U427 (N_427,In_561,In_3392);
or U428 (N_428,In_1015,In_784);
and U429 (N_429,In_2289,In_2260);
or U430 (N_430,In_1441,In_2364);
or U431 (N_431,In_2150,In_3056);
and U432 (N_432,In_4088,In_1449);
nor U433 (N_433,In_2109,In_2648);
or U434 (N_434,In_288,In_1795);
nor U435 (N_435,In_3513,In_4630);
xor U436 (N_436,In_112,In_525);
and U437 (N_437,In_3311,In_2444);
xor U438 (N_438,In_2422,In_4456);
or U439 (N_439,In_2694,In_3040);
nor U440 (N_440,In_83,In_2952);
or U441 (N_441,In_1374,In_2993);
xor U442 (N_442,In_1424,In_2766);
or U443 (N_443,In_3991,In_3396);
xor U444 (N_444,In_3037,In_3790);
or U445 (N_445,In_4589,In_4026);
xor U446 (N_446,In_4416,In_3948);
nor U447 (N_447,In_3405,In_4421);
nor U448 (N_448,In_184,In_2656);
nor U449 (N_449,In_256,In_2075);
xor U450 (N_450,In_2393,In_3966);
or U451 (N_451,In_4572,In_1733);
nand U452 (N_452,In_1582,In_4942);
and U453 (N_453,In_2379,In_3946);
or U454 (N_454,In_2201,In_4566);
or U455 (N_455,In_3463,In_4072);
xnor U456 (N_456,In_4377,In_3793);
or U457 (N_457,In_3012,In_2008);
nor U458 (N_458,In_2099,In_78);
nand U459 (N_459,In_1822,In_1639);
nor U460 (N_460,In_162,In_1219);
xor U461 (N_461,In_3224,In_3113);
xnor U462 (N_462,In_2549,In_4);
xor U463 (N_463,In_1085,In_2911);
or U464 (N_464,In_3710,In_4627);
nor U465 (N_465,In_1629,In_3100);
nor U466 (N_466,In_3721,In_3109);
nand U467 (N_467,In_766,In_2189);
or U468 (N_468,In_2198,In_4426);
nand U469 (N_469,In_2710,In_1498);
nand U470 (N_470,In_2050,In_4867);
nor U471 (N_471,In_1866,In_3552);
or U472 (N_472,In_539,In_3362);
nand U473 (N_473,In_4678,In_4318);
xnor U474 (N_474,In_2049,In_4317);
xor U475 (N_475,In_1533,In_593);
nand U476 (N_476,In_4173,In_604);
xnor U477 (N_477,In_2825,In_1152);
or U478 (N_478,In_4521,In_1973);
or U479 (N_479,In_3155,In_1522);
and U480 (N_480,In_2852,In_3785);
nand U481 (N_481,In_2148,In_266);
or U482 (N_482,In_3950,In_1948);
nand U483 (N_483,In_3361,In_1438);
nor U484 (N_484,In_4403,In_3218);
nand U485 (N_485,In_2363,In_2905);
nand U486 (N_486,In_1770,In_1626);
nand U487 (N_487,In_1598,In_4919);
nor U488 (N_488,In_2533,In_1744);
nor U489 (N_489,In_1826,In_7);
nand U490 (N_490,In_4420,In_2073);
or U491 (N_491,In_1538,In_90);
or U492 (N_492,In_1539,In_2717);
or U493 (N_493,In_3182,In_2672);
or U494 (N_494,In_1101,In_4001);
nand U495 (N_495,In_4672,In_2888);
nor U496 (N_496,In_4023,In_999);
nor U497 (N_497,In_4084,In_996);
nand U498 (N_498,In_4772,In_3096);
xor U499 (N_499,In_3545,In_1815);
and U500 (N_500,In_159,In_2197);
xor U501 (N_501,In_892,In_3384);
and U502 (N_502,In_2003,In_602);
nor U503 (N_503,In_152,In_941);
or U504 (N_504,In_608,In_4599);
and U505 (N_505,In_3586,In_3448);
xnor U506 (N_506,In_410,In_2651);
nor U507 (N_507,In_3912,In_4239);
and U508 (N_508,In_2622,In_4977);
nor U509 (N_509,In_3789,In_1968);
nor U510 (N_510,In_1187,In_3712);
nor U511 (N_511,In_929,In_4492);
and U512 (N_512,In_472,In_2402);
nand U513 (N_513,In_174,In_3604);
and U514 (N_514,In_2335,In_635);
xnor U515 (N_515,In_3763,In_2849);
and U516 (N_516,In_4171,In_4835);
nor U517 (N_517,In_1280,In_2111);
nand U518 (N_518,In_3588,In_4817);
and U519 (N_519,In_821,In_3149);
and U520 (N_520,In_2832,In_2959);
and U521 (N_521,In_1174,In_943);
xnor U522 (N_522,In_413,In_2640);
nor U523 (N_523,In_2347,In_3067);
nand U524 (N_524,In_1319,In_4111);
nor U525 (N_525,In_229,In_1403);
xnor U526 (N_526,In_2745,In_3690);
nor U527 (N_527,In_1277,In_598);
xor U528 (N_528,In_987,In_4771);
and U529 (N_529,In_3741,In_4155);
nor U530 (N_530,In_1630,In_4151);
nand U531 (N_531,In_3846,In_2509);
nor U532 (N_532,In_3815,In_1042);
xnor U533 (N_533,In_4537,In_82);
nand U534 (N_534,In_590,In_4646);
and U535 (N_535,In_1662,In_4357);
and U536 (N_536,In_250,In_1517);
and U537 (N_537,In_1956,In_236);
nand U538 (N_538,In_1620,In_3101);
or U539 (N_539,In_3986,In_2196);
nor U540 (N_540,In_952,In_2782);
nand U541 (N_541,In_1224,In_1621);
and U542 (N_542,In_977,In_1262);
xor U543 (N_543,In_3479,In_1969);
or U544 (N_544,In_332,In_3114);
or U545 (N_545,In_3029,In_1300);
xor U546 (N_546,In_3377,In_2418);
nor U547 (N_547,In_1525,In_4267);
nand U548 (N_548,In_4198,In_690);
and U549 (N_549,In_4592,In_1480);
xnor U550 (N_550,In_3769,In_1252);
nand U551 (N_551,In_2361,In_4802);
nand U552 (N_552,In_1873,In_2843);
nand U553 (N_553,In_205,In_226);
and U554 (N_554,In_1809,In_2676);
or U555 (N_555,In_1907,In_2370);
or U556 (N_556,In_1811,In_232);
xor U557 (N_557,In_4531,In_754);
nand U558 (N_558,In_4756,In_1667);
and U559 (N_559,In_4020,In_3021);
xnor U560 (N_560,In_2876,In_4585);
nand U561 (N_561,In_308,In_985);
xor U562 (N_562,In_523,In_3576);
xor U563 (N_563,In_4723,In_895);
xor U564 (N_564,In_4657,In_584);
nand U565 (N_565,In_1454,In_4105);
and U566 (N_566,In_391,In_4983);
or U567 (N_567,In_1436,In_1927);
nor U568 (N_568,In_1904,In_1588);
or U569 (N_569,In_501,In_4329);
and U570 (N_570,In_2854,In_123);
or U571 (N_571,In_622,In_839);
xor U572 (N_572,In_2714,In_3571);
nand U573 (N_573,In_3730,In_842);
and U574 (N_574,In_4052,In_662);
nand U575 (N_575,In_503,In_2748);
xnor U576 (N_576,In_2664,In_4808);
and U577 (N_577,In_3167,In_2115);
or U578 (N_578,In_661,In_4484);
and U579 (N_579,In_4733,In_2132);
and U580 (N_580,In_133,In_3982);
and U581 (N_581,In_4066,In_2338);
or U582 (N_582,In_4294,In_2407);
or U583 (N_583,In_1716,In_4460);
nand U584 (N_584,In_4936,In_4949);
or U585 (N_585,In_4064,In_2847);
nor U586 (N_586,In_4540,In_4882);
nand U587 (N_587,In_2467,In_917);
nand U588 (N_588,In_419,In_4188);
xnor U589 (N_589,In_317,In_1754);
xnor U590 (N_590,In_3447,In_1358);
xor U591 (N_591,In_1599,In_2312);
and U592 (N_592,In_3075,In_772);
and U593 (N_593,In_897,In_3242);
or U594 (N_594,In_1225,In_923);
or U595 (N_595,In_1885,In_2004);
or U596 (N_596,In_3504,In_621);
nor U597 (N_597,In_4796,In_2211);
nand U598 (N_598,In_522,In_4612);
nand U599 (N_599,In_2853,In_3136);
nor U600 (N_600,In_3599,In_2517);
or U601 (N_601,In_4780,In_2587);
or U602 (N_602,In_3120,In_1912);
nor U603 (N_603,In_4679,In_2414);
nand U604 (N_604,In_3882,In_4168);
xor U605 (N_605,In_4122,In_2998);
nor U606 (N_606,In_4074,In_4236);
or U607 (N_607,In_3403,In_2346);
nor U608 (N_608,In_4933,In_3255);
nor U609 (N_609,In_2623,In_1958);
and U610 (N_610,In_130,In_555);
and U611 (N_611,In_4159,In_1934);
nor U612 (N_612,In_2562,In_3965);
or U613 (N_613,In_475,In_60);
nand U614 (N_614,In_4387,In_4289);
or U615 (N_615,In_439,In_2425);
nand U616 (N_616,In_3154,In_3205);
or U617 (N_617,In_2958,In_1316);
and U618 (N_618,In_358,In_4883);
nor U619 (N_619,In_2801,In_4163);
nand U620 (N_620,In_3919,In_4730);
nor U621 (N_621,In_4706,In_1710);
or U622 (N_622,In_4276,In_1595);
xnor U623 (N_623,In_4245,In_4174);
and U624 (N_624,In_696,In_3104);
or U625 (N_625,In_1431,In_3402);
xnor U626 (N_626,In_2877,In_3934);
xnor U627 (N_627,In_3883,In_2091);
xnor U628 (N_628,In_4439,In_538);
nor U629 (N_629,In_1711,In_1818);
and U630 (N_630,In_1670,In_4988);
xnor U631 (N_631,In_2009,In_4099);
xor U632 (N_632,In_1704,In_535);
and U633 (N_633,In_599,In_4610);
xor U634 (N_634,In_3908,In_2705);
nand U635 (N_635,In_3547,In_1750);
and U636 (N_636,In_4459,In_4901);
and U637 (N_637,In_1730,In_2496);
or U638 (N_638,In_1854,In_2977);
xnor U639 (N_639,In_404,In_1964);
nor U640 (N_640,In_13,In_3283);
or U641 (N_641,In_2518,In_3);
xor U642 (N_642,In_1335,In_1981);
nand U643 (N_643,In_1823,In_4021);
and U644 (N_644,In_4553,In_2572);
and U645 (N_645,In_4311,In_3653);
and U646 (N_646,In_3413,In_1576);
nand U647 (N_647,In_2535,In_1401);
nor U648 (N_648,In_708,In_1257);
and U649 (N_649,In_4594,In_880);
or U650 (N_650,In_4255,In_1184);
xor U651 (N_651,In_267,In_2458);
or U652 (N_652,In_77,In_4162);
nor U653 (N_653,In_962,In_1740);
and U654 (N_654,In_3193,In_4164);
or U655 (N_655,In_3225,In_2308);
nor U656 (N_656,In_4282,In_4981);
nand U657 (N_657,In_3974,In_1832);
nor U658 (N_658,In_888,In_88);
and U659 (N_659,In_1398,In_4645);
and U660 (N_660,In_110,In_1136);
xor U661 (N_661,In_3353,In_1299);
nor U662 (N_662,In_3737,In_4569);
nor U663 (N_663,In_4197,In_2383);
xnor U664 (N_664,In_3145,In_4056);
and U665 (N_665,In_4079,In_63);
nand U666 (N_666,In_830,In_3566);
nand U667 (N_667,In_2139,In_4024);
and U668 (N_668,In_3091,In_3497);
xor U669 (N_669,In_1888,In_2910);
and U670 (N_670,In_325,In_4568);
nand U671 (N_671,In_251,In_3245);
or U672 (N_672,In_1248,In_886);
nand U673 (N_673,In_3826,In_805);
xor U674 (N_674,In_38,In_617);
xor U675 (N_675,In_2028,In_2309);
or U676 (N_676,In_1411,In_6);
and U677 (N_677,In_2126,In_883);
nand U678 (N_678,In_4342,In_2420);
nand U679 (N_679,In_4037,In_1891);
and U680 (N_680,In_4334,In_633);
or U681 (N_681,In_3063,In_24);
xnor U682 (N_682,In_64,In_436);
and U683 (N_683,In_2490,In_2744);
nand U684 (N_684,In_1095,In_2750);
or U685 (N_685,In_4252,In_4476);
xor U686 (N_686,In_813,In_3340);
nand U687 (N_687,In_3285,In_1058);
nor U688 (N_688,In_2159,In_714);
and U689 (N_689,In_579,In_1451);
or U690 (N_690,In_1607,In_904);
xor U691 (N_691,In_1725,In_3521);
nor U692 (N_692,In_1385,In_3438);
and U693 (N_693,In_2565,In_684);
nand U694 (N_694,In_1440,In_2678);
or U695 (N_695,In_729,In_3115);
or U696 (N_696,In_4616,In_1455);
and U697 (N_697,In_2006,In_1392);
and U698 (N_698,In_4838,In_1182);
and U699 (N_699,In_96,In_408);
nor U700 (N_700,In_2769,In_3484);
and U701 (N_701,In_443,In_3527);
or U702 (N_702,In_3942,In_371);
nand U703 (N_703,In_417,In_1264);
nand U704 (N_704,In_4012,In_4186);
or U705 (N_705,In_3695,In_4577);
nor U706 (N_706,In_1221,In_146);
nor U707 (N_707,In_299,In_4841);
xor U708 (N_708,In_3057,In_4398);
or U709 (N_709,In_4114,In_4031);
xnor U710 (N_710,In_129,In_4033);
and U711 (N_711,In_2824,In_4582);
and U712 (N_712,In_119,In_4804);
or U713 (N_713,In_1671,In_2253);
or U714 (N_714,In_1406,In_3537);
xor U715 (N_715,In_1243,In_2495);
or U716 (N_716,In_2380,In_2391);
xnor U717 (N_717,In_2220,In_1916);
nor U718 (N_718,In_2862,In_97);
nor U719 (N_719,In_4063,In_4992);
xor U720 (N_720,In_3162,In_788);
xnor U721 (N_721,In_2455,In_1077);
nand U722 (N_722,In_2229,In_2128);
and U723 (N_723,In_4243,In_3518);
or U724 (N_724,In_1999,In_1207);
or U725 (N_725,In_4716,In_4083);
xor U726 (N_726,In_2283,In_925);
nor U727 (N_727,In_748,In_3330);
and U728 (N_728,In_4002,In_3993);
nor U729 (N_729,In_945,In_1218);
or U730 (N_730,In_3290,In_1137);
or U731 (N_731,In_2469,In_882);
xnor U732 (N_732,In_4040,In_2011);
nor U733 (N_733,In_40,In_1373);
xor U734 (N_734,In_1978,In_183);
or U735 (N_735,In_3391,In_699);
nand U736 (N_736,In_4350,In_4671);
nor U737 (N_737,In_1357,In_4256);
nor U738 (N_738,In_2807,In_148);
nor U739 (N_739,In_2398,In_1256);
or U740 (N_740,In_434,In_3273);
and U741 (N_741,In_4890,In_969);
nand U742 (N_742,In_1022,In_258);
nand U743 (N_743,In_1573,In_1156);
nor U744 (N_744,In_4560,In_2423);
xnor U745 (N_745,In_3797,In_259);
or U746 (N_746,In_4641,In_3800);
and U747 (N_747,In_4604,In_1035);
nor U748 (N_748,In_3806,In_4880);
nand U749 (N_749,In_992,In_4465);
and U750 (N_750,In_4120,In_2321);
or U751 (N_751,In_2147,In_643);
nor U752 (N_752,In_4286,In_2204);
xor U753 (N_753,In_281,In_4918);
nor U754 (N_754,In_1163,In_4068);
or U755 (N_755,In_965,In_4681);
xor U756 (N_756,In_4986,In_2588);
or U757 (N_757,In_4104,In_3068);
and U758 (N_758,In_468,In_1752);
and U759 (N_759,In_2250,In_2005);
nor U760 (N_760,In_422,In_3042);
and U761 (N_761,In_2100,In_2523);
xnor U762 (N_762,In_1416,In_2409);
nand U763 (N_763,In_1773,In_2626);
or U764 (N_764,In_2316,In_782);
xnor U765 (N_765,In_1370,In_4389);
nor U766 (N_766,In_2921,In_4310);
xor U767 (N_767,In_3036,In_75);
or U768 (N_768,In_1170,In_1734);
nand U769 (N_769,In_1861,In_2792);
nand U770 (N_770,In_2311,In_323);
nor U771 (N_771,In_2770,In_2631);
or U772 (N_772,In_2352,In_4515);
xor U773 (N_773,In_3280,In_2720);
or U774 (N_774,In_285,In_2046);
and U775 (N_775,In_3319,In_1038);
and U776 (N_776,In_1199,In_3970);
and U777 (N_777,In_140,In_4445);
nor U778 (N_778,In_2908,In_4270);
nor U779 (N_779,In_4461,In_2231);
nor U780 (N_780,In_2874,In_4574);
xnor U781 (N_781,In_1166,In_2528);
nor U782 (N_782,In_1017,In_520);
nand U783 (N_783,In_3926,In_2679);
and U784 (N_784,In_4046,In_1390);
or U785 (N_785,In_3125,In_1507);
nor U786 (N_786,In_1846,In_4866);
xor U787 (N_787,In_4859,In_2081);
nor U788 (N_788,In_2410,In_3652);
nor U789 (N_789,In_2484,In_2154);
nor U790 (N_790,In_1980,In_536);
or U791 (N_791,In_3903,In_854);
or U792 (N_792,In_1606,In_2175);
and U793 (N_793,In_3001,In_3517);
and U794 (N_794,In_2892,In_2546);
xnor U795 (N_795,In_1983,In_3316);
and U796 (N_796,In_4076,In_2343);
nand U797 (N_797,In_204,In_107);
xnor U798 (N_798,In_212,In_1514);
or U799 (N_799,In_1301,In_3809);
nor U800 (N_800,In_2891,In_2406);
xor U801 (N_801,In_921,In_2505);
xor U802 (N_802,In_3076,In_4720);
or U803 (N_803,In_2653,In_780);
nand U804 (N_804,In_1941,In_2582);
or U805 (N_805,In_4315,In_1139);
nor U806 (N_806,In_4769,In_4953);
nand U807 (N_807,In_151,In_1658);
or U808 (N_808,In_809,In_2187);
and U809 (N_809,In_1775,In_182);
nand U810 (N_810,In_1393,In_127);
and U811 (N_811,In_4695,In_993);
or U812 (N_812,In_298,In_3520);
nor U813 (N_813,In_2296,In_1687);
nor U814 (N_814,In_3247,In_679);
nor U815 (N_815,In_4674,In_3969);
xnor U816 (N_816,In_282,In_1747);
nand U817 (N_817,In_720,In_3818);
nor U818 (N_818,In_4128,In_1727);
and U819 (N_819,In_1186,In_4161);
or U820 (N_820,In_1394,In_4964);
or U821 (N_821,In_2314,In_1932);
xor U822 (N_822,In_2436,In_2433);
xor U823 (N_823,In_3562,In_785);
or U824 (N_824,In_858,In_2898);
or U825 (N_825,In_4367,In_2485);
nor U826 (N_826,In_1557,In_3563);
or U827 (N_827,In_2621,In_4062);
nor U828 (N_828,In_4994,In_4495);
and U829 (N_829,In_1580,In_2885);
or U830 (N_830,In_1327,In_2597);
nand U831 (N_831,In_4702,In_2025);
or U832 (N_832,In_145,In_2491);
and U833 (N_833,In_1612,In_1082);
and U834 (N_834,In_2680,In_510);
nand U835 (N_835,In_783,In_3146);
or U836 (N_836,In_4575,In_2145);
nor U837 (N_837,In_2256,In_3975);
nand U838 (N_838,In_933,In_2884);
xor U839 (N_839,In_351,In_1903);
and U840 (N_840,In_4941,In_2340);
nand U841 (N_841,In_956,In_4777);
and U842 (N_842,In_3460,In_1864);
xnor U843 (N_843,In_3185,In_1060);
nand U844 (N_844,In_1192,In_2654);
nor U845 (N_845,In_4738,In_948);
xor U846 (N_846,In_4330,In_1475);
nor U847 (N_847,In_3138,In_3419);
nand U848 (N_848,In_1081,In_243);
and U849 (N_849,In_4284,In_311);
nor U850 (N_850,In_2324,In_3770);
nor U851 (N_851,In_249,In_1408);
and U852 (N_852,In_3174,In_1064);
nor U853 (N_853,In_1816,In_3444);
or U854 (N_854,In_3191,In_4648);
xnor U855 (N_855,In_1326,In_3246);
and U856 (N_856,In_1078,In_828);
nand U857 (N_857,In_3746,In_1304);
nand U858 (N_858,In_3979,In_2541);
or U859 (N_859,In_2815,In_844);
xnor U860 (N_860,In_0,In_2007);
and U861 (N_861,In_48,In_4424);
nand U862 (N_862,In_4544,In_2971);
xnor U863 (N_863,In_3306,In_4595);
or U864 (N_864,In_3675,In_1245);
nor U865 (N_865,In_4381,In_4663);
xor U866 (N_866,In_4996,In_2761);
nor U867 (N_867,In_244,In_1287);
and U868 (N_868,In_3898,In_2368);
xnor U869 (N_869,In_3568,In_4191);
nor U870 (N_870,In_3901,In_2944);
and U871 (N_871,In_3794,In_1321);
xnor U872 (N_872,In_1213,In_1021);
xor U873 (N_873,In_3976,In_586);
xor U874 (N_874,In_4957,In_4140);
nand U875 (N_875,In_4661,In_4607);
xnor U876 (N_876,In_3376,In_2447);
nor U877 (N_877,In_1817,In_4927);
nand U878 (N_878,In_4274,In_4551);
nand U879 (N_879,In_275,In_1062);
xnor U880 (N_880,In_428,In_2929);
and U881 (N_881,In_1331,In_2395);
or U882 (N_882,In_1413,In_1571);
or U883 (N_883,In_2756,In_2327);
xor U884 (N_884,In_3879,In_2970);
xnor U885 (N_885,In_1676,In_3229);
nor U886 (N_886,In_3700,In_4509);
or U887 (N_887,In_2094,In_2610);
xor U888 (N_888,In_2700,In_2448);
nor U889 (N_889,In_3176,In_1737);
nor U890 (N_890,In_1359,In_1590);
xnor U891 (N_891,In_3788,In_1602);
nand U892 (N_892,In_2721,In_2983);
nand U893 (N_893,In_2166,In_2930);
nand U894 (N_894,In_4615,In_4879);
nand U895 (N_895,In_2121,In_2827);
nand U896 (N_896,In_1518,In_4968);
nand U897 (N_897,In_1283,In_4199);
and U898 (N_898,In_4382,In_1988);
xnor U899 (N_899,In_564,In_2329);
or U900 (N_900,In_1342,In_1387);
nand U901 (N_901,In_3236,In_3929);
xnor U902 (N_902,In_2954,In_3079);
nor U903 (N_903,In_2339,In_736);
xnor U904 (N_904,In_3677,In_4081);
or U905 (N_905,In_3394,In_2507);
and U906 (N_906,In_3265,In_4467);
xor U907 (N_907,In_4413,In_2104);
or U908 (N_908,In_4268,In_3015);
xor U909 (N_909,In_3222,In_382);
or U910 (N_910,In_3720,In_398);
nor U911 (N_911,In_450,In_2472);
nand U912 (N_912,In_3874,In_2445);
or U913 (N_913,In_3004,In_811);
or U914 (N_914,In_406,In_1881);
and U915 (N_915,In_3804,In_344);
or U916 (N_916,In_4840,In_1332);
nand U917 (N_917,In_2096,In_407);
and U918 (N_918,In_1505,In_2351);
nor U919 (N_919,In_3107,In_264);
and U920 (N_920,In_3610,In_2624);
nor U921 (N_921,In_2924,In_967);
and U922 (N_922,In_1312,In_4961);
or U923 (N_923,In_4689,In_2837);
nor U924 (N_924,In_2468,In_4813);
nor U925 (N_925,In_4345,In_3918);
or U926 (N_926,In_1633,In_3382);
nand U927 (N_927,In_1859,In_2711);
nor U928 (N_928,In_3983,In_4785);
or U929 (N_929,In_101,In_4471);
and U930 (N_930,In_3792,In_2394);
nand U931 (N_931,In_1375,In_4325);
and U932 (N_932,In_3896,In_2986);
and U933 (N_933,In_4045,In_2337);
nor U934 (N_934,In_2746,In_618);
and U935 (N_935,In_1645,In_4394);
or U936 (N_936,In_3594,In_3089);
xor U937 (N_937,In_2598,In_4232);
nor U938 (N_938,In_3631,In_2772);
and U939 (N_939,In_3178,In_3461);
or U940 (N_940,In_3723,In_1002);
xnor U941 (N_941,In_1519,In_3296);
nor U942 (N_942,In_154,In_728);
xor U943 (N_943,In_3889,In_4365);
and U944 (N_944,In_3899,In_2786);
and U945 (N_945,In_1173,In_4593);
nor U946 (N_946,In_3077,In_2299);
and U947 (N_947,In_216,In_911);
or U948 (N_948,In_2511,In_1506);
nor U949 (N_949,In_3234,In_2939);
xor U950 (N_950,In_4436,In_2909);
or U951 (N_951,In_1399,In_2593);
nor U952 (N_952,In_3681,In_2251);
or U953 (N_953,In_3870,In_2180);
nor U954 (N_954,In_4240,In_4843);
nand U955 (N_955,In_3750,In_2817);
xnor U956 (N_956,In_4014,In_4972);
and U957 (N_957,In_3727,In_1627);
xor U958 (N_958,In_2072,In_3452);
nand U959 (N_959,In_2302,In_801);
and U960 (N_960,In_4422,In_2985);
and U961 (N_961,In_3728,In_2160);
nand U962 (N_962,In_2857,In_2514);
and U963 (N_963,In_3698,In_2031);
nor U964 (N_964,In_713,In_1986);
or U965 (N_965,In_2743,In_2297);
nor U966 (N_966,In_3602,In_284);
nor U967 (N_967,In_1466,In_2063);
xnor U968 (N_968,In_4614,In_3474);
nor U969 (N_969,In_4588,In_541);
nor U970 (N_970,In_4153,In_2334);
or U971 (N_971,In_283,In_1657);
or U972 (N_972,In_4906,In_4909);
and U973 (N_973,In_4185,In_698);
nor U974 (N_974,In_3716,In_263);
or U975 (N_975,In_4878,In_4704);
and U976 (N_976,In_4856,In_1282);
nand U977 (N_977,In_4201,In_552);
nand U978 (N_978,In_292,In_4488);
nand U979 (N_979,In_352,In_2538);
xnor U980 (N_980,In_4501,In_1141);
xor U981 (N_981,In_1405,In_1943);
nand U982 (N_982,In_1209,In_3337);
xor U983 (N_983,In_4109,In_497);
or U984 (N_984,In_3747,In_1933);
or U985 (N_985,In_3778,In_3890);
xor U986 (N_986,In_1143,In_3252);
xor U987 (N_987,In_2788,In_3002);
or U988 (N_988,In_2365,In_3219);
and U989 (N_989,In_2453,In_4842);
and U990 (N_990,In_1742,In_540);
nand U991 (N_991,In_1628,In_2629);
xnor U992 (N_992,In_3268,In_4179);
or U993 (N_993,In_3493,In_105);
or U994 (N_994,In_3200,In_1259);
or U995 (N_995,In_1070,In_1235);
or U996 (N_996,In_4379,In_3410);
nand U997 (N_997,In_4212,In_61);
and U998 (N_998,In_293,In_4216);
nor U999 (N_999,In_4828,In_4489);
xnor U1000 (N_1000,In_1908,In_2632);
xor U1001 (N_1001,In_1805,In_2221);
xnor U1002 (N_1002,In_156,In_1320);
xnor U1003 (N_1003,In_4448,In_3608);
xnor U1004 (N_1004,In_2374,In_2636);
nor U1005 (N_1005,In_4510,In_3328);
nand U1006 (N_1006,In_1428,In_574);
xor U1007 (N_1007,In_2760,In_4718);
and U1008 (N_1008,In_4384,In_2836);
and U1009 (N_1009,In_3469,In_2350);
nor U1010 (N_1010,In_4565,In_3365);
nor U1011 (N_1011,In_3276,In_1721);
xor U1012 (N_1012,In_3907,In_1549);
nor U1013 (N_1013,In_4280,In_1018);
xnor U1014 (N_1014,In_2878,In_3672);
nor U1015 (N_1015,In_1692,In_4693);
nand U1016 (N_1016,In_1055,In_1766);
and U1017 (N_1017,In_3584,In_4196);
xor U1018 (N_1018,In_689,In_4713);
or U1019 (N_1019,In_2182,In_3287);
nand U1020 (N_1020,In_3288,In_3972);
nand U1021 (N_1021,In_2992,In_3468);
and U1022 (N_1022,In_208,In_791);
nand U1023 (N_1023,In_2989,In_3168);
nand U1024 (N_1024,In_372,In_542);
or U1025 (N_1025,In_4736,In_98);
or U1026 (N_1026,In_4204,In_2879);
xnor U1027 (N_1027,In_2475,In_106);
nand U1028 (N_1028,In_4847,In_2441);
or U1029 (N_1029,In_1157,In_1290);
nand U1030 (N_1030,In_3130,In_2431);
nand U1031 (N_1031,In_1753,In_1260);
xor U1032 (N_1032,In_3358,In_3416);
nand U1033 (N_1033,In_3956,In_2345);
and U1034 (N_1034,In_1210,In_3888);
nand U1035 (N_1035,In_2079,In_1989);
nand U1036 (N_1036,In_4511,In_178);
or U1037 (N_1037,In_1360,In_3127);
xor U1038 (N_1038,In_2524,In_3062);
xnor U1039 (N_1039,In_1982,In_3342);
nand U1040 (N_1040,In_2933,In_4119);
nor U1041 (N_1041,In_3536,In_2319);
xnor U1042 (N_1042,In_4078,In_2053);
nor U1043 (N_1043,In_738,In_1722);
nand U1044 (N_1044,In_3891,In_4784);
nand U1045 (N_1045,In_2531,In_4763);
nand U1046 (N_1046,In_2556,In_2203);
and U1047 (N_1047,In_955,In_1794);
nand U1048 (N_1048,In_1132,In_2539);
xor U1049 (N_1049,In_4712,In_3742);
xnor U1050 (N_1050,In_261,In_1079);
nor U1051 (N_1051,In_735,In_3614);
and U1052 (N_1052,In_3740,In_1465);
xnor U1053 (N_1053,In_4910,In_4154);
or U1054 (N_1054,In_3626,In_2554);
or U1055 (N_1055,In_3031,In_4670);
and U1056 (N_1056,In_269,In_1114);
and U1057 (N_1057,In_3118,In_1003);
or U1058 (N_1058,In_4288,In_669);
and U1059 (N_1059,In_1251,In_2438);
or U1060 (N_1060,In_1165,In_3994);
nor U1061 (N_1061,In_1696,In_3639);
nor U1062 (N_1062,In_4917,In_368);
and U1063 (N_1063,In_4322,In_2738);
and U1064 (N_1064,In_2568,In_578);
and U1065 (N_1065,In_756,In_3139);
xor U1066 (N_1066,In_963,In_4792);
or U1067 (N_1067,In_4409,In_2320);
nand U1068 (N_1068,In_995,In_1762);
or U1069 (N_1069,In_4721,In_3751);
and U1070 (N_1070,In_744,In_1389);
and U1071 (N_1071,In_3186,In_3250);
nand U1072 (N_1072,In_644,In_2353);
nor U1073 (N_1073,In_4117,In_4851);
xnor U1074 (N_1074,In_1532,In_966);
and U1075 (N_1075,In_166,In_4889);
and U1076 (N_1076,In_1807,In_1608);
nand U1077 (N_1077,In_4458,In_4955);
and U1078 (N_1078,In_2360,In_2493);
and U1079 (N_1079,In_2618,In_1748);
or U1080 (N_1080,In_383,In_252);
nor U1081 (N_1081,In_506,In_3863);
xor U1082 (N_1082,In_1348,In_2097);
and U1083 (N_1083,In_1648,In_2603);
or U1084 (N_1084,In_4858,In_1700);
nand U1085 (N_1085,In_884,In_33);
nor U1086 (N_1086,In_3261,In_270);
nand U1087 (N_1087,In_3098,In_4903);
nor U1088 (N_1088,In_1216,In_300);
and U1089 (N_1089,In_3387,In_3745);
and U1090 (N_1090,In_964,In_2595);
and U1091 (N_1091,In_4452,In_3995);
nand U1092 (N_1092,In_4231,In_4513);
and U1093 (N_1093,In_2557,In_4803);
or U1094 (N_1094,In_3709,In_2784);
nand U1095 (N_1095,In_287,In_879);
and U1096 (N_1096,In_4793,In_1640);
xor U1097 (N_1097,In_4638,In_4997);
xor U1098 (N_1098,In_3641,In_2871);
or U1099 (N_1099,In_4177,In_3049);
nand U1100 (N_1100,In_595,In_3558);
xnor U1101 (N_1101,In_1693,In_4178);
and U1102 (N_1102,In_3999,In_3756);
nor U1103 (N_1103,In_3406,In_2987);
nand U1104 (N_1104,In_660,In_3841);
nand U1105 (N_1105,In_1443,In_545);
xor U1106 (N_1106,In_4481,In_4740);
and U1107 (N_1107,In_1130,In_3642);
nor U1108 (N_1108,In_190,In_3519);
and U1109 (N_1109,In_2170,In_3916);
and U1110 (N_1110,In_4206,In_1202);
nand U1111 (N_1111,In_2781,In_4010);
and U1112 (N_1112,In_775,In_4562);
and U1113 (N_1113,In_639,In_3541);
and U1114 (N_1114,In_1844,In_4130);
nand U1115 (N_1115,In_823,In_1542);
or U1116 (N_1116,In_2117,In_3099);
nor U1117 (N_1117,In_1896,In_1276);
or U1118 (N_1118,In_659,In_2586);
and U1119 (N_1119,In_3308,In_4782);
nand U1120 (N_1120,In_2994,In_742);
or U1121 (N_1121,In_1073,In_4005);
nor U1122 (N_1122,In_1208,In_1432);
xnor U1123 (N_1123,In_3364,In_4635);
xor U1124 (N_1124,In_4754,In_1536);
or U1125 (N_1125,In_2076,In_2794);
nor U1126 (N_1126,In_1634,In_132);
xor U1127 (N_1127,In_4184,In_4830);
and U1128 (N_1128,In_4691,In_3900);
and U1129 (N_1129,In_2955,In_3302);
xor U1130 (N_1130,In_550,In_3133);
and U1131 (N_1131,In_2241,In_804);
and U1132 (N_1132,In_902,In_4984);
xnor U1133 (N_1133,In_2424,In_4881);
nand U1134 (N_1134,In_2034,In_647);
or U1135 (N_1135,In_4044,In_881);
or U1136 (N_1136,In_498,In_3159);
nor U1137 (N_1137,In_2176,In_838);
nor U1138 (N_1138,In_1429,In_2966);
or U1139 (N_1139,In_3620,In_3666);
nand U1140 (N_1140,In_2569,In_3482);
nor U1141 (N_1141,In_1112,In_3998);
nand U1142 (N_1142,In_1268,In_4850);
nand U1143 (N_1143,In_4809,In_2627);
nor U1144 (N_1144,In_2793,In_2195);
or U1145 (N_1145,In_1103,In_3429);
or U1146 (N_1146,In_518,In_4629);
nor U1147 (N_1147,In_473,In_2123);
or U1148 (N_1148,In_2388,In_715);
and U1149 (N_1149,In_3351,In_84);
nand U1150 (N_1150,In_2151,In_4013);
xnor U1151 (N_1151,In_4347,In_4067);
or U1152 (N_1152,In_4434,In_4134);
and U1153 (N_1153,In_2599,In_4998);
xnor U1154 (N_1154,In_887,In_1741);
nor U1155 (N_1155,In_2615,In_1140);
xor U1156 (N_1156,In_4303,In_2127);
nand U1157 (N_1157,In_3355,In_1562);
and U1158 (N_1158,In_2917,In_3635);
nand U1159 (N_1159,In_2205,In_3825);
or U1160 (N_1160,In_1563,In_322);
or U1161 (N_1161,In_1910,In_4029);
nor U1162 (N_1162,In_2734,In_32);
nand U1163 (N_1163,In_4292,In_3415);
or U1164 (N_1164,In_4034,In_465);
xor U1165 (N_1165,In_951,In_990);
nor U1166 (N_1166,In_2359,In_1685);
or U1167 (N_1167,In_2371,In_570);
or U1168 (N_1168,In_1247,In_2886);
nor U1169 (N_1169,In_1852,In_1698);
and U1170 (N_1170,In_2171,In_3344);
xnor U1171 (N_1171,In_612,In_3111);
nand U1172 (N_1172,In_1738,In_4483);
nor U1173 (N_1173,In_820,In_3550);
nand U1174 (N_1174,In_3834,In_2238);
or U1175 (N_1175,In_3603,In_947);
nand U1176 (N_1176,In_4103,In_4443);
and U1177 (N_1177,In_1254,In_4227);
or U1178 (N_1178,In_1976,In_841);
and U1179 (N_1179,In_1691,In_409);
and U1180 (N_1180,In_2732,In_4141);
or U1181 (N_1181,In_3449,In_916);
or U1182 (N_1182,In_1402,In_1979);
nor U1183 (N_1183,In_936,In_958);
and U1184 (N_1184,In_4077,In_3719);
and U1185 (N_1185,In_2881,In_4190);
nor U1186 (N_1186,In_2015,In_4597);
or U1187 (N_1187,In_2742,In_3606);
and U1188 (N_1188,In_778,In_4535);
and U1189 (N_1189,In_978,In_3930);
xnor U1190 (N_1190,In_3209,In_3996);
and U1191 (N_1191,In_706,In_4533);
or U1192 (N_1192,In_4655,In_1011);
xnor U1193 (N_1193,In_1020,In_59);
xor U1194 (N_1194,In_2974,In_1914);
xnor U1195 (N_1195,In_1528,In_723);
nor U1196 (N_1196,In_2301,In_2067);
nand U1197 (N_1197,In_528,In_3680);
and U1198 (N_1198,In_1092,In_502);
or U1199 (N_1199,In_3925,In_3322);
nand U1200 (N_1200,In_4563,In_3861);
nand U1201 (N_1201,In_3702,In_3583);
xnor U1202 (N_1202,In_4472,In_1499);
xor U1203 (N_1203,In_2013,In_1876);
xor U1204 (N_1204,In_4857,In_187);
or U1205 (N_1205,In_426,In_2155);
and U1206 (N_1206,In_193,In_4429);
and U1207 (N_1207,In_4665,In_3754);
nor U1208 (N_1208,In_4320,In_3239);
xor U1209 (N_1209,In_4741,In_2056);
xor U1210 (N_1210,In_932,In_4223);
nor U1211 (N_1211,In_716,In_3638);
and U1212 (N_1212,In_2277,In_1530);
xor U1213 (N_1213,In_3071,In_2778);
or U1214 (N_1214,In_3170,In_4608);
xor U1215 (N_1215,In_4257,In_4390);
xor U1216 (N_1216,In_3335,In_1712);
nand U1217 (N_1217,In_1371,In_280);
or U1218 (N_1218,In_1294,In_4969);
xnor U1219 (N_1219,In_2305,In_4653);
xnor U1220 (N_1220,In_1310,In_1768);
nor U1221 (N_1221,In_527,In_3478);
xnor U1222 (N_1222,In_1583,In_329);
and U1223 (N_1223,In_2405,In_872);
and U1224 (N_1224,In_1729,In_3997);
xnor U1225 (N_1225,In_547,In_961);
xor U1226 (N_1226,In_611,In_2579);
xor U1227 (N_1227,In_556,In_4516);
or U1228 (N_1228,In_1942,In_4370);
xor U1229 (N_1229,In_982,In_1965);
nor U1230 (N_1230,In_2577,In_1071);
xnor U1231 (N_1231,In_3459,In_296);
and U1232 (N_1232,In_1400,In_3323);
nor U1233 (N_1233,In_4814,In_711);
nand U1234 (N_1234,In_832,In_2948);
xor U1235 (N_1235,In_2055,In_4943);
xor U1236 (N_1236,In_863,In_3981);
nor U1237 (N_1237,In_3274,In_2161);
and U1238 (N_1238,In_3636,In_1592);
and U1239 (N_1239,In_954,In_1637);
and U1240 (N_1240,In_1472,In_421);
nand U1241 (N_1241,In_1476,In_362);
xnor U1242 (N_1242,In_802,In_4259);
and U1243 (N_1243,In_4450,In_4869);
nor U1244 (N_1244,In_3988,In_2731);
xor U1245 (N_1245,In_1056,In_2604);
nor U1246 (N_1246,In_4987,In_1609);
and U1247 (N_1247,In_3807,In_3445);
and U1248 (N_1248,In_214,In_4896);
and U1249 (N_1249,In_4208,In_3674);
or U1250 (N_1250,In_2691,In_2789);
nor U1251 (N_1251,In_1545,In_1723);
or U1252 (N_1252,In_3629,In_4517);
nand U1253 (N_1253,In_3984,In_1368);
nand U1254 (N_1254,In_1250,In_2730);
or U1255 (N_1255,In_2829,In_2280);
nor U1256 (N_1256,In_3673,In_1745);
and U1257 (N_1257,In_3548,In_425);
or U1258 (N_1258,In_4924,In_2661);
and U1259 (N_1259,In_3210,In_2997);
xor U1260 (N_1260,In_4262,In_4989);
or U1261 (N_1261,In_2225,In_2960);
and U1262 (N_1262,In_1521,In_1720);
nand U1263 (N_1263,In_2697,In_4688);
and U1264 (N_1264,In_3607,In_3436);
or U1265 (N_1265,In_4121,In_3658);
and U1266 (N_1266,In_2300,In_3755);
and U1267 (N_1267,In_1502,In_4351);
xor U1268 (N_1268,In_1452,In_195);
xnor U1269 (N_1269,In_2926,In_2157);
and U1270 (N_1270,In_3411,In_2589);
nor U1271 (N_1271,In_2848,In_1162);
nand U1272 (N_1272,In_3332,In_4794);
nand U1273 (N_1273,In_3026,In_3279);
nand U1274 (N_1274,In_1949,In_1570);
xor U1275 (N_1275,In_306,In_4902);
nor U1276 (N_1276,In_2961,In_4985);
and U1277 (N_1277,In_4220,In_2186);
nand U1278 (N_1278,In_4348,In_4639);
nand U1279 (N_1279,In_3987,In_681);
and U1280 (N_1280,In_3501,In_4502);
nor U1281 (N_1281,In_1054,In_365);
and U1282 (N_1282,In_1825,In_991);
and U1283 (N_1283,In_657,In_4441);
or U1284 (N_1284,In_4609,In_3313);
xor U1285 (N_1285,In_4503,In_2027);
nand U1286 (N_1286,In_4898,In_3508);
nand U1287 (N_1287,In_3230,In_430);
nor U1288 (N_1288,In_4451,In_4361);
nor U1289 (N_1289,In_2268,In_3892);
nand U1290 (N_1290,In_3851,In_2396);
and U1291 (N_1291,In_2143,In_2138);
nor U1292 (N_1292,In_3134,In_4339);
or U1293 (N_1293,In_4326,In_3347);
and U1294 (N_1294,In_1673,In_4278);
nor U1295 (N_1295,In_4296,In_3688);
xnor U1296 (N_1296,In_3110,In_4374);
xnor U1297 (N_1297,In_3069,In_642);
nor U1298 (N_1298,In_2465,In_849);
xor U1299 (N_1299,In_3241,In_4601);
or U1300 (N_1300,In_2643,In_3909);
nand U1301 (N_1301,In_3622,In_3078);
or U1302 (N_1302,In_4094,In_2816);
xnor U1303 (N_1303,In_707,In_1586);
nand U1304 (N_1304,In_2033,In_4225);
nand U1305 (N_1305,In_3171,In_3726);
and U1306 (N_1306,In_3315,In_1831);
or U1307 (N_1307,In_3289,In_3543);
or U1308 (N_1308,In_675,In_4328);
and U1309 (N_1309,In_3655,In_3106);
nand U1310 (N_1310,In_1728,In_610);
and U1311 (N_1311,In_517,In_47);
xor U1312 (N_1312,In_3238,In_3485);
nor U1313 (N_1313,In_3736,In_1855);
and U1314 (N_1314,In_2430,In_1684);
or U1315 (N_1315,In_2575,In_3823);
and U1316 (N_1316,In_3765,In_855);
or U1317 (N_1317,In_2102,In_1957);
nand U1318 (N_1318,In_4427,In_856);
nand U1319 (N_1319,In_2882,In_4400);
or U1320 (N_1320,In_1417,In_515);
and U1321 (N_1321,In_2887,In_4246);
and U1322 (N_1322,In_2010,In_1094);
xnor U1323 (N_1323,In_1096,In_2802);
nor U1324 (N_1324,In_1013,In_1688);
and U1325 (N_1325,In_504,In_3887);
and U1326 (N_1326,In_1535,In_734);
nor U1327 (N_1327,In_175,In_238);
or U1328 (N_1328,In_3375,In_833);
and U1329 (N_1329,In_3050,In_631);
nand U1330 (N_1330,In_4169,In_144);
and U1331 (N_1331,In_3937,In_2779);
xor U1332 (N_1332,In_636,In_3011);
nand U1333 (N_1333,In_1444,In_4466);
nand U1334 (N_1334,In_2602,In_875);
nor U1335 (N_1335,In_3935,In_3374);
and U1336 (N_1336,In_2681,In_4167);
nand U1337 (N_1337,In_1159,In_4536);
nor U1338 (N_1338,In_1554,In_1066);
nand U1339 (N_1339,In_2428,In_2753);
nor U1340 (N_1340,In_3839,In_1771);
nor U1341 (N_1341,In_983,In_3473);
and U1342 (N_1342,In_8,In_3421);
nand U1343 (N_1343,In_2698,In_3151);
xor U1344 (N_1344,In_641,In_1931);
and U1345 (N_1345,In_4444,In_378);
or U1346 (N_1346,In_3786,In_781);
xnor U1347 (N_1347,In_3634,In_1087);
nor U1348 (N_1348,In_4491,In_2249);
xor U1349 (N_1349,In_1829,In_1155);
nand U1350 (N_1350,In_4139,In_3957);
and U1351 (N_1351,In_909,In_4770);
or U1352 (N_1352,In_4591,In_257);
or U1353 (N_1353,In_4682,In_1635);
nor U1354 (N_1354,In_998,In_3400);
nor U1355 (N_1355,In_2041,In_960);
or U1356 (N_1356,In_4349,In_438);
xnor U1357 (N_1357,In_822,In_4061);
xnor U1358 (N_1358,In_357,In_1926);
or U1359 (N_1359,In_165,In_1782);
nand U1360 (N_1360,In_3591,In_2129);
xnor U1361 (N_1361,In_4564,In_1463);
or U1362 (N_1362,In_3053,In_2668);
xor U1363 (N_1363,In_2896,In_4928);
nand U1364 (N_1364,In_1707,In_1672);
xnor U1365 (N_1365,In_375,In_494);
nor U1366 (N_1366,In_1461,In_431);
nor U1367 (N_1367,In_1732,In_2609);
or U1368 (N_1368,In_4751,In_2336);
nor U1369 (N_1369,In_1951,In_1749);
nand U1370 (N_1370,In_3676,In_2401);
nor U1371 (N_1371,In_4490,In_1801);
nand U1372 (N_1372,In_548,In_4945);
nand U1373 (N_1373,In_3881,In_4586);
nor U1374 (N_1374,In_1709,In_3180);
xor U1375 (N_1375,In_4584,In_4108);
nor U1376 (N_1376,In_4960,In_304);
and U1377 (N_1377,In_3248,In_2583);
and U1378 (N_1378,In_4938,In_2103);
nand U1379 (N_1379,In_3949,In_4291);
and U1380 (N_1380,In_3352,In_2808);
or U1381 (N_1381,In_201,In_4853);
xor U1382 (N_1382,In_3625,In_1269);
or U1383 (N_1383,In_3033,In_4724);
nor U1384 (N_1384,In_3434,In_2095);
nand U1385 (N_1385,In_1229,In_1361);
nor U1386 (N_1386,In_1970,In_3801);
and U1387 (N_1387,In_3952,In_2432);
and U1388 (N_1388,In_613,In_234);
and U1389 (N_1389,In_2619,In_1295);
nand U1390 (N_1390,In_2216,In_2504);
or U1391 (N_1391,In_1142,In_4333);
and U1392 (N_1392,In_1862,In_4229);
and U1393 (N_1393,In_2071,In_2092);
or U1394 (N_1394,In_217,In_740);
or U1395 (N_1395,In_1391,In_626);
and U1396 (N_1396,In_3774,In_2105);
and U1397 (N_1397,In_3226,In_3161);
nor U1398 (N_1398,In_2638,In_3577);
or U1399 (N_1399,In_2584,In_2835);
xor U1400 (N_1400,In_4700,In_2701);
and U1401 (N_1401,In_2200,In_395);
and U1402 (N_1402,In_2726,In_2087);
or U1403 (N_1403,In_2270,In_4831);
xor U1404 (N_1404,In_4557,In_1717);
and U1405 (N_1405,In_2389,In_2677);
nand U1406 (N_1406,In_367,In_4766);
xor U1407 (N_1407,In_1074,In_230);
and U1408 (N_1408,In_2950,In_1503);
xnor U1409 (N_1409,In_3456,In_1007);
and U1410 (N_1410,In_656,In_1128);
nand U1411 (N_1411,In_1622,In_1778);
and U1412 (N_1412,In_2232,In_3523);
xor U1413 (N_1413,In_2611,In_615);
xor U1414 (N_1414,In_2596,In_1731);
nand U1415 (N_1415,In_4415,In_4649);
xnor U1416 (N_1416,In_2809,In_4930);
or U1417 (N_1417,In_340,In_3858);
and U1418 (N_1418,In_189,In_1820);
nand U1419 (N_1419,In_4399,In_2122);
or U1420 (N_1420,In_3487,In_1318);
xnor U1421 (N_1421,In_1275,In_986);
and U1422 (N_1422,In_2362,In_2767);
and U1423 (N_1423,In_225,In_3018);
or U1424 (N_1424,In_4408,In_831);
xnor U1425 (N_1425,In_1469,In_4567);
or U1426 (N_1426,In_141,In_4366);
or U1427 (N_1427,In_4894,In_4778);
nand U1428 (N_1428,In_94,In_4055);
or U1429 (N_1429,In_1041,In_99);
nor U1430 (N_1430,In_4932,In_339);
and U1431 (N_1431,In_1579,In_4152);
and U1432 (N_1432,In_3432,In_3043);
and U1433 (N_1433,In_2659,In_1075);
xnor U1434 (N_1434,In_4368,In_1382);
nand U1435 (N_1435,In_197,In_2002);
or U1436 (N_1436,In_442,In_1242);
xor U1437 (N_1437,In_3542,In_4820);
and U1438 (N_1438,In_1515,In_721);
xor U1439 (N_1439,In_1308,In_4757);
and U1440 (N_1440,In_2209,In_846);
xor U1441 (N_1441,In_3683,In_4497);
or U1442 (N_1442,In_2183,In_625);
and U1443 (N_1443,In_3017,In_1473);
or U1444 (N_1444,In_2988,In_1372);
and U1445 (N_1445,In_4110,In_2703);
and U1446 (N_1446,In_4485,In_297);
and U1447 (N_1447,In_3301,In_4011);
nor U1448 (N_1448,In_3258,In_17);
xnor U1449 (N_1449,In_4106,In_1045);
and U1450 (N_1450,In_4006,In_2199);
xnor U1451 (N_1451,In_4123,In_3574);
or U1452 (N_1452,In_524,In_1777);
xnor U1453 (N_1453,In_4507,In_866);
and U1454 (N_1454,In_4908,In_1780);
nand U1455 (N_1455,In_463,In_3047);
nor U1456 (N_1456,In_2315,In_3811);
nand U1457 (N_1457,In_3694,In_1313);
nor U1458 (N_1458,In_653,In_4865);
and U1459 (N_1459,In_918,In_337);
or U1460 (N_1460,In_4819,In_3843);
and U1461 (N_1461,In_3201,In_2957);
and U1462 (N_1462,In_4327,In_2267);
nor U1463 (N_1463,In_4341,In_2536);
nand U1464 (N_1464,In_489,In_2688);
or U1465 (N_1465,In_2563,In_2519);
nor U1466 (N_1466,In_4260,In_1122);
xor U1467 (N_1467,In_1388,In_1090);
nand U1468 (N_1468,In_2724,In_3044);
nor U1469 (N_1469,In_3179,In_1072);
nand U1470 (N_1470,In_3835,In_2845);
xor U1471 (N_1471,In_1383,In_135);
or U1472 (N_1472,In_2856,In_2039);
xnor U1473 (N_1473,In_979,In_1284);
nand U1474 (N_1474,In_4454,In_2451);
and U1475 (N_1475,In_4053,In_2042);
and U1476 (N_1476,In_697,In_192);
nor U1477 (N_1477,In_4085,In_2776);
or U1478 (N_1478,In_1222,In_11);
nor U1479 (N_1479,In_2605,In_1603);
and U1480 (N_1480,In_4767,In_862);
and U1481 (N_1481,In_203,In_2064);
nand U1482 (N_1482,In_4337,In_4939);
nor U1483 (N_1483,In_4980,In_2551);
xor U1484 (N_1484,In_3020,In_3703);
xor U1485 (N_1485,In_3816,In_4958);
and U1486 (N_1486,In_1364,In_3761);
nand U1487 (N_1487,In_701,In_4948);
or U1488 (N_1488,In_4714,In_480);
xor U1489 (N_1489,In_3612,In_2515);
and U1490 (N_1490,In_338,In_931);
and U1491 (N_1491,In_3092,In_3032);
xnor U1492 (N_1492,In_837,In_109);
nor U1493 (N_1493,In_26,In_2142);
and U1494 (N_1494,In_16,In_161);
nand U1495 (N_1495,In_1705,In_2764);
xnor U1496 (N_1496,In_1023,In_2915);
nor U1497 (N_1497,In_4432,In_4437);
nor U1498 (N_1498,In_850,In_1792);
xor U1499 (N_1499,In_1126,In_864);
or U1500 (N_1500,In_1975,In_2647);
or U1501 (N_1501,In_2566,In_320);
nand U1502 (N_1502,In_4254,In_2120);
xor U1503 (N_1503,In_4355,In_4293);
xor U1504 (N_1504,In_2771,In_4016);
or U1505 (N_1505,In_3773,In_3657);
xor U1506 (N_1506,In_2044,In_467);
nand U1507 (N_1507,In_1228,In_3293);
or U1508 (N_1508,In_3555,In_150);
nor U1509 (N_1509,In_4070,In_685);
nand U1510 (N_1510,In_4275,In_492);
xor U1511 (N_1511,In_3490,In_4783);
or U1512 (N_1512,In_2281,In_765);
nand U1513 (N_1513,In_730,In_975);
or U1514 (N_1514,In_423,In_1297);
and U1515 (N_1515,In_3701,In_486);
and U1516 (N_1516,In_12,In_1453);
xnor U1517 (N_1517,In_4505,In_2810);
nand U1518 (N_1518,In_563,In_4258);
or U1519 (N_1519,In_2673,In_2666);
nand U1520 (N_1520,In_3678,In_1513);
nor U1521 (N_1521,In_1044,In_2790);
nor U1522 (N_1522,In_3348,In_1746);
and U1523 (N_1523,In_4999,In_1006);
nand U1524 (N_1524,In_2174,In_4093);
and U1525 (N_1525,In_3525,In_2797);
xnor U1526 (N_1526,In_2130,In_900);
nand U1527 (N_1527,In_3502,In_478);
nand U1528 (N_1528,In_3729,In_2774);
nor U1529 (N_1529,In_2228,In_3124);
or U1530 (N_1530,In_1821,In_1119);
xnor U1531 (N_1531,In_2550,In_4753);
and U1532 (N_1532,In_4526,In_2516);
or U1533 (N_1533,In_3281,In_3441);
xor U1534 (N_1534,In_582,In_3921);
xor U1535 (N_1535,In_1151,In_565);
nor U1536 (N_1536,In_3088,In_4952);
nor U1537 (N_1537,In_330,In_1412);
nor U1538 (N_1538,In_470,In_1196);
nor U1539 (N_1539,In_1061,In_3123);
nand U1540 (N_1540,In_1651,In_4338);
xor U1541 (N_1541,In_4886,In_1110);
or U1542 (N_1542,In_3087,In_4474);
xnor U1543 (N_1543,In_25,In_397);
and U1544 (N_1544,In_1037,In_4737);
nand U1545 (N_1545,In_3028,In_1850);
or U1546 (N_1546,In_2045,In_3483);
and U1547 (N_1547,In_988,In_3962);
and U1548 (N_1548,In_2454,In_4967);
nand U1549 (N_1549,In_3708,In_2303);
xnor U1550 (N_1550,In_667,In_194);
nand U1551 (N_1551,In_3880,In_1337);
and U1552 (N_1552,In_3776,In_4625);
or U1553 (N_1553,In_4176,In_3827);
and U1554 (N_1554,In_3693,In_4209);
or U1555 (N_1555,In_2326,In_4089);
nor U1556 (N_1556,In_31,In_674);
nand U1557 (N_1557,In_2674,In_1255);
nand U1558 (N_1558,In_85,In_4271);
and U1559 (N_1559,In_3227,In_1824);
xnor U1560 (N_1560,In_3579,In_3472);
nand U1561 (N_1561,In_4727,In_3961);
nand U1562 (N_1562,In_4375,In_364);
nand U1563 (N_1563,In_3917,In_3660);
or U1564 (N_1564,In_3292,In_1947);
and U1565 (N_1565,In_326,In_1615);
or U1566 (N_1566,In_4558,In_168);
xor U1567 (N_1567,In_1819,In_2313);
nand U1568 (N_1568,In_2146,In_331);
nand U1569 (N_1569,In_4872,In_361);
or U1570 (N_1570,In_4701,In_1053);
xnor U1571 (N_1571,In_2500,In_1407);
nor U1572 (N_1572,In_4332,In_4290);
xnor U1573 (N_1573,In_1918,In_920);
nor U1574 (N_1574,In_2548,In_2473);
nand U1575 (N_1575,In_4935,In_4309);
or U1576 (N_1576,In_1220,In_946);
xor U1577 (N_1577,In_1857,In_1099);
nand U1578 (N_1578,In_1482,In_1967);
or U1579 (N_1579,In_4036,In_218);
or U1580 (N_1580,In_1739,In_3724);
xnor U1581 (N_1581,In_1153,In_2462);
nand U1582 (N_1582,In_3336,In_4321);
nand U1583 (N_1583,In_239,In_2968);
nor U1584 (N_1584,In_2918,In_4124);
nor U1585 (N_1585,In_2795,In_1939);
nand U1586 (N_1586,In_2625,In_3744);
or U1587 (N_1587,In_3553,In_2085);
or U1588 (N_1588,In_603,In_1194);
nand U1589 (N_1589,In_1414,In_3314);
nand U1590 (N_1590,In_1641,In_3670);
or U1591 (N_1591,In_3277,In_973);
and U1592 (N_1592,In_1030,In_2269);
or U1593 (N_1593,In_4552,In_71);
or U1594 (N_1594,In_453,In_1971);
or U1595 (N_1595,In_2069,In_52);
or U1596 (N_1596,In_451,In_4273);
nor U1597 (N_1597,In_4019,In_461);
nor U1598 (N_1598,In_808,In_2331);
or U1599 (N_1599,In_4050,In_4410);
and U1600 (N_1600,In_4993,In_4618);
nor U1601 (N_1601,In_1632,In_3321);
and U1602 (N_1602,In_449,In_66);
and U1603 (N_1603,In_2864,In_637);
and U1604 (N_1604,In_2580,In_1678);
or U1605 (N_1605,In_3616,In_4266);
xor U1606 (N_1606,In_3324,In_34);
or U1607 (N_1607,In_1048,In_4360);
xnor U1608 (N_1608,In_1575,In_3260);
and U1609 (N_1609,In_389,In_4827);
nand U1610 (N_1610,In_3370,In_4187);
or U1611 (N_1611,In_3175,In_3158);
nand U1612 (N_1612,In_693,In_4090);
or U1613 (N_1613,In_890,In_2119);
nor U1614 (N_1614,In_704,In_1100);
or U1615 (N_1615,In_2570,In_4694);
xor U1616 (N_1616,In_2765,In_2070);
nor U1617 (N_1617,In_58,In_3059);
and U1618 (N_1618,In_3199,In_558);
nand U1619 (N_1619,In_913,In_3194);
xor U1620 (N_1620,In_3598,In_4414);
xnor U1621 (N_1621,In_3305,In_3567);
nand U1622 (N_1622,In_1439,In_2922);
or U1623 (N_1623,In_95,In_1031);
nor U1624 (N_1624,In_3476,In_529);
xnor U1625 (N_1625,In_2419,In_286);
xnor U1626 (N_1626,In_3007,In_1865);
nand U1627 (N_1627,In_3423,In_4739);
xnor U1628 (N_1628,In_2110,In_2416);
nor U1629 (N_1629,In_4698,In_117);
nand U1630 (N_1630,In_2408,In_1116);
and U1631 (N_1631,In_2083,In_4082);
nor U1632 (N_1632,In_718,In_3561);
or U1633 (N_1633,In_1230,In_4684);
or U1634 (N_1634,In_334,In_658);
xnor U1635 (N_1635,In_1446,In_4696);
and U1636 (N_1636,In_4829,In_4101);
nand U1637 (N_1637,In_1610,In_2452);
and U1638 (N_1638,In_1164,In_2290);
or U1639 (N_1639,In_2573,In_1005);
xnor U1640 (N_1640,In_2474,In_2354);
xor U1641 (N_1641,In_4514,In_1027);
nand U1642 (N_1642,In_3426,In_4200);
or U1643 (N_1643,In_575,In_4482);
nor U1644 (N_1644,In_2571,In_1185);
nand U1645 (N_1645,In_2903,In_4677);
and U1646 (N_1646,In_3488,In_4893);
and U1647 (N_1647,In_1674,In_585);
nor U1648 (N_1648,In_2149,In_4189);
nand U1649 (N_1649,In_207,In_4852);
nand U1650 (N_1650,In_1706,In_4049);
and U1651 (N_1651,In_3836,In_1487);
and U1652 (N_1652,In_2369,In_2357);
nor U1653 (N_1653,In_3803,In_1339);
xor U1654 (N_1654,In_2665,In_291);
nor U1655 (N_1655,In_4500,In_4904);
and U1656 (N_1656,In_3197,In_3054);
or U1657 (N_1657,In_1559,In_537);
and U1658 (N_1658,In_1024,In_3831);
xor U1659 (N_1659,In_179,In_1847);
nand U1660 (N_1660,In_2826,In_861);
xor U1661 (N_1661,In_4632,In_1423);
nand U1662 (N_1662,In_2946,In_3064);
xnor U1663 (N_1663,In_1148,In_3160);
nand U1664 (N_1664,In_456,In_1874);
xor U1665 (N_1665,In_3354,In_4004);
or U1666 (N_1666,In_1984,In_1464);
or U1667 (N_1667,In_1135,In_4499);
xnor U1668 (N_1668,In_3005,In_4570);
nor U1669 (N_1669,In_2062,In_1445);
nand U1670 (N_1670,In_3257,In_1869);
nand U1671 (N_1671,In_2022,In_228);
or U1672 (N_1672,In_2916,In_1810);
xnor U1673 (N_1673,In_4768,In_1395);
nand U1674 (N_1674,In_3131,In_420);
xnor U1675 (N_1675,In_1930,In_526);
or U1676 (N_1676,In_3805,In_2306);
and U1677 (N_1677,In_554,In_629);
xnor U1678 (N_1678,In_3963,In_3630);
nand U1679 (N_1679,In_1597,In_3457);
xor U1680 (N_1680,In_2657,In_191);
xor U1681 (N_1681,In_878,In_4870);
nand U1682 (N_1682,In_3535,In_2540);
nand U1683 (N_1683,In_3855,In_1922);
nor U1684 (N_1684,In_4600,In_1540);
nand U1685 (N_1685,In_447,In_905);
nor U1686 (N_1686,In_3373,In_583);
or U1687 (N_1687,In_2457,In_2956);
nand U1688 (N_1688,In_508,In_2534);
nor U1689 (N_1689,In_4352,In_2118);
nor U1690 (N_1690,In_4875,In_102);
or U1691 (N_1691,In_3466,In_390);
or U1692 (N_1692,In_4528,In_3886);
nor U1693 (N_1693,In_4971,In_1197);
and U1694 (N_1694,In_1241,In_1311);
or U1695 (N_1695,In_683,In_1779);
nor U1696 (N_1696,In_1016,In_2082);
nand U1697 (N_1697,In_1479,In_1430);
or U1698 (N_1698,In_3137,In_2024);
and U1699 (N_1699,In_1489,In_79);
nor U1700 (N_1700,In_4146,In_219);
or U1701 (N_1701,In_4868,In_3848);
and U1702 (N_1702,In_2893,In_3684);
nand U1703 (N_1703,In_4554,In_601);
and U1704 (N_1704,In_3443,In_1991);
nand U1705 (N_1705,In_2456,In_1198);
and U1706 (N_1706,In_2561,In_2137);
or U1707 (N_1707,In_202,In_3954);
xor U1708 (N_1708,In_2762,In_1123);
nand U1709 (N_1709,In_799,In_2152);
nor U1710 (N_1710,In_3086,In_1477);
or U1711 (N_1711,In_588,In_1713);
xor U1712 (N_1712,In_3269,In_3731);
nor U1713 (N_1713,In_3587,In_2494);
nor U1714 (N_1714,In_1759,In_1328);
xor U1715 (N_1715,In_2715,In_1952);
or U1716 (N_1716,In_3360,In_4406);
xor U1717 (N_1717,In_898,In_4673);
nand U1718 (N_1718,In_1057,In_2116);
nor U1719 (N_1719,In_3711,In_3649);
nand U1720 (N_1720,In_4891,In_2263);
nor U1721 (N_1721,In_4885,In_167);
nor U1722 (N_1722,In_2233,In_4172);
xor U1723 (N_1723,In_2317,In_2543);
nand U1724 (N_1724,In_3034,In_1334);
or U1725 (N_1725,In_1568,In_3713);
nor U1726 (N_1726,In_4132,In_4479);
or U1727 (N_1727,In_1996,In_2242);
xor U1728 (N_1728,In_2310,In_3897);
nand U1729 (N_1729,In_459,In_3282);
or U1730 (N_1730,In_3633,In_1756);
nand U1731 (N_1731,In_1134,In_1467);
nor U1732 (N_1732,In_4038,In_481);
nor U1733 (N_1733,In_3329,In_2940);
xor U1734 (N_1734,In_1726,In_1649);
and U1735 (N_1735,In_3102,In_4144);
nor U1736 (N_1736,In_1813,In_3664);
nand U1737 (N_1737,In_65,In_4726);
nor U1738 (N_1738,In_3386,In_1366);
or U1739 (N_1739,In_516,In_4662);
and U1740 (N_1740,In_695,In_553);
xnor U1741 (N_1741,In_1447,In_4207);
xnor U1742 (N_1742,In_1839,In_3849);
or U1743 (N_1743,In_726,In_3480);
nand U1744 (N_1744,In_3442,In_2278);
or U1745 (N_1745,In_4664,In_2868);
nor U1746 (N_1746,In_1365,In_1894);
xor U1747 (N_1747,In_747,In_957);
or U1748 (N_1748,In_668,In_3023);
xnor U1749 (N_1749,In_3539,In_868);
or U1750 (N_1750,In_247,In_1679);
or U1751 (N_1751,In_632,In_1345);
or U1752 (N_1752,In_4316,In_2125);
nor U1753 (N_1753,In_366,In_373);
nor U1754 (N_1754,In_4805,In_3142);
xor U1755 (N_1755,In_1421,In_2463);
nor U1756 (N_1756,In_2163,In_1669);
or U1757 (N_1757,In_1203,In_2642);
and U1758 (N_1758,In_2259,In_2366);
nand U1759 (N_1759,In_136,In_2141);
or U1760 (N_1760,In_160,In_532);
nor U1761 (N_1761,In_1039,In_3532);
xnor U1762 (N_1762,In_2434,In_1124);
nor U1763 (N_1763,In_2020,In_1564);
xor U1764 (N_1764,In_3964,In_224);
nand U1765 (N_1765,In_3847,In_3905);
or U1766 (N_1766,In_789,In_3771);
or U1767 (N_1767,In_3235,In_4340);
nand U1768 (N_1768,In_3119,In_3052);
xnor U1769 (N_1769,In_2722,In_126);
nand U1770 (N_1770,In_592,In_609);
nor U1771 (N_1771,In_1736,In_654);
or U1772 (N_1772,In_4855,In_4581);
or U1773 (N_1773,In_3534,In_3397);
and U1774 (N_1774,In_2763,In_3767);
nand U1775 (N_1775,In_1990,In_4265);
xnor U1776 (N_1776,In_4900,In_3367);
or U1777 (N_1777,In_45,In_544);
nor U1778 (N_1778,In_3854,In_3733);
nor U1779 (N_1779,In_301,In_3157);
xor U1780 (N_1780,In_4473,In_1214);
or U1781 (N_1781,In_2399,In_483);
and U1782 (N_1782,In_845,In_4642);
and U1783 (N_1783,In_2276,In_1644);
xor U1784 (N_1784,In_3085,In_2164);
xnor U1785 (N_1785,In_237,In_4652);
and U1786 (N_1786,In_1897,In_3528);
nor U1787 (N_1787,In_3270,In_566);
xor U1788 (N_1788,In_1010,In_4861);
nand U1789 (N_1789,In_3163,In_3757);
nand U1790 (N_1790,In_3450,In_3947);
and U1791 (N_1791,In_3524,In_4759);
nor U1792 (N_1792,In_2328,In_3379);
and U1793 (N_1793,In_3924,In_3560);
xnor U1794 (N_1794,In_108,In_4973);
and U1795 (N_1795,In_2134,In_2545);
nor U1796 (N_1796,In_4669,In_1409);
xor U1797 (N_1797,In_4354,In_2866);
nor U1798 (N_1798,In_2089,In_464);
xnor U1799 (N_1799,In_4131,In_2907);
and U1800 (N_1800,In_1508,In_4463);
nor U1801 (N_1801,In_2168,In_3628);
nand U1802 (N_1802,In_4219,In_115);
or U1803 (N_1803,In_3759,In_692);
nand U1804 (N_1804,In_2224,In_316);
xnor U1805 (N_1805,In_386,In_3692);
or U1806 (N_1806,In_1084,In_3796);
xor U1807 (N_1807,In_2173,In_1377);
nand U1808 (N_1808,In_912,In_3072);
and U1809 (N_1809,In_2068,In_2178);
nor U1810 (N_1810,In_28,In_997);
or U1811 (N_1811,In_2963,In_4680);
and U1812 (N_1812,In_877,In_2449);
xor U1813 (N_1813,In_3345,In_4746);
and U1814 (N_1814,In_477,In_3958);
xor U1815 (N_1815,In_3326,In_2234);
or U1816 (N_1816,In_3187,In_4675);
and U1817 (N_1817,In_1798,In_2675);
nor U1818 (N_1818,In_2052,In_4359);
nand U1819 (N_1819,In_1652,In_100);
and U1820 (N_1820,In_533,In_3978);
nand U1821 (N_1821,In_1593,In_500);
or U1822 (N_1822,In_2800,In_4009);
nand U1823 (N_1823,In_3148,In_121);
and U1824 (N_1824,In_4455,In_620);
xnor U1825 (N_1825,In_4224,In_1105);
nand U1826 (N_1826,In_169,In_4773);
nor U1827 (N_1827,In_1548,In_818);
or U1828 (N_1828,In_910,In_1883);
and U1829 (N_1829,In_4205,In_255);
nand U1830 (N_1830,In_1690,In_2113);
or U1831 (N_1831,In_2996,In_867);
nor U1832 (N_1832,In_4775,In_1459);
nor U1833 (N_1833,In_3147,In_2246);
xnor U1834 (N_1834,In_4423,In_253);
xor U1835 (N_1835,In_4407,In_4285);
nand U1836 (N_1836,In_3338,In_1149);
nand U1837 (N_1837,In_2964,In_1993);
and U1838 (N_1838,In_3783,In_3931);
or U1839 (N_1839,In_1893,In_3648);
nand U1840 (N_1840,In_2614,In_369);
and U1841 (N_1841,In_1263,In_3221);
nand U1842 (N_1842,In_2883,In_4925);
nor U1843 (N_1843,In_2135,In_2080);
and U1844 (N_1844,In_507,In_3097);
nand U1845 (N_1845,In_2032,In_2880);
nor U1846 (N_1846,In_2901,In_3232);
nand U1847 (N_1847,In_2747,In_2759);
nor U1848 (N_1848,In_2600,In_302);
xnor U1849 (N_1849,In_4725,In_2612);
xor U1850 (N_1850,In_1267,In_86);
xor U1851 (N_1851,In_1086,In_2213);
and U1852 (N_1852,In_4269,In_2489);
or U1853 (N_1853,In_4705,In_343);
xnor U1854 (N_1854,In_188,In_2850);
nand U1855 (N_1855,In_2757,In_2480);
or U1856 (N_1856,In_3943,In_1972);
xor U1857 (N_1857,In_1654,In_414);
nand U1858 (N_1858,In_4047,In_1682);
nand U1859 (N_1859,In_2838,In_724);
xnor U1860 (N_1860,In_2530,In_4686);
nand U1861 (N_1861,In_3395,In_3777);
or U1862 (N_1862,In_4166,In_186);
xnor U1863 (N_1863,In_4362,In_3417);
and U1864 (N_1864,In_3401,In_2012);
and U1865 (N_1865,In_2048,In_1764);
nor U1866 (N_1866,In_874,In_199);
or U1867 (N_1867,In_2261,In_3734);
and U1868 (N_1868,In_4762,In_295);
or U1869 (N_1869,In_4728,In_953);
xnor U1870 (N_1870,In_4180,In_1787);
nand U1871 (N_1871,In_4798,In_3331);
or U1872 (N_1872,In_1680,In_3334);
or U1873 (N_1873,In_1793,In_1578);
nor U1874 (N_1874,In_4619,In_1330);
nand U1875 (N_1875,In_514,In_530);
nand U1876 (N_1876,In_3844,In_1171);
or U1877 (N_1877,In_4397,In_1594);
nor U1878 (N_1878,In_4624,In_2526);
nand U1879 (N_1879,In_4042,In_4864);
nand U1880 (N_1880,In_3914,In_4837);
and U1881 (N_1881,In_1204,In_4895);
nor U1882 (N_1882,In_3357,In_3217);
xor U1883 (N_1883,In_3378,In_3689);
nor U1884 (N_1884,In_4000,In_3959);
and U1885 (N_1885,In_448,In_2223);
nand U1886 (N_1886,In_1565,In_1828);
or U1887 (N_1887,In_1797,In_2990);
xor U1888 (N_1888,In_1868,In_2979);
xnor U1889 (N_1889,In_2212,In_231);
nand U1890 (N_1890,In_4404,In_703);
nand U1891 (N_1891,In_3990,In_4442);
nand U1892 (N_1892,In_118,In_4970);
nor U1893 (N_1893,In_3735,In_3618);
nor U1894 (N_1894,In_446,In_4545);
or U1895 (N_1895,In_1581,In_3725);
or U1896 (N_1896,In_671,In_1483);
xor U1897 (N_1897,In_4025,In_440);
nor U1898 (N_1898,In_3465,In_840);
xor U1899 (N_1899,In_4324,In_2477);
nand U1900 (N_1900,In_745,In_3039);
nand U1901 (N_1901,In_2245,In_1497);
or U1902 (N_1902,In_3203,In_4228);
and U1903 (N_1903,In_495,In_3531);
xor U1904 (N_1904,In_3105,In_2244);
xor U1905 (N_1905,In_277,In_594);
nand U1906 (N_1906,In_1437,In_1426);
nand U1907 (N_1907,In_4892,In_1574);
or U1908 (N_1908,In_4578,In_3817);
and U1909 (N_1909,In_687,In_2689);
nand U1910 (N_1910,In_50,In_2973);
nand U1911 (N_1911,In_1266,In_4573);
xor U1912 (N_1912,In_2435,In_1663);
nand U1913 (N_1913,In_4175,In_750);
nor U1914 (N_1914,In_143,In_1355);
nand U1915 (N_1915,In_4606,In_4008);
nor U1916 (N_1916,In_3505,In_4884);
nand U1917 (N_1917,In_753,In_4965);
or U1918 (N_1918,In_4899,In_2090);
and U1919 (N_1919,In_3286,In_1806);
xnor U1920 (N_1920,In_4449,In_1584);
xor U1921 (N_1921,In_1898,In_551);
nand U1922 (N_1922,In_2775,In_2777);
or U1923 (N_1923,In_562,In_2796);
nor U1924 (N_1924,In_3705,In_3152);
nand U1925 (N_1925,In_3832,In_3095);
or U1926 (N_1926,In_1133,In_2214);
and U1927 (N_1927,In_488,In_1350);
nand U1928 (N_1928,In_3498,In_4071);
nor U1929 (N_1929,In_4202,In_3842);
nor U1930 (N_1930,In_3910,In_3762);
nand U1931 (N_1931,In_4822,In_2367);
or U1932 (N_1932,In_2650,In_2559);
nor U1933 (N_1933,In_790,In_3714);
nor U1934 (N_1934,In_3732,In_1083);
nand U1935 (N_1935,In_2450,In_1067);
or U1936 (N_1936,In_51,In_1178);
or U1937 (N_1937,In_815,In_1246);
xnor U1938 (N_1938,In_1034,In_3760);
xor U1939 (N_1939,In_3904,In_819);
and U1940 (N_1940,In_1233,In_4385);
nor U1941 (N_1941,In_2047,In_3196);
or U1942 (N_1942,In_731,In_573);
nand U1943 (N_1943,In_4915,In_3779);
or U1944 (N_1944,In_4750,In_3530);
nor U1945 (N_1945,In_3297,In_4690);
and U1946 (N_1946,In_1191,In_926);
xor U1947 (N_1947,In_4035,In_2591);
nor U1948 (N_1948,In_3066,In_2460);
nor U1949 (N_1949,In_403,In_4192);
nand U1950 (N_1950,In_1938,In_2645);
or U1951 (N_1951,In_2527,In_1962);
xor U1952 (N_1952,In_3317,In_1333);
or U1953 (N_1953,In_3206,In_4486);
xnor U1954 (N_1954,In_1227,In_572);
nand U1955 (N_1955,In_1604,In_49);
or U1956 (N_1956,In_2381,In_1167);
or U1957 (N_1957,In_2248,In_1814);
or U1958 (N_1958,In_1511,In_1623);
and U1959 (N_1959,In_3927,In_571);
xor U1960 (N_1960,In_3198,In_2140);
or U1961 (N_1961,In_826,In_73);
xnor U1962 (N_1962,In_2133,In_3010);
or U1963 (N_1963,In_1205,In_2440);
xor U1964 (N_1964,In_1961,In_2529);
nand U1965 (N_1965,In_1751,In_4611);
and U1966 (N_1966,In_4048,In_1102);
and U1967 (N_1967,In_4546,In_4976);
nor U1968 (N_1968,In_2254,In_2628);
nor U1969 (N_1969,In_2914,In_200);
and U1970 (N_1970,In_4658,In_2699);
nand U1971 (N_1971,In_1743,In_2375);
nand U1972 (N_1972,In_2036,In_1526);
nor U1973 (N_1973,In_3103,In_1274);
xnor U1974 (N_1974,In_2652,In_4181);
xnor U1975 (N_1975,In_1664,In_2323);
nor U1976 (N_1976,In_2923,In_278);
and U1977 (N_1977,In_1619,In_2503);
or U1978 (N_1978,In_3609,In_1650);
or U1979 (N_1979,In_124,In_2931);
nand U1980 (N_1980,In_760,In_2646);
nor U1981 (N_1981,In_37,In_4818);
or U1982 (N_1982,In_1799,In_3014);
xor U1983 (N_1983,In_487,In_3188);
nand U1984 (N_1984,In_1127,In_2413);
nor U1985 (N_1985,In_3753,In_3893);
or U1986 (N_1986,In_3393,In_663);
nand U1987 (N_1987,In_3575,In_2291);
nor U1988 (N_1988,In_2707,In_1789);
xnor U1989 (N_1989,In_350,In_1724);
nand U1990 (N_1990,In_3875,In_2294);
and U1991 (N_1991,In_4634,In_4799);
and U1992 (N_1992,In_3108,In_2937);
nor U1993 (N_1993,In_3775,In_3425);
and U1994 (N_1994,In_4149,In_732);
nor U1995 (N_1995,In_3595,In_2060);
nand U1996 (N_1996,In_2038,In_2384);
and U1997 (N_1997,In_3589,In_546);
nor U1998 (N_1998,In_1715,In_4742);
or U1999 (N_1999,In_4059,In_3529);
xor U2000 (N_2000,In_4707,In_2813);
nand U2001 (N_2001,In_76,In_4477);
or U2002 (N_2002,In_1341,In_3596);
xor U2003 (N_2003,In_4446,In_81);
and U2004 (N_2004,In_2897,In_3046);
or U2005 (N_2005,In_4412,In_4527);
and U2006 (N_2006,In_4931,In_1098);
nand U2007 (N_2007,In_638,In_4238);
nor U2008 (N_2008,In_4863,In_2397);
xnor U2009 (N_2009,In_313,In_4129);
nor U2010 (N_2010,In_2236,In_1212);
and U2011 (N_2011,In_3884,In_3822);
nor U2012 (N_2012,In_2023,In_870);
xor U2013 (N_2013,In_4920,In_814);
xnor U2014 (N_2014,In_4054,In_4849);
nor U2015 (N_2015,In_1708,In_3477);
nor U2016 (N_2016,In_345,In_220);
or U2017 (N_2017,In_499,In_3388);
and U2018 (N_2018,In_4277,In_14);
and U2019 (N_2019,In_3971,In_3181);
nand U2020 (N_2020,In_3911,In_180);
nor U2021 (N_2021,In_3933,In_2984);
xor U2022 (N_2022,In_2719,In_1804);
and U2023 (N_2023,In_3940,In_1524);
xnor U2024 (N_2024,In_1997,In_2403);
nor U2025 (N_2025,In_1899,In_1457);
nor U2026 (N_2026,In_2304,In_1776);
or U2027 (N_2027,In_3369,In_3192);
and U2028 (N_2028,In_346,In_3207);
xor U2029 (N_2029,In_2508,In_1481);
and U2030 (N_2030,In_2967,In_3135);
xnor U2031 (N_2031,In_370,In_3651);
or U2032 (N_2032,In_4810,In_2037);
nand U2033 (N_2033,In_1572,In_2735);
nor U2034 (N_2034,In_1929,In_1179);
nand U2035 (N_2035,In_1353,In_4127);
nand U2036 (N_2036,In_3090,In_1872);
nor U2037 (N_2037,In_4250,In_1495);
xnor U2038 (N_2038,In_2634,In_1238);
or U2039 (N_2039,In_4982,In_272);
nand U2040 (N_2040,In_128,In_2889);
or U2041 (N_2041,In_399,In_1946);
and U2042 (N_2042,In_4708,In_3083);
nand U2043 (N_2043,In_307,In_3383);
xnor U2044 (N_2044,In_989,In_2969);
and U2045 (N_2045,In_321,In_4743);
nand U2046 (N_2046,In_3718,In_1494);
nor U2047 (N_2047,In_1211,In_3060);
or U2048 (N_2048,In_648,In_1158);
nand U2049 (N_2049,In_279,In_559);
or U2050 (N_2050,In_2978,In_2243);
or U2051 (N_2051,In_1638,In_2754);
nand U2052 (N_2052,In_2798,In_4978);
nand U2053 (N_2053,In_1349,In_549);
nor U2054 (N_2054,In_222,In_1323);
nand U2055 (N_2055,In_2819,In_4761);
xnor U2056 (N_2056,In_2867,In_3687);
or U2057 (N_2057,In_3850,In_387);
or U2058 (N_2058,In_4666,In_2991);
xor U2059 (N_2059,In_437,In_1541);
xnor U2060 (N_2060,In_614,In_3398);
and U2061 (N_2061,In_2202,In_4383);
nor U2062 (N_2062,In_1052,In_3385);
or U2063 (N_2063,In_4613,In_3333);
or U2064 (N_2064,In_2635,In_4776);
nand U2065 (N_2065,In_2608,In_2065);
nand U2066 (N_2066,In_3573,In_3008);
and U2067 (N_2067,In_1088,In_271);
nor U2068 (N_2068,In_4522,In_1625);
nand U2069 (N_2069,In_380,In_4816);
xnor U2070 (N_2070,In_3717,In_1108);
xor U2071 (N_2071,In_1552,In_2016);
nand U2072 (N_2072,In_3418,In_2000);
and U2073 (N_2073,In_2333,In_1765);
and U2074 (N_2074,In_2858,In_394);
nor U2075 (N_2075,In_2581,In_4251);
xor U2076 (N_2076,In_3799,In_737);
nand U2077 (N_2077,In_4846,In_3122);
xnor U2078 (N_2078,In_1351,In_1125);
nor U2079 (N_2079,In_3240,In_1534);
xnor U2080 (N_2080,In_4874,In_694);
or U2081 (N_2081,In_3471,In_4297);
xor U2082 (N_2082,In_806,In_688);
nand U2083 (N_2083,In_3968,In_30);
nand U2084 (N_2084,In_591,In_1278);
xor U2085 (N_2085,In_2459,In_4715);
and U2086 (N_2086,In_3637,In_3749);
xnor U2087 (N_2087,In_2415,In_4241);
or U2088 (N_2088,In_1512,In_1689);
or U2089 (N_2089,In_4080,In_1921);
and U2090 (N_2090,In_646,In_274);
xor U2091 (N_2091,In_4732,In_3195);
nand U2092 (N_2092,In_2101,In_1892);
xor U2093 (N_2093,In_1065,In_672);
or U2094 (N_2094,In_3864,In_1172);
nor U2095 (N_2095,In_560,In_4242);
nor U2096 (N_2096,In_241,In_2288);
xnor U2097 (N_2097,In_2190,In_577);
and U2098 (N_2098,In_354,In_4417);
and U2099 (N_2099,In_4654,In_1234);
and U2100 (N_2100,In_1569,In_1833);
and U2101 (N_2101,In_4710,In_4877);
or U2102 (N_2102,In_4137,In_2727);
or U2103 (N_2103,In_3704,In_2712);
nand U2104 (N_2104,In_4790,In_4839);
or U2105 (N_2105,In_2001,In_3491);
nand U2106 (N_2106,In_834,In_2378);
and U2107 (N_2107,In_1181,In_1161);
or U2108 (N_2108,In_1960,In_1683);
and U2109 (N_2109,In_441,In_576);
and U2110 (N_2110,In_424,In_859);
xor U2111 (N_2111,In_1384,In_922);
nor U2112 (N_2112,In_4378,In_645);
nor U2113 (N_2113,In_1206,In_4640);
or U2114 (N_2114,In_2172,In_1781);
or U2115 (N_2115,In_655,In_3237);
nand U2116 (N_2116,In_3722,In_2252);
nor U2117 (N_2117,In_1701,In_1915);
and U2118 (N_2118,In_4559,In_4095);
nor U2119 (N_2119,In_2574,In_3503);
or U2120 (N_2120,In_1600,In_318);
nand U2121 (N_2121,In_751,In_3868);
nand U2122 (N_2122,In_4755,In_795);
and U2123 (N_2123,In_4926,In_1329);
or U2124 (N_2124,In_3656,In_1520);
nor U2125 (N_2125,In_980,In_1253);
nor U2126 (N_2126,In_3869,In_3390);
nor U2127 (N_2127,In_412,In_3685);
and U2128 (N_2128,In_944,In_2613);
and U2129 (N_2129,In_4396,In_758);
or U2130 (N_2130,In_3169,In_4580);
nand U2131 (N_2131,In_3144,In_4911);
xnor U2132 (N_2132,In_971,In_4815);
xnor U2133 (N_2133,In_4734,In_1317);
and U2134 (N_2134,In_4304,In_3644);
or U2135 (N_2135,In_3768,In_4211);
nand U2136 (N_2136,In_1889,In_764);
nand U2137 (N_2137,In_1763,In_770);
nand U2138 (N_2138,In_984,In_937);
nand U2139 (N_2139,In_3065,In_3973);
nand U2140 (N_2140,In_1790,In_589);
nand U2141 (N_2141,In_4102,In_2758);
and U2142 (N_2142,In_134,In_2780);
or U2143 (N_2143,In_894,In_4617);
xnor U2144 (N_2144,In_1758,In_2412);
or U2145 (N_2145,In_4380,In_1240);
nor U2146 (N_2146,In_4126,In_3024);
nor U2147 (N_2147,In_1769,In_4493);
xor U2148 (N_2148,In_3650,In_3143);
nor U2149 (N_2149,In_3938,In_2057);
nand U2150 (N_2150,In_4457,In_4344);
nand U2151 (N_2151,In_2387,In_23);
nand U2152 (N_2152,In_903,In_2194);
and U2153 (N_2153,In_4237,In_3605);
nor U2154 (N_2154,In_4402,In_1000);
xnor U2155 (N_2155,In_774,In_2279);
and U2156 (N_2156,In_3177,In_111);
and U2157 (N_2157,In_2318,In_1937);
xor U2158 (N_2158,In_4158,In_4529);
nand U2159 (N_2159,In_1309,In_976);
or U2160 (N_2160,In_1695,In_587);
nand U2161 (N_2161,In_4160,In_2443);
or U2162 (N_2162,In_4876,In_2783);
xor U2163 (N_2163,In_2112,In_757);
xor U2164 (N_2164,In_3422,In_2392);
and U2165 (N_2165,In_3643,In_2018);
or U2166 (N_2166,In_3821,In_4508);
nor U2167 (N_2167,In_2207,In_1419);
and U2168 (N_2168,In_314,In_4478);
and U2169 (N_2169,In_935,In_1895);
nand U2170 (N_2170,In_181,In_1129);
xnor U2171 (N_2171,In_3795,In_2417);
nor U2172 (N_2172,In_896,In_4703);
or U2173 (N_2173,In_2669,In_959);
xor U2174 (N_2174,In_4287,In_1215);
xor U2175 (N_2175,In_1919,In_3980);
nor U2176 (N_2176,In_4091,In_836);
xor U2177 (N_2177,In_4922,In_1905);
nand U2178 (N_2178,In_4395,In_4430);
nand U2179 (N_2179,In_3022,In_1033);
or U2180 (N_2180,In_3977,In_44);
xnor U2181 (N_2181,In_1653,In_3481);
and U2182 (N_2182,In_3593,In_4069);
xor U2183 (N_2183,In_3256,In_363);
and U2184 (N_2184,In_4369,In_3781);
and U2185 (N_2185,In_4092,In_3051);
and U2186 (N_2186,In_2486,In_755);
or U2187 (N_2187,In_1381,In_379);
xor U2188 (N_2188,In_131,In_4539);
nor U2189 (N_2189,In_393,In_4523);
nand U2190 (N_2190,In_303,In_1953);
nand U2191 (N_2191,In_2481,In_1379);
xor U2192 (N_2192,In_4222,In_1111);
nand U2193 (N_2193,In_2426,In_3074);
and U2194 (N_2194,In_4518,In_4030);
or U2195 (N_2195,In_4683,In_1702);
nor U2196 (N_2196,In_2040,In_1347);
and U2197 (N_2197,In_3132,In_2912);
nand U2198 (N_2198,In_377,In_315);
nand U2199 (N_2199,In_1504,In_1767);
or U2200 (N_2200,In_3951,In_606);
nor U2201 (N_2201,In_3856,In_3464);
xor U2202 (N_2202,In_649,In_1656);
nor U2203 (N_2203,In_3791,In_2685);
nand U2204 (N_2204,In_116,In_1314);
xnor U2205 (N_2205,In_3499,In_21);
nand U2206 (N_2206,In_2074,In_41);
nor U2207 (N_2207,In_2752,In_1840);
xnor U2208 (N_2208,In_4147,In_1537);
nor U2209 (N_2209,In_2325,In_1490);
xor U2210 (N_2210,In_4032,In_3183);
xor U2211 (N_2211,In_2181,In_619);
and U2212 (N_2212,In_1906,In_2400);
nand U2213 (N_2213,In_1614,In_673);
xnor U2214 (N_2214,In_1577,In_427);
or U2215 (N_2215,In_4636,In_2564);
and U2216 (N_2216,In_4788,In_1049);
nand U2217 (N_2217,In_3939,In_1757);
nand U2218 (N_2218,In_3128,In_1012);
and U2219 (N_2219,In_1677,In_2271);
nor U2220 (N_2220,In_2059,In_3211);
nand U2221 (N_2221,In_2512,In_2660);
or U2222 (N_2222,In_1177,In_4183);
or U2223 (N_2223,In_4194,In_2713);
nand U2224 (N_2224,In_2812,In_2217);
and U2225 (N_2225,In_974,In_4836);
xor U2226 (N_2226,In_484,In_2552);
nand U2227 (N_2227,In_3862,In_4548);
and U2228 (N_2228,In_2461,In_1613);
nor U2229 (N_2229,In_381,In_1686);
nor U2230 (N_2230,In_1448,In_2839);
nand U2231 (N_2231,In_3829,In_2768);
or U2232 (N_2232,In_1298,In_1589);
xor U2233 (N_2233,In_710,In_567);
nor U2234 (N_2234,In_1008,In_4203);
or U2235 (N_2235,In_42,In_2728);
or U2236 (N_2236,In_3758,In_3866);
nand U2237 (N_2237,In_1346,In_3025);
and U2238 (N_2238,In_664,In_1928);
nor U2239 (N_2239,In_215,In_171);
and U2240 (N_2240,In_768,In_3557);
nand U2241 (N_2241,In_1117,In_476);
and U2242 (N_2242,In_120,In_3894);
and U2243 (N_2243,In_1138,In_3533);
and U2244 (N_2244,In_18,In_4626);
nand U2245 (N_2245,In_2644,In_4934);
or U2246 (N_2246,In_1936,In_2131);
nand U2247 (N_2247,In_3932,In_2684);
nand U2248 (N_2248,In_1491,In_376);
or U2249 (N_2249,In_1994,In_149);
nor U2250 (N_2250,In_3070,In_3895);
xnor U2251 (N_2251,In_4015,In_2641);
or U2252 (N_2252,In_1397,In_4487);
or U2253 (N_2253,In_4579,In_2733);
and U2254 (N_2254,In_4940,In_4975);
and U2255 (N_2255,In_3857,In_2177);
nor U2256 (N_2256,In_857,In_901);
nand U2257 (N_2257,In_485,In_2739);
nand U2258 (N_2258,In_1488,In_676);
nor U2259 (N_2259,In_860,In_2851);
nor U2260 (N_2260,In_2695,In_3592);
nor U2261 (N_2261,In_3253,In_4795);
nor U2262 (N_2262,In_1617,In_1080);
and U2263 (N_2263,In_686,In_312);
nor U2264 (N_2264,In_3611,In_4647);
nor U2265 (N_2265,In_1867,In_1802);
nor U2266 (N_2266,In_2590,In_3944);
nor U2267 (N_2267,In_3509,In_3941);
nand U2268 (N_2268,In_2470,In_670);
and U2269 (N_2269,In_1863,In_2607);
or U2270 (N_2270,In_392,In_3420);
nand U2271 (N_2271,In_3339,In_4758);
nor U2272 (N_2272,In_3661,In_827);
or U2273 (N_2273,In_2555,In_2014);
nand U2274 (N_2274,In_385,In_3291);
and U2275 (N_2275,In_1882,In_2165);
and U2276 (N_2276,In_4075,In_3409);
or U2277 (N_2277,In_4475,In_3372);
and U2278 (N_2278,In_3082,In_3621);
xnor U2279 (N_2279,In_2017,In_142);
nand U2280 (N_2280,In_4097,In_968);
or U2281 (N_2281,In_1886,In_1131);
or U2282 (N_2282,In_3294,In_4959);
or U2283 (N_2283,In_2058,In_1344);
nor U2284 (N_2284,In_246,In_22);
nor U2285 (N_2285,In_3787,In_147);
nor U2286 (N_2286,In_3624,In_4308);
xnor U2287 (N_2287,In_2671,In_1591);
xor U2288 (N_2288,In_616,In_1834);
nand U2289 (N_2289,In_1544,In_3691);
nor U2290 (N_2290,In_3080,In_3318);
and U2291 (N_2291,In_2029,In_4950);
nor U2292 (N_2292,In_359,In_3837);
and U2293 (N_2293,In_4832,In_4170);
and U2294 (N_2294,In_2736,In_4530);
or U2295 (N_2295,In_2030,In_1755);
xnor U2296 (N_2296,In_1471,In_4376);
nand U2297 (N_2297,In_3030,In_691);
nand U2298 (N_2298,In_4017,In_3707);
or U2299 (N_2299,In_2702,In_2834);
or U2300 (N_2300,In_2061,In_3019);
or U2301 (N_2301,In_2035,In_1004);
xor U2302 (N_2302,In_1560,In_3554);
nand U2303 (N_2303,In_157,In_2376);
xor U2304 (N_2304,In_4512,In_1900);
or U2305 (N_2305,In_4393,In_4392);
or U2306 (N_2306,In_1838,In_2872);
xnor U2307 (N_2307,In_2,In_3126);
and U2308 (N_2308,In_2501,In_3812);
nor U2309 (N_2309,In_1302,In_2828);
or U2310 (N_2310,In_4966,In_2429);
or U2311 (N_2311,In_3312,In_1118);
or U2312 (N_2312,In_3590,In_2938);
xor U2313 (N_2313,In_4887,In_1180);
nor U2314 (N_2314,In_4418,In_1553);
nand U2315 (N_2315,In_2820,In_103);
or U2316 (N_2316,In_2498,In_1386);
or U2317 (N_2317,In_1853,In_493);
and U2318 (N_2318,In_4631,In_4826);
nor U2319 (N_2319,In_2805,In_2158);
xor U2320 (N_2320,In_2975,In_3985);
nor U2321 (N_2321,In_223,In_1959);
nand U2322 (N_2322,In_3343,In_2179);
and U2323 (N_2323,In_1636,In_2136);
nand U2324 (N_2324,In_3549,In_873);
and U2325 (N_2325,In_1842,In_384);
nand U2326 (N_2326,In_1659,In_4470);
xor U2327 (N_2327,In_4462,In_1877);
and U2328 (N_2328,In_3915,In_3243);
xnor U2329 (N_2329,In_2293,In_1418);
nor U2330 (N_2330,In_2567,In_4125);
nor U2331 (N_2331,In_3885,In_3601);
and U2332 (N_2332,In_4371,In_906);
and U2333 (N_2333,In_3259,In_2341);
and U2334 (N_2334,In_2696,In_847);
xor U2335 (N_2335,In_2785,In_2492);
or U2336 (N_2336,In_2869,In_455);
and U2337 (N_2337,In_3112,In_1237);
xor U2338 (N_2338,In_1026,In_4165);
and U2339 (N_2339,In_4538,In_482);
xnor U2340 (N_2340,In_4644,In_3659);
xnor U2341 (N_2341,In_39,In_852);
nand U2342 (N_2342,In_3249,In_4660);
nand U2343 (N_2343,In_2846,In_1924);
nand U2344 (N_2344,In_3431,In_4213);
nand U2345 (N_2345,In_3356,In_717);
nor U2346 (N_2346,In_4148,In_1410);
nor U2347 (N_2347,In_3298,In_3646);
or U2348 (N_2348,In_2617,In_1270);
or U2349 (N_2349,In_3506,In_807);
nor U2350 (N_2350,In_2295,In_2483);
nor U2351 (N_2351,In_348,In_2066);
xor U2352 (N_2352,In_4628,In_3458);
and U2353 (N_2353,In_628,In_682);
xnor U2354 (N_2354,In_4779,In_2709);
xor U2355 (N_2355,In_4115,In_1193);
nor U2356 (N_2356,In_733,In_2773);
nor U2357 (N_2357,In_336,In_4305);
nor U2358 (N_2358,In_1596,In_4118);
and U2359 (N_2359,In_2861,In_3368);
nor U2360 (N_2360,In_600,In_2532);
or U2361 (N_2361,In_4912,In_1352);
xor U2362 (N_2362,In_1433,In_3564);
and U2363 (N_2363,In_2822,In_209);
nor U2364 (N_2364,In_4157,In_1935);
nor U2365 (N_2365,In_1697,In_4065);
nor U2366 (N_2366,In_3819,In_2466);
nor U2367 (N_2367,In_3840,In_3462);
and U2368 (N_2368,In_2934,In_1646);
xor U2369 (N_2369,In_356,In_3813);
nand U2370 (N_2370,In_2348,In_3381);
or U2371 (N_2371,In_3486,In_2499);
nor U2372 (N_2372,In_1427,In_1195);
or U2373 (N_2373,In_1029,In_3623);
xnor U2374 (N_2374,In_2439,In_466);
and U2375 (N_2375,In_2755,In_650);
nor U2376 (N_2376,In_4954,In_3859);
nor U2377 (N_2377,In_1183,In_779);
nand U2378 (N_2378,In_1909,In_972);
nor U2379 (N_2379,In_1050,In_3665);
and U2380 (N_2380,In_1261,In_1201);
and U2381 (N_2381,In_4833,In_1047);
xnor U2382 (N_2382,In_4729,In_57);
nor U2383 (N_2383,In_4711,In_4764);
and U2384 (N_2384,In_1009,In_3045);
nor U2385 (N_2385,In_72,In_2188);
xor U2386 (N_2386,In_1880,In_416);
or U2387 (N_2387,In_91,In_2107);
or U2388 (N_2388,In_3820,In_3093);
xor U2389 (N_2389,In_3190,In_568);
xor U2390 (N_2390,In_2476,In_3121);
nor U2391 (N_2391,In_776,In_3551);
nor U2392 (N_2392,In_4041,In_3494);
nand U2393 (N_2393,In_122,In_1837);
and U2394 (N_2394,In_2976,In_2920);
xnor U2395 (N_2395,In_1974,In_1624);
nor U2396 (N_2396,In_1069,In_994);
xnor U2397 (N_2397,In_3451,In_163);
or U2398 (N_2398,In_1760,In_2215);
nand U2399 (N_2399,In_173,In_4498);
xor U2400 (N_2400,In_3437,In_848);
and U2401 (N_2401,In_1239,In_4343);
xnor U2402 (N_2402,In_4364,In_1492);
nand U2403 (N_2403,In_3556,In_3228);
nor U2404 (N_2404,In_2655,In_3233);
xnor U2405 (N_2405,In_3522,In_4897);
nand U2406 (N_2406,In_1830,In_4825);
and U2407 (N_2407,In_1788,In_534);
nand U2408 (N_2408,In_496,In_1369);
nor U2409 (N_2409,In_1289,In_938);
nand U2410 (N_2410,In_889,In_1169);
xor U2411 (N_2411,In_1232,In_3055);
or U2412 (N_2412,In_114,In_1442);
nor U2413 (N_2413,In_1977,In_3341);
nor U2414 (N_2414,In_4116,In_1954);
xnor U2415 (N_2415,In_113,In_1378);
nor U2416 (N_2416,In_970,In_4234);
nor U2417 (N_2417,In_1315,In_4261);
xor U2418 (N_2418,In_4789,In_4298);
nor U2419 (N_2419,In_69,In_940);
nand U2420 (N_2420,In_2206,In_2332);
nand U2421 (N_2421,In_1791,In_2227);
or U2422 (N_2422,In_327,In_3906);
xnor U2423 (N_2423,In_1051,In_4620);
xnor U2424 (N_2424,In_1884,In_3960);
nand U2425 (N_2425,In_513,In_491);
nor U2426 (N_2426,In_1887,In_4824);
xnor U2427 (N_2427,In_3540,In_1367);
and U2428 (N_2428,In_680,In_4431);
xor U2429 (N_2429,In_221,In_1);
or U2430 (N_2430,In_3428,In_1032);
and U2431 (N_2431,In_3600,In_2553);
and U2432 (N_2432,In_265,In_355);
nand U2433 (N_2433,In_4319,In_2751);
nand U2434 (N_2434,In_4440,In_1786);
xor U2435 (N_2435,In_3212,In_1354);
xnor U2436 (N_2436,In_4692,In_2169);
or U2437 (N_2437,In_2687,In_1851);
and U2438 (N_2438,In_1146,In_4419);
nand U2439 (N_2439,In_1631,In_2054);
nand U2440 (N_2440,In_3878,In_1516);
nor U2441 (N_2441,In_1281,In_1493);
nand U2442 (N_2442,In_1849,In_2108);
or U2443 (N_2443,In_10,In_4425);
nor U2444 (N_2444,In_4133,In_1188);
nor U2445 (N_2445,In_3013,In_4787);
and U2446 (N_2446,In_4812,In_1456);
nand U2447 (N_2447,In_907,In_1468);
or U2448 (N_2448,In_46,In_2980);
nand U2449 (N_2449,In_1509,In_89);
nand U2450 (N_2450,In_4107,In_2247);
xor U2451 (N_2451,In_3094,In_273);
and U2452 (N_2452,In_777,In_4263);
xor U2453 (N_2453,In_4057,In_1735);
xor U2454 (N_2454,In_3084,In_2962);
nor U2455 (N_2455,In_2787,In_4556);
or U2456 (N_2456,In_70,In_2272);
xnor U2457 (N_2457,In_4774,In_4447);
nor U2458 (N_2458,In_797,In_899);
nand U2459 (N_2459,In_2544,In_3204);
nor U2460 (N_2460,In_2240,In_1200);
nand U2461 (N_2461,In_2144,In_3116);
and U2462 (N_2462,In_2193,In_4058);
or U2463 (N_2463,In_29,In_787);
or U2464 (N_2464,In_4043,In_4142);
xor U2465 (N_2465,In_2814,In_739);
nor U2466 (N_2466,In_3739,In_3433);
and U2467 (N_2467,In_4823,In_1661);
nor U2468 (N_2468,In_3715,In_1547);
and U2469 (N_2469,In_429,In_4233);
nor U2470 (N_2470,In_4249,In_2218);
nand U2471 (N_2471,In_4748,In_2191);
or U2472 (N_2472,In_2663,In_235);
nor U2473 (N_2473,In_4587,In_4962);
nand U2474 (N_2474,In_4401,In_1106);
or U2475 (N_2475,In_4921,In_2875);
nor U2476 (N_2476,In_2257,In_4845);
or U2477 (N_2477,In_1435,In_3489);
or U2478 (N_2478,In_2725,In_3654);
and U2479 (N_2479,In_4435,In_4913);
nor U2480 (N_2480,In_3156,In_2019);
nand U2481 (N_2481,In_1025,In_2385);
xor U2482 (N_2482,In_2740,In_798);
nand U2483 (N_2483,In_3581,In_2639);
xnor U2484 (N_2484,In_2741,In_1089);
or U2485 (N_2485,In_3865,In_1848);
and U2486 (N_2486,In_1812,In_2749);
xor U2487 (N_2487,In_4633,In_792);
xnor U2488 (N_2488,In_2806,In_3922);
nand U2489 (N_2489,In_1296,In_3412);
xor U2490 (N_2490,In_2842,In_2230);
nor U2491 (N_2491,In_702,In_835);
xor U2492 (N_2492,In_3511,In_2471);
xor U2493 (N_2493,In_1460,In_1843);
nor U2494 (N_2494,In_1510,In_3006);
and U2495 (N_2495,In_3663,In_4028);
nand U2496 (N_2496,In_1271,In_705);
or U2497 (N_2497,In_4576,In_4214);
and U2498 (N_2498,In_1761,In_761);
or U2499 (N_2499,In_4411,In_1940);
and U2500 (N_2500,N_1224,N_784);
nor U2501 (N_2501,N_2027,N_1652);
nand U2502 (N_2502,N_428,N_1598);
nor U2503 (N_2503,N_1143,N_373);
and U2504 (N_2504,N_934,N_1434);
and U2505 (N_2505,N_2210,N_1268);
or U2506 (N_2506,N_750,N_104);
or U2507 (N_2507,N_1527,N_254);
nand U2508 (N_2508,N_2085,N_1610);
xnor U2509 (N_2509,N_505,N_1428);
or U2510 (N_2510,N_344,N_128);
nand U2511 (N_2511,N_2443,N_1552);
xnor U2512 (N_2512,N_1666,N_1608);
or U2513 (N_2513,N_2097,N_1432);
xor U2514 (N_2514,N_674,N_2006);
nor U2515 (N_2515,N_285,N_1994);
or U2516 (N_2516,N_1635,N_2220);
or U2517 (N_2517,N_501,N_1489);
nand U2518 (N_2518,N_607,N_2264);
and U2519 (N_2519,N_2204,N_2284);
xor U2520 (N_2520,N_2378,N_1396);
or U2521 (N_2521,N_1450,N_882);
xnor U2522 (N_2522,N_54,N_2126);
xor U2523 (N_2523,N_1775,N_1648);
or U2524 (N_2524,N_166,N_1920);
nor U2525 (N_2525,N_2069,N_475);
xnor U2526 (N_2526,N_786,N_1096);
nor U2527 (N_2527,N_1237,N_4);
or U2528 (N_2528,N_358,N_2371);
and U2529 (N_2529,N_534,N_1746);
nand U2530 (N_2530,N_1874,N_1133);
or U2531 (N_2531,N_2002,N_2256);
nand U2532 (N_2532,N_504,N_1767);
or U2533 (N_2533,N_3,N_1938);
or U2534 (N_2534,N_1616,N_486);
or U2535 (N_2535,N_1711,N_1470);
nand U2536 (N_2536,N_1591,N_1424);
or U2537 (N_2537,N_1297,N_2376);
nor U2538 (N_2538,N_325,N_2295);
xor U2539 (N_2539,N_2334,N_1305);
nor U2540 (N_2540,N_2026,N_1828);
nor U2541 (N_2541,N_1100,N_223);
nor U2542 (N_2542,N_1731,N_1211);
nand U2543 (N_2543,N_457,N_1668);
xor U2544 (N_2544,N_2070,N_2494);
nand U2545 (N_2545,N_1600,N_2309);
nand U2546 (N_2546,N_935,N_1567);
xor U2547 (N_2547,N_617,N_1080);
or U2548 (N_2548,N_918,N_958);
or U2549 (N_2549,N_248,N_87);
and U2550 (N_2550,N_2177,N_310);
xor U2551 (N_2551,N_801,N_217);
and U2552 (N_2552,N_435,N_1864);
xor U2553 (N_2553,N_1893,N_1330);
or U2554 (N_2554,N_999,N_2161);
or U2555 (N_2555,N_814,N_1808);
xnor U2556 (N_2556,N_1634,N_239);
nand U2557 (N_2557,N_2482,N_1673);
nor U2558 (N_2558,N_1831,N_1482);
and U2559 (N_2559,N_1622,N_2294);
nand U2560 (N_2560,N_2231,N_2014);
nand U2561 (N_2561,N_2305,N_581);
xor U2562 (N_2562,N_1872,N_1197);
or U2563 (N_2563,N_1764,N_2184);
or U2564 (N_2564,N_1447,N_987);
nor U2565 (N_2565,N_1397,N_641);
nor U2566 (N_2566,N_2235,N_1459);
xor U2567 (N_2567,N_546,N_1559);
nor U2568 (N_2568,N_2083,N_920);
or U2569 (N_2569,N_410,N_1493);
xor U2570 (N_2570,N_2263,N_2268);
nand U2571 (N_2571,N_1366,N_1914);
and U2572 (N_2572,N_2078,N_2318);
nand U2573 (N_2573,N_589,N_1070);
and U2574 (N_2574,N_618,N_762);
xnor U2575 (N_2575,N_1276,N_744);
or U2576 (N_2576,N_1388,N_1431);
nor U2577 (N_2577,N_1316,N_917);
nand U2578 (N_2578,N_889,N_2476);
and U2579 (N_2579,N_694,N_1667);
xor U2580 (N_2580,N_88,N_499);
nor U2581 (N_2581,N_948,N_669);
nor U2582 (N_2582,N_1650,N_1823);
nand U2583 (N_2583,N_2456,N_1761);
and U2584 (N_2584,N_1149,N_594);
or U2585 (N_2585,N_214,N_1871);
nand U2586 (N_2586,N_2003,N_192);
xnor U2587 (N_2587,N_944,N_700);
xnor U2588 (N_2588,N_2306,N_320);
or U2589 (N_2589,N_271,N_1543);
xor U2590 (N_2590,N_2245,N_464);
nor U2591 (N_2591,N_1776,N_1658);
nor U2592 (N_2592,N_1359,N_1429);
nor U2593 (N_2593,N_616,N_2192);
nor U2594 (N_2594,N_2140,N_1346);
and U2595 (N_2595,N_2286,N_516);
and U2596 (N_2596,N_416,N_2466);
nand U2597 (N_2597,N_1819,N_870);
and U2598 (N_2598,N_1075,N_2211);
nor U2599 (N_2599,N_245,N_463);
nand U2600 (N_2600,N_1538,N_35);
and U2601 (N_2601,N_2200,N_562);
or U2602 (N_2602,N_555,N_693);
and U2603 (N_2603,N_2458,N_284);
xor U2604 (N_2604,N_1468,N_1333);
and U2605 (N_2605,N_343,N_429);
xnor U2606 (N_2606,N_1510,N_330);
or U2607 (N_2607,N_728,N_1247);
or U2608 (N_2608,N_129,N_2178);
nor U2609 (N_2609,N_2278,N_800);
and U2610 (N_2610,N_208,N_1354);
nand U2611 (N_2611,N_1970,N_630);
nor U2612 (N_2612,N_1594,N_1645);
and U2613 (N_2613,N_905,N_803);
nor U2614 (N_2614,N_431,N_1875);
or U2615 (N_2615,N_1483,N_1275);
or U2616 (N_2616,N_877,N_400);
or U2617 (N_2617,N_1981,N_1679);
and U2618 (N_2618,N_1602,N_1727);
nand U2619 (N_2619,N_1534,N_238);
xor U2620 (N_2620,N_1323,N_1974);
nor U2621 (N_2621,N_2137,N_2448);
and U2622 (N_2622,N_1671,N_422);
or U2623 (N_2623,N_1439,N_2179);
xor U2624 (N_2624,N_24,N_629);
nor U2625 (N_2625,N_591,N_2285);
xor U2626 (N_2626,N_1982,N_584);
nand U2627 (N_2627,N_676,N_985);
xnor U2628 (N_2628,N_2079,N_211);
nand U2629 (N_2629,N_1628,N_2118);
xor U2630 (N_2630,N_1709,N_717);
or U2631 (N_2631,N_765,N_2174);
and U2632 (N_2632,N_1633,N_1408);
nand U2633 (N_2633,N_368,N_462);
or U2634 (N_2634,N_1751,N_891);
nor U2635 (N_2635,N_2023,N_631);
xnor U2636 (N_2636,N_810,N_1314);
and U2637 (N_2637,N_222,N_646);
or U2638 (N_2638,N_268,N_926);
nand U2639 (N_2639,N_1183,N_157);
nor U2640 (N_2640,N_200,N_610);
nand U2641 (N_2641,N_950,N_1369);
or U2642 (N_2642,N_1490,N_116);
nor U2643 (N_2643,N_1554,N_2359);
xnor U2644 (N_2644,N_433,N_471);
and U2645 (N_2645,N_2410,N_311);
nor U2646 (N_2646,N_1399,N_852);
nor U2647 (N_2647,N_907,N_1094);
nor U2648 (N_2648,N_2317,N_1682);
nand U2649 (N_2649,N_2405,N_1619);
and U2650 (N_2650,N_472,N_409);
xnor U2651 (N_2651,N_2463,N_335);
and U2652 (N_2652,N_2187,N_123);
xor U2653 (N_2653,N_747,N_106);
or U2654 (N_2654,N_1331,N_1599);
nor U2655 (N_2655,N_2375,N_1350);
xor U2656 (N_2656,N_198,N_1206);
nor U2657 (N_2657,N_1843,N_2379);
nand U2658 (N_2658,N_565,N_888);
and U2659 (N_2659,N_841,N_353);
or U2660 (N_2660,N_1779,N_1248);
nor U2661 (N_2661,N_1072,N_59);
xnor U2662 (N_2662,N_533,N_967);
or U2663 (N_2663,N_2416,N_1234);
and U2664 (N_2664,N_390,N_1117);
nor U2665 (N_2665,N_1586,N_1549);
nand U2666 (N_2666,N_1908,N_28);
and U2667 (N_2667,N_2346,N_1945);
and U2668 (N_2668,N_1090,N_845);
nor U2669 (N_2669,N_1193,N_365);
xor U2670 (N_2670,N_1278,N_1896);
nand U2671 (N_2671,N_1380,N_1563);
and U2672 (N_2672,N_2325,N_10);
nand U2673 (N_2673,N_1939,N_1315);
and U2674 (N_2674,N_705,N_201);
nor U2675 (N_2675,N_957,N_708);
nand U2676 (N_2676,N_1318,N_2020);
xor U2677 (N_2677,N_122,N_113);
nor U2678 (N_2678,N_1150,N_1298);
xor U2679 (N_2679,N_58,N_1273);
and U2680 (N_2680,N_394,N_252);
xnor U2681 (N_2681,N_1110,N_178);
xor U2682 (N_2682,N_1400,N_1018);
xnor U2683 (N_2683,N_1593,N_1866);
xor U2684 (N_2684,N_996,N_9);
or U2685 (N_2685,N_1917,N_467);
or U2686 (N_2686,N_529,N_2216);
and U2687 (N_2687,N_1691,N_1925);
nand U2688 (N_2688,N_2066,N_1269);
and U2689 (N_2689,N_1686,N_71);
nand U2690 (N_2690,N_261,N_136);
nor U2691 (N_2691,N_836,N_1);
nand U2692 (N_2692,N_771,N_1267);
xnor U2693 (N_2693,N_1087,N_628);
and U2694 (N_2694,N_470,N_850);
xnor U2695 (N_2695,N_1029,N_1449);
nand U2696 (N_2696,N_2468,N_2195);
or U2697 (N_2697,N_678,N_726);
and U2698 (N_2698,N_1217,N_2253);
nor U2699 (N_2699,N_1550,N_1719);
xor U2700 (N_2700,N_2225,N_2241);
nand U2701 (N_2701,N_2290,N_2428);
or U2702 (N_2702,N_876,N_661);
nor U2703 (N_2703,N_2275,N_1985);
xor U2704 (N_2704,N_2365,N_685);
xnor U2705 (N_2705,N_799,N_234);
or U2706 (N_2706,N_2148,N_61);
or U2707 (N_2707,N_186,N_1791);
nand U2708 (N_2708,N_246,N_1123);
xor U2709 (N_2709,N_1415,N_972);
and U2710 (N_2710,N_2368,N_2158);
xor U2711 (N_2711,N_2064,N_2389);
xor U2712 (N_2712,N_1614,N_2000);
and U2713 (N_2713,N_823,N_2367);
or U2714 (N_2714,N_1730,N_1698);
or U2715 (N_2715,N_18,N_340);
or U2716 (N_2716,N_2121,N_1230);
nand U2717 (N_2717,N_1609,N_489);
nand U2718 (N_2718,N_866,N_2454);
xor U2719 (N_2719,N_1784,N_492);
xor U2720 (N_2720,N_328,N_2355);
nand U2721 (N_2721,N_2082,N_807);
or U2722 (N_2722,N_99,N_1533);
nor U2723 (N_2723,N_183,N_1627);
and U2724 (N_2724,N_449,N_1801);
and U2725 (N_2725,N_356,N_1846);
or U2726 (N_2726,N_1927,N_1502);
xnor U2727 (N_2727,N_1465,N_2009);
xor U2728 (N_2728,N_1371,N_1756);
nor U2729 (N_2729,N_2381,N_2144);
nor U2730 (N_2730,N_2270,N_847);
nand U2731 (N_2731,N_1332,N_176);
nor U2732 (N_2732,N_1855,N_502);
nand U2733 (N_2733,N_1820,N_493);
xnor U2734 (N_2734,N_436,N_1041);
and U2735 (N_2735,N_2203,N_2061);
nand U2736 (N_2736,N_1532,N_1638);
and U2737 (N_2737,N_1947,N_243);
nor U2738 (N_2738,N_2426,N_1888);
and U2739 (N_2739,N_1844,N_2434);
xor U2740 (N_2740,N_1291,N_291);
and U2741 (N_2741,N_1701,N_657);
or U2742 (N_2742,N_1902,N_614);
nand U2743 (N_2743,N_1051,N_2213);
and U2744 (N_2744,N_1969,N_180);
nand U2745 (N_2745,N_484,N_2163);
and U2746 (N_2746,N_709,N_1515);
nor U2747 (N_2747,N_1054,N_2030);
and U2748 (N_2748,N_992,N_1540);
or U2749 (N_2749,N_2304,N_2212);
xnor U2750 (N_2750,N_2360,N_1270);
nor U2751 (N_2751,N_933,N_44);
xnor U2752 (N_2752,N_49,N_2191);
nor U2753 (N_2753,N_1389,N_1996);
nor U2754 (N_2754,N_297,N_568);
or U2755 (N_2755,N_582,N_1977);
nand U2756 (N_2756,N_1215,N_111);
nand U2757 (N_2757,N_858,N_1246);
nand U2758 (N_2758,N_1735,N_542);
or U2759 (N_2759,N_1499,N_2419);
and U2760 (N_2760,N_1623,N_1368);
nand U2761 (N_2761,N_2157,N_2150);
xnor U2762 (N_2762,N_36,N_1148);
or U2763 (N_2763,N_244,N_2433);
nor U2764 (N_2764,N_792,N_830);
nor U2765 (N_2765,N_2234,N_1103);
xor U2766 (N_2766,N_1773,N_1028);
xnor U2767 (N_2767,N_366,N_156);
xnor U2768 (N_2768,N_608,N_417);
xor U2769 (N_2769,N_827,N_715);
or U2770 (N_2770,N_838,N_442);
xnor U2771 (N_2771,N_185,N_100);
and U2772 (N_2772,N_1639,N_622);
or U2773 (N_2773,N_1317,N_1906);
xnor U2774 (N_2774,N_1467,N_1281);
nor U2775 (N_2775,N_2065,N_1975);
and U2776 (N_2776,N_292,N_126);
or U2777 (N_2777,N_2141,N_1107);
nand U2778 (N_2778,N_643,N_1827);
xnor U2779 (N_2779,N_577,N_636);
nand U2780 (N_2780,N_1868,N_2337);
xnor U2781 (N_2781,N_711,N_1320);
nor U2782 (N_2782,N_1463,N_1955);
nand U2783 (N_2783,N_526,N_1363);
xor U2784 (N_2784,N_1976,N_1034);
nand U2785 (N_2785,N_1835,N_1055);
or U2786 (N_2786,N_840,N_307);
and U2787 (N_2787,N_1964,N_2237);
or U2788 (N_2788,N_863,N_1142);
nand U2789 (N_2789,N_357,N_808);
or U2790 (N_2790,N_434,N_1841);
nand U2791 (N_2791,N_2119,N_900);
xnor U2792 (N_2792,N_2228,N_2050);
and U2793 (N_2793,N_1007,N_386);
or U2794 (N_2794,N_655,N_714);
or U2795 (N_2795,N_1595,N_545);
xor U2796 (N_2796,N_1084,N_2138);
xor U2797 (N_2797,N_2056,N_1766);
xnor U2798 (N_2798,N_1024,N_1588);
or U2799 (N_2799,N_599,N_2094);
or U2800 (N_2800,N_488,N_2135);
nor U2801 (N_2801,N_2124,N_161);
xnor U2802 (N_2802,N_783,N_1729);
and U2803 (N_2803,N_1743,N_1294);
nand U2804 (N_2804,N_2394,N_1073);
and U2805 (N_2805,N_1319,N_978);
xor U2806 (N_2806,N_281,N_1857);
and U2807 (N_2807,N_2431,N_1484);
xor U2808 (N_2808,N_1741,N_778);
nor U2809 (N_2809,N_8,N_207);
and U2810 (N_2810,N_1777,N_1916);
xor U2811 (N_2811,N_1068,N_2287);
xor U2812 (N_2812,N_2193,N_602);
or U2813 (N_2813,N_1040,N_569);
and U2814 (N_2814,N_548,N_1264);
nor U2815 (N_2815,N_219,N_1740);
and U2816 (N_2816,N_1241,N_1724);
and U2817 (N_2817,N_773,N_203);
xor U2818 (N_2818,N_627,N_144);
xor U2819 (N_2819,N_1391,N_1834);
nor U2820 (N_2820,N_231,N_418);
and U2821 (N_2821,N_319,N_1462);
nand U2822 (N_2822,N_962,N_1414);
xor U2823 (N_2823,N_52,N_115);
and U2824 (N_2824,N_85,N_559);
and U2825 (N_2825,N_1243,N_202);
and U2826 (N_2826,N_339,N_1647);
xor U2827 (N_2827,N_206,N_984);
xnor U2828 (N_2828,N_495,N_2159);
nor U2829 (N_2829,N_1663,N_1214);
and U2830 (N_2830,N_1669,N_2414);
and U2831 (N_2831,N_2060,N_2139);
nand U2832 (N_2832,N_2156,N_2331);
xor U2833 (N_2833,N_986,N_1056);
nor U2834 (N_2834,N_1733,N_1487);
xnor U2835 (N_2835,N_1548,N_702);
nor U2836 (N_2836,N_1962,N_138);
or U2837 (N_2837,N_415,N_1010);
or U2838 (N_2838,N_2105,N_80);
or U2839 (N_2839,N_857,N_2430);
xnor U2840 (N_2840,N_1886,N_1122);
nor U2841 (N_2841,N_1525,N_2190);
nor U2842 (N_2842,N_1624,N_1002);
or U2843 (N_2843,N_619,N_1009);
and U2844 (N_2844,N_142,N_834);
nand U2845 (N_2845,N_1012,N_258);
or U2846 (N_2846,N_84,N_2199);
and U2847 (N_2847,N_33,N_1407);
xor U2848 (N_2848,N_1566,N_1889);
nor U2849 (N_2849,N_2122,N_1421);
and U2850 (N_2850,N_1046,N_1960);
or U2851 (N_2851,N_1426,N_2096);
nand U2852 (N_2852,N_1911,N_1180);
and U2853 (N_2853,N_898,N_2129);
xnor U2854 (N_2854,N_375,N_820);
nand U2855 (N_2855,N_2080,N_1477);
xor U2856 (N_2856,N_687,N_1876);
and U2857 (N_2857,N_324,N_420);
and U2858 (N_2858,N_532,N_1692);
or U2859 (N_2859,N_1696,N_1714);
xor U2860 (N_2860,N_355,N_2391);
nand U2861 (N_2861,N_27,N_259);
nand U2862 (N_2862,N_1725,N_518);
or U2863 (N_2863,N_1703,N_498);
or U2864 (N_2864,N_155,N_1192);
xor U2865 (N_2865,N_2266,N_556);
nand U2866 (N_2866,N_531,N_345);
nand U2867 (N_2867,N_1071,N_2173);
and U2868 (N_2868,N_322,N_2068);
or U2869 (N_2869,N_1514,N_131);
or U2870 (N_2870,N_197,N_2219);
xor U2871 (N_2871,N_1390,N_1349);
or U2872 (N_2872,N_2429,N_1959);
and U2873 (N_2873,N_2147,N_1812);
or U2874 (N_2874,N_1219,N_1047);
or U2875 (N_2875,N_485,N_1473);
and U2876 (N_2876,N_2320,N_1113);
or U2877 (N_2877,N_774,N_408);
xnor U2878 (N_2878,N_326,N_1615);
nand U2879 (N_2879,N_963,N_1677);
or U2880 (N_2880,N_1157,N_2073);
or U2881 (N_2881,N_1572,N_1901);
nor U2882 (N_2882,N_2473,N_1367);
and U2883 (N_2883,N_1971,N_327);
nor U2884 (N_2884,N_2108,N_1111);
and U2885 (N_2885,N_1718,N_2262);
and U2886 (N_2886,N_2182,N_110);
nor U2887 (N_2887,N_26,N_1092);
xor U2888 (N_2888,N_2267,N_817);
or U2889 (N_2889,N_2442,N_1444);
nor U2890 (N_2890,N_1995,N_181);
xor U2891 (N_2891,N_43,N_1941);
nand U2892 (N_2892,N_673,N_121);
xor U2893 (N_2893,N_1536,N_2090);
xor U2894 (N_2894,N_973,N_768);
and U2895 (N_2895,N_1233,N_2353);
and U2896 (N_2896,N_1220,N_2438);
nor U2897 (N_2897,N_1576,N_405);
nand U2898 (N_2898,N_64,N_2049);
xor U2899 (N_2899,N_2092,N_1675);
xor U2900 (N_2900,N_143,N_1023);
xnor U2901 (N_2901,N_1963,N_2288);
nor U2902 (N_2902,N_1937,N_1528);
and U2903 (N_2903,N_2397,N_103);
and U2904 (N_2904,N_1286,N_1457);
nand U2905 (N_2905,N_2497,N_2424);
nand U2906 (N_2906,N_404,N_1423);
nand U2907 (N_2907,N_242,N_1553);
nand U2908 (N_2908,N_1393,N_20);
nor U2909 (N_2909,N_1555,N_474);
xor U2910 (N_2910,N_98,N_440);
nand U2911 (N_2911,N_1951,N_1285);
and U2912 (N_2912,N_1762,N_1607);
nor U2913 (N_2913,N_437,N_510);
and U2914 (N_2914,N_1057,N_1585);
xnor U2915 (N_2915,N_380,N_848);
and U2916 (N_2916,N_797,N_2277);
nor U2917 (N_2917,N_1678,N_522);
or U2918 (N_2918,N_364,N_1155);
and U2919 (N_2919,N_1693,N_1817);
or U2920 (N_2920,N_2233,N_2418);
xnor U2921 (N_2921,N_1918,N_2180);
xor U2922 (N_2922,N_1999,N_1411);
and U2923 (N_2923,N_1038,N_511);
xnor U2924 (N_2924,N_2441,N_1605);
nor U2925 (N_2925,N_1385,N_1929);
nand U2926 (N_2926,N_2453,N_1509);
or U2927 (N_2927,N_1744,N_1562);
nand U2928 (N_2928,N_452,N_162);
or U2929 (N_2929,N_372,N_2462);
xor U2930 (N_2930,N_645,N_277);
nand U2931 (N_2931,N_300,N_301);
nor U2932 (N_2932,N_1209,N_1919);
xor U2933 (N_2933,N_1335,N_1341);
and U2934 (N_2934,N_249,N_1728);
nor U2935 (N_2935,N_1479,N_1300);
nor U2936 (N_2936,N_777,N_2425);
nand U2937 (N_2937,N_1485,N_1620);
nand U2938 (N_2938,N_47,N_1505);
nand U2939 (N_2939,N_1655,N_218);
or U2940 (N_2940,N_1636,N_2293);
or U2941 (N_2941,N_1398,N_854);
nand U2942 (N_2942,N_1419,N_412);
and U2943 (N_2943,N_1845,N_95);
or U2944 (N_2944,N_770,N_2062);
nor U2945 (N_2945,N_1991,N_1058);
or U2946 (N_2946,N_1076,N_215);
nor U2947 (N_2947,N_338,N_1089);
and U2948 (N_2948,N_590,N_2155);
and U2949 (N_2949,N_1461,N_1603);
and U2950 (N_2950,N_1182,N_1565);
xnor U2951 (N_2951,N_1494,N_1417);
xor U2952 (N_2952,N_561,N_699);
and U2953 (N_2953,N_1942,N_1880);
and U2954 (N_2954,N_818,N_583);
xnor U2955 (N_2955,N_2324,N_2340);
nor U2956 (N_2956,N_2384,N_1309);
xnor U2957 (N_2957,N_703,N_1687);
or U2958 (N_2958,N_2089,N_2036);
nand U2959 (N_2959,N_2127,N_735);
nand U2960 (N_2960,N_1228,N_868);
and U2961 (N_2961,N_109,N_753);
nor U2962 (N_2962,N_2004,N_1838);
nor U2963 (N_2963,N_633,N_459);
and U2964 (N_2964,N_939,N_2252);
nor U2965 (N_2965,N_1114,N_1749);
xor U2966 (N_2966,N_147,N_552);
nor U2967 (N_2967,N_781,N_1153);
and U2968 (N_2968,N_141,N_2205);
xnor U2969 (N_2969,N_2383,N_334);
xor U2970 (N_2970,N_2313,N_831);
or U2971 (N_2971,N_1587,N_1944);
nor U2972 (N_2972,N_273,N_1427);
and U2973 (N_2973,N_1859,N_153);
or U2974 (N_2974,N_875,N_1227);
nor U2975 (N_2975,N_13,N_824);
xnor U2976 (N_2976,N_2257,N_1934);
and U2977 (N_2977,N_160,N_1125);
nand U2978 (N_2978,N_1581,N_2274);
nor U2979 (N_2979,N_968,N_943);
xnor U2980 (N_2980,N_1033,N_289);
or U2981 (N_2981,N_253,N_1402);
xnor U2982 (N_2982,N_1795,N_294);
xnor U2983 (N_2983,N_1005,N_367);
nand U2984 (N_2984,N_25,N_974);
nor U2985 (N_2985,N_1558,N_1127);
or U2986 (N_2986,N_1672,N_2243);
xor U2987 (N_2987,N_2040,N_2186);
or U2988 (N_2988,N_1837,N_839);
or U2989 (N_2989,N_2168,N_554);
and U2990 (N_2990,N_887,N_893);
nor U2991 (N_2991,N_361,N_74);
nand U2992 (N_2992,N_2486,N_689);
nand U2993 (N_2993,N_132,N_1283);
xor U2994 (N_2994,N_212,N_829);
xor U2995 (N_2995,N_1334,N_1912);
or U2996 (N_2996,N_480,N_2250);
nand U2997 (N_2997,N_2460,N_309);
xor U2998 (N_2998,N_407,N_1524);
xnor U2999 (N_2999,N_2232,N_2133);
nand U3000 (N_3000,N_1832,N_154);
xor U3001 (N_3001,N_1966,N_1061);
nand U3002 (N_3002,N_787,N_2114);
nand U3003 (N_3003,N_2478,N_426);
and U3004 (N_3004,N_1077,N_563);
and U3005 (N_3005,N_906,N_1304);
xnor U3006 (N_3006,N_403,N_107);
or U3007 (N_3007,N_1685,N_2017);
nor U3008 (N_3008,N_2132,N_1265);
nand U3009 (N_3009,N_751,N_698);
xnor U3010 (N_3010,N_514,N_1203);
or U3011 (N_3011,N_587,N_826);
xnor U3012 (N_3012,N_1049,N_2055);
or U3013 (N_3013,N_1106,N_2103);
or U3014 (N_3014,N_2115,N_1858);
and U3015 (N_3015,N_1337,N_2308);
nor U3016 (N_3016,N_224,N_1611);
nand U3017 (N_3017,N_1852,N_660);
nand U3018 (N_3018,N_48,N_1850);
nand U3019 (N_3019,N_2393,N_979);
and U3020 (N_3020,N_1095,N_2314);
and U3021 (N_3021,N_1798,N_2330);
and U3022 (N_3022,N_1456,N_1438);
xor U3023 (N_3023,N_956,N_1646);
nand U3024 (N_3024,N_1568,N_479);
xor U3025 (N_3025,N_746,N_537);
and U3026 (N_3026,N_2423,N_67);
xor U3027 (N_3027,N_2104,N_72);
and U3028 (N_3028,N_1120,N_1644);
nor U3029 (N_3029,N_2217,N_1694);
or U3030 (N_3030,N_913,N_1877);
and U3031 (N_3031,N_2471,N_1252);
nor U3032 (N_3032,N_815,N_874);
nor U3033 (N_3033,N_1968,N_2189);
or U3034 (N_3034,N_881,N_1141);
or U3035 (N_3035,N_496,N_460);
and U3036 (N_3036,N_894,N_482);
xnor U3037 (N_3037,N_1516,N_2054);
nor U3038 (N_3038,N_1905,N_1519);
nand U3039 (N_3039,N_2053,N_11);
or U3040 (N_3040,N_789,N_1360);
and U3041 (N_3041,N_377,N_1043);
nor U3042 (N_3042,N_2008,N_1940);
and U3043 (N_3043,N_649,N_2215);
and U3044 (N_3044,N_1190,N_2154);
nand U3045 (N_3045,N_659,N_1355);
and U3046 (N_3046,N_1539,N_1452);
xnor U3047 (N_3047,N_2239,N_578);
and U3048 (N_3048,N_2197,N_1003);
and U3049 (N_3049,N_235,N_1121);
xnor U3050 (N_3050,N_2338,N_1723);
nor U3051 (N_3051,N_1307,N_527);
nor U3052 (N_3052,N_1736,N_29);
nand U3053 (N_3053,N_146,N_1664);
nor U3054 (N_3054,N_2319,N_1923);
and U3055 (N_3055,N_1261,N_1763);
and U3056 (N_3056,N_2296,N_1546);
and U3057 (N_3057,N_2439,N_1659);
nand U3058 (N_3058,N_1956,N_896);
nor U3059 (N_3059,N_118,N_2349);
xnor U3060 (N_3060,N_1684,N_164);
nor U3061 (N_3061,N_1474,N_1425);
or U3062 (N_3062,N_615,N_1979);
and U3063 (N_3063,N_2035,N_1198);
and U3064 (N_3064,N_1132,N_2136);
nor U3065 (N_3065,N_908,N_2072);
nand U3066 (N_3066,N_57,N_1258);
nor U3067 (N_3067,N_1027,N_2269);
nand U3068 (N_3068,N_1375,N_1151);
xor U3069 (N_3069,N_419,N_2450);
xor U3070 (N_3070,N_1287,N_886);
nand U3071 (N_3071,N_954,N_1204);
or U3072 (N_3072,N_1815,N_448);
or U3073 (N_3073,N_221,N_134);
and U3074 (N_3074,N_1471,N_860);
or U3075 (N_3075,N_736,N_1695);
xor U3076 (N_3076,N_988,N_1327);
xor U3077 (N_3077,N_1903,N_105);
and U3078 (N_3078,N_2093,N_1022);
and U3079 (N_3079,N_1881,N_662);
nand U3080 (N_3080,N_1582,N_233);
xnor U3081 (N_3081,N_1401,N_1469);
or U3082 (N_3082,N_1706,N_251);
nand U3083 (N_3083,N_1032,N_216);
xor U3084 (N_3084,N_272,N_7);
xnor U3085 (N_3085,N_1311,N_1322);
and U3086 (N_3086,N_1992,N_1935);
and U3087 (N_3087,N_758,N_177);
nor U3088 (N_3088,N_2160,N_696);
and U3089 (N_3089,N_864,N_2392);
nor U3090 (N_3090,N_299,N_2297);
and U3091 (N_3091,N_454,N_2445);
xor U3092 (N_3092,N_1455,N_1232);
or U3093 (N_3093,N_1313,N_1913);
and U3094 (N_3094,N_1171,N_269);
and U3095 (N_3095,N_575,N_2407);
nand U3096 (N_3096,N_1894,N_225);
xnor U3097 (N_3097,N_1816,N_2123);
and U3098 (N_3098,N_1755,N_387);
nor U3099 (N_3099,N_966,N_1892);
or U3100 (N_3100,N_928,N_2404);
xor U3101 (N_3101,N_2299,N_897);
or U3102 (N_3102,N_1067,N_278);
xor U3103 (N_3103,N_1272,N_2229);
nor U3104 (N_3104,N_293,N_1356);
or U3105 (N_3105,N_1422,N_1683);
and U3106 (N_3106,N_140,N_1606);
xor U3107 (N_3107,N_871,N_256);
and U3108 (N_3108,N_779,N_2492);
and U3109 (N_3109,N_539,N_82);
and U3110 (N_3110,N_949,N_1557);
nand U3111 (N_3111,N_2051,N_2432);
and U3112 (N_3112,N_1943,N_392);
nand U3113 (N_3113,N_804,N_1236);
and U3114 (N_3114,N_124,N_1653);
nor U3115 (N_3115,N_2348,N_2401);
or U3116 (N_3116,N_1365,N_2301);
xnor U3117 (N_3117,N_916,N_1822);
or U3118 (N_3118,N_1240,N_179);
nand U3119 (N_3119,N_1697,N_1099);
and U3120 (N_3120,N_302,N_30);
nand U3121 (N_3121,N_2013,N_363);
nor U3122 (N_3122,N_1172,N_1098);
nor U3123 (N_3123,N_718,N_2007);
or U3124 (N_3124,N_19,N_952);
nor U3125 (N_3125,N_31,N_1662);
xnor U3126 (N_3126,N_2447,N_2236);
xnor U3127 (N_3127,N_1184,N_1511);
and U3128 (N_3128,N_2125,N_209);
xnor U3129 (N_3129,N_1993,N_2045);
nand U3130 (N_3130,N_1921,N_686);
and U3131 (N_3131,N_666,N_805);
nand U3132 (N_3132,N_1904,N_1949);
or U3133 (N_3133,N_1804,N_1481);
or U3134 (N_3134,N_521,N_1329);
and U3135 (N_3135,N_2461,N_1464);
and U3136 (N_3136,N_1174,N_79);
xnor U3137 (N_3137,N_1048,N_304);
or U3138 (N_3138,N_2100,N_1613);
or U3139 (N_3139,N_550,N_1021);
nor U3140 (N_3140,N_2421,N_1175);
xnor U3141 (N_3141,N_1218,N_1440);
or U3142 (N_3142,N_66,N_1336);
nand U3143 (N_3143,N_1475,N_127);
xor U3144 (N_3144,N_1179,N_809);
nand U3145 (N_3145,N_1436,N_1409);
xnor U3146 (N_3146,N_535,N_2350);
nand U3147 (N_3147,N_2489,N_1556);
nor U3148 (N_3148,N_855,N_724);
nand U3149 (N_3149,N_145,N_1416);
nor U3150 (N_3150,N_1063,N_940);
or U3151 (N_3151,N_1310,N_2399);
and U3152 (N_3152,N_112,N_595);
xor U3153 (N_3153,N_169,N_1689);
and U3154 (N_3154,N_1164,N_1091);
nor U3155 (N_3155,N_86,N_1321);
nor U3156 (N_3156,N_1166,N_2395);
xnor U3157 (N_3157,N_1231,N_588);
or U3158 (N_3158,N_842,N_989);
and U3159 (N_3159,N_1074,N_232);
nand U3160 (N_3160,N_980,N_439);
xor U3161 (N_3161,N_664,N_2152);
or U3162 (N_3162,N_2106,N_453);
and U3163 (N_3163,N_2031,N_55);
nor U3164 (N_3164,N_1079,N_1025);
or U3165 (N_3165,N_2223,N_331);
nand U3166 (N_3166,N_316,N_1053);
xnor U3167 (N_3167,N_567,N_69);
and U3168 (N_3168,N_371,N_795);
xnor U3169 (N_3169,N_1069,N_228);
xnor U3170 (N_3170,N_2099,N_653);
nor U3171 (N_3171,N_295,N_890);
xor U3172 (N_3172,N_682,N_1742);
or U3173 (N_3173,N_1760,N_1458);
and U3174 (N_3174,N_1802,N_572);
nor U3175 (N_3175,N_1786,N_362);
nand U3176 (N_3176,N_2312,N_1083);
nand U3177 (N_3177,N_2091,N_930);
or U3178 (N_3178,N_1601,N_1825);
nor U3179 (N_3179,N_89,N_39);
nor U3180 (N_3180,N_92,N_6);
nand U3181 (N_3181,N_396,N_2498);
nor U3182 (N_3182,N_743,N_1328);
nand U3183 (N_3183,N_1097,N_2185);
xor U3184 (N_3184,N_1262,N_1177);
nor U3185 (N_3185,N_2333,N_263);
and U3186 (N_3186,N_276,N_1488);
xor U3187 (N_3187,N_1418,N_998);
and U3188 (N_3188,N_279,N_2339);
or U3189 (N_3189,N_1570,N_869);
nand U3190 (N_3190,N_1271,N_2409);
nand U3191 (N_3191,N_2449,N_1078);
and U3192 (N_3192,N_929,N_880);
nor U3193 (N_3193,N_1052,N_776);
nand U3194 (N_3194,N_2176,N_626);
and U3195 (N_3195,N_656,N_1898);
or U3196 (N_3196,N_1140,N_1681);
and U3197 (N_3197,N_187,N_2477);
xnor U3198 (N_3198,N_1376,N_1460);
and U3199 (N_3199,N_638,N_393);
xnor U3200 (N_3200,N_2075,N_904);
xor U3201 (N_3201,N_648,N_1961);
and U3202 (N_3202,N_650,N_378);
or U3203 (N_3203,N_706,N_547);
xnor U3204 (N_3204,N_1946,N_1035);
xor U3205 (N_3205,N_1101,N_257);
and U3206 (N_3206,N_2117,N_184);
and U3207 (N_3207,N_399,N_2012);
nand U3208 (N_3208,N_931,N_102);
nor U3209 (N_3209,N_598,N_1936);
or U3210 (N_3210,N_790,N_859);
or U3211 (N_3211,N_1560,N_1535);
and U3212 (N_3212,N_159,N_1710);
and U3213 (N_3213,N_229,N_2402);
nor U3214 (N_3214,N_1382,N_2248);
xor U3215 (N_3215,N_1520,N_1910);
and U3216 (N_3216,N_1042,N_959);
nand U3217 (N_3217,N_1930,N_2411);
nor U3218 (N_3218,N_321,N_2033);
xnor U3219 (N_3219,N_1102,N_2095);
and U3220 (N_3220,N_444,N_148);
nand U3221 (N_3221,N_2281,N_1144);
nand U3222 (N_3222,N_1308,N_476);
and U3223 (N_3223,N_960,N_1803);
or U3224 (N_3224,N_1170,N_704);
or U3225 (N_3225,N_2403,N_170);
xnor U3226 (N_3226,N_1242,N_658);
nand U3227 (N_3227,N_2029,N_837);
nand U3228 (N_3228,N_2321,N_2271);
or U3229 (N_3229,N_1435,N_2328);
or U3230 (N_3230,N_2088,N_1873);
nand U3231 (N_3231,N_1019,N_573);
and U3232 (N_3232,N_432,N_2081);
and U3233 (N_3233,N_2153,N_2345);
and U3234 (N_3234,N_873,N_2249);
nor U3235 (N_3235,N_1342,N_1497);
xnor U3236 (N_3236,N_1478,N_538);
nor U3237 (N_3237,N_1783,N_2172);
xor U3238 (N_3238,N_2194,N_351);
and U3239 (N_3239,N_600,N_2351);
and U3240 (N_3240,N_135,N_793);
xnor U3241 (N_3241,N_2261,N_2128);
and U3242 (N_3242,N_91,N_303);
and U3243 (N_3243,N_1299,N_849);
nand U3244 (N_3244,N_2071,N_305);
xor U3245 (N_3245,N_2221,N_1406);
and U3246 (N_3246,N_1990,N_1472);
nor U3247 (N_3247,N_1790,N_189);
and U3248 (N_3248,N_652,N_1357);
or U3249 (N_3249,N_1720,N_812);
and U3250 (N_3250,N_56,N_625);
nor U3251 (N_3251,N_942,N_1296);
nor U3252 (N_3252,N_1793,N_2043);
or U3253 (N_3253,N_16,N_1501);
nand U3254 (N_3254,N_759,N_1093);
nor U3255 (N_3255,N_270,N_283);
xor U3256 (N_3256,N_2452,N_1712);
or U3257 (N_3257,N_519,N_447);
and U3258 (N_3258,N_369,N_152);
xor U3259 (N_3259,N_1109,N_1173);
xor U3260 (N_3260,N_2107,N_1986);
and U3261 (N_3261,N_1661,N_149);
xnor U3262 (N_3262,N_1250,N_990);
nor U3263 (N_3263,N_503,N_597);
xnor U3264 (N_3264,N_1626,N_2015);
and U3265 (N_3265,N_1721,N_720);
or U3266 (N_3266,N_1748,N_60);
xor U3267 (N_3267,N_1163,N_508);
and U3268 (N_3268,N_2116,N_37);
nor U3269 (N_3269,N_34,N_909);
and U3270 (N_3270,N_1221,N_692);
or U3271 (N_3271,N_1290,N_2459);
nor U3272 (N_3272,N_1797,N_1708);
or U3273 (N_3273,N_1226,N_1448);
nor U3274 (N_3274,N_2005,N_425);
nand U3275 (N_3275,N_1280,N_346);
and U3276 (N_3276,N_2048,N_2214);
and U3277 (N_3277,N_1799,N_1772);
and U3278 (N_3278,N_1826,N_507);
nand U3279 (N_3279,N_2451,N_1840);
nor U3280 (N_3280,N_2039,N_195);
xnor U3281 (N_3281,N_438,N_1301);
nand U3282 (N_3282,N_729,N_1088);
and U3283 (N_3283,N_1351,N_1135);
xnor U3284 (N_3284,N_2362,N_1085);
or U3285 (N_3285,N_348,N_1138);
xor U3286 (N_3286,N_1118,N_2145);
nor U3287 (N_3287,N_483,N_450);
and U3288 (N_3288,N_382,N_846);
or U3289 (N_3289,N_1251,N_1394);
nor U3290 (N_3290,N_2188,N_308);
nand U3291 (N_3291,N_635,N_1000);
or U3292 (N_3292,N_468,N_1915);
nand U3293 (N_3293,N_2406,N_167);
and U3294 (N_3294,N_596,N_117);
and U3295 (N_3295,N_2224,N_2335);
nand U3296 (N_3296,N_2044,N_2170);
xnor U3297 (N_3297,N_2440,N_2332);
and U3298 (N_3298,N_632,N_1769);
xnor U3299 (N_3299,N_862,N_2242);
or U3300 (N_3300,N_1412,N_63);
or U3301 (N_3301,N_1632,N_1665);
and U3302 (N_3302,N_2,N_2260);
xnor U3303 (N_3303,N_1325,N_1324);
and U3304 (N_3304,N_199,N_2364);
and U3305 (N_3305,N_2427,N_1891);
and U3306 (N_3306,N_769,N_923);
and U3307 (N_3307,N_2455,N_323);
and U3308 (N_3308,N_2420,N_2283);
and U3309 (N_3309,N_668,N_722);
and U3310 (N_3310,N_1284,N_2254);
xnor U3311 (N_3311,N_1011,N_2142);
xor U3312 (N_3312,N_843,N_794);
xor U3313 (N_3313,N_1878,N_912);
xnor U3314 (N_3314,N_910,N_2098);
xor U3315 (N_3315,N_932,N_1529);
nor U3316 (N_3316,N_2206,N_1948);
nand U3317 (N_3317,N_477,N_509);
nor U3318 (N_3318,N_1199,N_1200);
nor U3319 (N_3319,N_2258,N_1617);
and U3320 (N_3320,N_2422,N_1115);
nand U3321 (N_3321,N_1154,N_1403);
nor U3322 (N_3322,N_2292,N_120);
and U3323 (N_3323,N_712,N_354);
and U3324 (N_3324,N_1386,N_642);
nor U3325 (N_3325,N_752,N_250);
or U3326 (N_3326,N_2315,N_915);
nand U3327 (N_3327,N_816,N_2181);
nor U3328 (N_3328,N_997,N_574);
nand U3329 (N_3329,N_756,N_766);
nor U3330 (N_3330,N_255,N_376);
nand U3331 (N_3331,N_1008,N_388);
or U3332 (N_3332,N_1800,N_1064);
nor U3333 (N_3333,N_634,N_899);
xor U3334 (N_3334,N_798,N_191);
nand U3335 (N_3335,N_1129,N_1781);
or U3336 (N_3336,N_1688,N_1523);
xor U3337 (N_3337,N_1805,N_1924);
nor U3338 (N_3338,N_515,N_1500);
nand U3339 (N_3339,N_733,N_188);
nor U3340 (N_3340,N_914,N_754);
or U3341 (N_3341,N_1378,N_2058);
nand U3342 (N_3342,N_1690,N_782);
nor U3343 (N_3343,N_740,N_32);
nor U3344 (N_3344,N_2479,N_730);
and U3345 (N_3345,N_23,N_517);
xnor U3346 (N_3346,N_1722,N_1732);
nor U3347 (N_3347,N_165,N_1105);
xor U3348 (N_3348,N_1235,N_1186);
nor U3349 (N_3349,N_760,N_329);
xnor U3350 (N_3350,N_1965,N_788);
or U3351 (N_3351,N_2109,N_697);
nand U3352 (N_3352,N_2323,N_2021);
or U3353 (N_3353,N_1383,N_1384);
nor U3354 (N_3354,N_2322,N_2481);
or U3355 (N_3355,N_1108,N_1128);
and U3356 (N_3356,N_780,N_609);
or U3357 (N_3357,N_1037,N_1124);
or U3358 (N_3358,N_947,N_1745);
xnor U3359 (N_3359,N_1578,N_1162);
nor U3360 (N_3360,N_951,N_1116);
or U3361 (N_3361,N_342,N_1806);
and U3362 (N_3362,N_1597,N_991);
nand U3363 (N_3363,N_1404,N_1774);
and U3364 (N_3364,N_901,N_2475);
and U3365 (N_3365,N_2276,N_2028);
and U3366 (N_3366,N_1702,N_1312);
nand U3367 (N_3367,N_551,N_1853);
or U3368 (N_3368,N_637,N_2162);
nand U3369 (N_3369,N_173,N_1674);
nor U3370 (N_3370,N_721,N_406);
and U3371 (N_3371,N_267,N_1569);
and U3372 (N_3372,N_1491,N_1641);
nand U3373 (N_3373,N_2342,N_671);
and U3374 (N_3374,N_644,N_2435);
xor U3375 (N_3375,N_576,N_1358);
nand U3376 (N_3376,N_1026,N_2025);
and U3377 (N_3377,N_349,N_2087);
nand U3378 (N_3378,N_2032,N_553);
and U3379 (N_3379,N_1338,N_1978);
nand U3380 (N_3380,N_1013,N_601);
nor U3381 (N_3381,N_2067,N_2474);
nor U3382 (N_3382,N_1890,N_1030);
xnor U3383 (N_3383,N_1860,N_1065);
nand U3384 (N_3384,N_1158,N_543);
nand U3385 (N_3385,N_1789,N_287);
nor U3386 (N_3386,N_266,N_70);
nor U3387 (N_3387,N_313,N_964);
and U3388 (N_3388,N_1020,N_158);
and U3389 (N_3389,N_612,N_2412);
nor U3390 (N_3390,N_902,N_1082);
nand U3391 (N_3391,N_220,N_1547);
or U3392 (N_3392,N_90,N_1495);
nor U3393 (N_3393,N_469,N_38);
nand U3394 (N_3394,N_1340,N_466);
nor U3395 (N_3395,N_336,N_1066);
nor U3396 (N_3396,N_2240,N_1134);
xnor U3397 (N_3397,N_1631,N_679);
and U3398 (N_3398,N_1196,N_2247);
xor U3399 (N_3399,N_879,N_1957);
xnor U3400 (N_3400,N_1583,N_1796);
nand U3401 (N_3401,N_1952,N_1517);
xor U3402 (N_3402,N_1201,N_1185);
and U3403 (N_3403,N_2207,N_22);
nor U3404 (N_3404,N_1289,N_2047);
and U3405 (N_3405,N_1637,N_314);
nor U3406 (N_3406,N_133,N_288);
nand U3407 (N_3407,N_2374,N_227);
xor U3408 (N_3408,N_395,N_2018);
or U3409 (N_3409,N_226,N_665);
xnor U3410 (N_3410,N_982,N_1551);
xor U3411 (N_3411,N_1207,N_2227);
nand U3412 (N_3412,N_1716,N_385);
nor U3413 (N_3413,N_620,N_1680);
and U3414 (N_3414,N_14,N_1160);
and U3415 (N_3415,N_707,N_2146);
nor U3416 (N_3416,N_2499,N_1754);
or U3417 (N_3417,N_995,N_1884);
nor U3418 (N_3418,N_757,N_1792);
nor U3419 (N_3419,N_1119,N_1577);
and U3420 (N_3420,N_1293,N_520);
nor U3421 (N_3421,N_1897,N_1542);
or U3422 (N_3422,N_825,N_1347);
nand U3423 (N_3423,N_45,N_2390);
nor U3424 (N_3424,N_884,N_1050);
nor U3425 (N_3425,N_1496,N_1787);
or U3426 (N_3426,N_512,N_75);
nor U3427 (N_3427,N_119,N_2464);
nand U3428 (N_3428,N_101,N_2001);
xor U3429 (N_3429,N_835,N_1480);
xnor U3430 (N_3430,N_684,N_236);
and U3431 (N_3431,N_1530,N_1446);
or U3432 (N_3432,N_1362,N_1466);
xnor U3433 (N_3433,N_2289,N_2046);
nor U3434 (N_3434,N_1205,N_802);
or U3435 (N_3435,N_772,N_2446);
nand U3436 (N_3436,N_1503,N_1654);
and U3437 (N_3437,N_374,N_1984);
nand U3438 (N_3438,N_204,N_1814);
or U3439 (N_3439,N_506,N_1112);
or U3440 (N_3440,N_1778,N_1381);
nor U3441 (N_3441,N_925,N_2372);
or U3442 (N_3442,N_603,N_993);
nand U3443 (N_3443,N_2291,N_981);
xnor U3444 (N_3444,N_40,N_883);
nand U3445 (N_3445,N_1997,N_1788);
and U3446 (N_3446,N_1571,N_15);
and U3447 (N_3447,N_481,N_1352);
nor U3448 (N_3448,N_639,N_961);
nor U3449 (N_3449,N_2165,N_163);
nor U3450 (N_3450,N_2310,N_1045);
nand U3451 (N_3451,N_491,N_1713);
xnor U3452 (N_3452,N_623,N_1295);
nor U3453 (N_3453,N_490,N_494);
nor U3454 (N_3454,N_359,N_1830);
or U3455 (N_3455,N_65,N_2316);
nor U3456 (N_3456,N_585,N_274);
nand U3457 (N_3457,N_2329,N_2396);
xnor U3458 (N_3458,N_1131,N_175);
nand U3459 (N_3459,N_333,N_1768);
or U3460 (N_3460,N_1782,N_1883);
nand U3461 (N_3461,N_821,N_1856);
and U3462 (N_3462,N_286,N_139);
nand U3463 (N_3463,N_1739,N_443);
or U3464 (N_3464,N_1345,N_384);
xor U3465 (N_3465,N_2120,N_247);
nor U3466 (N_3466,N_523,N_461);
xnor U3467 (N_3467,N_114,N_2273);
and U3468 (N_3468,N_1372,N_1590);
nand U3469 (N_3469,N_1303,N_1642);
nor U3470 (N_3470,N_1704,N_811);
xor U3471 (N_3471,N_2011,N_424);
or U3472 (N_3472,N_2496,N_193);
and U3473 (N_3473,N_1044,N_716);
and U3474 (N_3474,N_1392,N_1451);
and U3475 (N_3475,N_306,N_878);
or U3476 (N_3476,N_73,N_2467);
and U3477 (N_3477,N_2057,N_2495);
nor U3478 (N_3478,N_1031,N_1865);
xnor U3479 (N_3479,N_2111,N_1954);
and U3480 (N_3480,N_1810,N_861);
and U3481 (N_3481,N_813,N_1017);
nor U3482 (N_3482,N_911,N_2183);
or U3483 (N_3483,N_2298,N_1757);
xor U3484 (N_3484,N_2370,N_391);
or U3485 (N_3485,N_1001,N_1869);
or U3486 (N_3486,N_2246,N_755);
and U3487 (N_3487,N_2361,N_530);
and U3488 (N_3488,N_430,N_1062);
or U3489 (N_3489,N_2343,N_500);
or U3490 (N_3490,N_701,N_2307);
or U3491 (N_3491,N_1476,N_2373);
xor U3492 (N_3492,N_2485,N_1060);
xnor U3493 (N_3493,N_624,N_2244);
xnor U3494 (N_3494,N_741,N_130);
nor U3495 (N_3495,N_2388,N_540);
and U3496 (N_3496,N_579,N_2259);
nand U3497 (N_3497,N_2038,N_1454);
nand U3498 (N_3498,N_275,N_1580);
or U3499 (N_3499,N_2444,N_383);
xor U3500 (N_3500,N_1036,N_1973);
and U3501 (N_3501,N_260,N_2149);
xnor U3502 (N_3502,N_1437,N_1245);
or U3503 (N_3503,N_513,N_1807);
xnor U3504 (N_3504,N_2076,N_895);
nand U3505 (N_3505,N_2400,N_1145);
xnor U3506 (N_3506,N_1980,N_1506);
or U3507 (N_3507,N_977,N_265);
nor U3508 (N_3508,N_421,N_1836);
nor U3509 (N_3509,N_2490,N_1998);
or U3510 (N_3510,N_1191,N_1257);
and U3511 (N_3511,N_1441,N_2387);
and U3512 (N_3512,N_21,N_1589);
xnor U3513 (N_3513,N_2166,N_240);
nor U3514 (N_3514,N_1737,N_1526);
and U3515 (N_3515,N_1811,N_298);
nand U3516 (N_3516,N_1139,N_1387);
xor U3517 (N_3517,N_2037,N_1178);
or U3518 (N_3518,N_230,N_1933);
and U3519 (N_3519,N_414,N_1212);
or U3520 (N_3520,N_1705,N_592);
nand U3521 (N_3521,N_1453,N_719);
nor U3522 (N_3522,N_1707,N_663);
and U3523 (N_3523,N_856,N_68);
xnor U3524 (N_3524,N_1854,N_2300);
nand U3525 (N_3525,N_1442,N_1288);
nand U3526 (N_3526,N_1851,N_1900);
or U3527 (N_3527,N_2265,N_352);
nor U3528 (N_3528,N_402,N_945);
and U3529 (N_3529,N_1379,N_667);
xor U3530 (N_3530,N_725,N_1244);
or U3531 (N_3531,N_2251,N_946);
nand U3532 (N_3532,N_2302,N_941);
xnor U3533 (N_3533,N_557,N_53);
nand U3534 (N_3534,N_2209,N_1643);
or U3535 (N_3535,N_1625,N_1213);
nand U3536 (N_3536,N_1254,N_1136);
and U3537 (N_3537,N_1395,N_2326);
nand U3538 (N_3538,N_2413,N_478);
nor U3539 (N_3539,N_921,N_190);
and U3540 (N_3540,N_927,N_1015);
xnor U3541 (N_3541,N_2202,N_41);
nor U3542 (N_3542,N_822,N_1202);
nor U3543 (N_3543,N_955,N_1657);
xnor U3544 (N_3544,N_796,N_1238);
nor U3545 (N_3545,N_681,N_1545);
or U3546 (N_3546,N_1987,N_621);
xor U3547 (N_3547,N_381,N_604);
xor U3548 (N_3548,N_1518,N_194);
or U3549 (N_3549,N_2016,N_1405);
nand U3550 (N_3550,N_2347,N_1326);
xor U3551 (N_3551,N_1660,N_1833);
or U3552 (N_3552,N_1887,N_2024);
and U3553 (N_3553,N_2101,N_1229);
nor U3554 (N_3554,N_1717,N_1818);
xnor U3555 (N_3555,N_1907,N_1104);
nand U3556 (N_3556,N_806,N_541);
or U3557 (N_3557,N_171,N_2488);
nand U3558 (N_3558,N_290,N_446);
nor U3559 (N_3559,N_413,N_1374);
xor U3560 (N_3560,N_1771,N_1513);
xor U3561 (N_3561,N_2052,N_497);
or U3562 (N_3562,N_688,N_1137);
nor U3563 (N_3563,N_832,N_919);
nand U3564 (N_3564,N_1521,N_723);
or U3565 (N_3565,N_1839,N_544);
nand U3566 (N_3566,N_731,N_2131);
and U3567 (N_3567,N_571,N_1081);
nand U3568 (N_3568,N_280,N_672);
nand U3569 (N_3569,N_867,N_315);
or U3570 (N_3570,N_586,N_2386);
and U3571 (N_3571,N_196,N_205);
xnor U3572 (N_3572,N_2255,N_360);
xnor U3573 (N_3573,N_1189,N_965);
or U3574 (N_3574,N_1168,N_1187);
nand U3575 (N_3575,N_670,N_970);
nand U3576 (N_3576,N_1194,N_172);
xnor U3577 (N_3577,N_2218,N_1738);
and U3578 (N_3578,N_525,N_94);
and U3579 (N_3579,N_1339,N_1700);
or U3580 (N_3580,N_1758,N_2086);
or U3581 (N_3581,N_1169,N_566);
nand U3582 (N_3582,N_1879,N_455);
nor U3583 (N_3583,N_1039,N_1156);
xor U3584 (N_3584,N_2279,N_2143);
or U3585 (N_3585,N_1988,N_742);
nor U3586 (N_3586,N_1765,N_2226);
nand U3587 (N_3587,N_613,N_312);
nand U3588 (N_3588,N_1676,N_2208);
nor U3589 (N_3589,N_1370,N_2465);
and U3590 (N_3590,N_2113,N_2487);
and U3591 (N_3591,N_317,N_2457);
and U3592 (N_3592,N_549,N_125);
xnor U3593 (N_3593,N_737,N_1575);
nand U3594 (N_3594,N_282,N_1596);
xor U3595 (N_3595,N_1445,N_1592);
or U3596 (N_3596,N_558,N_337);
or U3597 (N_3597,N_1249,N_2102);
or U3598 (N_3598,N_1561,N_885);
or U3599 (N_3599,N_1579,N_1629);
nand U3600 (N_3600,N_2175,N_892);
nor U3601 (N_3601,N_1152,N_844);
xnor U3602 (N_3602,N_2436,N_1507);
and U3603 (N_3603,N_2415,N_1443);
and U3604 (N_3604,N_971,N_1147);
or U3605 (N_3605,N_1004,N_42);
nor U3606 (N_3606,N_1165,N_2336);
nand U3607 (N_3607,N_423,N_2382);
xor U3608 (N_3608,N_1926,N_936);
nand U3609 (N_3609,N_1302,N_713);
and U3610 (N_3610,N_1159,N_2084);
xnor U3611 (N_3611,N_2198,N_2327);
nand U3612 (N_3612,N_2238,N_1612);
or U3613 (N_3613,N_1263,N_739);
nor U3614 (N_3614,N_1849,N_922);
and U3615 (N_3615,N_150,N_2041);
nand U3616 (N_3616,N_456,N_745);
and U3617 (N_3617,N_1208,N_1780);
nor U3618 (N_3618,N_46,N_1006);
xor U3619 (N_3619,N_1726,N_398);
xor U3620 (N_3620,N_2272,N_1292);
or U3621 (N_3621,N_241,N_953);
nand U3622 (N_3622,N_2341,N_2356);
or U3623 (N_3623,N_1255,N_695);
or U3624 (N_3624,N_97,N_2303);
xor U3625 (N_3625,N_1824,N_1361);
xor U3626 (N_3626,N_2417,N_1544);
xor U3627 (N_3627,N_76,N_775);
and U3628 (N_3628,N_5,N_441);
nor U3629 (N_3629,N_2480,N_1574);
nor U3630 (N_3630,N_1433,N_2380);
and U3631 (N_3631,N_1512,N_1967);
and U3632 (N_3632,N_1343,N_1188);
nand U3633 (N_3633,N_1899,N_975);
nor U3634 (N_3634,N_1753,N_791);
nand U3635 (N_3635,N_710,N_1016);
nand U3636 (N_3636,N_677,N_1086);
and U3637 (N_3637,N_2034,N_1260);
nor U3638 (N_3638,N_2134,N_580);
and U3639 (N_3639,N_828,N_168);
xnor U3640 (N_3640,N_651,N_350);
nor U3641 (N_3641,N_2280,N_1344);
or U3642 (N_3642,N_2369,N_2222);
or U3643 (N_3643,N_2358,N_2042);
nor U3644 (N_3644,N_732,N_938);
or U3645 (N_3645,N_1649,N_1604);
and U3646 (N_3646,N_1922,N_1239);
nand U3647 (N_3647,N_734,N_1870);
or U3648 (N_3648,N_50,N_1863);
nor U3649 (N_3649,N_465,N_2169);
xor U3650 (N_3650,N_1508,N_2112);
nand U3651 (N_3651,N_0,N_524);
or U3652 (N_3652,N_1222,N_1928);
and U3653 (N_3653,N_1266,N_1348);
or U3654 (N_3654,N_570,N_1531);
nand U3655 (N_3655,N_1885,N_1670);
and U3656 (N_3656,N_1862,N_341);
nand U3657 (N_3657,N_819,N_593);
nand U3658 (N_3658,N_767,N_487);
xor U3659 (N_3659,N_2352,N_748);
nand U3660 (N_3660,N_1498,N_1715);
nor U3661 (N_3661,N_1059,N_749);
xnor U3662 (N_3662,N_2059,N_1640);
and U3663 (N_3663,N_451,N_237);
and U3664 (N_3664,N_401,N_2344);
or U3665 (N_3665,N_976,N_296);
xnor U3666 (N_3666,N_1847,N_1492);
or U3667 (N_3667,N_564,N_763);
or U3668 (N_3668,N_1420,N_1989);
nor U3669 (N_3669,N_182,N_2472);
and U3670 (N_3670,N_2484,N_683);
nor U3671 (N_3671,N_1794,N_903);
or U3672 (N_3672,N_1932,N_1785);
and U3673 (N_3673,N_1983,N_1972);
or U3674 (N_3674,N_411,N_1410);
xnor U3675 (N_3675,N_1747,N_389);
xnor U3676 (N_3676,N_81,N_2077);
nor U3677 (N_3677,N_2022,N_1931);
or U3678 (N_3678,N_1584,N_1413);
nand U3679 (N_3679,N_1161,N_2019);
xnor U3680 (N_3680,N_96,N_764);
nor U3681 (N_3681,N_1750,N_654);
nor U3682 (N_3682,N_1364,N_1895);
xnor U3683 (N_3683,N_370,N_1821);
xor U3684 (N_3684,N_2483,N_1259);
and U3685 (N_3685,N_1564,N_738);
and U3686 (N_3686,N_62,N_1216);
nor U3687 (N_3687,N_833,N_1277);
nor U3688 (N_3688,N_78,N_1486);
nor U3689 (N_3689,N_210,N_640);
nand U3690 (N_3690,N_1699,N_983);
or U3691 (N_3691,N_1656,N_536);
xnor U3692 (N_3692,N_1306,N_1848);
xnor U3693 (N_3693,N_853,N_1953);
xnor U3694 (N_3694,N_994,N_1651);
nand U3695 (N_3695,N_761,N_2469);
nor U3696 (N_3696,N_2130,N_83);
nand U3697 (N_3697,N_2151,N_872);
and U3698 (N_3698,N_379,N_1225);
nand U3699 (N_3699,N_1373,N_2282);
nor U3700 (N_3700,N_1842,N_17);
and U3701 (N_3701,N_2164,N_2063);
or U3702 (N_3702,N_1950,N_2171);
nor U3703 (N_3703,N_690,N_1882);
xnor U3704 (N_3704,N_1770,N_264);
xor U3705 (N_3705,N_969,N_675);
nand U3706 (N_3706,N_445,N_1867);
and U3707 (N_3707,N_528,N_2398);
or U3708 (N_3708,N_2010,N_77);
nor U3709 (N_3709,N_1541,N_2363);
or U3710 (N_3710,N_2196,N_108);
or U3711 (N_3711,N_1522,N_611);
nand U3712 (N_3712,N_318,N_1210);
and U3713 (N_3713,N_397,N_865);
xnor U3714 (N_3714,N_2311,N_1353);
or U3715 (N_3715,N_1253,N_1279);
or U3716 (N_3716,N_2366,N_1223);
and U3717 (N_3717,N_1126,N_924);
and U3718 (N_3718,N_1813,N_1274);
xor U3719 (N_3719,N_937,N_1809);
xnor U3720 (N_3720,N_727,N_1621);
xnor U3721 (N_3721,N_1504,N_137);
nand U3722 (N_3722,N_1130,N_1958);
nor U3723 (N_3723,N_560,N_2074);
and U3724 (N_3724,N_851,N_680);
nor U3725 (N_3725,N_174,N_262);
nand U3726 (N_3726,N_51,N_1377);
xor U3727 (N_3727,N_1829,N_2230);
and U3728 (N_3728,N_1014,N_606);
nand U3729 (N_3729,N_1430,N_1537);
and U3730 (N_3730,N_473,N_1573);
nand U3731 (N_3731,N_2493,N_605);
xnor U3732 (N_3732,N_1146,N_2377);
nand U3733 (N_3733,N_2385,N_2110);
nor U3734 (N_3734,N_2437,N_1909);
xor U3735 (N_3735,N_2167,N_2357);
xor U3736 (N_3736,N_458,N_427);
or U3737 (N_3737,N_1734,N_151);
nor U3738 (N_3738,N_2354,N_1181);
xor U3739 (N_3739,N_1195,N_1618);
and U3740 (N_3740,N_1759,N_347);
nor U3741 (N_3741,N_1752,N_1167);
nor U3742 (N_3742,N_213,N_93);
nor U3743 (N_3743,N_2470,N_647);
nor U3744 (N_3744,N_2201,N_1256);
xnor U3745 (N_3745,N_1176,N_691);
and U3746 (N_3746,N_1861,N_332);
and U3747 (N_3747,N_785,N_2408);
and U3748 (N_3748,N_1282,N_1630);
and U3749 (N_3749,N_2491,N_12);
nand U3750 (N_3750,N_331,N_2189);
nor U3751 (N_3751,N_884,N_899);
xor U3752 (N_3752,N_2032,N_520);
nand U3753 (N_3753,N_436,N_358);
and U3754 (N_3754,N_1319,N_2161);
or U3755 (N_3755,N_1513,N_618);
nor U3756 (N_3756,N_1489,N_1055);
or U3757 (N_3757,N_1339,N_1939);
and U3758 (N_3758,N_1028,N_1195);
or U3759 (N_3759,N_1379,N_904);
or U3760 (N_3760,N_1206,N_1312);
and U3761 (N_3761,N_1178,N_1144);
xnor U3762 (N_3762,N_832,N_2375);
or U3763 (N_3763,N_2000,N_2031);
nand U3764 (N_3764,N_1757,N_464);
xnor U3765 (N_3765,N_1370,N_1101);
xnor U3766 (N_3766,N_185,N_760);
or U3767 (N_3767,N_1373,N_1579);
nor U3768 (N_3768,N_368,N_727);
nand U3769 (N_3769,N_1261,N_925);
xnor U3770 (N_3770,N_2054,N_569);
or U3771 (N_3771,N_2471,N_362);
nor U3772 (N_3772,N_1323,N_226);
nor U3773 (N_3773,N_896,N_2322);
nor U3774 (N_3774,N_2043,N_1776);
and U3775 (N_3775,N_1289,N_2348);
nor U3776 (N_3776,N_1839,N_2434);
xnor U3777 (N_3777,N_1972,N_123);
xor U3778 (N_3778,N_2383,N_406);
and U3779 (N_3779,N_1816,N_1329);
or U3780 (N_3780,N_294,N_2098);
and U3781 (N_3781,N_2250,N_1499);
nand U3782 (N_3782,N_239,N_367);
and U3783 (N_3783,N_2211,N_79);
nand U3784 (N_3784,N_9,N_763);
and U3785 (N_3785,N_1136,N_422);
or U3786 (N_3786,N_944,N_350);
xor U3787 (N_3787,N_1038,N_1031);
and U3788 (N_3788,N_1343,N_1811);
and U3789 (N_3789,N_204,N_1698);
nor U3790 (N_3790,N_2038,N_1226);
nand U3791 (N_3791,N_434,N_620);
xor U3792 (N_3792,N_276,N_1052);
and U3793 (N_3793,N_1666,N_1585);
or U3794 (N_3794,N_339,N_1513);
nor U3795 (N_3795,N_1931,N_602);
nand U3796 (N_3796,N_2141,N_925);
nand U3797 (N_3797,N_116,N_2079);
and U3798 (N_3798,N_1427,N_2046);
xnor U3799 (N_3799,N_1265,N_151);
or U3800 (N_3800,N_2287,N_901);
nand U3801 (N_3801,N_2491,N_1951);
and U3802 (N_3802,N_1652,N_422);
xnor U3803 (N_3803,N_812,N_1227);
or U3804 (N_3804,N_735,N_1380);
and U3805 (N_3805,N_2428,N_2001);
or U3806 (N_3806,N_1762,N_1611);
nor U3807 (N_3807,N_2147,N_2426);
xnor U3808 (N_3808,N_664,N_1462);
and U3809 (N_3809,N_1559,N_987);
nand U3810 (N_3810,N_2170,N_1491);
xor U3811 (N_3811,N_2193,N_495);
or U3812 (N_3812,N_1171,N_811);
and U3813 (N_3813,N_847,N_994);
and U3814 (N_3814,N_432,N_653);
nor U3815 (N_3815,N_541,N_2213);
or U3816 (N_3816,N_542,N_815);
nor U3817 (N_3817,N_1714,N_2158);
or U3818 (N_3818,N_670,N_2427);
and U3819 (N_3819,N_1933,N_2465);
nor U3820 (N_3820,N_90,N_2291);
or U3821 (N_3821,N_909,N_1279);
nor U3822 (N_3822,N_1566,N_2237);
or U3823 (N_3823,N_1930,N_282);
xnor U3824 (N_3824,N_1948,N_1904);
or U3825 (N_3825,N_1787,N_608);
and U3826 (N_3826,N_1382,N_790);
xor U3827 (N_3827,N_1673,N_657);
nand U3828 (N_3828,N_1446,N_1927);
nor U3829 (N_3829,N_1096,N_1564);
xor U3830 (N_3830,N_2425,N_1505);
xnor U3831 (N_3831,N_1986,N_1205);
and U3832 (N_3832,N_1595,N_1073);
or U3833 (N_3833,N_1785,N_2265);
or U3834 (N_3834,N_1420,N_2276);
nand U3835 (N_3835,N_1865,N_2204);
nand U3836 (N_3836,N_764,N_1991);
or U3837 (N_3837,N_676,N_673);
nand U3838 (N_3838,N_1976,N_942);
nor U3839 (N_3839,N_896,N_2099);
xor U3840 (N_3840,N_1058,N_1345);
nor U3841 (N_3841,N_40,N_1667);
nor U3842 (N_3842,N_243,N_2278);
nand U3843 (N_3843,N_667,N_962);
nor U3844 (N_3844,N_2137,N_1305);
xnor U3845 (N_3845,N_121,N_1436);
nand U3846 (N_3846,N_2041,N_356);
nor U3847 (N_3847,N_1177,N_1178);
nor U3848 (N_3848,N_666,N_858);
xor U3849 (N_3849,N_2301,N_1804);
xor U3850 (N_3850,N_2089,N_1782);
nor U3851 (N_3851,N_1393,N_637);
or U3852 (N_3852,N_559,N_473);
nand U3853 (N_3853,N_2104,N_1364);
nor U3854 (N_3854,N_1266,N_1755);
and U3855 (N_3855,N_2195,N_2222);
or U3856 (N_3856,N_645,N_260);
or U3857 (N_3857,N_2177,N_1749);
nand U3858 (N_3858,N_561,N_2112);
and U3859 (N_3859,N_756,N_1645);
xnor U3860 (N_3860,N_1209,N_2074);
or U3861 (N_3861,N_2054,N_2042);
and U3862 (N_3862,N_954,N_1298);
and U3863 (N_3863,N_1561,N_915);
or U3864 (N_3864,N_119,N_77);
and U3865 (N_3865,N_323,N_1322);
and U3866 (N_3866,N_995,N_1990);
nor U3867 (N_3867,N_167,N_1072);
nor U3868 (N_3868,N_2356,N_1775);
nand U3869 (N_3869,N_1295,N_1002);
xnor U3870 (N_3870,N_1957,N_931);
or U3871 (N_3871,N_505,N_768);
or U3872 (N_3872,N_1272,N_2294);
nor U3873 (N_3873,N_1275,N_296);
and U3874 (N_3874,N_1015,N_1404);
nand U3875 (N_3875,N_1716,N_421);
and U3876 (N_3876,N_185,N_652);
or U3877 (N_3877,N_2161,N_1149);
nor U3878 (N_3878,N_166,N_1109);
or U3879 (N_3879,N_239,N_2359);
xor U3880 (N_3880,N_1216,N_1305);
and U3881 (N_3881,N_176,N_638);
nand U3882 (N_3882,N_487,N_818);
and U3883 (N_3883,N_1759,N_911);
nand U3884 (N_3884,N_1687,N_1183);
and U3885 (N_3885,N_77,N_2333);
nor U3886 (N_3886,N_2264,N_82);
xor U3887 (N_3887,N_1444,N_2194);
and U3888 (N_3888,N_607,N_837);
xor U3889 (N_3889,N_944,N_1278);
nor U3890 (N_3890,N_376,N_427);
and U3891 (N_3891,N_904,N_798);
or U3892 (N_3892,N_2067,N_450);
nor U3893 (N_3893,N_1918,N_1124);
and U3894 (N_3894,N_2139,N_73);
and U3895 (N_3895,N_1177,N_1238);
or U3896 (N_3896,N_1137,N_1944);
or U3897 (N_3897,N_1925,N_750);
nand U3898 (N_3898,N_1228,N_1200);
nand U3899 (N_3899,N_616,N_870);
nor U3900 (N_3900,N_2105,N_1993);
nand U3901 (N_3901,N_592,N_2105);
nor U3902 (N_3902,N_281,N_1457);
nor U3903 (N_3903,N_1670,N_2109);
nor U3904 (N_3904,N_593,N_250);
and U3905 (N_3905,N_2188,N_2430);
and U3906 (N_3906,N_2388,N_1431);
or U3907 (N_3907,N_740,N_2185);
nor U3908 (N_3908,N_1678,N_237);
nand U3909 (N_3909,N_2471,N_364);
and U3910 (N_3910,N_1668,N_1244);
and U3911 (N_3911,N_1105,N_72);
nor U3912 (N_3912,N_1595,N_393);
and U3913 (N_3913,N_1275,N_1348);
or U3914 (N_3914,N_353,N_2277);
nor U3915 (N_3915,N_1117,N_617);
and U3916 (N_3916,N_364,N_255);
nor U3917 (N_3917,N_1319,N_1535);
nand U3918 (N_3918,N_358,N_164);
nor U3919 (N_3919,N_1089,N_1524);
and U3920 (N_3920,N_435,N_1683);
and U3921 (N_3921,N_2324,N_468);
or U3922 (N_3922,N_1232,N_1761);
or U3923 (N_3923,N_1684,N_334);
nand U3924 (N_3924,N_827,N_2343);
xor U3925 (N_3925,N_641,N_1088);
nand U3926 (N_3926,N_2265,N_1249);
and U3927 (N_3927,N_1951,N_56);
nand U3928 (N_3928,N_2431,N_1264);
and U3929 (N_3929,N_966,N_2434);
or U3930 (N_3930,N_2254,N_1150);
xor U3931 (N_3931,N_474,N_2110);
and U3932 (N_3932,N_1844,N_1091);
xor U3933 (N_3933,N_2171,N_885);
nand U3934 (N_3934,N_2466,N_309);
and U3935 (N_3935,N_2295,N_197);
and U3936 (N_3936,N_1068,N_844);
and U3937 (N_3937,N_2236,N_1099);
xor U3938 (N_3938,N_1562,N_1348);
nand U3939 (N_3939,N_792,N_69);
and U3940 (N_3940,N_2006,N_893);
and U3941 (N_3941,N_2132,N_1968);
nor U3942 (N_3942,N_1815,N_1774);
or U3943 (N_3943,N_1278,N_776);
nor U3944 (N_3944,N_281,N_1405);
or U3945 (N_3945,N_411,N_317);
nor U3946 (N_3946,N_401,N_653);
nand U3947 (N_3947,N_16,N_436);
and U3948 (N_3948,N_2243,N_254);
or U3949 (N_3949,N_1388,N_196);
nor U3950 (N_3950,N_227,N_1540);
nor U3951 (N_3951,N_1548,N_537);
nor U3952 (N_3952,N_2100,N_920);
and U3953 (N_3953,N_1958,N_1522);
nor U3954 (N_3954,N_1597,N_2252);
and U3955 (N_3955,N_1112,N_1719);
nor U3956 (N_3956,N_2237,N_2082);
nand U3957 (N_3957,N_1675,N_627);
nand U3958 (N_3958,N_756,N_1243);
nand U3959 (N_3959,N_802,N_319);
nor U3960 (N_3960,N_2254,N_2188);
xor U3961 (N_3961,N_1041,N_2181);
nor U3962 (N_3962,N_770,N_876);
nor U3963 (N_3963,N_878,N_1031);
or U3964 (N_3964,N_835,N_1855);
nand U3965 (N_3965,N_2395,N_2248);
nor U3966 (N_3966,N_1037,N_1576);
xnor U3967 (N_3967,N_97,N_644);
nor U3968 (N_3968,N_2164,N_485);
and U3969 (N_3969,N_2093,N_1440);
nand U3970 (N_3970,N_74,N_2343);
or U3971 (N_3971,N_1112,N_2097);
nand U3972 (N_3972,N_667,N_1960);
and U3973 (N_3973,N_785,N_1378);
xnor U3974 (N_3974,N_247,N_1699);
xnor U3975 (N_3975,N_733,N_2333);
nand U3976 (N_3976,N_696,N_1724);
and U3977 (N_3977,N_1301,N_1036);
nor U3978 (N_3978,N_4,N_1152);
nor U3979 (N_3979,N_1447,N_1553);
or U3980 (N_3980,N_1888,N_2009);
xnor U3981 (N_3981,N_2122,N_1946);
nand U3982 (N_3982,N_325,N_1464);
or U3983 (N_3983,N_1088,N_1978);
xnor U3984 (N_3984,N_1003,N_396);
and U3985 (N_3985,N_45,N_403);
and U3986 (N_3986,N_2094,N_453);
and U3987 (N_3987,N_2345,N_1882);
nor U3988 (N_3988,N_1971,N_2396);
and U3989 (N_3989,N_323,N_956);
or U3990 (N_3990,N_706,N_1243);
and U3991 (N_3991,N_1073,N_809);
or U3992 (N_3992,N_626,N_2399);
or U3993 (N_3993,N_838,N_918);
nand U3994 (N_3994,N_993,N_726);
xor U3995 (N_3995,N_11,N_2361);
nand U3996 (N_3996,N_2136,N_241);
nor U3997 (N_3997,N_2012,N_1923);
and U3998 (N_3998,N_862,N_225);
nand U3999 (N_3999,N_1406,N_2132);
xor U4000 (N_4000,N_462,N_2184);
nor U4001 (N_4001,N_1388,N_1345);
nor U4002 (N_4002,N_1461,N_39);
nand U4003 (N_4003,N_330,N_2095);
nor U4004 (N_4004,N_2133,N_2254);
nor U4005 (N_4005,N_1101,N_1055);
nor U4006 (N_4006,N_646,N_321);
nand U4007 (N_4007,N_1015,N_1749);
nor U4008 (N_4008,N_1811,N_1705);
or U4009 (N_4009,N_873,N_255);
xor U4010 (N_4010,N_2060,N_1075);
or U4011 (N_4011,N_222,N_334);
xor U4012 (N_4012,N_1679,N_616);
or U4013 (N_4013,N_2077,N_945);
nand U4014 (N_4014,N_698,N_1289);
xor U4015 (N_4015,N_2399,N_594);
or U4016 (N_4016,N_1930,N_1582);
xnor U4017 (N_4017,N_1589,N_516);
or U4018 (N_4018,N_705,N_819);
and U4019 (N_4019,N_1795,N_1859);
nor U4020 (N_4020,N_906,N_1849);
xnor U4021 (N_4021,N_993,N_2037);
and U4022 (N_4022,N_45,N_360);
or U4023 (N_4023,N_1134,N_1182);
and U4024 (N_4024,N_806,N_1582);
and U4025 (N_4025,N_1593,N_797);
or U4026 (N_4026,N_780,N_672);
nor U4027 (N_4027,N_578,N_2273);
xor U4028 (N_4028,N_1387,N_1230);
xnor U4029 (N_4029,N_776,N_1274);
and U4030 (N_4030,N_2038,N_1014);
and U4031 (N_4031,N_1824,N_682);
xnor U4032 (N_4032,N_506,N_1589);
xnor U4033 (N_4033,N_886,N_305);
or U4034 (N_4034,N_693,N_2311);
xor U4035 (N_4035,N_801,N_148);
nor U4036 (N_4036,N_858,N_1998);
and U4037 (N_4037,N_1248,N_647);
nor U4038 (N_4038,N_2100,N_2392);
xor U4039 (N_4039,N_2321,N_1147);
or U4040 (N_4040,N_1839,N_1168);
or U4041 (N_4041,N_1309,N_1042);
nor U4042 (N_4042,N_350,N_1737);
nand U4043 (N_4043,N_2315,N_1935);
nand U4044 (N_4044,N_1414,N_2391);
and U4045 (N_4045,N_548,N_2068);
nor U4046 (N_4046,N_462,N_972);
xor U4047 (N_4047,N_2095,N_1033);
and U4048 (N_4048,N_534,N_1564);
nor U4049 (N_4049,N_1357,N_666);
xor U4050 (N_4050,N_88,N_1239);
nor U4051 (N_4051,N_1729,N_2043);
nor U4052 (N_4052,N_2345,N_380);
nand U4053 (N_4053,N_850,N_348);
and U4054 (N_4054,N_1067,N_229);
nand U4055 (N_4055,N_409,N_2048);
xor U4056 (N_4056,N_370,N_2234);
nor U4057 (N_4057,N_263,N_1728);
and U4058 (N_4058,N_1278,N_165);
xor U4059 (N_4059,N_1575,N_1170);
and U4060 (N_4060,N_1436,N_1470);
nor U4061 (N_4061,N_126,N_924);
and U4062 (N_4062,N_947,N_2071);
xnor U4063 (N_4063,N_131,N_352);
xor U4064 (N_4064,N_946,N_1989);
nand U4065 (N_4065,N_1434,N_2359);
and U4066 (N_4066,N_1493,N_560);
nor U4067 (N_4067,N_2010,N_1626);
or U4068 (N_4068,N_2159,N_2383);
nand U4069 (N_4069,N_769,N_1567);
and U4070 (N_4070,N_2475,N_967);
xor U4071 (N_4071,N_86,N_2131);
nand U4072 (N_4072,N_1034,N_891);
or U4073 (N_4073,N_702,N_2424);
or U4074 (N_4074,N_207,N_728);
nor U4075 (N_4075,N_1952,N_901);
and U4076 (N_4076,N_948,N_1474);
or U4077 (N_4077,N_840,N_607);
and U4078 (N_4078,N_1674,N_380);
and U4079 (N_4079,N_373,N_2468);
and U4080 (N_4080,N_1453,N_139);
nor U4081 (N_4081,N_1366,N_2169);
nand U4082 (N_4082,N_39,N_1469);
or U4083 (N_4083,N_459,N_387);
or U4084 (N_4084,N_502,N_1499);
nor U4085 (N_4085,N_2294,N_475);
nor U4086 (N_4086,N_2473,N_2182);
and U4087 (N_4087,N_26,N_1829);
nand U4088 (N_4088,N_121,N_2183);
nor U4089 (N_4089,N_232,N_558);
nand U4090 (N_4090,N_804,N_833);
or U4091 (N_4091,N_2062,N_2016);
nand U4092 (N_4092,N_2142,N_1229);
or U4093 (N_4093,N_538,N_173);
or U4094 (N_4094,N_1588,N_200);
nand U4095 (N_4095,N_1235,N_396);
and U4096 (N_4096,N_134,N_1637);
and U4097 (N_4097,N_721,N_1102);
and U4098 (N_4098,N_341,N_975);
xnor U4099 (N_4099,N_921,N_1710);
xnor U4100 (N_4100,N_745,N_1096);
and U4101 (N_4101,N_1973,N_810);
or U4102 (N_4102,N_1325,N_2332);
nand U4103 (N_4103,N_570,N_177);
or U4104 (N_4104,N_2266,N_632);
or U4105 (N_4105,N_2398,N_473);
xnor U4106 (N_4106,N_2101,N_1951);
or U4107 (N_4107,N_2270,N_1940);
or U4108 (N_4108,N_848,N_2232);
or U4109 (N_4109,N_2089,N_189);
and U4110 (N_4110,N_1887,N_276);
and U4111 (N_4111,N_1496,N_1894);
xnor U4112 (N_4112,N_2271,N_1897);
or U4113 (N_4113,N_246,N_236);
and U4114 (N_4114,N_933,N_896);
nand U4115 (N_4115,N_1502,N_1626);
nand U4116 (N_4116,N_179,N_585);
xnor U4117 (N_4117,N_1702,N_2198);
nand U4118 (N_4118,N_272,N_1681);
nand U4119 (N_4119,N_2085,N_2292);
xnor U4120 (N_4120,N_309,N_2018);
nor U4121 (N_4121,N_2025,N_527);
and U4122 (N_4122,N_2060,N_553);
or U4123 (N_4123,N_2151,N_1684);
or U4124 (N_4124,N_2032,N_88);
nand U4125 (N_4125,N_1158,N_1333);
nor U4126 (N_4126,N_1795,N_714);
or U4127 (N_4127,N_2193,N_1844);
and U4128 (N_4128,N_1432,N_115);
and U4129 (N_4129,N_1988,N_473);
and U4130 (N_4130,N_1811,N_708);
nand U4131 (N_4131,N_2205,N_635);
and U4132 (N_4132,N_376,N_1681);
xor U4133 (N_4133,N_1158,N_961);
xor U4134 (N_4134,N_1498,N_1153);
nand U4135 (N_4135,N_660,N_548);
xor U4136 (N_4136,N_1368,N_2161);
and U4137 (N_4137,N_1498,N_1666);
or U4138 (N_4138,N_2328,N_540);
or U4139 (N_4139,N_1979,N_2296);
and U4140 (N_4140,N_101,N_501);
nand U4141 (N_4141,N_1853,N_2356);
or U4142 (N_4142,N_551,N_2006);
nor U4143 (N_4143,N_783,N_319);
and U4144 (N_4144,N_83,N_1340);
and U4145 (N_4145,N_1785,N_1362);
or U4146 (N_4146,N_791,N_1200);
nand U4147 (N_4147,N_318,N_724);
or U4148 (N_4148,N_1858,N_2306);
nor U4149 (N_4149,N_2371,N_2276);
and U4150 (N_4150,N_1523,N_502);
nand U4151 (N_4151,N_1449,N_1565);
or U4152 (N_4152,N_395,N_522);
nor U4153 (N_4153,N_46,N_1138);
nand U4154 (N_4154,N_329,N_962);
or U4155 (N_4155,N_1047,N_233);
nand U4156 (N_4156,N_2011,N_695);
and U4157 (N_4157,N_1150,N_660);
xnor U4158 (N_4158,N_224,N_1252);
nand U4159 (N_4159,N_902,N_919);
xnor U4160 (N_4160,N_1723,N_2139);
nor U4161 (N_4161,N_1495,N_177);
and U4162 (N_4162,N_1006,N_2097);
nand U4163 (N_4163,N_1371,N_380);
and U4164 (N_4164,N_1351,N_317);
nor U4165 (N_4165,N_47,N_1757);
and U4166 (N_4166,N_900,N_1040);
or U4167 (N_4167,N_1938,N_1772);
xnor U4168 (N_4168,N_346,N_225);
nor U4169 (N_4169,N_826,N_767);
or U4170 (N_4170,N_599,N_2308);
nor U4171 (N_4171,N_914,N_1922);
or U4172 (N_4172,N_1587,N_779);
xor U4173 (N_4173,N_888,N_2080);
xor U4174 (N_4174,N_1788,N_599);
nor U4175 (N_4175,N_316,N_764);
or U4176 (N_4176,N_1270,N_1619);
nand U4177 (N_4177,N_1361,N_325);
nor U4178 (N_4178,N_2402,N_1054);
or U4179 (N_4179,N_338,N_927);
nand U4180 (N_4180,N_280,N_1344);
or U4181 (N_4181,N_747,N_2410);
nor U4182 (N_4182,N_2148,N_321);
xor U4183 (N_4183,N_1683,N_1852);
or U4184 (N_4184,N_1249,N_520);
or U4185 (N_4185,N_2220,N_1985);
and U4186 (N_4186,N_800,N_1062);
nor U4187 (N_4187,N_722,N_1377);
or U4188 (N_4188,N_820,N_2465);
or U4189 (N_4189,N_624,N_1191);
and U4190 (N_4190,N_1520,N_643);
nor U4191 (N_4191,N_28,N_274);
nor U4192 (N_4192,N_1211,N_1879);
and U4193 (N_4193,N_538,N_1851);
nor U4194 (N_4194,N_1803,N_430);
and U4195 (N_4195,N_2237,N_946);
or U4196 (N_4196,N_2443,N_1594);
nor U4197 (N_4197,N_1598,N_230);
and U4198 (N_4198,N_45,N_690);
xnor U4199 (N_4199,N_508,N_43);
or U4200 (N_4200,N_2019,N_683);
xor U4201 (N_4201,N_638,N_1212);
xor U4202 (N_4202,N_683,N_2298);
nor U4203 (N_4203,N_609,N_1516);
or U4204 (N_4204,N_1754,N_1271);
or U4205 (N_4205,N_1783,N_476);
nor U4206 (N_4206,N_2153,N_1400);
nand U4207 (N_4207,N_1890,N_188);
or U4208 (N_4208,N_1174,N_1729);
or U4209 (N_4209,N_69,N_851);
and U4210 (N_4210,N_1437,N_79);
nand U4211 (N_4211,N_1334,N_1016);
nand U4212 (N_4212,N_1479,N_643);
and U4213 (N_4213,N_100,N_2298);
and U4214 (N_4214,N_1473,N_1509);
and U4215 (N_4215,N_1406,N_2291);
nor U4216 (N_4216,N_2439,N_2433);
nand U4217 (N_4217,N_1091,N_238);
xnor U4218 (N_4218,N_733,N_75);
nand U4219 (N_4219,N_1395,N_1573);
nand U4220 (N_4220,N_2186,N_522);
nand U4221 (N_4221,N_531,N_83);
or U4222 (N_4222,N_1142,N_1247);
and U4223 (N_4223,N_42,N_558);
or U4224 (N_4224,N_1332,N_467);
nand U4225 (N_4225,N_1670,N_1759);
or U4226 (N_4226,N_1927,N_2173);
nor U4227 (N_4227,N_77,N_733);
nor U4228 (N_4228,N_1596,N_53);
and U4229 (N_4229,N_1426,N_1846);
nor U4230 (N_4230,N_456,N_782);
nand U4231 (N_4231,N_1111,N_668);
xnor U4232 (N_4232,N_878,N_812);
or U4233 (N_4233,N_180,N_978);
and U4234 (N_4234,N_595,N_660);
and U4235 (N_4235,N_477,N_1694);
nor U4236 (N_4236,N_153,N_599);
nand U4237 (N_4237,N_1730,N_2084);
nand U4238 (N_4238,N_510,N_619);
nor U4239 (N_4239,N_1922,N_691);
and U4240 (N_4240,N_1689,N_942);
or U4241 (N_4241,N_2275,N_2399);
or U4242 (N_4242,N_2432,N_1369);
or U4243 (N_4243,N_2436,N_1807);
xor U4244 (N_4244,N_1971,N_1771);
or U4245 (N_4245,N_458,N_2467);
and U4246 (N_4246,N_552,N_644);
and U4247 (N_4247,N_1142,N_695);
nor U4248 (N_4248,N_1038,N_792);
xnor U4249 (N_4249,N_382,N_990);
nand U4250 (N_4250,N_1034,N_675);
nor U4251 (N_4251,N_2479,N_245);
nand U4252 (N_4252,N_163,N_261);
and U4253 (N_4253,N_2196,N_1583);
nand U4254 (N_4254,N_2405,N_1819);
nand U4255 (N_4255,N_62,N_177);
xor U4256 (N_4256,N_1053,N_541);
or U4257 (N_4257,N_1432,N_1271);
xnor U4258 (N_4258,N_2155,N_1967);
or U4259 (N_4259,N_1292,N_2271);
xnor U4260 (N_4260,N_93,N_1667);
nor U4261 (N_4261,N_1883,N_2133);
nand U4262 (N_4262,N_214,N_221);
nor U4263 (N_4263,N_876,N_1681);
and U4264 (N_4264,N_39,N_1751);
and U4265 (N_4265,N_2137,N_472);
and U4266 (N_4266,N_437,N_61);
or U4267 (N_4267,N_819,N_512);
nor U4268 (N_4268,N_2181,N_596);
nor U4269 (N_4269,N_2187,N_1288);
and U4270 (N_4270,N_1074,N_49);
nand U4271 (N_4271,N_240,N_1614);
nand U4272 (N_4272,N_1528,N_2415);
nand U4273 (N_4273,N_1748,N_243);
or U4274 (N_4274,N_1454,N_194);
and U4275 (N_4275,N_1086,N_600);
or U4276 (N_4276,N_651,N_1758);
and U4277 (N_4277,N_1338,N_296);
or U4278 (N_4278,N_2012,N_549);
or U4279 (N_4279,N_538,N_2160);
and U4280 (N_4280,N_493,N_1929);
nand U4281 (N_4281,N_487,N_1756);
nor U4282 (N_4282,N_1434,N_80);
nor U4283 (N_4283,N_1817,N_732);
nor U4284 (N_4284,N_424,N_311);
or U4285 (N_4285,N_1427,N_205);
nor U4286 (N_4286,N_1359,N_1858);
and U4287 (N_4287,N_1109,N_1212);
xnor U4288 (N_4288,N_2479,N_1074);
nand U4289 (N_4289,N_2025,N_1529);
xor U4290 (N_4290,N_1957,N_912);
and U4291 (N_4291,N_2391,N_61);
or U4292 (N_4292,N_803,N_2098);
nand U4293 (N_4293,N_824,N_2463);
and U4294 (N_4294,N_1667,N_1741);
or U4295 (N_4295,N_2484,N_1055);
nor U4296 (N_4296,N_1155,N_737);
and U4297 (N_4297,N_1252,N_1173);
and U4298 (N_4298,N_1289,N_479);
or U4299 (N_4299,N_312,N_585);
nand U4300 (N_4300,N_1192,N_543);
or U4301 (N_4301,N_1913,N_1694);
and U4302 (N_4302,N_536,N_1221);
xor U4303 (N_4303,N_2445,N_896);
nor U4304 (N_4304,N_2427,N_1858);
nor U4305 (N_4305,N_283,N_2391);
nor U4306 (N_4306,N_2210,N_706);
nand U4307 (N_4307,N_57,N_519);
nor U4308 (N_4308,N_1367,N_2358);
or U4309 (N_4309,N_1350,N_2021);
nand U4310 (N_4310,N_1744,N_2255);
nand U4311 (N_4311,N_378,N_1634);
xnor U4312 (N_4312,N_1749,N_834);
or U4313 (N_4313,N_174,N_2101);
xor U4314 (N_4314,N_2428,N_1392);
nor U4315 (N_4315,N_2385,N_198);
and U4316 (N_4316,N_1999,N_450);
nor U4317 (N_4317,N_1,N_406);
xor U4318 (N_4318,N_597,N_2354);
or U4319 (N_4319,N_2071,N_168);
nand U4320 (N_4320,N_377,N_19);
nor U4321 (N_4321,N_448,N_466);
xnor U4322 (N_4322,N_2387,N_1652);
and U4323 (N_4323,N_1525,N_1331);
xnor U4324 (N_4324,N_712,N_381);
and U4325 (N_4325,N_971,N_1710);
nor U4326 (N_4326,N_1571,N_385);
nor U4327 (N_4327,N_1823,N_243);
or U4328 (N_4328,N_1365,N_2355);
xnor U4329 (N_4329,N_1038,N_1351);
or U4330 (N_4330,N_132,N_860);
nand U4331 (N_4331,N_855,N_565);
or U4332 (N_4332,N_228,N_733);
xor U4333 (N_4333,N_1054,N_1482);
or U4334 (N_4334,N_765,N_78);
nor U4335 (N_4335,N_188,N_997);
nand U4336 (N_4336,N_2006,N_413);
nor U4337 (N_4337,N_2125,N_50);
or U4338 (N_4338,N_2179,N_2177);
or U4339 (N_4339,N_48,N_74);
or U4340 (N_4340,N_4,N_2016);
nor U4341 (N_4341,N_1626,N_404);
and U4342 (N_4342,N_948,N_288);
nand U4343 (N_4343,N_1579,N_1545);
nand U4344 (N_4344,N_1907,N_1245);
or U4345 (N_4345,N_2269,N_412);
nor U4346 (N_4346,N_1572,N_239);
and U4347 (N_4347,N_639,N_287);
and U4348 (N_4348,N_2258,N_634);
or U4349 (N_4349,N_582,N_1625);
xnor U4350 (N_4350,N_984,N_210);
or U4351 (N_4351,N_242,N_37);
nand U4352 (N_4352,N_372,N_2153);
xor U4353 (N_4353,N_2033,N_1985);
nor U4354 (N_4354,N_54,N_1642);
or U4355 (N_4355,N_1791,N_1498);
and U4356 (N_4356,N_606,N_2052);
and U4357 (N_4357,N_435,N_1971);
nand U4358 (N_4358,N_1153,N_582);
nand U4359 (N_4359,N_2434,N_226);
or U4360 (N_4360,N_104,N_2408);
xor U4361 (N_4361,N_1365,N_400);
nor U4362 (N_4362,N_2488,N_1362);
nand U4363 (N_4363,N_1276,N_1318);
or U4364 (N_4364,N_90,N_2460);
nor U4365 (N_4365,N_2439,N_1291);
nand U4366 (N_4366,N_1169,N_1332);
or U4367 (N_4367,N_2472,N_264);
nand U4368 (N_4368,N_2218,N_718);
nor U4369 (N_4369,N_353,N_1487);
and U4370 (N_4370,N_1816,N_0);
nand U4371 (N_4371,N_93,N_1150);
nor U4372 (N_4372,N_1162,N_145);
nand U4373 (N_4373,N_984,N_1465);
nand U4374 (N_4374,N_1417,N_799);
xor U4375 (N_4375,N_629,N_1684);
xnor U4376 (N_4376,N_1510,N_422);
and U4377 (N_4377,N_2467,N_424);
xor U4378 (N_4378,N_1172,N_2094);
or U4379 (N_4379,N_1462,N_1997);
nand U4380 (N_4380,N_1355,N_726);
xor U4381 (N_4381,N_837,N_810);
and U4382 (N_4382,N_1853,N_132);
nand U4383 (N_4383,N_1470,N_2337);
nand U4384 (N_4384,N_303,N_62);
or U4385 (N_4385,N_234,N_1935);
and U4386 (N_4386,N_2119,N_2256);
nand U4387 (N_4387,N_1995,N_1389);
and U4388 (N_4388,N_540,N_454);
and U4389 (N_4389,N_495,N_2099);
and U4390 (N_4390,N_1714,N_2433);
or U4391 (N_4391,N_2089,N_2319);
and U4392 (N_4392,N_671,N_2249);
and U4393 (N_4393,N_577,N_407);
nor U4394 (N_4394,N_1097,N_1581);
nor U4395 (N_4395,N_1999,N_2230);
and U4396 (N_4396,N_2378,N_1289);
nand U4397 (N_4397,N_1558,N_1311);
nor U4398 (N_4398,N_545,N_338);
nand U4399 (N_4399,N_371,N_1063);
nor U4400 (N_4400,N_985,N_1795);
and U4401 (N_4401,N_1025,N_561);
and U4402 (N_4402,N_1379,N_1027);
and U4403 (N_4403,N_667,N_2017);
xor U4404 (N_4404,N_386,N_741);
or U4405 (N_4405,N_1615,N_2417);
nor U4406 (N_4406,N_2477,N_364);
xnor U4407 (N_4407,N_1992,N_753);
xnor U4408 (N_4408,N_1020,N_548);
nor U4409 (N_4409,N_1366,N_13);
or U4410 (N_4410,N_2475,N_1948);
and U4411 (N_4411,N_1436,N_2033);
or U4412 (N_4412,N_1502,N_308);
nor U4413 (N_4413,N_1960,N_29);
nor U4414 (N_4414,N_1510,N_1369);
nor U4415 (N_4415,N_664,N_343);
nor U4416 (N_4416,N_1392,N_2276);
or U4417 (N_4417,N_377,N_1008);
nor U4418 (N_4418,N_2373,N_1574);
nand U4419 (N_4419,N_292,N_1800);
and U4420 (N_4420,N_634,N_457);
xor U4421 (N_4421,N_1618,N_1639);
and U4422 (N_4422,N_1867,N_807);
xor U4423 (N_4423,N_28,N_698);
nor U4424 (N_4424,N_2473,N_1728);
xor U4425 (N_4425,N_1270,N_250);
nor U4426 (N_4426,N_950,N_2069);
nand U4427 (N_4427,N_942,N_1881);
or U4428 (N_4428,N_2000,N_2019);
nor U4429 (N_4429,N_1197,N_487);
xor U4430 (N_4430,N_695,N_665);
or U4431 (N_4431,N_1618,N_2493);
nor U4432 (N_4432,N_2227,N_1175);
xor U4433 (N_4433,N_1210,N_854);
nand U4434 (N_4434,N_2155,N_541);
and U4435 (N_4435,N_2182,N_2196);
xnor U4436 (N_4436,N_1159,N_1861);
nor U4437 (N_4437,N_1821,N_506);
and U4438 (N_4438,N_2364,N_1874);
or U4439 (N_4439,N_2037,N_697);
xnor U4440 (N_4440,N_1448,N_560);
or U4441 (N_4441,N_1233,N_1689);
nor U4442 (N_4442,N_896,N_2412);
nor U4443 (N_4443,N_1915,N_2492);
and U4444 (N_4444,N_793,N_1717);
nand U4445 (N_4445,N_491,N_35);
and U4446 (N_4446,N_546,N_1480);
nor U4447 (N_4447,N_609,N_1102);
xnor U4448 (N_4448,N_1983,N_294);
nor U4449 (N_4449,N_1850,N_368);
nand U4450 (N_4450,N_1796,N_790);
and U4451 (N_4451,N_1800,N_985);
xor U4452 (N_4452,N_744,N_2288);
nor U4453 (N_4453,N_2297,N_701);
nor U4454 (N_4454,N_1887,N_2394);
and U4455 (N_4455,N_772,N_1134);
or U4456 (N_4456,N_2299,N_1017);
and U4457 (N_4457,N_1570,N_111);
or U4458 (N_4458,N_2466,N_2076);
xnor U4459 (N_4459,N_752,N_2220);
nand U4460 (N_4460,N_656,N_1801);
or U4461 (N_4461,N_2288,N_1611);
and U4462 (N_4462,N_2492,N_1626);
nor U4463 (N_4463,N_1177,N_1940);
or U4464 (N_4464,N_1131,N_403);
nor U4465 (N_4465,N_2024,N_1080);
nor U4466 (N_4466,N_186,N_240);
and U4467 (N_4467,N_2058,N_240);
nor U4468 (N_4468,N_82,N_623);
and U4469 (N_4469,N_2053,N_1347);
nand U4470 (N_4470,N_2335,N_1566);
xnor U4471 (N_4471,N_836,N_2248);
nor U4472 (N_4472,N_793,N_1477);
or U4473 (N_4473,N_1692,N_1402);
nor U4474 (N_4474,N_953,N_756);
or U4475 (N_4475,N_1886,N_389);
xor U4476 (N_4476,N_166,N_1754);
xor U4477 (N_4477,N_738,N_1449);
and U4478 (N_4478,N_2305,N_2075);
and U4479 (N_4479,N_2427,N_2117);
and U4480 (N_4480,N_1520,N_2024);
or U4481 (N_4481,N_1489,N_1019);
xnor U4482 (N_4482,N_390,N_1019);
nor U4483 (N_4483,N_1610,N_740);
xnor U4484 (N_4484,N_1814,N_2339);
and U4485 (N_4485,N_2119,N_2030);
and U4486 (N_4486,N_995,N_2145);
nor U4487 (N_4487,N_24,N_81);
and U4488 (N_4488,N_255,N_2308);
nand U4489 (N_4489,N_1067,N_1887);
xor U4490 (N_4490,N_362,N_2459);
xor U4491 (N_4491,N_2144,N_1835);
nor U4492 (N_4492,N_2383,N_22);
nand U4493 (N_4493,N_964,N_1309);
and U4494 (N_4494,N_2373,N_286);
and U4495 (N_4495,N_1559,N_2355);
and U4496 (N_4496,N_215,N_2334);
nor U4497 (N_4497,N_285,N_1106);
nor U4498 (N_4498,N_643,N_1599);
or U4499 (N_4499,N_575,N_1794);
or U4500 (N_4500,N_2326,N_2336);
nand U4501 (N_4501,N_2428,N_2414);
nor U4502 (N_4502,N_1469,N_2303);
nor U4503 (N_4503,N_459,N_411);
or U4504 (N_4504,N_474,N_1607);
nand U4505 (N_4505,N_1486,N_722);
nand U4506 (N_4506,N_1596,N_962);
xor U4507 (N_4507,N_1746,N_1821);
nand U4508 (N_4508,N_2196,N_920);
nor U4509 (N_4509,N_2095,N_2482);
and U4510 (N_4510,N_536,N_1346);
nand U4511 (N_4511,N_1186,N_1804);
xor U4512 (N_4512,N_714,N_1881);
or U4513 (N_4513,N_1939,N_127);
and U4514 (N_4514,N_1368,N_115);
nor U4515 (N_4515,N_1023,N_1563);
nand U4516 (N_4516,N_1980,N_1153);
and U4517 (N_4517,N_579,N_587);
or U4518 (N_4518,N_95,N_1777);
xor U4519 (N_4519,N_831,N_1574);
or U4520 (N_4520,N_2271,N_650);
xnor U4521 (N_4521,N_1296,N_2021);
nor U4522 (N_4522,N_1721,N_1411);
xnor U4523 (N_4523,N_1724,N_1741);
or U4524 (N_4524,N_415,N_2372);
or U4525 (N_4525,N_1422,N_2111);
or U4526 (N_4526,N_273,N_605);
and U4527 (N_4527,N_2073,N_104);
nand U4528 (N_4528,N_2496,N_927);
xor U4529 (N_4529,N_2009,N_232);
nor U4530 (N_4530,N_278,N_269);
and U4531 (N_4531,N_345,N_95);
nand U4532 (N_4532,N_1808,N_2289);
or U4533 (N_4533,N_1370,N_1544);
and U4534 (N_4534,N_1681,N_97);
nor U4535 (N_4535,N_902,N_1675);
or U4536 (N_4536,N_1155,N_2260);
and U4537 (N_4537,N_1411,N_2485);
and U4538 (N_4538,N_943,N_2280);
nand U4539 (N_4539,N_818,N_598);
nand U4540 (N_4540,N_193,N_1206);
or U4541 (N_4541,N_1976,N_1323);
xnor U4542 (N_4542,N_2287,N_1186);
xnor U4543 (N_4543,N_1913,N_1749);
xnor U4544 (N_4544,N_1588,N_1475);
nand U4545 (N_4545,N_1235,N_1204);
and U4546 (N_4546,N_2481,N_2430);
xor U4547 (N_4547,N_449,N_1407);
or U4548 (N_4548,N_2264,N_2167);
nor U4549 (N_4549,N_2370,N_457);
and U4550 (N_4550,N_1795,N_1556);
nand U4551 (N_4551,N_858,N_935);
xor U4552 (N_4552,N_591,N_58);
nor U4553 (N_4553,N_1538,N_63);
or U4554 (N_4554,N_1620,N_1135);
nand U4555 (N_4555,N_1488,N_1020);
and U4556 (N_4556,N_609,N_242);
nand U4557 (N_4557,N_1956,N_1039);
nand U4558 (N_4558,N_339,N_2428);
and U4559 (N_4559,N_1309,N_1100);
or U4560 (N_4560,N_2057,N_334);
or U4561 (N_4561,N_1212,N_2324);
and U4562 (N_4562,N_1876,N_459);
nor U4563 (N_4563,N_2115,N_879);
nand U4564 (N_4564,N_1244,N_1188);
or U4565 (N_4565,N_1784,N_770);
and U4566 (N_4566,N_1335,N_1399);
or U4567 (N_4567,N_119,N_1939);
nor U4568 (N_4568,N_2478,N_2138);
xnor U4569 (N_4569,N_516,N_153);
or U4570 (N_4570,N_1251,N_2253);
or U4571 (N_4571,N_532,N_1517);
nand U4572 (N_4572,N_2319,N_1761);
nor U4573 (N_4573,N_218,N_22);
nand U4574 (N_4574,N_674,N_2338);
nand U4575 (N_4575,N_1057,N_2001);
or U4576 (N_4576,N_1089,N_926);
nand U4577 (N_4577,N_989,N_2471);
nand U4578 (N_4578,N_640,N_319);
or U4579 (N_4579,N_345,N_715);
and U4580 (N_4580,N_1038,N_740);
xor U4581 (N_4581,N_2225,N_2184);
nor U4582 (N_4582,N_1088,N_436);
and U4583 (N_4583,N_1074,N_2130);
xnor U4584 (N_4584,N_882,N_540);
nor U4585 (N_4585,N_2053,N_1706);
xor U4586 (N_4586,N_143,N_1429);
nand U4587 (N_4587,N_1424,N_1783);
nand U4588 (N_4588,N_756,N_870);
xor U4589 (N_4589,N_2342,N_1410);
nor U4590 (N_4590,N_1528,N_290);
nand U4591 (N_4591,N_2498,N_623);
and U4592 (N_4592,N_2087,N_58);
or U4593 (N_4593,N_2346,N_1226);
xnor U4594 (N_4594,N_1984,N_398);
nand U4595 (N_4595,N_638,N_1198);
nand U4596 (N_4596,N_412,N_819);
nand U4597 (N_4597,N_1824,N_1652);
nor U4598 (N_4598,N_1542,N_1232);
nor U4599 (N_4599,N_1413,N_1134);
or U4600 (N_4600,N_1994,N_2213);
nand U4601 (N_4601,N_2299,N_2239);
or U4602 (N_4602,N_1948,N_243);
or U4603 (N_4603,N_1629,N_822);
or U4604 (N_4604,N_54,N_1286);
and U4605 (N_4605,N_1833,N_1788);
and U4606 (N_4606,N_948,N_2348);
nor U4607 (N_4607,N_1832,N_748);
and U4608 (N_4608,N_1724,N_1352);
and U4609 (N_4609,N_520,N_1986);
or U4610 (N_4610,N_2214,N_263);
nand U4611 (N_4611,N_1307,N_1497);
xnor U4612 (N_4612,N_2110,N_649);
nor U4613 (N_4613,N_2178,N_416);
nor U4614 (N_4614,N_852,N_1879);
xnor U4615 (N_4615,N_947,N_2050);
or U4616 (N_4616,N_2402,N_42);
nor U4617 (N_4617,N_1800,N_142);
xnor U4618 (N_4618,N_1246,N_745);
nand U4619 (N_4619,N_1020,N_570);
and U4620 (N_4620,N_2373,N_1662);
xor U4621 (N_4621,N_1121,N_1598);
xnor U4622 (N_4622,N_771,N_1245);
nand U4623 (N_4623,N_806,N_1973);
and U4624 (N_4624,N_1340,N_2477);
nand U4625 (N_4625,N_1748,N_2065);
or U4626 (N_4626,N_347,N_2387);
or U4627 (N_4627,N_2020,N_36);
nand U4628 (N_4628,N_392,N_1642);
nor U4629 (N_4629,N_2343,N_2230);
nor U4630 (N_4630,N_366,N_65);
nand U4631 (N_4631,N_831,N_1779);
nor U4632 (N_4632,N_233,N_180);
and U4633 (N_4633,N_1673,N_2492);
nand U4634 (N_4634,N_511,N_747);
nor U4635 (N_4635,N_2172,N_663);
xor U4636 (N_4636,N_1302,N_2202);
and U4637 (N_4637,N_1564,N_899);
or U4638 (N_4638,N_1428,N_2018);
or U4639 (N_4639,N_1516,N_1422);
and U4640 (N_4640,N_1217,N_2226);
xnor U4641 (N_4641,N_942,N_1230);
nand U4642 (N_4642,N_1204,N_1296);
or U4643 (N_4643,N_281,N_927);
xnor U4644 (N_4644,N_2334,N_1584);
nor U4645 (N_4645,N_1071,N_1999);
nand U4646 (N_4646,N_449,N_2331);
and U4647 (N_4647,N_1870,N_1190);
nand U4648 (N_4648,N_1202,N_2191);
and U4649 (N_4649,N_698,N_1131);
xor U4650 (N_4650,N_4,N_168);
nand U4651 (N_4651,N_490,N_1574);
or U4652 (N_4652,N_1821,N_811);
xor U4653 (N_4653,N_1735,N_733);
xor U4654 (N_4654,N_1467,N_1800);
xnor U4655 (N_4655,N_1676,N_1952);
and U4656 (N_4656,N_576,N_473);
xor U4657 (N_4657,N_661,N_1767);
nor U4658 (N_4658,N_1421,N_176);
or U4659 (N_4659,N_1344,N_881);
or U4660 (N_4660,N_179,N_628);
nor U4661 (N_4661,N_1244,N_1640);
xor U4662 (N_4662,N_1879,N_1941);
or U4663 (N_4663,N_290,N_1845);
and U4664 (N_4664,N_1266,N_1251);
or U4665 (N_4665,N_31,N_2109);
and U4666 (N_4666,N_469,N_26);
and U4667 (N_4667,N_2401,N_1546);
nor U4668 (N_4668,N_1900,N_1559);
nand U4669 (N_4669,N_1693,N_1386);
and U4670 (N_4670,N_211,N_401);
nor U4671 (N_4671,N_469,N_1123);
and U4672 (N_4672,N_2430,N_432);
xor U4673 (N_4673,N_1619,N_1411);
or U4674 (N_4674,N_1167,N_2277);
and U4675 (N_4675,N_337,N_2253);
xnor U4676 (N_4676,N_1874,N_2439);
and U4677 (N_4677,N_1518,N_1852);
xnor U4678 (N_4678,N_2334,N_581);
nand U4679 (N_4679,N_1113,N_1583);
or U4680 (N_4680,N_1112,N_376);
xnor U4681 (N_4681,N_273,N_1002);
and U4682 (N_4682,N_1115,N_744);
xor U4683 (N_4683,N_1116,N_1882);
nand U4684 (N_4684,N_1458,N_341);
nand U4685 (N_4685,N_1317,N_2448);
and U4686 (N_4686,N_2038,N_1294);
or U4687 (N_4687,N_133,N_572);
nor U4688 (N_4688,N_334,N_560);
nor U4689 (N_4689,N_2247,N_1906);
nand U4690 (N_4690,N_1241,N_1273);
nand U4691 (N_4691,N_955,N_123);
nand U4692 (N_4692,N_1407,N_2401);
and U4693 (N_4693,N_393,N_1379);
xnor U4694 (N_4694,N_357,N_649);
and U4695 (N_4695,N_913,N_1576);
and U4696 (N_4696,N_376,N_934);
nand U4697 (N_4697,N_729,N_1379);
nand U4698 (N_4698,N_1581,N_1336);
xor U4699 (N_4699,N_1198,N_1432);
and U4700 (N_4700,N_2247,N_1277);
nor U4701 (N_4701,N_610,N_1544);
nand U4702 (N_4702,N_2094,N_1325);
nor U4703 (N_4703,N_992,N_2088);
nand U4704 (N_4704,N_103,N_1569);
and U4705 (N_4705,N_1963,N_1563);
or U4706 (N_4706,N_1717,N_1143);
nand U4707 (N_4707,N_78,N_859);
nor U4708 (N_4708,N_1939,N_495);
or U4709 (N_4709,N_54,N_1224);
nand U4710 (N_4710,N_883,N_1429);
or U4711 (N_4711,N_1612,N_165);
nor U4712 (N_4712,N_878,N_961);
nor U4713 (N_4713,N_1286,N_2171);
and U4714 (N_4714,N_2268,N_258);
nand U4715 (N_4715,N_96,N_359);
xnor U4716 (N_4716,N_1635,N_1584);
nand U4717 (N_4717,N_464,N_511);
and U4718 (N_4718,N_1997,N_2249);
xnor U4719 (N_4719,N_1992,N_2271);
or U4720 (N_4720,N_2393,N_1967);
xor U4721 (N_4721,N_919,N_770);
or U4722 (N_4722,N_2033,N_353);
xor U4723 (N_4723,N_1412,N_769);
and U4724 (N_4724,N_1262,N_353);
xnor U4725 (N_4725,N_1680,N_1614);
nand U4726 (N_4726,N_2372,N_2479);
xnor U4727 (N_4727,N_413,N_1571);
or U4728 (N_4728,N_1920,N_1876);
and U4729 (N_4729,N_489,N_208);
and U4730 (N_4730,N_2366,N_1696);
xnor U4731 (N_4731,N_577,N_638);
nand U4732 (N_4732,N_2299,N_2089);
or U4733 (N_4733,N_1340,N_1448);
or U4734 (N_4734,N_1415,N_2476);
xor U4735 (N_4735,N_23,N_647);
xnor U4736 (N_4736,N_618,N_1947);
nand U4737 (N_4737,N_1895,N_298);
nor U4738 (N_4738,N_1471,N_1280);
or U4739 (N_4739,N_902,N_2385);
nor U4740 (N_4740,N_1442,N_1798);
xor U4741 (N_4741,N_1941,N_1972);
nor U4742 (N_4742,N_141,N_1942);
and U4743 (N_4743,N_1787,N_258);
and U4744 (N_4744,N_248,N_2211);
nand U4745 (N_4745,N_1530,N_1546);
xnor U4746 (N_4746,N_39,N_2121);
and U4747 (N_4747,N_980,N_278);
nand U4748 (N_4748,N_144,N_535);
xor U4749 (N_4749,N_2001,N_1206);
nand U4750 (N_4750,N_1316,N_1409);
and U4751 (N_4751,N_2306,N_1907);
nor U4752 (N_4752,N_169,N_1601);
xnor U4753 (N_4753,N_1567,N_1765);
xnor U4754 (N_4754,N_338,N_2293);
nor U4755 (N_4755,N_2376,N_1480);
and U4756 (N_4756,N_2351,N_1708);
or U4757 (N_4757,N_556,N_2190);
or U4758 (N_4758,N_1387,N_72);
nor U4759 (N_4759,N_76,N_933);
or U4760 (N_4760,N_352,N_1695);
nand U4761 (N_4761,N_1732,N_2339);
or U4762 (N_4762,N_1123,N_2038);
and U4763 (N_4763,N_1193,N_2022);
or U4764 (N_4764,N_2387,N_885);
and U4765 (N_4765,N_4,N_145);
and U4766 (N_4766,N_1689,N_64);
or U4767 (N_4767,N_2352,N_1507);
nor U4768 (N_4768,N_1302,N_1670);
and U4769 (N_4769,N_952,N_2234);
xor U4770 (N_4770,N_658,N_1138);
or U4771 (N_4771,N_120,N_1832);
nor U4772 (N_4772,N_1005,N_160);
nor U4773 (N_4773,N_642,N_92);
xnor U4774 (N_4774,N_2175,N_331);
or U4775 (N_4775,N_928,N_1068);
and U4776 (N_4776,N_1036,N_1513);
xor U4777 (N_4777,N_2003,N_1488);
and U4778 (N_4778,N_1214,N_1121);
nor U4779 (N_4779,N_2214,N_486);
xnor U4780 (N_4780,N_252,N_1947);
nand U4781 (N_4781,N_1477,N_1579);
or U4782 (N_4782,N_620,N_1399);
or U4783 (N_4783,N_1971,N_367);
nor U4784 (N_4784,N_399,N_1718);
or U4785 (N_4785,N_1567,N_445);
nor U4786 (N_4786,N_939,N_2240);
and U4787 (N_4787,N_954,N_943);
and U4788 (N_4788,N_1962,N_442);
xnor U4789 (N_4789,N_136,N_2229);
nor U4790 (N_4790,N_1936,N_1561);
nand U4791 (N_4791,N_1620,N_1535);
nor U4792 (N_4792,N_2448,N_2159);
and U4793 (N_4793,N_1814,N_117);
or U4794 (N_4794,N_2272,N_50);
nand U4795 (N_4795,N_743,N_224);
or U4796 (N_4796,N_2336,N_1169);
xor U4797 (N_4797,N_1700,N_736);
nand U4798 (N_4798,N_1028,N_1579);
and U4799 (N_4799,N_1522,N_928);
xor U4800 (N_4800,N_835,N_67);
nor U4801 (N_4801,N_1241,N_600);
xor U4802 (N_4802,N_32,N_1035);
or U4803 (N_4803,N_1938,N_138);
and U4804 (N_4804,N_206,N_2294);
or U4805 (N_4805,N_1360,N_1667);
nand U4806 (N_4806,N_2255,N_958);
and U4807 (N_4807,N_418,N_937);
nand U4808 (N_4808,N_1622,N_1893);
or U4809 (N_4809,N_1234,N_2144);
xor U4810 (N_4810,N_333,N_1793);
nand U4811 (N_4811,N_376,N_1564);
xnor U4812 (N_4812,N_1020,N_1537);
and U4813 (N_4813,N_1509,N_1556);
nand U4814 (N_4814,N_2088,N_1148);
or U4815 (N_4815,N_34,N_2172);
nand U4816 (N_4816,N_942,N_1981);
nand U4817 (N_4817,N_2159,N_1574);
and U4818 (N_4818,N_1474,N_1681);
xnor U4819 (N_4819,N_38,N_764);
nor U4820 (N_4820,N_758,N_1033);
xnor U4821 (N_4821,N_1928,N_219);
nand U4822 (N_4822,N_550,N_1473);
or U4823 (N_4823,N_545,N_326);
nand U4824 (N_4824,N_2490,N_1177);
nand U4825 (N_4825,N_2191,N_268);
xor U4826 (N_4826,N_1546,N_243);
nand U4827 (N_4827,N_638,N_673);
and U4828 (N_4828,N_429,N_2000);
nand U4829 (N_4829,N_1245,N_225);
nor U4830 (N_4830,N_528,N_826);
nand U4831 (N_4831,N_1306,N_1604);
and U4832 (N_4832,N_1284,N_2395);
and U4833 (N_4833,N_119,N_122);
xor U4834 (N_4834,N_324,N_1583);
or U4835 (N_4835,N_450,N_879);
xor U4836 (N_4836,N_2233,N_1300);
nor U4837 (N_4837,N_225,N_1022);
nor U4838 (N_4838,N_316,N_25);
xnor U4839 (N_4839,N_1056,N_2300);
nand U4840 (N_4840,N_446,N_24);
and U4841 (N_4841,N_1163,N_59);
nand U4842 (N_4842,N_851,N_2030);
nand U4843 (N_4843,N_628,N_1381);
nor U4844 (N_4844,N_874,N_1537);
nand U4845 (N_4845,N_941,N_1719);
nor U4846 (N_4846,N_2256,N_1400);
xnor U4847 (N_4847,N_355,N_2428);
xor U4848 (N_4848,N_935,N_674);
or U4849 (N_4849,N_29,N_597);
and U4850 (N_4850,N_2222,N_2240);
xor U4851 (N_4851,N_2188,N_2400);
xnor U4852 (N_4852,N_194,N_422);
nand U4853 (N_4853,N_11,N_1343);
and U4854 (N_4854,N_2296,N_2303);
xnor U4855 (N_4855,N_1641,N_1272);
xor U4856 (N_4856,N_503,N_589);
xnor U4857 (N_4857,N_2343,N_313);
nand U4858 (N_4858,N_1871,N_2309);
or U4859 (N_4859,N_437,N_2303);
nor U4860 (N_4860,N_629,N_236);
and U4861 (N_4861,N_1297,N_1075);
and U4862 (N_4862,N_2108,N_1035);
nor U4863 (N_4863,N_2051,N_1033);
nor U4864 (N_4864,N_765,N_229);
nand U4865 (N_4865,N_1706,N_1460);
and U4866 (N_4866,N_87,N_423);
xnor U4867 (N_4867,N_1189,N_704);
nand U4868 (N_4868,N_592,N_550);
xor U4869 (N_4869,N_60,N_1950);
nor U4870 (N_4870,N_1507,N_2338);
or U4871 (N_4871,N_83,N_1998);
or U4872 (N_4872,N_2378,N_1478);
xor U4873 (N_4873,N_1257,N_1846);
nor U4874 (N_4874,N_309,N_705);
xor U4875 (N_4875,N_1361,N_289);
and U4876 (N_4876,N_1024,N_1865);
or U4877 (N_4877,N_2045,N_2321);
nand U4878 (N_4878,N_647,N_1856);
or U4879 (N_4879,N_1435,N_56);
or U4880 (N_4880,N_455,N_2147);
nor U4881 (N_4881,N_1553,N_1292);
nor U4882 (N_4882,N_1211,N_2054);
nor U4883 (N_4883,N_151,N_2453);
and U4884 (N_4884,N_1007,N_1165);
nand U4885 (N_4885,N_332,N_1478);
or U4886 (N_4886,N_328,N_1988);
nor U4887 (N_4887,N_2153,N_1393);
and U4888 (N_4888,N_836,N_1914);
nor U4889 (N_4889,N_474,N_1084);
and U4890 (N_4890,N_1656,N_400);
nor U4891 (N_4891,N_1581,N_503);
nand U4892 (N_4892,N_1676,N_1452);
nand U4893 (N_4893,N_2357,N_1386);
nor U4894 (N_4894,N_409,N_590);
and U4895 (N_4895,N_1338,N_251);
nor U4896 (N_4896,N_2075,N_668);
and U4897 (N_4897,N_1041,N_2051);
nand U4898 (N_4898,N_1163,N_384);
nor U4899 (N_4899,N_2062,N_864);
or U4900 (N_4900,N_975,N_2125);
nand U4901 (N_4901,N_2134,N_1929);
and U4902 (N_4902,N_2190,N_798);
nand U4903 (N_4903,N_998,N_1463);
or U4904 (N_4904,N_324,N_673);
xor U4905 (N_4905,N_1678,N_2006);
nand U4906 (N_4906,N_924,N_52);
nor U4907 (N_4907,N_693,N_2273);
or U4908 (N_4908,N_572,N_1787);
and U4909 (N_4909,N_1461,N_2140);
nor U4910 (N_4910,N_298,N_2084);
xnor U4911 (N_4911,N_192,N_1707);
and U4912 (N_4912,N_1673,N_1900);
and U4913 (N_4913,N_1511,N_1791);
or U4914 (N_4914,N_1955,N_1674);
xnor U4915 (N_4915,N_797,N_2067);
nand U4916 (N_4916,N_1711,N_1171);
nor U4917 (N_4917,N_1998,N_1280);
or U4918 (N_4918,N_2486,N_407);
nor U4919 (N_4919,N_1934,N_1468);
or U4920 (N_4920,N_512,N_2408);
or U4921 (N_4921,N_391,N_126);
nor U4922 (N_4922,N_2472,N_1630);
xnor U4923 (N_4923,N_711,N_64);
nand U4924 (N_4924,N_1465,N_1864);
nand U4925 (N_4925,N_460,N_1251);
or U4926 (N_4926,N_522,N_13);
xor U4927 (N_4927,N_688,N_1069);
or U4928 (N_4928,N_1450,N_1813);
xor U4929 (N_4929,N_1197,N_2102);
nor U4930 (N_4930,N_1805,N_1655);
nor U4931 (N_4931,N_2169,N_458);
xnor U4932 (N_4932,N_1249,N_417);
nand U4933 (N_4933,N_2210,N_843);
or U4934 (N_4934,N_12,N_2071);
and U4935 (N_4935,N_1477,N_1862);
and U4936 (N_4936,N_1527,N_2388);
xnor U4937 (N_4937,N_1777,N_68);
nor U4938 (N_4938,N_1693,N_488);
and U4939 (N_4939,N_160,N_775);
xnor U4940 (N_4940,N_653,N_709);
or U4941 (N_4941,N_882,N_148);
nand U4942 (N_4942,N_955,N_1816);
xor U4943 (N_4943,N_461,N_1932);
or U4944 (N_4944,N_1208,N_2160);
and U4945 (N_4945,N_1323,N_744);
nand U4946 (N_4946,N_2290,N_268);
nor U4947 (N_4947,N_150,N_87);
nand U4948 (N_4948,N_2209,N_919);
or U4949 (N_4949,N_1905,N_425);
nand U4950 (N_4950,N_578,N_948);
nor U4951 (N_4951,N_2054,N_705);
or U4952 (N_4952,N_333,N_2250);
nor U4953 (N_4953,N_2137,N_1139);
xor U4954 (N_4954,N_1021,N_1466);
nand U4955 (N_4955,N_16,N_1430);
and U4956 (N_4956,N_576,N_2217);
and U4957 (N_4957,N_2177,N_2420);
and U4958 (N_4958,N_557,N_1502);
or U4959 (N_4959,N_995,N_2316);
xor U4960 (N_4960,N_2267,N_2402);
and U4961 (N_4961,N_905,N_1698);
xor U4962 (N_4962,N_1282,N_1281);
xnor U4963 (N_4963,N_2107,N_785);
or U4964 (N_4964,N_2148,N_445);
or U4965 (N_4965,N_102,N_2035);
xnor U4966 (N_4966,N_2348,N_1814);
nand U4967 (N_4967,N_1075,N_2378);
nor U4968 (N_4968,N_2152,N_630);
xor U4969 (N_4969,N_1102,N_538);
nor U4970 (N_4970,N_2178,N_2238);
nor U4971 (N_4971,N_1381,N_1043);
nor U4972 (N_4972,N_916,N_1928);
or U4973 (N_4973,N_1615,N_2353);
xor U4974 (N_4974,N_2306,N_2393);
nor U4975 (N_4975,N_1387,N_97);
nand U4976 (N_4976,N_23,N_32);
and U4977 (N_4977,N_234,N_1570);
or U4978 (N_4978,N_1706,N_1526);
and U4979 (N_4979,N_212,N_1834);
or U4980 (N_4980,N_545,N_527);
xnor U4981 (N_4981,N_1058,N_1489);
nand U4982 (N_4982,N_1291,N_798);
nand U4983 (N_4983,N_668,N_479);
xor U4984 (N_4984,N_987,N_593);
and U4985 (N_4985,N_483,N_287);
and U4986 (N_4986,N_1368,N_421);
and U4987 (N_4987,N_1783,N_1472);
nor U4988 (N_4988,N_1176,N_1165);
xor U4989 (N_4989,N_747,N_9);
and U4990 (N_4990,N_942,N_319);
nand U4991 (N_4991,N_1102,N_1988);
xnor U4992 (N_4992,N_700,N_1036);
nand U4993 (N_4993,N_1191,N_936);
and U4994 (N_4994,N_339,N_979);
and U4995 (N_4995,N_491,N_2480);
and U4996 (N_4996,N_1919,N_76);
xnor U4997 (N_4997,N_197,N_2447);
nor U4998 (N_4998,N_2371,N_1933);
xnor U4999 (N_4999,N_1138,N_1080);
xnor U5000 (N_5000,N_3027,N_4777);
and U5001 (N_5001,N_3811,N_2642);
or U5002 (N_5002,N_2934,N_3461);
nand U5003 (N_5003,N_3255,N_2897);
xnor U5004 (N_5004,N_3242,N_4206);
and U5005 (N_5005,N_2846,N_4231);
or U5006 (N_5006,N_3573,N_4120);
and U5007 (N_5007,N_3231,N_3591);
or U5008 (N_5008,N_4057,N_2673);
nor U5009 (N_5009,N_2838,N_3551);
xnor U5010 (N_5010,N_3252,N_4640);
xor U5011 (N_5011,N_4028,N_2827);
or U5012 (N_5012,N_3767,N_3297);
xnor U5013 (N_5013,N_3257,N_4821);
nand U5014 (N_5014,N_3971,N_2848);
nand U5015 (N_5015,N_4114,N_4862);
nand U5016 (N_5016,N_3195,N_4778);
and U5017 (N_5017,N_2582,N_4944);
or U5018 (N_5018,N_3812,N_3922);
xnor U5019 (N_5019,N_2512,N_3208);
and U5020 (N_5020,N_2812,N_4567);
nand U5021 (N_5021,N_4017,N_3694);
xnor U5022 (N_5022,N_2730,N_2938);
and U5023 (N_5023,N_4527,N_4771);
or U5024 (N_5024,N_4358,N_2698);
nand U5025 (N_5025,N_4662,N_3025);
and U5026 (N_5026,N_4015,N_2920);
nor U5027 (N_5027,N_4915,N_3783);
nor U5028 (N_5028,N_4882,N_3589);
or U5029 (N_5029,N_2940,N_4804);
nand U5030 (N_5030,N_3251,N_4994);
nor U5031 (N_5031,N_4996,N_3369);
or U5032 (N_5032,N_3705,N_4556);
nor U5033 (N_5033,N_4395,N_4728);
nand U5034 (N_5034,N_3840,N_4024);
nor U5035 (N_5035,N_3608,N_3264);
nand U5036 (N_5036,N_2667,N_3809);
xnor U5037 (N_5037,N_4968,N_4569);
xor U5038 (N_5038,N_4229,N_4455);
and U5039 (N_5039,N_4923,N_3951);
or U5040 (N_5040,N_4310,N_4265);
nor U5041 (N_5041,N_3194,N_4051);
xor U5042 (N_5042,N_2945,N_3082);
xor U5043 (N_5043,N_4195,N_4444);
nor U5044 (N_5044,N_3782,N_4703);
nor U5045 (N_5045,N_4440,N_3053);
and U5046 (N_5046,N_3584,N_4926);
and U5047 (N_5047,N_3201,N_4130);
nor U5048 (N_5048,N_3590,N_2779);
and U5049 (N_5049,N_3096,N_3943);
or U5050 (N_5050,N_4006,N_3068);
or U5051 (N_5051,N_4184,N_4725);
nand U5052 (N_5052,N_2861,N_3736);
xnor U5053 (N_5053,N_4502,N_4039);
nand U5054 (N_5054,N_3556,N_3755);
or U5055 (N_5055,N_3666,N_4881);
nand U5056 (N_5056,N_3581,N_2620);
and U5057 (N_5057,N_2629,N_3651);
or U5058 (N_5058,N_3126,N_3462);
nand U5059 (N_5059,N_2553,N_4718);
nor U5060 (N_5060,N_4489,N_3683);
nor U5061 (N_5061,N_3475,N_3883);
nand U5062 (N_5062,N_4408,N_3348);
and U5063 (N_5063,N_3919,N_3160);
or U5064 (N_5064,N_4940,N_3289);
or U5065 (N_5065,N_4371,N_3704);
and U5066 (N_5066,N_2649,N_4370);
and U5067 (N_5067,N_2648,N_4917);
nor U5068 (N_5068,N_3265,N_3328);
xnor U5069 (N_5069,N_3725,N_4207);
nand U5070 (N_5070,N_3769,N_2533);
xnor U5071 (N_5071,N_4244,N_4951);
xnor U5072 (N_5072,N_3456,N_3031);
or U5073 (N_5073,N_3978,N_4794);
xor U5074 (N_5074,N_3534,N_4507);
and U5075 (N_5075,N_2614,N_4360);
and U5076 (N_5076,N_3794,N_3948);
xor U5077 (N_5077,N_4529,N_4009);
and U5078 (N_5078,N_4619,N_2768);
or U5079 (N_5079,N_4390,N_4989);
nor U5080 (N_5080,N_3513,N_3610);
xor U5081 (N_5081,N_4941,N_4400);
nand U5082 (N_5082,N_3775,N_3323);
or U5083 (N_5083,N_4956,N_4344);
or U5084 (N_5084,N_3277,N_4425);
nand U5085 (N_5085,N_4406,N_3990);
nor U5086 (N_5086,N_4791,N_4337);
or U5087 (N_5087,N_3431,N_4072);
nand U5088 (N_5088,N_4572,N_3463);
xor U5089 (N_5089,N_4167,N_4945);
or U5090 (N_5090,N_4014,N_4822);
and U5091 (N_5091,N_3844,N_4590);
nand U5092 (N_5092,N_4318,N_3597);
xnor U5093 (N_5093,N_3485,N_3223);
nor U5094 (N_5094,N_4171,N_3715);
and U5095 (N_5095,N_2637,N_3123);
nand U5096 (N_5096,N_4029,N_4885);
or U5097 (N_5097,N_2993,N_4078);
or U5098 (N_5098,N_4317,N_3253);
nor U5099 (N_5099,N_4116,N_4185);
or U5100 (N_5100,N_3390,N_3508);
nor U5101 (N_5101,N_3383,N_3301);
and U5102 (N_5102,N_3890,N_3713);
and U5103 (N_5103,N_4332,N_3550);
nand U5104 (N_5104,N_4403,N_2966);
nand U5105 (N_5105,N_3532,N_2815);
nand U5106 (N_5106,N_4659,N_4924);
nand U5107 (N_5107,N_4525,N_3702);
or U5108 (N_5108,N_4046,N_4271);
nor U5109 (N_5109,N_4002,N_4495);
nand U5110 (N_5110,N_4255,N_3607);
and U5111 (N_5111,N_2894,N_2801);
xor U5112 (N_5112,N_2803,N_3181);
xnor U5113 (N_5113,N_2932,N_4049);
and U5114 (N_5114,N_4324,N_2933);
nand U5115 (N_5115,N_3384,N_4075);
or U5116 (N_5116,N_4824,N_4779);
or U5117 (N_5117,N_2685,N_3529);
and U5118 (N_5118,N_2645,N_3215);
nor U5119 (N_5119,N_4892,N_3227);
or U5120 (N_5120,N_4736,N_3452);
nand U5121 (N_5121,N_3499,N_3299);
nand U5122 (N_5122,N_3362,N_4521);
nand U5123 (N_5123,N_3980,N_3973);
xor U5124 (N_5124,N_4099,N_3744);
nand U5125 (N_5125,N_4478,N_3266);
nor U5126 (N_5126,N_3555,N_2747);
xor U5127 (N_5127,N_2719,N_4452);
nor U5128 (N_5128,N_3742,N_3337);
nand U5129 (N_5129,N_4712,N_4580);
or U5130 (N_5130,N_3386,N_3806);
and U5131 (N_5131,N_2592,N_3930);
xor U5132 (N_5132,N_4136,N_3032);
nand U5133 (N_5133,N_4341,N_3070);
and U5134 (N_5134,N_4362,N_2744);
nand U5135 (N_5135,N_3292,N_4987);
nor U5136 (N_5136,N_4998,N_2962);
and U5137 (N_5137,N_2657,N_4252);
nand U5138 (N_5138,N_4069,N_3909);
and U5139 (N_5139,N_2559,N_3984);
and U5140 (N_5140,N_4971,N_2893);
nor U5141 (N_5141,N_2856,N_3088);
nor U5142 (N_5142,N_2599,N_3043);
nor U5143 (N_5143,N_3199,N_2900);
nand U5144 (N_5144,N_3056,N_4316);
nor U5145 (N_5145,N_2769,N_4559);
or U5146 (N_5146,N_4418,N_2824);
and U5147 (N_5147,N_3979,N_4067);
or U5148 (N_5148,N_3611,N_3049);
or U5149 (N_5149,N_4638,N_3450);
nor U5150 (N_5150,N_2729,N_3949);
nor U5151 (N_5151,N_3011,N_4304);
and U5152 (N_5152,N_3953,N_2712);
nand U5153 (N_5153,N_3515,N_4102);
nor U5154 (N_5154,N_2888,N_2628);
xnor U5155 (N_5155,N_3445,N_3073);
nor U5156 (N_5156,N_2575,N_4745);
and U5157 (N_5157,N_2640,N_4157);
nand U5158 (N_5158,N_3213,N_3024);
nand U5159 (N_5159,N_4850,N_4367);
nand U5160 (N_5160,N_4274,N_4674);
and U5161 (N_5161,N_3633,N_4472);
nand U5162 (N_5162,N_2626,N_3838);
xnor U5163 (N_5163,N_3240,N_4172);
nor U5164 (N_5164,N_3531,N_4933);
nor U5165 (N_5165,N_4284,N_3727);
and U5166 (N_5166,N_2583,N_3685);
nor U5167 (N_5167,N_3481,N_4701);
xnor U5168 (N_5168,N_3756,N_3764);
and U5169 (N_5169,N_3745,N_3465);
or U5170 (N_5170,N_3247,N_3500);
nand U5171 (N_5171,N_2806,N_2631);
and U5172 (N_5172,N_4857,N_3678);
and U5173 (N_5173,N_4710,N_3587);
nor U5174 (N_5174,N_2758,N_4177);
nand U5175 (N_5175,N_4147,N_2728);
nand U5176 (N_5176,N_2802,N_3224);
and U5177 (N_5177,N_4330,N_3220);
nor U5178 (N_5178,N_3030,N_4286);
nor U5179 (N_5179,N_4744,N_2689);
and U5180 (N_5180,N_2664,N_4614);
and U5181 (N_5181,N_4315,N_3144);
xor U5182 (N_5182,N_3720,N_4869);
xor U5183 (N_5183,N_3051,N_3853);
nand U5184 (N_5184,N_4333,N_4162);
xor U5185 (N_5185,N_4826,N_2763);
nand U5186 (N_5186,N_2942,N_4957);
and U5187 (N_5187,N_4380,N_4625);
or U5188 (N_5188,N_4133,N_4805);
or U5189 (N_5189,N_4482,N_2505);
xor U5190 (N_5190,N_4348,N_3879);
nor U5191 (N_5191,N_4212,N_4415);
or U5192 (N_5192,N_2594,N_4123);
xnor U5193 (N_5193,N_4410,N_3969);
nor U5194 (N_5194,N_3205,N_4591);
nand U5195 (N_5195,N_3609,N_3161);
and U5196 (N_5196,N_4325,N_2694);
and U5197 (N_5197,N_4173,N_3966);
or U5198 (N_5198,N_4799,N_4488);
and U5199 (N_5199,N_3770,N_4769);
nand U5200 (N_5200,N_3864,N_3230);
and U5201 (N_5201,N_3855,N_2950);
or U5202 (N_5202,N_3668,N_4128);
or U5203 (N_5203,N_2767,N_4241);
or U5204 (N_5204,N_2836,N_3287);
nand U5205 (N_5205,N_3333,N_2672);
nand U5206 (N_5206,N_2654,N_2952);
or U5207 (N_5207,N_4907,N_2574);
and U5208 (N_5208,N_4776,N_4209);
or U5209 (N_5209,N_2743,N_3002);
nor U5210 (N_5210,N_3428,N_2896);
and U5211 (N_5211,N_3547,N_4909);
xor U5212 (N_5212,N_4563,N_2713);
xnor U5213 (N_5213,N_3340,N_4044);
or U5214 (N_5214,N_2562,N_3413);
nor U5215 (N_5215,N_2907,N_3276);
xnor U5216 (N_5216,N_4752,N_2556);
or U5217 (N_5217,N_3075,N_4010);
and U5218 (N_5218,N_3069,N_3376);
xor U5219 (N_5219,N_4842,N_4812);
or U5220 (N_5220,N_3779,N_3457);
and U5221 (N_5221,N_4503,N_4218);
nand U5222 (N_5222,N_3799,N_4442);
or U5223 (N_5223,N_4129,N_3006);
or U5224 (N_5224,N_4124,N_3878);
nor U5225 (N_5225,N_4511,N_3303);
and U5226 (N_5226,N_3378,N_3814);
or U5227 (N_5227,N_3646,N_4679);
or U5228 (N_5228,N_2825,N_3886);
xor U5229 (N_5229,N_3471,N_3837);
xor U5230 (N_5230,N_4815,N_4609);
nor U5231 (N_5231,N_4545,N_2847);
and U5232 (N_5232,N_4031,N_4743);
or U5233 (N_5233,N_4523,N_4880);
nand U5234 (N_5234,N_4107,N_4758);
nand U5235 (N_5235,N_3425,N_4890);
and U5236 (N_5236,N_4033,N_3202);
nor U5237 (N_5237,N_3158,N_3548);
nand U5238 (N_5238,N_3817,N_4616);
and U5239 (N_5239,N_2524,N_4677);
xor U5240 (N_5240,N_2568,N_3080);
and U5241 (N_5241,N_3526,N_2604);
and U5242 (N_5242,N_3959,N_4458);
or U5243 (N_5243,N_2760,N_3661);
nand U5244 (N_5244,N_4308,N_3647);
nor U5245 (N_5245,N_3674,N_2548);
xnor U5246 (N_5246,N_2884,N_3753);
nor U5247 (N_5247,N_3870,N_3539);
and U5248 (N_5248,N_2726,N_4093);
and U5249 (N_5249,N_2883,N_3955);
nand U5250 (N_5250,N_4810,N_4118);
xnor U5251 (N_5251,N_3179,N_3407);
and U5252 (N_5252,N_3822,N_2761);
xnor U5253 (N_5253,N_2697,N_3843);
or U5254 (N_5254,N_4746,N_4657);
nand U5255 (N_5255,N_3325,N_3660);
and U5256 (N_5256,N_4524,N_2809);
or U5257 (N_5257,N_4997,N_3697);
or U5258 (N_5258,N_4025,N_4424);
nor U5259 (N_5259,N_3188,N_3899);
nor U5260 (N_5260,N_4647,N_2578);
and U5261 (N_5261,N_4827,N_2717);
nor U5262 (N_5262,N_4401,N_4603);
nand U5263 (N_5263,N_4686,N_4240);
or U5264 (N_5264,N_3576,N_4861);
nor U5265 (N_5265,N_3695,N_2869);
and U5266 (N_5266,N_3352,N_2804);
nand U5267 (N_5267,N_4379,N_3574);
xnor U5268 (N_5268,N_2701,N_2970);
xnor U5269 (N_5269,N_3423,N_2532);
nand U5270 (N_5270,N_4141,N_2590);
nor U5271 (N_5271,N_4943,N_4179);
nand U5272 (N_5272,N_2676,N_3285);
xor U5273 (N_5273,N_3818,N_3165);
and U5274 (N_5274,N_2585,N_4327);
nand U5275 (N_5275,N_2774,N_3245);
or U5276 (N_5276,N_3987,N_4279);
and U5277 (N_5277,N_3374,N_3832);
and U5278 (N_5278,N_4194,N_2880);
xor U5279 (N_5279,N_3093,N_4874);
xnor U5280 (N_5280,N_4801,N_4236);
or U5281 (N_5281,N_3599,N_4076);
nor U5282 (N_5282,N_4699,N_3913);
xor U5283 (N_5283,N_3875,N_4516);
nand U5284 (N_5284,N_4397,N_3774);
nor U5285 (N_5285,N_3440,N_2875);
or U5286 (N_5286,N_2563,N_3732);
nor U5287 (N_5287,N_4034,N_2611);
nor U5288 (N_5288,N_4906,N_2500);
nor U5289 (N_5289,N_3766,N_3677);
xor U5290 (N_5290,N_4465,N_4307);
xor U5291 (N_5291,N_3901,N_3825);
nand U5292 (N_5292,N_4431,N_2659);
and U5293 (N_5293,N_3358,N_4192);
nand U5294 (N_5294,N_4306,N_4865);
xnor U5295 (N_5295,N_2683,N_3468);
nand U5296 (N_5296,N_3616,N_3841);
nand U5297 (N_5297,N_4052,N_2733);
nand U5298 (N_5298,N_4412,N_3330);
nor U5299 (N_5299,N_2855,N_3592);
nor U5300 (N_5300,N_3022,N_2877);
or U5301 (N_5301,N_4226,N_3829);
nand U5302 (N_5302,N_2851,N_3882);
nor U5303 (N_5303,N_2885,N_3327);
xor U5304 (N_5304,N_4878,N_3846);
and U5305 (N_5305,N_3918,N_3411);
nor U5306 (N_5306,N_2864,N_3669);
nor U5307 (N_5307,N_2765,N_4303);
nand U5308 (N_5308,N_2876,N_3561);
nor U5309 (N_5309,N_4018,N_2634);
nor U5310 (N_5310,N_2951,N_3896);
nor U5311 (N_5311,N_3293,N_3520);
xnor U5312 (N_5312,N_4095,N_4553);
xnor U5313 (N_5313,N_3460,N_3653);
or U5314 (N_5314,N_4479,N_3115);
and U5315 (N_5315,N_4407,N_4931);
or U5316 (N_5316,N_3162,N_4973);
nor U5317 (N_5317,N_2899,N_4237);
nand U5318 (N_5318,N_3149,N_4264);
and U5319 (N_5319,N_4338,N_3638);
or U5320 (N_5320,N_4643,N_4328);
xnor U5321 (N_5321,N_3035,N_3020);
nand U5322 (N_5322,N_3887,N_4087);
nand U5323 (N_5323,N_4276,N_4929);
and U5324 (N_5324,N_3459,N_3672);
xnor U5325 (N_5325,N_3209,N_3739);
nor U5326 (N_5326,N_4653,N_3780);
or U5327 (N_5327,N_3938,N_4427);
and U5328 (N_5328,N_3409,N_3418);
xnor U5329 (N_5329,N_2721,N_2636);
nand U5330 (N_5330,N_4221,N_3946);
or U5331 (N_5331,N_2598,N_4660);
xor U5332 (N_5332,N_3124,N_3700);
nand U5333 (N_5333,N_4731,N_4454);
and U5334 (N_5334,N_2707,N_2773);
nor U5335 (N_5335,N_4655,N_3795);
and U5336 (N_5336,N_3466,N_4707);
or U5337 (N_5337,N_4916,N_4835);
xnor U5338 (N_5338,N_3003,N_2929);
or U5339 (N_5339,N_2718,N_3153);
or U5340 (N_5340,N_3826,N_4708);
or U5341 (N_5341,N_4690,N_3007);
or U5342 (N_5342,N_2982,N_3860);
nor U5343 (N_5343,N_4834,N_2745);
nor U5344 (N_5344,N_2587,N_3687);
or U5345 (N_5345,N_4611,N_3273);
and U5346 (N_5346,N_3368,N_4356);
nand U5347 (N_5347,N_2845,N_4975);
nand U5348 (N_5348,N_3914,N_3436);
nor U5349 (N_5349,N_3952,N_3396);
nand U5350 (N_5350,N_3698,N_4174);
or U5351 (N_5351,N_3797,N_4352);
nand U5352 (N_5352,N_4430,N_4484);
xor U5353 (N_5353,N_2817,N_4579);
or U5354 (N_5354,N_4673,N_3842);
nand U5355 (N_5355,N_4974,N_4990);
nand U5356 (N_5356,N_3308,N_4692);
nand U5357 (N_5357,N_2786,N_4098);
nor U5358 (N_5358,N_3239,N_2946);
and U5359 (N_5359,N_3467,N_2757);
nor U5360 (N_5360,N_3570,N_3198);
xnor U5361 (N_5361,N_2749,N_3639);
nand U5362 (N_5362,N_2709,N_4938);
and U5363 (N_5363,N_4150,N_4620);
xnor U5364 (N_5364,N_3291,N_2573);
and U5365 (N_5365,N_3229,N_3477);
or U5366 (N_5366,N_4574,N_2520);
and U5367 (N_5367,N_3986,N_4186);
nor U5368 (N_5368,N_4460,N_4622);
nor U5369 (N_5369,N_3120,N_4627);
nor U5370 (N_5370,N_3988,N_4409);
xnor U5371 (N_5371,N_4387,N_2503);
nand U5372 (N_5372,N_3146,N_3868);
or U5373 (N_5373,N_4369,N_4080);
and U5374 (N_5374,N_3164,N_2787);
nor U5375 (N_5375,N_4381,N_4831);
nor U5376 (N_5376,N_2919,N_3370);
xor U5377 (N_5377,N_4152,N_2770);
nand U5378 (N_5378,N_3422,N_3975);
and U5379 (N_5379,N_3884,N_3816);
xnor U5380 (N_5380,N_2704,N_4282);
nor U5381 (N_5381,N_2660,N_2783);
and U5382 (N_5382,N_4663,N_4565);
nor U5383 (N_5383,N_4526,N_3081);
or U5384 (N_5384,N_4920,N_4334);
and U5385 (N_5385,N_4723,N_4512);
nand U5386 (N_5386,N_4054,N_4092);
or U5387 (N_5387,N_2669,N_3286);
xor U5388 (N_5388,N_4800,N_3320);
and U5389 (N_5389,N_3496,N_4966);
nor U5390 (N_5390,N_4349,N_3156);
nor U5391 (N_5391,N_3319,N_3933);
nand U5392 (N_5392,N_3912,N_2510);
or U5393 (N_5393,N_3079,N_4426);
or U5394 (N_5394,N_3334,N_4168);
nor U5395 (N_5395,N_3606,N_4654);
nand U5396 (N_5396,N_4669,N_4722);
nand U5397 (N_5397,N_3077,N_4323);
or U5398 (N_5398,N_4269,N_4499);
nor U5399 (N_5399,N_3446,N_2901);
and U5400 (N_5400,N_3708,N_4199);
nand U5401 (N_5401,N_2850,N_3116);
nand U5402 (N_5402,N_3925,N_4645);
nor U5403 (N_5403,N_3100,N_3222);
xor U5404 (N_5404,N_2677,N_3511);
nand U5405 (N_5405,N_4873,N_3349);
nand U5406 (N_5406,N_3628,N_2523);
xnor U5407 (N_5407,N_2853,N_3306);
or U5408 (N_5408,N_4615,N_4903);
nor U5409 (N_5409,N_3540,N_4963);
and U5410 (N_5410,N_2561,N_3784);
or U5411 (N_5411,N_2990,N_2678);
or U5412 (N_5412,N_3166,N_3614);
nand U5413 (N_5413,N_3112,N_3059);
or U5414 (N_5414,N_4038,N_4059);
nand U5415 (N_5415,N_3618,N_4202);
and U5416 (N_5416,N_3743,N_3619);
xor U5417 (N_5417,N_4058,N_3092);
nand U5418 (N_5418,N_4366,N_4583);
or U5419 (N_5419,N_2979,N_4661);
nand U5420 (N_5420,N_4983,N_4871);
or U5421 (N_5421,N_3354,N_4290);
or U5422 (N_5422,N_3524,N_3302);
nand U5423 (N_5423,N_4416,N_2814);
nor U5424 (N_5424,N_2684,N_3917);
and U5425 (N_5425,N_3125,N_4977);
xor U5426 (N_5426,N_4630,N_4927);
or U5427 (N_5427,N_2606,N_4012);
nor U5428 (N_5428,N_4109,N_3877);
nor U5429 (N_5429,N_3037,N_3852);
or U5430 (N_5430,N_4508,N_4176);
xor U5431 (N_5431,N_3437,N_2756);
nand U5432 (N_5432,N_4036,N_4721);
or U5433 (N_5433,N_4091,N_4446);
nor U5434 (N_5434,N_3226,N_4449);
xnor U5435 (N_5435,N_3356,N_3665);
nand U5436 (N_5436,N_2916,N_3000);
nor U5437 (N_5437,N_4952,N_3071);
or U5438 (N_5438,N_3109,N_4434);
and U5439 (N_5439,N_3193,N_3084);
xor U5440 (N_5440,N_2540,N_3398);
or U5441 (N_5441,N_4106,N_3183);
or U5442 (N_5442,N_2589,N_4585);
or U5443 (N_5443,N_2507,N_4339);
nor U5444 (N_5444,N_4519,N_2633);
xnor U5445 (N_5445,N_3342,N_3225);
or U5446 (N_5446,N_3136,N_4258);
xnor U5447 (N_5447,N_4773,N_4396);
xor U5448 (N_5448,N_4027,N_2764);
and U5449 (N_5449,N_2715,N_2601);
xnor U5450 (N_5450,N_4477,N_3013);
nor U5451 (N_5451,N_3424,N_2619);
nand U5452 (N_5452,N_3671,N_3267);
xor U5453 (N_5453,N_3985,N_4793);
and U5454 (N_5454,N_4414,N_4902);
and U5455 (N_5455,N_2531,N_2518);
xnor U5456 (N_5456,N_4262,N_4550);
xor U5457 (N_5457,N_4509,N_4011);
or U5458 (N_5458,N_3235,N_3902);
nand U5459 (N_5459,N_4101,N_3553);
nand U5460 (N_5460,N_3620,N_4249);
or U5461 (N_5461,N_4817,N_4535);
nand U5462 (N_5462,N_4113,N_4589);
or U5463 (N_5463,N_2777,N_4671);
xnor U5464 (N_5464,N_2904,N_2800);
nor U5465 (N_5465,N_3190,N_3042);
nor U5466 (N_5466,N_4605,N_3121);
xor U5467 (N_5467,N_4658,N_2610);
and U5468 (N_5468,N_3174,N_2666);
and U5469 (N_5469,N_4470,N_3344);
and U5470 (N_5470,N_4086,N_3528);
xnor U5471 (N_5471,N_2688,N_3406);
xnor U5472 (N_5472,N_4081,N_3249);
or U5473 (N_5473,N_3676,N_4300);
nor U5474 (N_5474,N_4964,N_4844);
xnor U5475 (N_5475,N_3693,N_4928);
xnor U5476 (N_5476,N_4079,N_3004);
nand U5477 (N_5477,N_2546,N_4775);
xnor U5478 (N_5478,N_4532,N_4937);
or U5479 (N_5479,N_4198,N_3216);
or U5480 (N_5480,N_4243,N_3430);
nor U5481 (N_5481,N_4908,N_4680);
nor U5482 (N_5482,N_3168,N_3941);
nor U5483 (N_5483,N_2504,N_2665);
and U5484 (N_5484,N_2964,N_2723);
and U5485 (N_5485,N_3012,N_4547);
nor U5486 (N_5486,N_4540,N_4646);
nor U5487 (N_5487,N_4498,N_3039);
or U5488 (N_5488,N_3892,N_3733);
and U5489 (N_5489,N_3150,N_3351);
or U5490 (N_5490,N_2731,N_4691);
and U5491 (N_5491,N_2608,N_2714);
nor U5492 (N_5492,N_3151,N_2949);
nand U5493 (N_5493,N_4139,N_4715);
and U5494 (N_5494,N_2644,N_3598);
nand U5495 (N_5495,N_4441,N_4108);
xor U5496 (N_5496,N_2506,N_4223);
nand U5497 (N_5497,N_3757,N_4515);
or U5498 (N_5498,N_3064,N_3028);
xor U5499 (N_5499,N_3572,N_2927);
and U5500 (N_5500,N_2748,N_4056);
nand U5501 (N_5501,N_2898,N_3976);
nor U5502 (N_5502,N_3097,N_3439);
xor U5503 (N_5503,N_3706,N_2558);
xnor U5504 (N_5504,N_4950,N_4760);
nand U5505 (N_5505,N_2857,N_2552);
nor U5506 (N_5506,N_3113,N_4687);
or U5507 (N_5507,N_3167,N_4122);
or U5508 (N_5508,N_2565,N_3617);
nor U5509 (N_5509,N_3800,N_3549);
nor U5510 (N_5510,N_4656,N_2740);
xor U5511 (N_5511,N_3861,N_3891);
nor U5512 (N_5512,N_2843,N_2530);
or U5513 (N_5513,N_4901,N_3670);
nand U5514 (N_5514,N_4879,N_3562);
and U5515 (N_5515,N_4321,N_4541);
xor U5516 (N_5516,N_4007,N_4000);
and U5517 (N_5517,N_3805,N_3426);
or U5518 (N_5518,N_4261,N_3648);
nor U5519 (N_5519,N_3382,N_4239);
and U5520 (N_5520,N_3833,N_4232);
nand U5521 (N_5521,N_2502,N_3545);
and U5522 (N_5522,N_4787,N_3737);
nand U5523 (N_5523,N_2973,N_3360);
nor U5524 (N_5524,N_2895,N_4864);
and U5525 (N_5525,N_3129,N_3900);
xor U5526 (N_5526,N_3629,N_4331);
xor U5527 (N_5527,N_3813,N_4642);
nor U5528 (N_5528,N_3719,N_2622);
xor U5529 (N_5529,N_3014,N_3041);
or U5530 (N_5530,N_3787,N_4716);
nor U5531 (N_5531,N_3140,N_2708);
nor U5532 (N_5532,N_3414,N_3128);
or U5533 (N_5533,N_3557,N_3350);
nand U5534 (N_5534,N_4277,N_3537);
and U5535 (N_5535,N_2528,N_4610);
nand U5536 (N_5536,N_3785,N_4738);
or U5537 (N_5537,N_3964,N_3936);
nand U5538 (N_5538,N_2621,N_2858);
nor U5539 (N_5539,N_3505,N_4437);
and U5540 (N_5540,N_4189,N_4637);
xor U5541 (N_5541,N_3400,N_3595);
xor U5542 (N_5542,N_4022,N_4768);
xor U5543 (N_5543,N_4984,N_4125);
and U5544 (N_5544,N_3105,N_3313);
nor U5545 (N_5545,N_2706,N_4705);
nor U5546 (N_5546,N_2988,N_3995);
nand U5547 (N_5547,N_4432,N_3881);
nor U5548 (N_5548,N_3801,N_3391);
and U5549 (N_5549,N_4420,N_3543);
or U5550 (N_5550,N_4551,N_2955);
nor U5551 (N_5551,N_2651,N_3517);
or U5552 (N_5552,N_2868,N_2742);
nor U5553 (N_5553,N_3565,N_3824);
or U5554 (N_5554,N_4624,N_2782);
and U5555 (N_5555,N_3569,N_4040);
xor U5556 (N_5556,N_3530,N_2600);
and U5557 (N_5557,N_3221,N_2944);
or U5558 (N_5558,N_4486,N_2519);
or U5559 (N_5559,N_4632,N_3679);
or U5560 (N_5560,N_4245,N_4008);
or U5561 (N_5561,N_3268,N_4720);
or U5562 (N_5562,N_3214,N_3403);
nand U5563 (N_5563,N_3680,N_4368);
nand U5564 (N_5564,N_3148,N_2960);
nor U5565 (N_5565,N_3626,N_4795);
or U5566 (N_5566,N_2947,N_3937);
nor U5567 (N_5567,N_3399,N_3586);
or U5568 (N_5568,N_4398,N_3604);
or U5569 (N_5569,N_3304,N_4248);
xor U5570 (N_5570,N_4825,N_4084);
nor U5571 (N_5571,N_4345,N_3170);
xnor U5572 (N_5572,N_2596,N_3178);
nor U5573 (N_5573,N_3790,N_2516);
and U5574 (N_5574,N_3566,N_4757);
or U5575 (N_5575,N_3060,N_4517);
xnor U5576 (N_5576,N_4786,N_3991);
nand U5577 (N_5577,N_3332,N_2795);
and U5578 (N_5578,N_2921,N_4298);
xnor U5579 (N_5579,N_4856,N_3746);
nor U5580 (N_5580,N_3331,N_3535);
xnor U5581 (N_5581,N_4257,N_2741);
and U5582 (N_5582,N_2863,N_2569);
and U5583 (N_5583,N_4492,N_3641);
or U5584 (N_5584,N_2612,N_4082);
or U5585 (N_5585,N_4702,N_4392);
nand U5586 (N_5586,N_3579,N_4510);
xnor U5587 (N_5587,N_2732,N_4062);
nand U5588 (N_5588,N_3491,N_3375);
or U5589 (N_5589,N_3114,N_3939);
nor U5590 (N_5590,N_3834,N_4263);
nor U5591 (N_5591,N_4225,N_3196);
or U5592 (N_5592,N_2823,N_4913);
nor U5593 (N_5593,N_3578,N_4291);
nor U5594 (N_5594,N_4270,N_4513);
xnor U5595 (N_5595,N_4383,N_4621);
or U5596 (N_5596,N_4595,N_2866);
nand U5597 (N_5597,N_3029,N_4772);
and U5598 (N_5598,N_4105,N_4413);
nor U5599 (N_5599,N_4675,N_2886);
xnor U5600 (N_5600,N_3904,N_3270);
xnor U5601 (N_5601,N_2974,N_2870);
xnor U5602 (N_5602,N_4796,N_2910);
xnor U5603 (N_5603,N_2859,N_3992);
or U5604 (N_5604,N_2892,N_3065);
and U5605 (N_5605,N_3663,N_3173);
and U5606 (N_5606,N_3147,N_3810);
and U5607 (N_5607,N_2794,N_4073);
or U5608 (N_5608,N_3504,N_3915);
nand U5609 (N_5609,N_4001,N_4782);
and U5610 (N_5610,N_4846,N_2906);
or U5611 (N_5611,N_3191,N_4190);
or U5612 (N_5612,N_2643,N_3091);
nor U5613 (N_5613,N_3684,N_2681);
nor U5614 (N_5614,N_2954,N_3486);
and U5615 (N_5615,N_2554,N_3217);
or U5616 (N_5616,N_4089,N_2820);
xor U5617 (N_5617,N_3280,N_3974);
nand U5618 (N_5618,N_3412,N_4774);
or U5619 (N_5619,N_3625,N_3982);
nand U5620 (N_5620,N_2724,N_2778);
xnor U5621 (N_5621,N_2792,N_4755);
and U5622 (N_5622,N_4137,N_4693);
xnor U5623 (N_5623,N_2605,N_3441);
or U5624 (N_5624,N_4026,N_4305);
nor U5625 (N_5625,N_3387,N_3759);
xor U5626 (N_5626,N_4247,N_2890);
xnor U5627 (N_5627,N_4314,N_4436);
or U5628 (N_5628,N_3152,N_4104);
nand U5629 (N_5629,N_2867,N_2881);
and U5630 (N_5630,N_4765,N_4053);
or U5631 (N_5631,N_2785,N_4897);
nor U5632 (N_5632,N_3726,N_4910);
xnor U5633 (N_5633,N_4238,N_3963);
xnor U5634 (N_5634,N_4342,N_2961);
nand U5635 (N_5635,N_4613,N_3052);
nand U5636 (N_5636,N_3204,N_4730);
nor U5637 (N_5637,N_2658,N_2579);
and U5638 (N_5638,N_4134,N_4048);
xnor U5639 (N_5639,N_3282,N_2525);
or U5640 (N_5640,N_3142,N_4188);
or U5641 (N_5641,N_4808,N_2544);
nor U5642 (N_5642,N_3389,N_4644);
nor U5643 (N_5643,N_4411,N_3636);
xnor U5644 (N_5644,N_4685,N_4494);
nor U5645 (N_5645,N_4160,N_3750);
or U5646 (N_5646,N_3256,N_3311);
or U5647 (N_5647,N_4530,N_3262);
nand U5648 (N_5648,N_4766,N_2511);
nand U5649 (N_5649,N_3583,N_3171);
or U5650 (N_5650,N_3339,N_4224);
nand U5651 (N_5651,N_3741,N_3005);
nor U5652 (N_5652,N_3640,N_3972);
nor U5653 (N_5653,N_3021,N_4993);
xnor U5654 (N_5654,N_3366,N_2996);
nor U5655 (N_5655,N_4178,N_3815);
xor U5656 (N_5656,N_2662,N_2545);
or U5657 (N_5657,N_4422,N_4756);
nand U5658 (N_5658,N_3099,N_2826);
xnor U5659 (N_5659,N_3315,N_4578);
or U5660 (N_5660,N_4568,N_4623);
nand U5661 (N_5661,N_2849,N_4148);
nor U5662 (N_5662,N_4891,N_3729);
or U5663 (N_5663,N_4855,N_3728);
xnor U5664 (N_5664,N_3206,N_3497);
nor U5665 (N_5665,N_3575,N_4083);
nor U5666 (N_5666,N_3310,N_3871);
nand U5667 (N_5667,N_2873,N_3897);
nor U5668 (N_5668,N_3823,N_2922);
and U5669 (N_5669,N_4807,N_3076);
nand U5670 (N_5670,N_3001,N_4949);
or U5671 (N_5671,N_3710,N_3089);
or U5672 (N_5672,N_3119,N_4970);
or U5673 (N_5673,N_3696,N_2959);
and U5674 (N_5674,N_4103,N_3098);
or U5675 (N_5675,N_3954,N_4814);
xor U5676 (N_5676,N_3664,N_4982);
nor U5677 (N_5677,N_2840,N_4467);
or U5678 (N_5678,N_3849,N_4650);
nor U5679 (N_5679,N_3279,N_3243);
nor U5680 (N_5680,N_4853,N_4648);
nor U5681 (N_5681,N_4528,N_2810);
xnor U5682 (N_5682,N_3288,N_4364);
nand U5683 (N_5683,N_2539,N_4904);
xnor U5684 (N_5684,N_4785,N_4858);
nor U5685 (N_5685,N_3427,N_2632);
and U5686 (N_5686,N_4820,N_3630);
or U5687 (N_5687,N_2638,N_3219);
and U5688 (N_5688,N_3654,N_4165);
xnor U5689 (N_5689,N_3544,N_4149);
nor U5690 (N_5690,N_3416,N_2534);
nand U5691 (N_5691,N_2860,N_4534);
nor U5692 (N_5692,N_3627,N_3015);
nor U5693 (N_5693,N_4112,N_2725);
xnor U5694 (N_5694,N_2987,N_4948);
xor U5695 (N_5695,N_4711,N_4683);
nand U5696 (N_5696,N_4992,N_4876);
xor U5697 (N_5697,N_3563,N_3103);
nand U5698 (N_5698,N_3650,N_4428);
nor U5699 (N_5699,N_4155,N_4740);
and U5700 (N_5700,N_2641,N_3498);
xor U5701 (N_5701,N_3525,N_4641);
nand U5702 (N_5702,N_4604,N_3872);
nor U5703 (N_5703,N_4158,N_4753);
or U5704 (N_5704,N_4839,N_4665);
and U5705 (N_5705,N_3261,N_3923);
nand U5706 (N_5706,N_4386,N_4346);
nand U5707 (N_5707,N_2570,N_4849);
nor U5708 (N_5708,N_3845,N_4608);
xnor U5709 (N_5709,N_3458,N_3410);
and U5710 (N_5710,N_3957,N_3749);
xor U5711 (N_5711,N_2828,N_2887);
nand U5712 (N_5712,N_3269,N_3786);
or U5713 (N_5713,N_3960,N_2754);
nor U5714 (N_5714,N_4593,N_2529);
nand U5715 (N_5715,N_3177,N_4169);
and U5716 (N_5716,N_2871,N_3415);
nand U5717 (N_5717,N_3250,N_4518);
xor U5718 (N_5718,N_2509,N_3649);
nor U5719 (N_5719,N_3246,N_3701);
or U5720 (N_5720,N_2668,N_3659);
and U5721 (N_5721,N_2816,N_3488);
nand U5722 (N_5722,N_3237,N_2635);
xnor U5723 (N_5723,N_2593,N_2624);
and U5724 (N_5724,N_4464,N_3585);
xnor U5725 (N_5725,N_3106,N_2994);
xnor U5726 (N_5726,N_4961,N_4003);
nor U5727 (N_5727,N_4995,N_3200);
or U5728 (N_5728,N_4617,N_4061);
and U5729 (N_5729,N_4170,N_3363);
and U5730 (N_5730,N_4889,N_3519);
and U5731 (N_5731,N_4233,N_2716);
or U5732 (N_5732,N_2591,N_2909);
xnor U5733 (N_5733,N_4900,N_2762);
or U5734 (N_5734,N_2702,N_2788);
nor U5735 (N_5735,N_4877,N_4309);
or U5736 (N_5736,N_4135,N_2586);
and U5737 (N_5737,N_3894,N_3796);
nand U5738 (N_5738,N_3278,N_3712);
and U5739 (N_5739,N_4382,N_4735);
nand U5740 (N_5740,N_2799,N_3803);
nand U5741 (N_5741,N_4986,N_3848);
nor U5742 (N_5742,N_3983,N_2941);
or U5743 (N_5743,N_4626,N_4828);
or U5744 (N_5744,N_4919,N_4159);
xnor U5745 (N_5745,N_4848,N_3087);
and U5746 (N_5746,N_3395,N_3429);
and U5747 (N_5747,N_4197,N_2541);
xnor U5748 (N_5748,N_4761,N_3055);
nor U5749 (N_5749,N_3130,N_3699);
nand U5750 (N_5750,N_3197,N_4667);
nor U5751 (N_5751,N_4088,N_3483);
xor U5752 (N_5752,N_4421,N_4533);
and U5753 (N_5753,N_2646,N_4164);
nor U5754 (N_5754,N_4750,N_4063);
nand U5755 (N_5755,N_3298,N_3343);
and U5756 (N_5756,N_3792,N_4520);
nand U5757 (N_5757,N_4500,N_3274);
xnor U5758 (N_5758,N_4077,N_3876);
nand U5759 (N_5759,N_3442,N_4343);
nand U5760 (N_5760,N_4602,N_3248);
nor U5761 (N_5761,N_3066,N_4905);
nand U5762 (N_5762,N_3835,N_4374);
and U5763 (N_5763,N_3305,N_2829);
and U5764 (N_5764,N_3862,N_4064);
nand U5765 (N_5765,N_4205,N_4289);
or U5766 (N_5766,N_2550,N_3388);
and U5767 (N_5767,N_3667,N_3281);
xor U5768 (N_5768,N_3258,N_3104);
and U5769 (N_5769,N_4490,N_4748);
xor U5770 (N_5770,N_4402,N_4965);
or U5771 (N_5771,N_3336,N_2998);
or U5772 (N_5772,N_3722,N_4047);
xor U5773 (N_5773,N_2674,N_4127);
and U5774 (N_5774,N_4816,N_2736);
nand U5775 (N_5775,N_2752,N_4476);
nor U5776 (N_5776,N_4639,N_4071);
xor U5777 (N_5777,N_4466,N_3689);
or U5778 (N_5778,N_2675,N_3489);
nor U5779 (N_5779,N_2967,N_3476);
xor U5780 (N_5780,N_3111,N_3394);
nor U5781 (N_5781,N_3730,N_3364);
nand U5782 (N_5782,N_3044,N_3347);
or U5783 (N_5783,N_3433,N_4600);
nand U5784 (N_5784,N_3326,N_3341);
nor U5785 (N_5785,N_2997,N_2517);
or U5786 (N_5786,N_4404,N_3856);
nand U5787 (N_5787,N_4297,N_4893);
or U5788 (N_5788,N_4783,N_4035);
and U5789 (N_5789,N_3571,N_2983);
nor U5790 (N_5790,N_2535,N_3272);
xor U5791 (N_5791,N_2936,N_3472);
nand U5792 (N_5792,N_4110,N_4388);
xnor U5793 (N_5793,N_4376,N_4888);
or U5794 (N_5794,N_3944,N_3516);
nand U5795 (N_5795,N_3716,N_3642);
nand U5796 (N_5796,N_2891,N_2751);
nor U5797 (N_5797,N_3023,N_4201);
nand U5798 (N_5798,N_3807,N_2639);
or U5799 (N_5799,N_3622,N_3965);
nand U5800 (N_5800,N_4803,N_2521);
nand U5801 (N_5801,N_3888,N_3981);
or U5802 (N_5802,N_4911,N_3063);
or U5803 (N_5803,N_3402,N_3122);
xor U5804 (N_5804,N_4558,N_4976);
xor U5805 (N_5805,N_4586,N_2695);
or U5806 (N_5806,N_4055,N_4097);
and U5807 (N_5807,N_4759,N_2618);
xnor U5808 (N_5808,N_4504,N_4784);
xnor U5809 (N_5809,N_3464,N_4234);
nor U5810 (N_5810,N_3132,N_3762);
or U5811 (N_5811,N_2526,N_4597);
or U5812 (N_5812,N_2854,N_4066);
and U5813 (N_5813,N_3163,N_2939);
and U5814 (N_5814,N_4714,N_4021);
xnor U5815 (N_5815,N_3085,N_4219);
or U5816 (N_5816,N_3603,N_4980);
xor U5817 (N_5817,N_2911,N_4115);
nand U5818 (N_5818,N_4042,N_3228);
or U5819 (N_5819,N_3397,N_3373);
xnor U5820 (N_5820,N_2555,N_3321);
xnor U5821 (N_5821,N_4819,N_4435);
xnor U5822 (N_5822,N_4764,N_3624);
or U5823 (N_5823,N_4689,N_4487);
xnor U5824 (N_5824,N_2722,N_3738);
xor U5825 (N_5825,N_2789,N_3612);
xor U5826 (N_5826,N_3644,N_4319);
and U5827 (N_5827,N_2832,N_3506);
nand U5828 (N_5828,N_2703,N_4294);
nor U5829 (N_5829,N_4299,N_2931);
nand U5830 (N_5830,N_3906,N_3962);
nand U5831 (N_5831,N_3533,N_4399);
and U5832 (N_5832,N_4561,N_3033);
and U5833 (N_5833,N_2700,N_4393);
nor U5834 (N_5834,N_2822,N_4514);
xor U5835 (N_5835,N_3798,N_4859);
xor U5836 (N_5836,N_3686,N_2971);
or U5837 (N_5837,N_3703,N_4474);
nand U5838 (N_5838,N_4313,N_3102);
and U5839 (N_5839,N_3911,N_4361);
nand U5840 (N_5840,N_3275,N_3454);
xnor U5841 (N_5841,N_4729,N_4050);
nor U5842 (N_5842,N_4899,N_4830);
nor U5843 (N_5843,N_4969,N_4811);
or U5844 (N_5844,N_3873,N_4564);
or U5845 (N_5845,N_3717,N_3724);
nor U5846 (N_5846,N_3444,N_3631);
or U5847 (N_5847,N_3993,N_4433);
xnor U5848 (N_5848,N_4144,N_4896);
or U5849 (N_5849,N_4215,N_4958);
and U5850 (N_5850,N_3159,N_4700);
or U5851 (N_5851,N_3045,N_2879);
nand U5852 (N_5852,N_2930,N_2976);
xor U5853 (N_5853,N_3898,N_4020);
nand U5854 (N_5854,N_3836,N_4023);
xor U5855 (N_5855,N_3507,N_3040);
nor U5856 (N_5856,N_4599,N_3931);
and U5857 (N_5857,N_4180,N_3184);
and U5858 (N_5858,N_3643,N_2515);
nand U5859 (N_5859,N_2953,N_3131);
or U5860 (N_5860,N_3509,N_4246);
xnor U5861 (N_5861,N_3772,N_3740);
xor U5862 (N_5862,N_3294,N_2680);
xnor U5863 (N_5863,N_3233,N_3502);
and U5864 (N_5864,N_4480,N_3470);
nand U5865 (N_5865,N_4253,N_3776);
nand U5866 (N_5866,N_3996,N_4895);
nor U5867 (N_5867,N_3026,N_3359);
xor U5868 (N_5868,N_3942,N_3711);
or U5869 (N_5869,N_4468,N_3300);
nand U5870 (N_5870,N_3688,N_4004);
nand U5871 (N_5871,N_3771,N_2609);
nand U5872 (N_5872,N_3318,N_4823);
and U5873 (N_5873,N_4539,N_4475);
and U5874 (N_5874,N_3234,N_2581);
or U5875 (N_5875,N_4672,N_3956);
or U5876 (N_5876,N_2734,N_3921);
nor U5877 (N_5877,N_4111,N_4942);
or U5878 (N_5878,N_3175,N_3432);
xor U5879 (N_5879,N_3777,N_4832);
or U5880 (N_5880,N_4496,N_2917);
nor U5881 (N_5881,N_4222,N_3312);
and U5882 (N_5882,N_3182,N_2522);
xor U5883 (N_5883,N_3718,N_2560);
and U5884 (N_5884,N_4988,N_3192);
nand U5885 (N_5885,N_4019,N_3155);
nand U5886 (N_5886,N_4463,N_4742);
xnor U5887 (N_5887,N_3058,N_4727);
xor U5888 (N_5888,N_3503,N_3094);
xor U5889 (N_5889,N_2830,N_3379);
xor U5890 (N_5890,N_2537,N_3353);
or U5891 (N_5891,N_3404,N_3945);
xor U5892 (N_5892,N_4385,N_2705);
nand U5893 (N_5893,N_3494,N_3046);
nor U5894 (N_5894,N_2999,N_4922);
and U5895 (N_5895,N_2682,N_4981);
or U5896 (N_5896,N_4979,N_4340);
or U5897 (N_5897,N_4932,N_4934);
nand U5898 (N_5898,N_4596,N_2991);
xnor U5899 (N_5899,N_4797,N_3259);
nand U5900 (N_5900,N_4405,N_2831);
nor U5901 (N_5901,N_2905,N_3419);
nand U5902 (N_5902,N_4747,N_4154);
or U5903 (N_5903,N_4292,N_4560);
xnor U5904 (N_5904,N_3656,N_3582);
or U5905 (N_5905,N_4840,N_4573);
nand U5906 (N_5906,N_4070,N_4175);
nand U5907 (N_5907,N_4912,N_3657);
nand U5908 (N_5908,N_2995,N_4497);
nor U5909 (N_5909,N_4570,N_2956);
xor U5910 (N_5910,N_3435,N_4493);
nor U5911 (N_5911,N_2776,N_4142);
nand U5912 (N_5912,N_4581,N_2797);
and U5913 (N_5913,N_4273,N_4936);
nor U5914 (N_5914,N_3940,N_3487);
nand U5915 (N_5915,N_2844,N_2811);
or U5916 (N_5916,N_3380,N_3317);
nor U5917 (N_5917,N_2992,N_4151);
or U5918 (N_5918,N_2793,N_3637);
xnor U5919 (N_5919,N_4065,N_4954);
xor U5920 (N_5920,N_3036,N_4272);
xor U5921 (N_5921,N_3361,N_3480);
nor U5922 (N_5922,N_3723,N_3999);
nor U5923 (N_5923,N_3791,N_3934);
and U5924 (N_5924,N_4163,N_4394);
or U5925 (N_5925,N_3078,N_3596);
nand U5926 (N_5926,N_4925,N_4417);
or U5927 (N_5927,N_3673,N_4554);
nand U5928 (N_5928,N_3751,N_4302);
xor U5929 (N_5929,N_4733,N_3417);
nand U5930 (N_5930,N_4918,N_2872);
nor U5931 (N_5931,N_4280,N_4781);
nor U5932 (N_5932,N_3009,N_3474);
nand U5933 (N_5933,N_3613,N_4536);
nand U5934 (N_5934,N_4322,N_4090);
or U5935 (N_5935,N_3634,N_2965);
nand U5936 (N_5936,N_4183,N_3580);
or U5937 (N_5937,N_4156,N_4960);
xor U5938 (N_5938,N_3372,N_3947);
or U5939 (N_5939,N_4870,N_3692);
nor U5940 (N_5940,N_2613,N_4612);
or U5941 (N_5941,N_4531,N_4350);
nand U5942 (N_5942,N_4719,N_3137);
or U5943 (N_5943,N_3405,N_3994);
nor U5944 (N_5944,N_3819,N_3420);
and U5945 (N_5945,N_3885,N_3839);
xnor U5946 (N_5946,N_4668,N_4914);
nor U5947 (N_5947,N_3316,N_3176);
and U5948 (N_5948,N_4256,N_4363);
xor U5949 (N_5949,N_3355,N_2935);
or U5950 (N_5950,N_3932,N_2710);
nor U5951 (N_5951,N_2687,N_2630);
or U5952 (N_5952,N_2862,N_3910);
and U5953 (N_5953,N_4780,N_4838);
xnor U5954 (N_5954,N_2699,N_3169);
nand U5955 (N_5955,N_3284,N_4978);
xor U5956 (N_5956,N_2808,N_3926);
or U5957 (N_5957,N_4126,N_3748);
or U5958 (N_5958,N_3600,N_4886);
nor U5959 (N_5959,N_4682,N_3521);
xor U5960 (N_5960,N_4461,N_2501);
xor U5961 (N_5961,N_2557,N_4732);
nand U5962 (N_5962,N_3083,N_4068);
and U5963 (N_5963,N_4230,N_4867);
nand U5964 (N_5964,N_4866,N_3232);
or U5965 (N_5965,N_4094,N_4538);
nor U5966 (N_5966,N_4546,N_4153);
and U5967 (N_5967,N_4696,N_2969);
or U5968 (N_5968,N_3139,N_4193);
or U5969 (N_5969,N_3236,N_3820);
xor U5970 (N_5970,N_3827,N_2874);
or U5971 (N_5971,N_3605,N_4887);
or U5972 (N_5972,N_3998,N_4117);
xor U5973 (N_5973,N_2903,N_3117);
nor U5974 (N_5974,N_4359,N_4287);
nand U5975 (N_5975,N_2913,N_3260);
xor U5976 (N_5976,N_4351,N_4096);
or U5977 (N_5977,N_3523,N_3559);
or U5978 (N_5978,N_3054,N_4544);
nor U5979 (N_5979,N_4818,N_2690);
nand U5980 (N_5980,N_3789,N_4275);
xor U5981 (N_5981,N_4211,N_2661);
or U5982 (N_5982,N_4666,N_2625);
xor U5983 (N_5983,N_4852,N_4930);
and U5984 (N_5984,N_4704,N_2753);
nand U5985 (N_5985,N_4355,N_3451);
and U5986 (N_5986,N_4471,N_4372);
nor U5987 (N_5987,N_3479,N_4813);
nand U5988 (N_5988,N_3095,N_4391);
or U5989 (N_5989,N_2975,N_4227);
nand U5990 (N_5990,N_4868,N_4389);
nor U5991 (N_5991,N_2577,N_4863);
and U5992 (N_5992,N_2958,N_2696);
nor U5993 (N_5993,N_2538,N_3212);
and U5994 (N_5994,N_2746,N_4767);
nor U5995 (N_5995,N_2784,N_3335);
nor U5996 (N_5996,N_4443,N_2650);
xor U5997 (N_5997,N_4336,N_2835);
xnor U5998 (N_5998,N_3271,N_3874);
nand U5999 (N_5999,N_4267,N_4883);
xor U6000 (N_6000,N_3621,N_3889);
and U6001 (N_6001,N_4191,N_2549);
or U6002 (N_6002,N_2670,N_3514);
or U6003 (N_6003,N_3189,N_2567);
nand U6004 (N_6004,N_4037,N_4469);
and U6005 (N_6005,N_2616,N_2989);
nor U6006 (N_6006,N_3958,N_4354);
nor U6007 (N_6007,N_2584,N_3967);
xor U6008 (N_6008,N_3577,N_4357);
xor U6009 (N_6009,N_2595,N_3492);
nand U6010 (N_6010,N_4260,N_3768);
xnor U6011 (N_6011,N_3050,N_3385);
or U6012 (N_6012,N_3141,N_4552);
or U6013 (N_6013,N_4854,N_4898);
or U6014 (N_6014,N_2615,N_3567);
nor U6015 (N_6015,N_3473,N_2839);
nor U6016 (N_6016,N_2943,N_2928);
nand U6017 (N_6017,N_3453,N_4283);
nand U6018 (N_6018,N_3865,N_2914);
and U6019 (N_6019,N_3802,N_3804);
and U6020 (N_6020,N_4713,N_4790);
xor U6021 (N_6021,N_4138,N_4829);
xor U6022 (N_6022,N_4584,N_2547);
nor U6023 (N_6023,N_4429,N_4213);
xor U6024 (N_6024,N_4836,N_4254);
or U6025 (N_6025,N_3207,N_4737);
xnor U6026 (N_6026,N_4439,N_3110);
and U6027 (N_6027,N_3615,N_3709);
nor U6028 (N_6028,N_3546,N_2663);
nand U6029 (N_6029,N_3793,N_3854);
xnor U6030 (N_6030,N_2551,N_2566);
nand U6031 (N_6031,N_2948,N_3623);
or U6032 (N_6032,N_3490,N_3662);
xnor U6033 (N_6033,N_2514,N_3185);
xnor U6034 (N_6034,N_3482,N_2671);
nand U6035 (N_6035,N_4203,N_2790);
nor U6036 (N_6036,N_4618,N_2771);
or U6037 (N_6037,N_4636,N_3346);
and U6038 (N_6038,N_2513,N_3731);
or U6039 (N_6039,N_4562,N_4582);
nor U6040 (N_6040,N_4161,N_4598);
and U6041 (N_6041,N_4016,N_4145);
nand U6042 (N_6042,N_4837,N_4875);
nor U6043 (N_6043,N_3134,N_4664);
xnor U6044 (N_6044,N_4770,N_3828);
nand U6045 (N_6045,N_4166,N_4259);
xnor U6046 (N_6046,N_4678,N_4763);
xor U6047 (N_6047,N_4762,N_3345);
and U6048 (N_6048,N_3478,N_4542);
xnor U6049 (N_6049,N_2607,N_3601);
and U6050 (N_6050,N_4592,N_3138);
xor U6051 (N_6051,N_4217,N_2711);
nand U6052 (N_6052,N_4684,N_3858);
nor U6053 (N_6053,N_4967,N_3541);
xnor U6054 (N_6054,N_3850,N_4894);
nor U6055 (N_6055,N_4384,N_4375);
or U6056 (N_6056,N_4575,N_4296);
and U6057 (N_6057,N_4935,N_2738);
and U6058 (N_6058,N_4955,N_3421);
nand U6059 (N_6059,N_4250,N_4845);
nor U6060 (N_6060,N_3016,N_4242);
nor U6061 (N_6061,N_3443,N_3072);
and U6062 (N_6062,N_3916,N_4268);
or U6063 (N_6063,N_4140,N_4450);
nand U6064 (N_6064,N_4633,N_4634);
and U6065 (N_6065,N_4991,N_2603);
xor U6066 (N_6066,N_3961,N_2834);
nand U6067 (N_6067,N_3867,N_3448);
or U6068 (N_6068,N_2923,N_4196);
xor U6069 (N_6069,N_3365,N_4045);
nand U6070 (N_6070,N_3863,N_4281);
and U6071 (N_6071,N_3324,N_3536);
nor U6072 (N_6072,N_2902,N_4288);
nor U6073 (N_6073,N_4377,N_3568);
nand U6074 (N_6074,N_4726,N_3329);
nand U6075 (N_6075,N_3929,N_4032);
nor U6076 (N_6076,N_4557,N_4485);
xnor U6077 (N_6077,N_3295,N_3781);
xor U6078 (N_6078,N_3880,N_4754);
nor U6079 (N_6079,N_3924,N_3062);
and U6080 (N_6080,N_4548,N_3658);
nor U6081 (N_6081,N_3455,N_4606);
nor U6082 (N_6082,N_3935,N_4119);
or U6083 (N_6083,N_3908,N_4451);
nand U6084 (N_6084,N_4457,N_3157);
xor U6085 (N_6085,N_4751,N_3763);
xor U6086 (N_6086,N_3133,N_2821);
and U6087 (N_6087,N_4635,N_4181);
xnor U6088 (N_6088,N_4447,N_3392);
or U6089 (N_6089,N_2597,N_4695);
nor U6090 (N_6090,N_4419,N_3017);
or U6091 (N_6091,N_3447,N_3538);
and U6092 (N_6092,N_3367,N_3501);
nor U6093 (N_6093,N_4734,N_3143);
nand U6094 (N_6094,N_2977,N_4353);
nand U6095 (N_6095,N_3322,N_4549);
xnor U6096 (N_6096,N_3314,N_3187);
and U6097 (N_6097,N_4872,N_2865);
and U6098 (N_6098,N_2588,N_4792);
or U6099 (N_6099,N_3338,N_2852);
nor U6100 (N_6100,N_4953,N_2602);
xnor U6101 (N_6101,N_4999,N_2926);
or U6102 (N_6102,N_2727,N_4555);
nand U6103 (N_6103,N_4833,N_3357);
xnor U6104 (N_6104,N_4013,N_2572);
nand U6105 (N_6105,N_3859,N_2735);
nor U6106 (N_6106,N_3210,N_4335);
and U6107 (N_6107,N_3067,N_2819);
nand U6108 (N_6108,N_2882,N_4587);
nand U6109 (N_6109,N_2791,N_4543);
nand U6110 (N_6110,N_3773,N_4506);
and U6111 (N_6111,N_2984,N_3086);
nor U6112 (N_6112,N_3211,N_3542);
xnor U6113 (N_6113,N_3752,N_4235);
and U6114 (N_6114,N_3675,N_3655);
and U6115 (N_6115,N_3681,N_2842);
or U6116 (N_6116,N_4577,N_2655);
or U6117 (N_6117,N_2580,N_4187);
nand U6118 (N_6118,N_3180,N_3145);
nand U6119 (N_6119,N_4132,N_3434);
xor U6120 (N_6120,N_4607,N_4285);
xor U6121 (N_6121,N_3560,N_2527);
or U6122 (N_6122,N_2656,N_3635);
xnor U6123 (N_6123,N_4438,N_2508);
and U6124 (N_6124,N_4030,N_4462);
nand U6125 (N_6125,N_2652,N_4959);
nor U6126 (N_6126,N_3495,N_3977);
nand U6127 (N_6127,N_3735,N_3034);
nor U6128 (N_6128,N_4214,N_4652);
nor U6129 (N_6129,N_4373,N_3263);
and U6130 (N_6130,N_2693,N_3241);
nand U6131 (N_6131,N_3866,N_4100);
or U6132 (N_6132,N_3135,N_2691);
nand U6133 (N_6133,N_4698,N_4594);
nor U6134 (N_6134,N_2978,N_3747);
and U6135 (N_6135,N_3851,N_4798);
and U6136 (N_6136,N_4724,N_3047);
nor U6137 (N_6137,N_3118,N_4456);
and U6138 (N_6138,N_4788,N_4266);
nand U6139 (N_6139,N_2775,N_4445);
xor U6140 (N_6140,N_2766,N_4802);
xor U6141 (N_6141,N_3950,N_3970);
xnor U6142 (N_6142,N_4681,N_4709);
xor U6143 (N_6143,N_4843,N_3989);
or U6144 (N_6144,N_3857,N_2837);
nor U6145 (N_6145,N_4278,N_2878);
or U6146 (N_6146,N_2841,N_4631);
nand U6147 (N_6147,N_2536,N_3927);
xnor U6148 (N_6148,N_3808,N_4228);
nand U6149 (N_6149,N_3512,N_3903);
xor U6150 (N_6150,N_2759,N_4473);
nor U6151 (N_6151,N_3632,N_3008);
nor U6152 (N_6152,N_3778,N_4851);
xor U6153 (N_6153,N_3438,N_4448);
nor U6154 (N_6154,N_3690,N_3090);
nand U6155 (N_6155,N_3469,N_3554);
and U6156 (N_6156,N_2889,N_3101);
and U6157 (N_6157,N_3588,N_3254);
nor U6158 (N_6158,N_3682,N_3010);
nand U6159 (N_6159,N_3203,N_3172);
or U6160 (N_6160,N_4200,N_4210);
and U6161 (N_6161,N_2571,N_4717);
or U6162 (N_6162,N_2805,N_4841);
nand U6163 (N_6163,N_4459,N_4005);
or U6164 (N_6164,N_4182,N_3788);
nand U6165 (N_6165,N_4329,N_4301);
or U6166 (N_6166,N_3758,N_4749);
and U6167 (N_6167,N_4311,N_4588);
and U6168 (N_6168,N_2925,N_3831);
nand U6169 (N_6169,N_4143,N_4628);
nand U6170 (N_6170,N_2937,N_4809);
xor U6171 (N_6171,N_2623,N_3830);
nand U6172 (N_6172,N_2543,N_4043);
and U6173 (N_6173,N_3244,N_4697);
and U6174 (N_6174,N_4041,N_2750);
nand U6175 (N_6175,N_4365,N_2542);
or U6176 (N_6176,N_4884,N_2957);
nor U6177 (N_6177,N_2912,N_3522);
nor U6178 (N_6178,N_2564,N_4651);
nor U6179 (N_6179,N_2833,N_2807);
xor U6180 (N_6180,N_4085,N_3493);
and U6181 (N_6181,N_3707,N_2915);
nand U6182 (N_6182,N_2813,N_3754);
nand U6183 (N_6183,N_4146,N_2798);
nand U6184 (N_6184,N_4676,N_2755);
nor U6185 (N_6185,N_3449,N_3558);
or U6186 (N_6186,N_2739,N_4220);
or U6187 (N_6187,N_2924,N_2908);
or U6188 (N_6188,N_3074,N_3907);
and U6189 (N_6189,N_3928,N_3127);
nand U6190 (N_6190,N_4789,N_3283);
xnor U6191 (N_6191,N_3393,N_2972);
or U6192 (N_6192,N_3218,N_3510);
and U6193 (N_6193,N_3107,N_3484);
and U6194 (N_6194,N_3645,N_2647);
and U6195 (N_6195,N_2627,N_3527);
and U6196 (N_6196,N_2780,N_4501);
or U6197 (N_6197,N_2576,N_2985);
nor U6198 (N_6198,N_4481,N_2737);
or U6199 (N_6199,N_3564,N_2963);
xnor U6200 (N_6200,N_2679,N_4453);
nor U6201 (N_6201,N_3296,N_3869);
nor U6202 (N_6202,N_3401,N_4312);
or U6203 (N_6203,N_3108,N_3381);
xnor U6204 (N_6204,N_2818,N_4121);
nor U6205 (N_6205,N_3154,N_3821);
nand U6206 (N_6206,N_3371,N_3594);
xnor U6207 (N_6207,N_4251,N_4847);
and U6208 (N_6208,N_2686,N_2781);
nand U6209 (N_6209,N_3238,N_3691);
nand U6210 (N_6210,N_4688,N_2981);
or U6211 (N_6211,N_4985,N_4131);
nor U6212 (N_6212,N_2720,N_3518);
xor U6213 (N_6213,N_4295,N_3920);
xor U6214 (N_6214,N_3038,N_4576);
nor U6215 (N_6215,N_4423,N_2986);
or U6216 (N_6216,N_4921,N_3290);
nor U6217 (N_6217,N_3018,N_4972);
and U6218 (N_6218,N_3893,N_4208);
and U6219 (N_6219,N_4649,N_3765);
and U6220 (N_6220,N_4962,N_2617);
and U6221 (N_6221,N_4505,N_3377);
and U6222 (N_6222,N_3048,N_4566);
or U6223 (N_6223,N_4326,N_3057);
nor U6224 (N_6224,N_2692,N_4537);
or U6225 (N_6225,N_2968,N_2918);
and U6226 (N_6226,N_3905,N_4571);
and U6227 (N_6227,N_4629,N_3652);
and U6228 (N_6228,N_3602,N_4347);
nor U6229 (N_6229,N_4806,N_2796);
xnor U6230 (N_6230,N_4947,N_4060);
or U6231 (N_6231,N_4670,N_3061);
and U6232 (N_6232,N_4706,N_3847);
and U6233 (N_6233,N_3552,N_3760);
xnor U6234 (N_6234,N_4320,N_4216);
and U6235 (N_6235,N_4939,N_3309);
xor U6236 (N_6236,N_4522,N_3714);
and U6237 (N_6237,N_3186,N_4074);
xnor U6238 (N_6238,N_4204,N_3968);
nor U6239 (N_6239,N_4293,N_2653);
or U6240 (N_6240,N_4378,N_3408);
and U6241 (N_6241,N_4860,N_2772);
and U6242 (N_6242,N_4694,N_2980);
and U6243 (N_6243,N_3997,N_3721);
or U6244 (N_6244,N_4739,N_4491);
xnor U6245 (N_6245,N_3895,N_3019);
nand U6246 (N_6246,N_4946,N_3734);
or U6247 (N_6247,N_4741,N_3593);
or U6248 (N_6248,N_4483,N_3307);
nor U6249 (N_6249,N_4601,N_3761);
xor U6250 (N_6250,N_3028,N_4957);
xnor U6251 (N_6251,N_3442,N_3640);
xnor U6252 (N_6252,N_2958,N_4017);
nand U6253 (N_6253,N_2512,N_3543);
nor U6254 (N_6254,N_4356,N_4841);
xor U6255 (N_6255,N_4771,N_2918);
nand U6256 (N_6256,N_4762,N_4760);
or U6257 (N_6257,N_2579,N_2653);
xnor U6258 (N_6258,N_2799,N_3086);
or U6259 (N_6259,N_3374,N_3987);
or U6260 (N_6260,N_3252,N_3871);
and U6261 (N_6261,N_2525,N_2739);
and U6262 (N_6262,N_4820,N_4921);
nand U6263 (N_6263,N_2873,N_2579);
and U6264 (N_6264,N_4926,N_3859);
and U6265 (N_6265,N_4967,N_3967);
or U6266 (N_6266,N_4260,N_3407);
xnor U6267 (N_6267,N_3297,N_4093);
nor U6268 (N_6268,N_3515,N_3037);
xnor U6269 (N_6269,N_4872,N_3079);
nor U6270 (N_6270,N_3478,N_4336);
or U6271 (N_6271,N_4951,N_3955);
or U6272 (N_6272,N_4487,N_3051);
nor U6273 (N_6273,N_2591,N_3607);
and U6274 (N_6274,N_4311,N_3360);
nor U6275 (N_6275,N_3397,N_4332);
or U6276 (N_6276,N_3055,N_4857);
nor U6277 (N_6277,N_2649,N_3718);
xnor U6278 (N_6278,N_3073,N_3438);
nor U6279 (N_6279,N_4282,N_4458);
xnor U6280 (N_6280,N_2994,N_2620);
and U6281 (N_6281,N_4968,N_4019);
nand U6282 (N_6282,N_2697,N_3984);
and U6283 (N_6283,N_3252,N_4917);
nand U6284 (N_6284,N_3814,N_2777);
nor U6285 (N_6285,N_3463,N_4550);
and U6286 (N_6286,N_3332,N_4150);
nand U6287 (N_6287,N_3080,N_3339);
xor U6288 (N_6288,N_4829,N_3957);
or U6289 (N_6289,N_3199,N_3575);
nand U6290 (N_6290,N_4056,N_3817);
or U6291 (N_6291,N_3336,N_2965);
xnor U6292 (N_6292,N_4669,N_4639);
and U6293 (N_6293,N_4775,N_3181);
nand U6294 (N_6294,N_4351,N_3224);
xor U6295 (N_6295,N_4596,N_4649);
or U6296 (N_6296,N_4857,N_4041);
or U6297 (N_6297,N_2621,N_2670);
or U6298 (N_6298,N_2892,N_3482);
and U6299 (N_6299,N_3211,N_4498);
nand U6300 (N_6300,N_4593,N_3475);
or U6301 (N_6301,N_4132,N_4617);
xor U6302 (N_6302,N_4985,N_3739);
nand U6303 (N_6303,N_2926,N_2792);
and U6304 (N_6304,N_2805,N_4415);
and U6305 (N_6305,N_3669,N_4640);
nor U6306 (N_6306,N_4459,N_4724);
nand U6307 (N_6307,N_4734,N_3268);
xnor U6308 (N_6308,N_4496,N_4656);
xor U6309 (N_6309,N_3622,N_4791);
nand U6310 (N_6310,N_2565,N_4792);
and U6311 (N_6311,N_2525,N_2973);
or U6312 (N_6312,N_4252,N_2859);
and U6313 (N_6313,N_3988,N_3853);
or U6314 (N_6314,N_4893,N_4842);
xnor U6315 (N_6315,N_3523,N_2762);
and U6316 (N_6316,N_3618,N_3237);
or U6317 (N_6317,N_2583,N_3535);
or U6318 (N_6318,N_2674,N_3917);
nor U6319 (N_6319,N_3494,N_3974);
nand U6320 (N_6320,N_2921,N_3494);
or U6321 (N_6321,N_2931,N_3576);
xnor U6322 (N_6322,N_2839,N_4083);
nor U6323 (N_6323,N_2663,N_3349);
or U6324 (N_6324,N_3010,N_3439);
and U6325 (N_6325,N_4865,N_4712);
or U6326 (N_6326,N_3140,N_3047);
nand U6327 (N_6327,N_2600,N_2520);
nand U6328 (N_6328,N_3825,N_4381);
nand U6329 (N_6329,N_4820,N_3154);
and U6330 (N_6330,N_4320,N_2521);
xnor U6331 (N_6331,N_4874,N_2964);
xor U6332 (N_6332,N_2698,N_3197);
and U6333 (N_6333,N_4624,N_4238);
nor U6334 (N_6334,N_4092,N_4498);
nor U6335 (N_6335,N_2968,N_4642);
xnor U6336 (N_6336,N_4896,N_4701);
nor U6337 (N_6337,N_2658,N_2552);
nor U6338 (N_6338,N_4175,N_4789);
or U6339 (N_6339,N_3244,N_3422);
nor U6340 (N_6340,N_4641,N_2530);
or U6341 (N_6341,N_3966,N_4239);
nand U6342 (N_6342,N_4981,N_3169);
xnor U6343 (N_6343,N_4990,N_4705);
nand U6344 (N_6344,N_4930,N_2923);
or U6345 (N_6345,N_4329,N_4082);
and U6346 (N_6346,N_4071,N_3164);
and U6347 (N_6347,N_2946,N_4551);
and U6348 (N_6348,N_4954,N_4274);
and U6349 (N_6349,N_4337,N_3745);
xor U6350 (N_6350,N_2725,N_4292);
and U6351 (N_6351,N_4645,N_2782);
or U6352 (N_6352,N_3377,N_3538);
and U6353 (N_6353,N_3463,N_4185);
nand U6354 (N_6354,N_3687,N_3148);
and U6355 (N_6355,N_3675,N_4387);
and U6356 (N_6356,N_3286,N_4221);
nor U6357 (N_6357,N_4569,N_3905);
nand U6358 (N_6358,N_4334,N_4429);
and U6359 (N_6359,N_4934,N_2868);
nand U6360 (N_6360,N_3930,N_3906);
and U6361 (N_6361,N_3804,N_3521);
or U6362 (N_6362,N_3331,N_3655);
nor U6363 (N_6363,N_3607,N_3534);
and U6364 (N_6364,N_2818,N_2655);
xor U6365 (N_6365,N_2846,N_3909);
nor U6366 (N_6366,N_3897,N_2954);
or U6367 (N_6367,N_4973,N_4497);
or U6368 (N_6368,N_3559,N_3743);
xnor U6369 (N_6369,N_4780,N_3768);
nor U6370 (N_6370,N_3908,N_2535);
or U6371 (N_6371,N_3961,N_4754);
nor U6372 (N_6372,N_4150,N_3574);
nand U6373 (N_6373,N_3957,N_2785);
xnor U6374 (N_6374,N_3515,N_4863);
and U6375 (N_6375,N_4510,N_3032);
nand U6376 (N_6376,N_3132,N_2562);
xnor U6377 (N_6377,N_3578,N_4899);
nand U6378 (N_6378,N_3063,N_4124);
xnor U6379 (N_6379,N_3521,N_2549);
nand U6380 (N_6380,N_2642,N_3472);
nor U6381 (N_6381,N_4754,N_4617);
or U6382 (N_6382,N_3638,N_2504);
nor U6383 (N_6383,N_4433,N_4717);
xnor U6384 (N_6384,N_4769,N_3981);
and U6385 (N_6385,N_3080,N_4235);
nand U6386 (N_6386,N_4792,N_4242);
nand U6387 (N_6387,N_3772,N_4276);
nor U6388 (N_6388,N_3098,N_4262);
and U6389 (N_6389,N_4818,N_3663);
nor U6390 (N_6390,N_3027,N_4880);
xor U6391 (N_6391,N_4060,N_2519);
and U6392 (N_6392,N_2764,N_3133);
or U6393 (N_6393,N_4975,N_3823);
nand U6394 (N_6394,N_4676,N_3336);
xor U6395 (N_6395,N_3726,N_3478);
or U6396 (N_6396,N_4014,N_3350);
nor U6397 (N_6397,N_3095,N_3540);
nand U6398 (N_6398,N_3783,N_3795);
and U6399 (N_6399,N_4482,N_4617);
nor U6400 (N_6400,N_3509,N_2598);
nor U6401 (N_6401,N_4056,N_4406);
nand U6402 (N_6402,N_3622,N_4876);
and U6403 (N_6403,N_4987,N_3331);
and U6404 (N_6404,N_3859,N_3118);
xnor U6405 (N_6405,N_3053,N_4801);
nor U6406 (N_6406,N_3089,N_3319);
nand U6407 (N_6407,N_2940,N_4224);
nand U6408 (N_6408,N_4871,N_3777);
nand U6409 (N_6409,N_2703,N_3426);
and U6410 (N_6410,N_4758,N_3222);
nand U6411 (N_6411,N_3685,N_4211);
and U6412 (N_6412,N_2972,N_4223);
nor U6413 (N_6413,N_4544,N_2539);
xnor U6414 (N_6414,N_4577,N_4371);
nor U6415 (N_6415,N_3205,N_4053);
and U6416 (N_6416,N_3222,N_3060);
and U6417 (N_6417,N_3557,N_2973);
or U6418 (N_6418,N_4251,N_4524);
or U6419 (N_6419,N_2610,N_3916);
and U6420 (N_6420,N_4357,N_4033);
nand U6421 (N_6421,N_4248,N_2693);
xor U6422 (N_6422,N_4947,N_4283);
nor U6423 (N_6423,N_4390,N_2507);
and U6424 (N_6424,N_4980,N_3974);
or U6425 (N_6425,N_3296,N_3643);
and U6426 (N_6426,N_4756,N_3794);
nand U6427 (N_6427,N_3307,N_3270);
and U6428 (N_6428,N_3143,N_3306);
nor U6429 (N_6429,N_4724,N_4910);
or U6430 (N_6430,N_4062,N_4212);
nor U6431 (N_6431,N_2867,N_4815);
or U6432 (N_6432,N_3664,N_2900);
and U6433 (N_6433,N_3310,N_3332);
xnor U6434 (N_6434,N_4287,N_2582);
or U6435 (N_6435,N_4766,N_2875);
nor U6436 (N_6436,N_4640,N_2507);
nor U6437 (N_6437,N_3067,N_2984);
or U6438 (N_6438,N_3471,N_4821);
xor U6439 (N_6439,N_4854,N_3035);
or U6440 (N_6440,N_2898,N_2821);
and U6441 (N_6441,N_4896,N_2811);
nor U6442 (N_6442,N_4111,N_4445);
nor U6443 (N_6443,N_4023,N_3290);
and U6444 (N_6444,N_3162,N_3487);
and U6445 (N_6445,N_4033,N_3552);
nor U6446 (N_6446,N_2822,N_4079);
xnor U6447 (N_6447,N_3171,N_4221);
nor U6448 (N_6448,N_3645,N_2754);
nor U6449 (N_6449,N_4436,N_4724);
and U6450 (N_6450,N_2510,N_4335);
and U6451 (N_6451,N_3429,N_2808);
or U6452 (N_6452,N_4388,N_4580);
xnor U6453 (N_6453,N_3838,N_4992);
nand U6454 (N_6454,N_3261,N_4301);
nor U6455 (N_6455,N_3868,N_3744);
nor U6456 (N_6456,N_3956,N_3713);
xnor U6457 (N_6457,N_3596,N_4688);
xnor U6458 (N_6458,N_3037,N_2576);
nor U6459 (N_6459,N_2898,N_4486);
or U6460 (N_6460,N_2546,N_4829);
and U6461 (N_6461,N_4514,N_4090);
or U6462 (N_6462,N_3526,N_3535);
xor U6463 (N_6463,N_2646,N_4557);
or U6464 (N_6464,N_3531,N_4752);
xnor U6465 (N_6465,N_2923,N_2726);
xnor U6466 (N_6466,N_4822,N_3808);
nand U6467 (N_6467,N_3243,N_2879);
nand U6468 (N_6468,N_4961,N_4783);
nor U6469 (N_6469,N_4077,N_2742);
or U6470 (N_6470,N_3584,N_4313);
nand U6471 (N_6471,N_3765,N_4087);
xor U6472 (N_6472,N_3153,N_3803);
nand U6473 (N_6473,N_4525,N_3486);
xnor U6474 (N_6474,N_4450,N_4865);
or U6475 (N_6475,N_3531,N_3493);
xor U6476 (N_6476,N_3889,N_4259);
or U6477 (N_6477,N_2644,N_4697);
and U6478 (N_6478,N_4994,N_2647);
xnor U6479 (N_6479,N_3767,N_2729);
xor U6480 (N_6480,N_3475,N_4351);
or U6481 (N_6481,N_2790,N_4072);
and U6482 (N_6482,N_4648,N_3328);
nor U6483 (N_6483,N_4180,N_4456);
xor U6484 (N_6484,N_3887,N_4113);
nor U6485 (N_6485,N_3243,N_3443);
nand U6486 (N_6486,N_3255,N_4962);
xor U6487 (N_6487,N_3790,N_4776);
nand U6488 (N_6488,N_4330,N_4293);
and U6489 (N_6489,N_4753,N_2969);
and U6490 (N_6490,N_4492,N_2820);
nor U6491 (N_6491,N_4704,N_3168);
and U6492 (N_6492,N_3536,N_4599);
nand U6493 (N_6493,N_3443,N_3592);
xnor U6494 (N_6494,N_4172,N_2987);
nor U6495 (N_6495,N_2818,N_4136);
xor U6496 (N_6496,N_3808,N_4173);
nor U6497 (N_6497,N_4678,N_3205);
nor U6498 (N_6498,N_2553,N_4184);
xor U6499 (N_6499,N_4736,N_3966);
xnor U6500 (N_6500,N_4005,N_4565);
nand U6501 (N_6501,N_4292,N_3061);
nand U6502 (N_6502,N_3600,N_3748);
nor U6503 (N_6503,N_4027,N_4711);
and U6504 (N_6504,N_3629,N_3084);
and U6505 (N_6505,N_2758,N_4934);
and U6506 (N_6506,N_4846,N_4651);
xor U6507 (N_6507,N_4774,N_3569);
or U6508 (N_6508,N_3351,N_3444);
or U6509 (N_6509,N_2559,N_3897);
xnor U6510 (N_6510,N_4630,N_4121);
and U6511 (N_6511,N_2926,N_4853);
nor U6512 (N_6512,N_2642,N_3266);
or U6513 (N_6513,N_3754,N_4589);
nand U6514 (N_6514,N_4163,N_3741);
nor U6515 (N_6515,N_4851,N_3478);
nand U6516 (N_6516,N_4136,N_4352);
and U6517 (N_6517,N_3840,N_4165);
nand U6518 (N_6518,N_4359,N_3667);
xor U6519 (N_6519,N_3523,N_3669);
xor U6520 (N_6520,N_3764,N_2691);
nor U6521 (N_6521,N_3300,N_2694);
nor U6522 (N_6522,N_4390,N_3856);
and U6523 (N_6523,N_4049,N_4923);
xnor U6524 (N_6524,N_4732,N_3246);
nand U6525 (N_6525,N_4758,N_3620);
xnor U6526 (N_6526,N_4818,N_2720);
or U6527 (N_6527,N_3436,N_4243);
and U6528 (N_6528,N_2927,N_3148);
or U6529 (N_6529,N_4347,N_3238);
xnor U6530 (N_6530,N_3152,N_3896);
and U6531 (N_6531,N_3789,N_3397);
nand U6532 (N_6532,N_4917,N_3753);
xnor U6533 (N_6533,N_4109,N_4694);
and U6534 (N_6534,N_2500,N_4749);
and U6535 (N_6535,N_3362,N_4187);
nand U6536 (N_6536,N_2820,N_2883);
nand U6537 (N_6537,N_3661,N_4172);
xnor U6538 (N_6538,N_2814,N_3993);
xnor U6539 (N_6539,N_3424,N_2526);
and U6540 (N_6540,N_3821,N_4911);
or U6541 (N_6541,N_3732,N_3071);
and U6542 (N_6542,N_2890,N_3760);
nor U6543 (N_6543,N_3363,N_4946);
or U6544 (N_6544,N_3422,N_4311);
and U6545 (N_6545,N_3725,N_2735);
xnor U6546 (N_6546,N_2919,N_2768);
or U6547 (N_6547,N_4860,N_4611);
or U6548 (N_6548,N_4530,N_2964);
nand U6549 (N_6549,N_2609,N_2927);
xor U6550 (N_6550,N_2570,N_4049);
nor U6551 (N_6551,N_2950,N_2652);
xor U6552 (N_6552,N_4254,N_3855);
xor U6553 (N_6553,N_4801,N_2618);
or U6554 (N_6554,N_2599,N_3491);
and U6555 (N_6555,N_3807,N_4659);
xnor U6556 (N_6556,N_4305,N_2644);
or U6557 (N_6557,N_4607,N_4371);
nor U6558 (N_6558,N_3298,N_4978);
and U6559 (N_6559,N_2617,N_3692);
nor U6560 (N_6560,N_3847,N_4724);
nand U6561 (N_6561,N_3387,N_4521);
and U6562 (N_6562,N_4798,N_4096);
xor U6563 (N_6563,N_4111,N_3847);
and U6564 (N_6564,N_4871,N_4005);
and U6565 (N_6565,N_4025,N_3007);
or U6566 (N_6566,N_4910,N_4093);
or U6567 (N_6567,N_4829,N_4967);
or U6568 (N_6568,N_4808,N_4718);
nor U6569 (N_6569,N_4691,N_2810);
nor U6570 (N_6570,N_4571,N_4713);
and U6571 (N_6571,N_4963,N_4224);
and U6572 (N_6572,N_4611,N_4082);
nand U6573 (N_6573,N_3554,N_4467);
or U6574 (N_6574,N_3899,N_2963);
xnor U6575 (N_6575,N_3784,N_3476);
nor U6576 (N_6576,N_2837,N_3505);
nand U6577 (N_6577,N_4770,N_3902);
nor U6578 (N_6578,N_4686,N_2610);
nand U6579 (N_6579,N_4251,N_3650);
nor U6580 (N_6580,N_4676,N_4913);
and U6581 (N_6581,N_2985,N_2698);
or U6582 (N_6582,N_3797,N_4147);
nand U6583 (N_6583,N_2674,N_3441);
and U6584 (N_6584,N_3284,N_2888);
and U6585 (N_6585,N_2675,N_4828);
and U6586 (N_6586,N_4866,N_2898);
xor U6587 (N_6587,N_4017,N_3855);
nand U6588 (N_6588,N_4121,N_4489);
nand U6589 (N_6589,N_3885,N_3968);
nand U6590 (N_6590,N_4327,N_2658);
or U6591 (N_6591,N_4918,N_3116);
or U6592 (N_6592,N_4192,N_3773);
xor U6593 (N_6593,N_4307,N_3027);
xor U6594 (N_6594,N_4779,N_3641);
xor U6595 (N_6595,N_3219,N_2552);
nand U6596 (N_6596,N_4563,N_3651);
xnor U6597 (N_6597,N_2566,N_4329);
and U6598 (N_6598,N_3215,N_2838);
and U6599 (N_6599,N_4616,N_4059);
xnor U6600 (N_6600,N_3612,N_2644);
nand U6601 (N_6601,N_2602,N_2527);
or U6602 (N_6602,N_3058,N_4554);
or U6603 (N_6603,N_2919,N_4185);
xor U6604 (N_6604,N_3580,N_4520);
nor U6605 (N_6605,N_4693,N_3098);
nor U6606 (N_6606,N_3222,N_4400);
nand U6607 (N_6607,N_2748,N_2669);
or U6608 (N_6608,N_3265,N_2800);
or U6609 (N_6609,N_2830,N_4788);
nand U6610 (N_6610,N_4984,N_3452);
nand U6611 (N_6611,N_2942,N_3406);
or U6612 (N_6612,N_3501,N_4782);
nand U6613 (N_6613,N_3720,N_2506);
and U6614 (N_6614,N_2894,N_3570);
nand U6615 (N_6615,N_4970,N_4608);
nor U6616 (N_6616,N_3832,N_4440);
nor U6617 (N_6617,N_3333,N_3403);
nand U6618 (N_6618,N_3162,N_3109);
nor U6619 (N_6619,N_4538,N_3716);
and U6620 (N_6620,N_3917,N_3278);
or U6621 (N_6621,N_3273,N_2815);
xor U6622 (N_6622,N_4416,N_4413);
and U6623 (N_6623,N_4941,N_3765);
nor U6624 (N_6624,N_4288,N_4339);
or U6625 (N_6625,N_4790,N_4231);
xnor U6626 (N_6626,N_4160,N_3970);
or U6627 (N_6627,N_3608,N_3164);
nor U6628 (N_6628,N_4406,N_3057);
xor U6629 (N_6629,N_2807,N_3132);
nor U6630 (N_6630,N_3952,N_4064);
xor U6631 (N_6631,N_3976,N_2676);
nand U6632 (N_6632,N_4092,N_2695);
or U6633 (N_6633,N_2868,N_3993);
nor U6634 (N_6634,N_2690,N_3122);
or U6635 (N_6635,N_2720,N_4363);
and U6636 (N_6636,N_3530,N_2904);
and U6637 (N_6637,N_3011,N_4303);
or U6638 (N_6638,N_4543,N_3682);
nor U6639 (N_6639,N_3690,N_3213);
nand U6640 (N_6640,N_3694,N_3844);
nand U6641 (N_6641,N_4781,N_4982);
nor U6642 (N_6642,N_3767,N_4012);
and U6643 (N_6643,N_3164,N_3236);
and U6644 (N_6644,N_4335,N_4356);
or U6645 (N_6645,N_3778,N_4886);
and U6646 (N_6646,N_4741,N_3295);
nor U6647 (N_6647,N_4566,N_3870);
nand U6648 (N_6648,N_2663,N_2741);
nor U6649 (N_6649,N_4541,N_4281);
nor U6650 (N_6650,N_3629,N_3347);
or U6651 (N_6651,N_3151,N_4761);
and U6652 (N_6652,N_3378,N_4865);
nand U6653 (N_6653,N_3270,N_4022);
nor U6654 (N_6654,N_4975,N_4406);
or U6655 (N_6655,N_4967,N_4114);
nor U6656 (N_6656,N_2904,N_2891);
and U6657 (N_6657,N_2709,N_3216);
nor U6658 (N_6658,N_2616,N_4012);
and U6659 (N_6659,N_4917,N_3499);
and U6660 (N_6660,N_3603,N_3884);
xnor U6661 (N_6661,N_3323,N_3748);
and U6662 (N_6662,N_3875,N_4576);
or U6663 (N_6663,N_4612,N_2545);
xor U6664 (N_6664,N_3629,N_2641);
xor U6665 (N_6665,N_3890,N_3035);
nor U6666 (N_6666,N_4550,N_2801);
nand U6667 (N_6667,N_4701,N_3227);
and U6668 (N_6668,N_4762,N_3739);
nand U6669 (N_6669,N_2644,N_3270);
or U6670 (N_6670,N_2703,N_4321);
xor U6671 (N_6671,N_3526,N_3258);
xnor U6672 (N_6672,N_4836,N_3498);
xnor U6673 (N_6673,N_4967,N_3955);
and U6674 (N_6674,N_4740,N_3573);
nor U6675 (N_6675,N_4677,N_3058);
xnor U6676 (N_6676,N_3398,N_3898);
xor U6677 (N_6677,N_2935,N_4816);
or U6678 (N_6678,N_3777,N_3448);
nand U6679 (N_6679,N_2525,N_2933);
or U6680 (N_6680,N_3197,N_4379);
nand U6681 (N_6681,N_4244,N_3139);
nand U6682 (N_6682,N_4295,N_2818);
xor U6683 (N_6683,N_3523,N_3555);
nor U6684 (N_6684,N_3680,N_4344);
nand U6685 (N_6685,N_4520,N_3354);
nand U6686 (N_6686,N_2839,N_2718);
or U6687 (N_6687,N_4774,N_4275);
xor U6688 (N_6688,N_2769,N_3771);
nand U6689 (N_6689,N_4497,N_3925);
nand U6690 (N_6690,N_3849,N_3327);
nand U6691 (N_6691,N_3977,N_4291);
nand U6692 (N_6692,N_4463,N_3377);
or U6693 (N_6693,N_2702,N_3779);
nor U6694 (N_6694,N_4335,N_3238);
xor U6695 (N_6695,N_3167,N_3822);
or U6696 (N_6696,N_4075,N_3937);
nor U6697 (N_6697,N_4723,N_3057);
xnor U6698 (N_6698,N_2588,N_3796);
and U6699 (N_6699,N_4421,N_3006);
xor U6700 (N_6700,N_3778,N_3133);
nand U6701 (N_6701,N_2880,N_3908);
or U6702 (N_6702,N_4594,N_3420);
nor U6703 (N_6703,N_3061,N_3638);
nand U6704 (N_6704,N_3909,N_4440);
nand U6705 (N_6705,N_4972,N_3164);
and U6706 (N_6706,N_4637,N_3827);
or U6707 (N_6707,N_4843,N_4571);
nand U6708 (N_6708,N_3702,N_3316);
nor U6709 (N_6709,N_4272,N_3269);
and U6710 (N_6710,N_4632,N_4643);
nor U6711 (N_6711,N_3738,N_2923);
xnor U6712 (N_6712,N_3204,N_4678);
and U6713 (N_6713,N_3770,N_4877);
and U6714 (N_6714,N_4065,N_2906);
or U6715 (N_6715,N_4051,N_4095);
nand U6716 (N_6716,N_3125,N_4326);
or U6717 (N_6717,N_3685,N_4247);
nand U6718 (N_6718,N_2674,N_3221);
nand U6719 (N_6719,N_3442,N_4609);
or U6720 (N_6720,N_4108,N_2797);
nand U6721 (N_6721,N_4166,N_4571);
or U6722 (N_6722,N_4949,N_4130);
and U6723 (N_6723,N_3033,N_3940);
nor U6724 (N_6724,N_2921,N_4313);
xnor U6725 (N_6725,N_2902,N_2783);
and U6726 (N_6726,N_3070,N_4254);
nor U6727 (N_6727,N_4552,N_4566);
nand U6728 (N_6728,N_4122,N_3859);
nand U6729 (N_6729,N_3212,N_3727);
and U6730 (N_6730,N_2889,N_3275);
and U6731 (N_6731,N_4067,N_4837);
or U6732 (N_6732,N_2678,N_4191);
nand U6733 (N_6733,N_3640,N_4733);
and U6734 (N_6734,N_2650,N_3080);
or U6735 (N_6735,N_2661,N_2592);
nand U6736 (N_6736,N_3593,N_4110);
xnor U6737 (N_6737,N_3275,N_3471);
nor U6738 (N_6738,N_3605,N_3504);
xnor U6739 (N_6739,N_4475,N_4810);
and U6740 (N_6740,N_3354,N_3619);
xnor U6741 (N_6741,N_3720,N_4104);
or U6742 (N_6742,N_3477,N_2625);
or U6743 (N_6743,N_2747,N_3032);
nand U6744 (N_6744,N_2774,N_2691);
xor U6745 (N_6745,N_4349,N_3707);
and U6746 (N_6746,N_3367,N_2755);
nand U6747 (N_6747,N_2548,N_2675);
or U6748 (N_6748,N_2500,N_4427);
and U6749 (N_6749,N_3557,N_4986);
nor U6750 (N_6750,N_2690,N_4886);
or U6751 (N_6751,N_3522,N_3145);
or U6752 (N_6752,N_4821,N_4807);
xor U6753 (N_6753,N_3905,N_4465);
or U6754 (N_6754,N_2738,N_2969);
nand U6755 (N_6755,N_2727,N_2678);
and U6756 (N_6756,N_4408,N_4279);
and U6757 (N_6757,N_3370,N_3227);
or U6758 (N_6758,N_3828,N_3115);
nand U6759 (N_6759,N_4051,N_3581);
nand U6760 (N_6760,N_2600,N_4138);
nor U6761 (N_6761,N_2923,N_3706);
xor U6762 (N_6762,N_2739,N_2571);
nand U6763 (N_6763,N_3840,N_3010);
nor U6764 (N_6764,N_3571,N_3186);
xor U6765 (N_6765,N_3000,N_3186);
and U6766 (N_6766,N_3323,N_4089);
or U6767 (N_6767,N_2992,N_2908);
nor U6768 (N_6768,N_4656,N_4488);
and U6769 (N_6769,N_4484,N_4490);
nand U6770 (N_6770,N_3065,N_3917);
nand U6771 (N_6771,N_3816,N_3025);
nor U6772 (N_6772,N_2966,N_3959);
or U6773 (N_6773,N_2544,N_4043);
nor U6774 (N_6774,N_4427,N_4210);
nor U6775 (N_6775,N_3821,N_4040);
xor U6776 (N_6776,N_2684,N_4063);
and U6777 (N_6777,N_3955,N_3245);
nor U6778 (N_6778,N_4248,N_3873);
nand U6779 (N_6779,N_2855,N_3430);
nor U6780 (N_6780,N_4636,N_4178);
or U6781 (N_6781,N_3190,N_3791);
xor U6782 (N_6782,N_2923,N_2869);
or U6783 (N_6783,N_3120,N_4313);
nor U6784 (N_6784,N_3238,N_4589);
and U6785 (N_6785,N_4702,N_3880);
xnor U6786 (N_6786,N_4757,N_4821);
nand U6787 (N_6787,N_3326,N_2974);
nand U6788 (N_6788,N_4265,N_2853);
and U6789 (N_6789,N_3572,N_2971);
nor U6790 (N_6790,N_3614,N_3282);
nand U6791 (N_6791,N_4266,N_4689);
and U6792 (N_6792,N_4059,N_4022);
and U6793 (N_6793,N_3987,N_3225);
or U6794 (N_6794,N_3562,N_3783);
xnor U6795 (N_6795,N_4815,N_4789);
and U6796 (N_6796,N_3737,N_3281);
and U6797 (N_6797,N_4272,N_2685);
xnor U6798 (N_6798,N_3793,N_3209);
nor U6799 (N_6799,N_4753,N_2738);
xnor U6800 (N_6800,N_3616,N_3622);
nor U6801 (N_6801,N_3802,N_3808);
nor U6802 (N_6802,N_4565,N_3939);
nand U6803 (N_6803,N_3225,N_3961);
and U6804 (N_6804,N_4504,N_2712);
and U6805 (N_6805,N_3602,N_4733);
or U6806 (N_6806,N_2660,N_4931);
nor U6807 (N_6807,N_4192,N_3688);
and U6808 (N_6808,N_3541,N_3496);
and U6809 (N_6809,N_3025,N_4730);
nand U6810 (N_6810,N_3358,N_4772);
nand U6811 (N_6811,N_2867,N_2845);
xnor U6812 (N_6812,N_4091,N_2623);
nand U6813 (N_6813,N_2515,N_2594);
or U6814 (N_6814,N_4327,N_3070);
nor U6815 (N_6815,N_4732,N_3422);
xor U6816 (N_6816,N_3236,N_4718);
xor U6817 (N_6817,N_2727,N_4551);
and U6818 (N_6818,N_3215,N_2881);
or U6819 (N_6819,N_4400,N_2545);
and U6820 (N_6820,N_4065,N_4265);
nor U6821 (N_6821,N_4898,N_4530);
or U6822 (N_6822,N_4958,N_3939);
nor U6823 (N_6823,N_3028,N_4064);
nor U6824 (N_6824,N_4293,N_3510);
xnor U6825 (N_6825,N_3567,N_4044);
and U6826 (N_6826,N_4132,N_3090);
xor U6827 (N_6827,N_4612,N_4244);
nor U6828 (N_6828,N_4377,N_4482);
nand U6829 (N_6829,N_4834,N_3317);
nand U6830 (N_6830,N_2513,N_2960);
or U6831 (N_6831,N_4020,N_3458);
nor U6832 (N_6832,N_3038,N_4231);
and U6833 (N_6833,N_2595,N_4362);
xnor U6834 (N_6834,N_3302,N_4946);
nand U6835 (N_6835,N_4357,N_3593);
or U6836 (N_6836,N_4696,N_2529);
nor U6837 (N_6837,N_4865,N_3553);
nand U6838 (N_6838,N_4761,N_2832);
nor U6839 (N_6839,N_2832,N_4922);
nor U6840 (N_6840,N_2762,N_3897);
nand U6841 (N_6841,N_4909,N_4772);
or U6842 (N_6842,N_4040,N_4823);
xnor U6843 (N_6843,N_3166,N_3740);
xor U6844 (N_6844,N_3324,N_3951);
nand U6845 (N_6845,N_3732,N_2654);
and U6846 (N_6846,N_3259,N_4745);
nor U6847 (N_6847,N_2774,N_3687);
nand U6848 (N_6848,N_4200,N_3873);
nor U6849 (N_6849,N_4427,N_4080);
nand U6850 (N_6850,N_2537,N_3917);
xnor U6851 (N_6851,N_3610,N_3131);
or U6852 (N_6852,N_3698,N_4292);
or U6853 (N_6853,N_3928,N_3011);
nand U6854 (N_6854,N_4317,N_3249);
xnor U6855 (N_6855,N_4028,N_4992);
and U6856 (N_6856,N_3659,N_4799);
xor U6857 (N_6857,N_3757,N_4545);
nor U6858 (N_6858,N_2620,N_2890);
xnor U6859 (N_6859,N_4338,N_2542);
or U6860 (N_6860,N_3881,N_4700);
or U6861 (N_6861,N_2645,N_4987);
or U6862 (N_6862,N_4633,N_2513);
nand U6863 (N_6863,N_3654,N_4479);
and U6864 (N_6864,N_3389,N_2739);
and U6865 (N_6865,N_4523,N_3944);
or U6866 (N_6866,N_4405,N_4005);
nand U6867 (N_6867,N_2537,N_3886);
nand U6868 (N_6868,N_3972,N_3250);
xor U6869 (N_6869,N_3540,N_4925);
and U6870 (N_6870,N_3805,N_3882);
nor U6871 (N_6871,N_3368,N_3034);
nand U6872 (N_6872,N_2818,N_4340);
nor U6873 (N_6873,N_4890,N_3292);
nand U6874 (N_6874,N_2534,N_3712);
xor U6875 (N_6875,N_3623,N_2867);
and U6876 (N_6876,N_4234,N_3244);
or U6877 (N_6877,N_4862,N_4861);
xor U6878 (N_6878,N_4926,N_2573);
and U6879 (N_6879,N_2979,N_4373);
and U6880 (N_6880,N_3815,N_4461);
or U6881 (N_6881,N_3683,N_3181);
nor U6882 (N_6882,N_3910,N_3000);
or U6883 (N_6883,N_4630,N_3127);
and U6884 (N_6884,N_3218,N_3297);
or U6885 (N_6885,N_4834,N_3469);
nand U6886 (N_6886,N_3015,N_4131);
nor U6887 (N_6887,N_4483,N_3573);
nand U6888 (N_6888,N_3639,N_3388);
nor U6889 (N_6889,N_4161,N_3550);
or U6890 (N_6890,N_4071,N_3986);
xor U6891 (N_6891,N_3758,N_3726);
and U6892 (N_6892,N_3903,N_3729);
or U6893 (N_6893,N_2689,N_3350);
and U6894 (N_6894,N_4325,N_3533);
xor U6895 (N_6895,N_4106,N_4933);
nor U6896 (N_6896,N_3238,N_4912);
nand U6897 (N_6897,N_3759,N_4595);
nand U6898 (N_6898,N_3794,N_2772);
xor U6899 (N_6899,N_2769,N_4349);
nand U6900 (N_6900,N_4478,N_4096);
or U6901 (N_6901,N_3319,N_4621);
nor U6902 (N_6902,N_2606,N_4619);
xnor U6903 (N_6903,N_4829,N_2860);
xor U6904 (N_6904,N_3518,N_4546);
or U6905 (N_6905,N_3124,N_2700);
nand U6906 (N_6906,N_4442,N_3743);
nand U6907 (N_6907,N_2789,N_4814);
nor U6908 (N_6908,N_2802,N_2830);
or U6909 (N_6909,N_4931,N_4246);
or U6910 (N_6910,N_2784,N_4415);
xor U6911 (N_6911,N_4330,N_4264);
nand U6912 (N_6912,N_4885,N_2559);
or U6913 (N_6913,N_3993,N_2678);
or U6914 (N_6914,N_3389,N_3148);
and U6915 (N_6915,N_3140,N_3655);
xor U6916 (N_6916,N_2832,N_3531);
and U6917 (N_6917,N_4179,N_3107);
xnor U6918 (N_6918,N_2979,N_4512);
and U6919 (N_6919,N_3395,N_2599);
nor U6920 (N_6920,N_3938,N_4013);
xor U6921 (N_6921,N_2902,N_4259);
nand U6922 (N_6922,N_2503,N_3747);
xor U6923 (N_6923,N_4806,N_4829);
and U6924 (N_6924,N_3354,N_4232);
and U6925 (N_6925,N_4431,N_3160);
nor U6926 (N_6926,N_4882,N_4966);
nand U6927 (N_6927,N_3376,N_4830);
nor U6928 (N_6928,N_3862,N_4332);
nand U6929 (N_6929,N_3479,N_4660);
nor U6930 (N_6930,N_4558,N_4853);
and U6931 (N_6931,N_3417,N_2907);
and U6932 (N_6932,N_4895,N_4473);
nand U6933 (N_6933,N_3971,N_4809);
or U6934 (N_6934,N_2975,N_3484);
nand U6935 (N_6935,N_2705,N_3751);
xor U6936 (N_6936,N_2823,N_3806);
xnor U6937 (N_6937,N_3753,N_4366);
xnor U6938 (N_6938,N_2752,N_3262);
xor U6939 (N_6939,N_4298,N_4981);
nand U6940 (N_6940,N_3002,N_3975);
and U6941 (N_6941,N_3289,N_4738);
nor U6942 (N_6942,N_3280,N_2841);
nand U6943 (N_6943,N_4271,N_3342);
and U6944 (N_6944,N_2539,N_2533);
nor U6945 (N_6945,N_4819,N_2555);
nand U6946 (N_6946,N_3824,N_3136);
nand U6947 (N_6947,N_3093,N_3643);
nor U6948 (N_6948,N_2751,N_4323);
or U6949 (N_6949,N_3761,N_4886);
nand U6950 (N_6950,N_4492,N_2973);
nor U6951 (N_6951,N_4152,N_4112);
and U6952 (N_6952,N_4085,N_2545);
nand U6953 (N_6953,N_3418,N_4572);
or U6954 (N_6954,N_3130,N_3821);
nand U6955 (N_6955,N_2745,N_2998);
nand U6956 (N_6956,N_4328,N_3783);
xnor U6957 (N_6957,N_4458,N_3958);
nor U6958 (N_6958,N_3775,N_2888);
nand U6959 (N_6959,N_3723,N_2852);
and U6960 (N_6960,N_3472,N_3766);
and U6961 (N_6961,N_3219,N_3906);
xnor U6962 (N_6962,N_2882,N_3178);
nand U6963 (N_6963,N_3971,N_4921);
xor U6964 (N_6964,N_3659,N_2509);
nor U6965 (N_6965,N_4119,N_3264);
xnor U6966 (N_6966,N_3404,N_4147);
nand U6967 (N_6967,N_4538,N_4370);
or U6968 (N_6968,N_3030,N_2909);
or U6969 (N_6969,N_2993,N_3839);
and U6970 (N_6970,N_3621,N_3646);
xnor U6971 (N_6971,N_4568,N_4861);
or U6972 (N_6972,N_2681,N_3380);
xnor U6973 (N_6973,N_3131,N_4683);
and U6974 (N_6974,N_4577,N_4372);
or U6975 (N_6975,N_3968,N_2695);
xnor U6976 (N_6976,N_4122,N_4906);
and U6977 (N_6977,N_2508,N_3990);
nor U6978 (N_6978,N_2788,N_4478);
or U6979 (N_6979,N_3823,N_4773);
and U6980 (N_6980,N_4620,N_3073);
nor U6981 (N_6981,N_3729,N_4270);
or U6982 (N_6982,N_4696,N_3929);
nor U6983 (N_6983,N_4475,N_2574);
nor U6984 (N_6984,N_2703,N_3656);
nor U6985 (N_6985,N_3764,N_3079);
nand U6986 (N_6986,N_2953,N_2515);
xor U6987 (N_6987,N_4032,N_3876);
nor U6988 (N_6988,N_3731,N_2880);
or U6989 (N_6989,N_3975,N_2663);
and U6990 (N_6990,N_2952,N_4175);
or U6991 (N_6991,N_2893,N_3590);
nand U6992 (N_6992,N_2889,N_2879);
xor U6993 (N_6993,N_3285,N_2837);
nand U6994 (N_6994,N_3101,N_3282);
nor U6995 (N_6995,N_4026,N_4418);
or U6996 (N_6996,N_4583,N_3704);
or U6997 (N_6997,N_4843,N_4583);
nand U6998 (N_6998,N_2724,N_2509);
or U6999 (N_6999,N_3272,N_3862);
xor U7000 (N_7000,N_4147,N_2843);
nor U7001 (N_7001,N_3918,N_4000);
xnor U7002 (N_7002,N_3677,N_3722);
nand U7003 (N_7003,N_3775,N_4192);
xnor U7004 (N_7004,N_4431,N_3826);
xor U7005 (N_7005,N_3334,N_2781);
or U7006 (N_7006,N_3284,N_3796);
xor U7007 (N_7007,N_3037,N_4233);
nand U7008 (N_7008,N_2936,N_3602);
nor U7009 (N_7009,N_2551,N_4629);
xor U7010 (N_7010,N_2931,N_4442);
and U7011 (N_7011,N_3393,N_2848);
or U7012 (N_7012,N_4135,N_4775);
nor U7013 (N_7013,N_4080,N_4708);
or U7014 (N_7014,N_3675,N_4917);
nor U7015 (N_7015,N_4933,N_2653);
and U7016 (N_7016,N_4472,N_3682);
and U7017 (N_7017,N_4186,N_3885);
xnor U7018 (N_7018,N_2565,N_3110);
or U7019 (N_7019,N_2500,N_2997);
or U7020 (N_7020,N_2962,N_3902);
nor U7021 (N_7021,N_4972,N_3302);
nor U7022 (N_7022,N_3828,N_3610);
xnor U7023 (N_7023,N_4406,N_3171);
or U7024 (N_7024,N_4739,N_2815);
and U7025 (N_7025,N_3636,N_4419);
nor U7026 (N_7026,N_4264,N_4909);
nand U7027 (N_7027,N_4256,N_4575);
and U7028 (N_7028,N_3704,N_3952);
or U7029 (N_7029,N_3156,N_3155);
or U7030 (N_7030,N_4112,N_3745);
and U7031 (N_7031,N_3095,N_3293);
and U7032 (N_7032,N_2717,N_4188);
and U7033 (N_7033,N_2604,N_4802);
and U7034 (N_7034,N_4821,N_4690);
nor U7035 (N_7035,N_3008,N_4399);
xnor U7036 (N_7036,N_3957,N_3443);
nand U7037 (N_7037,N_4558,N_3767);
nor U7038 (N_7038,N_4954,N_4314);
nor U7039 (N_7039,N_3563,N_4607);
nor U7040 (N_7040,N_2765,N_4907);
nor U7041 (N_7041,N_3475,N_4127);
and U7042 (N_7042,N_2805,N_3438);
nand U7043 (N_7043,N_3640,N_2909);
or U7044 (N_7044,N_3255,N_4863);
nor U7045 (N_7045,N_4469,N_3666);
nand U7046 (N_7046,N_3877,N_2727);
or U7047 (N_7047,N_3757,N_4191);
nand U7048 (N_7048,N_2587,N_2545);
nand U7049 (N_7049,N_4617,N_3600);
xnor U7050 (N_7050,N_4698,N_4913);
nor U7051 (N_7051,N_3973,N_4872);
nor U7052 (N_7052,N_4380,N_3175);
xor U7053 (N_7053,N_4538,N_4462);
nor U7054 (N_7054,N_4584,N_3227);
nor U7055 (N_7055,N_3599,N_3087);
nor U7056 (N_7056,N_3657,N_3876);
and U7057 (N_7057,N_2932,N_4287);
or U7058 (N_7058,N_3344,N_4914);
or U7059 (N_7059,N_3531,N_2940);
nand U7060 (N_7060,N_3491,N_4910);
xnor U7061 (N_7061,N_3705,N_3012);
xnor U7062 (N_7062,N_4324,N_2918);
nand U7063 (N_7063,N_2629,N_3608);
nor U7064 (N_7064,N_3282,N_2738);
nor U7065 (N_7065,N_2731,N_2606);
and U7066 (N_7066,N_4276,N_2772);
xnor U7067 (N_7067,N_3153,N_4614);
and U7068 (N_7068,N_2613,N_3740);
xnor U7069 (N_7069,N_3344,N_4637);
and U7070 (N_7070,N_4818,N_4961);
nor U7071 (N_7071,N_4141,N_3219);
and U7072 (N_7072,N_4760,N_3180);
and U7073 (N_7073,N_4164,N_3123);
nor U7074 (N_7074,N_2941,N_3462);
nand U7075 (N_7075,N_2999,N_2585);
or U7076 (N_7076,N_3909,N_2635);
nor U7077 (N_7077,N_3609,N_3200);
xor U7078 (N_7078,N_3464,N_3251);
and U7079 (N_7079,N_3217,N_3189);
nor U7080 (N_7080,N_4822,N_4167);
or U7081 (N_7081,N_4470,N_4563);
nor U7082 (N_7082,N_4774,N_4650);
and U7083 (N_7083,N_3277,N_4375);
xor U7084 (N_7084,N_2726,N_3201);
xor U7085 (N_7085,N_4121,N_4907);
or U7086 (N_7086,N_3332,N_3277);
nand U7087 (N_7087,N_4884,N_4659);
and U7088 (N_7088,N_3320,N_2788);
xor U7089 (N_7089,N_2719,N_4253);
nor U7090 (N_7090,N_3377,N_3218);
or U7091 (N_7091,N_3403,N_3004);
xnor U7092 (N_7092,N_2850,N_3262);
xor U7093 (N_7093,N_4982,N_4408);
xor U7094 (N_7094,N_3335,N_2537);
nand U7095 (N_7095,N_2741,N_3561);
and U7096 (N_7096,N_4477,N_3956);
and U7097 (N_7097,N_4616,N_4742);
nor U7098 (N_7098,N_3316,N_2666);
nand U7099 (N_7099,N_4159,N_3990);
xnor U7100 (N_7100,N_4947,N_3010);
xor U7101 (N_7101,N_3939,N_4539);
and U7102 (N_7102,N_3334,N_4717);
nor U7103 (N_7103,N_4911,N_4205);
xor U7104 (N_7104,N_2901,N_4526);
xnor U7105 (N_7105,N_3621,N_4059);
nor U7106 (N_7106,N_4193,N_4832);
nor U7107 (N_7107,N_4897,N_3306);
nand U7108 (N_7108,N_4669,N_4295);
or U7109 (N_7109,N_4634,N_2689);
nor U7110 (N_7110,N_3377,N_3926);
xnor U7111 (N_7111,N_4619,N_3297);
xnor U7112 (N_7112,N_4776,N_3663);
or U7113 (N_7113,N_3636,N_4630);
nor U7114 (N_7114,N_4536,N_3539);
nand U7115 (N_7115,N_3746,N_3889);
and U7116 (N_7116,N_3811,N_4182);
xnor U7117 (N_7117,N_3923,N_3231);
nor U7118 (N_7118,N_4126,N_4409);
and U7119 (N_7119,N_3669,N_4532);
xnor U7120 (N_7120,N_3944,N_4243);
and U7121 (N_7121,N_2544,N_3775);
nor U7122 (N_7122,N_4784,N_3059);
nor U7123 (N_7123,N_4701,N_4519);
xor U7124 (N_7124,N_4286,N_3409);
xnor U7125 (N_7125,N_2741,N_2896);
nor U7126 (N_7126,N_4606,N_3880);
xnor U7127 (N_7127,N_2851,N_3333);
or U7128 (N_7128,N_3672,N_4022);
xor U7129 (N_7129,N_4856,N_4574);
xnor U7130 (N_7130,N_3871,N_4778);
or U7131 (N_7131,N_4546,N_4617);
nor U7132 (N_7132,N_4176,N_3156);
or U7133 (N_7133,N_3807,N_4201);
and U7134 (N_7134,N_3272,N_3163);
and U7135 (N_7135,N_2763,N_4949);
xor U7136 (N_7136,N_4373,N_3880);
or U7137 (N_7137,N_3864,N_4834);
nor U7138 (N_7138,N_2776,N_4153);
nand U7139 (N_7139,N_4694,N_3517);
nand U7140 (N_7140,N_2820,N_2611);
nor U7141 (N_7141,N_3379,N_4824);
or U7142 (N_7142,N_2931,N_3375);
or U7143 (N_7143,N_4096,N_3613);
nor U7144 (N_7144,N_4900,N_3612);
nand U7145 (N_7145,N_4497,N_3763);
nand U7146 (N_7146,N_4504,N_4073);
nor U7147 (N_7147,N_4572,N_2619);
and U7148 (N_7148,N_4067,N_2788);
or U7149 (N_7149,N_3380,N_4462);
xor U7150 (N_7150,N_3138,N_4482);
or U7151 (N_7151,N_4017,N_3605);
and U7152 (N_7152,N_4583,N_4947);
and U7153 (N_7153,N_2752,N_2971);
nor U7154 (N_7154,N_4684,N_4297);
xor U7155 (N_7155,N_4322,N_2875);
xnor U7156 (N_7156,N_3071,N_4598);
nand U7157 (N_7157,N_4947,N_2566);
or U7158 (N_7158,N_3483,N_4738);
xor U7159 (N_7159,N_3329,N_3185);
and U7160 (N_7160,N_4004,N_4755);
and U7161 (N_7161,N_3145,N_4732);
or U7162 (N_7162,N_4557,N_3330);
nor U7163 (N_7163,N_3412,N_4728);
nor U7164 (N_7164,N_2628,N_4379);
and U7165 (N_7165,N_4653,N_4145);
and U7166 (N_7166,N_4240,N_4704);
or U7167 (N_7167,N_4453,N_3383);
nor U7168 (N_7168,N_2938,N_4983);
and U7169 (N_7169,N_4354,N_3418);
xnor U7170 (N_7170,N_4487,N_3295);
and U7171 (N_7171,N_3328,N_3141);
or U7172 (N_7172,N_3873,N_4526);
xor U7173 (N_7173,N_3055,N_3772);
or U7174 (N_7174,N_2546,N_4184);
nand U7175 (N_7175,N_3978,N_2847);
nor U7176 (N_7176,N_4284,N_3800);
nand U7177 (N_7177,N_3180,N_2934);
nand U7178 (N_7178,N_3944,N_3748);
xor U7179 (N_7179,N_3189,N_4446);
and U7180 (N_7180,N_4877,N_4732);
xor U7181 (N_7181,N_4443,N_4617);
or U7182 (N_7182,N_2614,N_3753);
nand U7183 (N_7183,N_4515,N_3209);
or U7184 (N_7184,N_4525,N_4937);
nor U7185 (N_7185,N_3838,N_2883);
nor U7186 (N_7186,N_3026,N_3632);
nand U7187 (N_7187,N_2689,N_3726);
nand U7188 (N_7188,N_4047,N_2766);
xnor U7189 (N_7189,N_3888,N_2848);
nand U7190 (N_7190,N_4406,N_3625);
or U7191 (N_7191,N_3935,N_4650);
and U7192 (N_7192,N_4915,N_4562);
nand U7193 (N_7193,N_2874,N_3268);
and U7194 (N_7194,N_3660,N_3231);
nand U7195 (N_7195,N_3024,N_2593);
nor U7196 (N_7196,N_2817,N_4812);
nor U7197 (N_7197,N_3963,N_4391);
xnor U7198 (N_7198,N_4170,N_4978);
or U7199 (N_7199,N_2643,N_4409);
and U7200 (N_7200,N_3991,N_4450);
or U7201 (N_7201,N_4835,N_3478);
xnor U7202 (N_7202,N_4384,N_4295);
xnor U7203 (N_7203,N_4105,N_2767);
nor U7204 (N_7204,N_3829,N_4094);
or U7205 (N_7205,N_4953,N_3420);
nand U7206 (N_7206,N_3171,N_3798);
and U7207 (N_7207,N_3581,N_4258);
or U7208 (N_7208,N_2829,N_4986);
nor U7209 (N_7209,N_4158,N_2824);
nor U7210 (N_7210,N_4697,N_4299);
or U7211 (N_7211,N_4822,N_4667);
xnor U7212 (N_7212,N_3790,N_4351);
xor U7213 (N_7213,N_2759,N_4123);
and U7214 (N_7214,N_3698,N_3856);
xnor U7215 (N_7215,N_3533,N_3928);
nor U7216 (N_7216,N_4756,N_2809);
or U7217 (N_7217,N_4030,N_2903);
xnor U7218 (N_7218,N_3417,N_4624);
and U7219 (N_7219,N_3703,N_3020);
or U7220 (N_7220,N_4961,N_4599);
nor U7221 (N_7221,N_3564,N_4584);
and U7222 (N_7222,N_2621,N_4806);
or U7223 (N_7223,N_3514,N_4963);
xor U7224 (N_7224,N_3525,N_3448);
nand U7225 (N_7225,N_4074,N_2742);
or U7226 (N_7226,N_3510,N_4884);
or U7227 (N_7227,N_3479,N_4161);
nor U7228 (N_7228,N_2651,N_2833);
nor U7229 (N_7229,N_4672,N_3737);
nor U7230 (N_7230,N_2759,N_2817);
xor U7231 (N_7231,N_3744,N_4544);
nand U7232 (N_7232,N_4606,N_3612);
xnor U7233 (N_7233,N_3830,N_3466);
and U7234 (N_7234,N_4160,N_3918);
nor U7235 (N_7235,N_3732,N_2791);
nand U7236 (N_7236,N_4956,N_3625);
nor U7237 (N_7237,N_2623,N_2697);
nand U7238 (N_7238,N_4929,N_4316);
or U7239 (N_7239,N_4933,N_3366);
or U7240 (N_7240,N_3716,N_3428);
or U7241 (N_7241,N_2788,N_3383);
xnor U7242 (N_7242,N_3882,N_3976);
nand U7243 (N_7243,N_4682,N_2974);
or U7244 (N_7244,N_4832,N_4323);
or U7245 (N_7245,N_3924,N_3224);
xor U7246 (N_7246,N_4134,N_3588);
nand U7247 (N_7247,N_2502,N_3110);
and U7248 (N_7248,N_4643,N_3053);
nor U7249 (N_7249,N_3329,N_3766);
xnor U7250 (N_7250,N_2870,N_3124);
xor U7251 (N_7251,N_2553,N_3699);
xor U7252 (N_7252,N_3496,N_3037);
or U7253 (N_7253,N_3479,N_3156);
nand U7254 (N_7254,N_2853,N_3141);
nor U7255 (N_7255,N_4966,N_4689);
nor U7256 (N_7256,N_4109,N_4792);
xnor U7257 (N_7257,N_4465,N_4522);
xor U7258 (N_7258,N_3150,N_3047);
and U7259 (N_7259,N_4331,N_2633);
nor U7260 (N_7260,N_2619,N_2816);
or U7261 (N_7261,N_3392,N_4642);
nor U7262 (N_7262,N_2966,N_3217);
nand U7263 (N_7263,N_4653,N_3818);
xnor U7264 (N_7264,N_3507,N_4061);
xor U7265 (N_7265,N_2931,N_4465);
nand U7266 (N_7266,N_3089,N_4672);
nand U7267 (N_7267,N_2513,N_4586);
and U7268 (N_7268,N_3451,N_4177);
xnor U7269 (N_7269,N_3919,N_3257);
and U7270 (N_7270,N_2796,N_2557);
or U7271 (N_7271,N_3410,N_3204);
xor U7272 (N_7272,N_4164,N_4409);
xor U7273 (N_7273,N_3116,N_4865);
and U7274 (N_7274,N_4979,N_4243);
nand U7275 (N_7275,N_4283,N_2799);
xnor U7276 (N_7276,N_2558,N_3402);
and U7277 (N_7277,N_4771,N_4055);
or U7278 (N_7278,N_4554,N_3236);
or U7279 (N_7279,N_4541,N_3828);
and U7280 (N_7280,N_3760,N_2889);
nand U7281 (N_7281,N_3986,N_3569);
or U7282 (N_7282,N_4281,N_2761);
nor U7283 (N_7283,N_3903,N_3437);
and U7284 (N_7284,N_3841,N_3856);
xor U7285 (N_7285,N_3055,N_3926);
or U7286 (N_7286,N_4837,N_3673);
or U7287 (N_7287,N_3491,N_4741);
and U7288 (N_7288,N_4174,N_3315);
or U7289 (N_7289,N_4958,N_4508);
and U7290 (N_7290,N_3364,N_2738);
nand U7291 (N_7291,N_3763,N_3987);
xnor U7292 (N_7292,N_3948,N_4301);
and U7293 (N_7293,N_2667,N_3647);
nand U7294 (N_7294,N_4366,N_4683);
nor U7295 (N_7295,N_4191,N_4730);
nor U7296 (N_7296,N_3916,N_4128);
and U7297 (N_7297,N_4354,N_3519);
and U7298 (N_7298,N_2985,N_3201);
and U7299 (N_7299,N_3514,N_4945);
or U7300 (N_7300,N_3957,N_4092);
or U7301 (N_7301,N_3893,N_4667);
nand U7302 (N_7302,N_4427,N_3069);
nand U7303 (N_7303,N_4827,N_4373);
or U7304 (N_7304,N_3684,N_3141);
and U7305 (N_7305,N_4217,N_4529);
xnor U7306 (N_7306,N_2786,N_2634);
xor U7307 (N_7307,N_4533,N_2960);
and U7308 (N_7308,N_3368,N_4771);
and U7309 (N_7309,N_2747,N_3325);
and U7310 (N_7310,N_4238,N_2977);
nand U7311 (N_7311,N_3923,N_3152);
or U7312 (N_7312,N_4493,N_4285);
and U7313 (N_7313,N_3070,N_3483);
nand U7314 (N_7314,N_3591,N_3636);
and U7315 (N_7315,N_4481,N_2918);
xor U7316 (N_7316,N_3092,N_4958);
and U7317 (N_7317,N_3099,N_2674);
xnor U7318 (N_7318,N_4195,N_4346);
nor U7319 (N_7319,N_4219,N_4593);
nor U7320 (N_7320,N_3489,N_3728);
or U7321 (N_7321,N_4086,N_4771);
or U7322 (N_7322,N_2786,N_2665);
nor U7323 (N_7323,N_3142,N_3555);
or U7324 (N_7324,N_2942,N_4854);
nand U7325 (N_7325,N_3666,N_2674);
or U7326 (N_7326,N_4372,N_4898);
xor U7327 (N_7327,N_3259,N_3995);
nand U7328 (N_7328,N_3329,N_4303);
xnor U7329 (N_7329,N_4661,N_3085);
and U7330 (N_7330,N_3807,N_4283);
nor U7331 (N_7331,N_4905,N_4972);
and U7332 (N_7332,N_4520,N_4528);
nor U7333 (N_7333,N_4373,N_2719);
nand U7334 (N_7334,N_3734,N_2703);
nor U7335 (N_7335,N_3267,N_2537);
xor U7336 (N_7336,N_4017,N_4754);
nand U7337 (N_7337,N_2753,N_3287);
nor U7338 (N_7338,N_2924,N_3960);
and U7339 (N_7339,N_2856,N_4946);
nor U7340 (N_7340,N_2676,N_3790);
and U7341 (N_7341,N_2865,N_2989);
nand U7342 (N_7342,N_3331,N_3728);
nand U7343 (N_7343,N_2801,N_2574);
or U7344 (N_7344,N_2617,N_3833);
nand U7345 (N_7345,N_3485,N_3069);
xnor U7346 (N_7346,N_4450,N_4894);
xor U7347 (N_7347,N_2568,N_4172);
nand U7348 (N_7348,N_3513,N_4634);
and U7349 (N_7349,N_4905,N_3902);
nand U7350 (N_7350,N_2739,N_3974);
nor U7351 (N_7351,N_4587,N_3247);
and U7352 (N_7352,N_4226,N_3948);
and U7353 (N_7353,N_4068,N_2670);
nand U7354 (N_7354,N_4652,N_2743);
and U7355 (N_7355,N_4025,N_4290);
nor U7356 (N_7356,N_4640,N_3157);
nand U7357 (N_7357,N_2982,N_3238);
xor U7358 (N_7358,N_2991,N_4430);
xor U7359 (N_7359,N_3353,N_4981);
and U7360 (N_7360,N_2585,N_2727);
nor U7361 (N_7361,N_3529,N_2615);
and U7362 (N_7362,N_4332,N_3453);
nand U7363 (N_7363,N_4607,N_3390);
nand U7364 (N_7364,N_4539,N_3572);
nand U7365 (N_7365,N_2967,N_2532);
xor U7366 (N_7366,N_2657,N_4727);
and U7367 (N_7367,N_4499,N_2922);
nor U7368 (N_7368,N_3026,N_4219);
nor U7369 (N_7369,N_2601,N_2639);
nand U7370 (N_7370,N_3386,N_3813);
nor U7371 (N_7371,N_4500,N_4245);
and U7372 (N_7372,N_4803,N_4786);
nor U7373 (N_7373,N_2851,N_4813);
nor U7374 (N_7374,N_2708,N_3113);
nand U7375 (N_7375,N_4810,N_3650);
xnor U7376 (N_7376,N_2522,N_4691);
or U7377 (N_7377,N_4639,N_3081);
and U7378 (N_7378,N_2610,N_3675);
xor U7379 (N_7379,N_3960,N_3433);
nand U7380 (N_7380,N_4049,N_3037);
or U7381 (N_7381,N_3585,N_3672);
or U7382 (N_7382,N_3431,N_3620);
xor U7383 (N_7383,N_4121,N_3038);
or U7384 (N_7384,N_2870,N_3612);
nand U7385 (N_7385,N_3837,N_4850);
nand U7386 (N_7386,N_4553,N_2701);
xnor U7387 (N_7387,N_3741,N_4691);
or U7388 (N_7388,N_3506,N_2626);
xnor U7389 (N_7389,N_3214,N_4550);
and U7390 (N_7390,N_2848,N_4793);
nor U7391 (N_7391,N_3181,N_3764);
and U7392 (N_7392,N_3381,N_2672);
nor U7393 (N_7393,N_4598,N_2800);
nand U7394 (N_7394,N_2633,N_2528);
nand U7395 (N_7395,N_2946,N_4251);
nor U7396 (N_7396,N_4858,N_3553);
nor U7397 (N_7397,N_4560,N_4476);
nand U7398 (N_7398,N_3685,N_4037);
or U7399 (N_7399,N_4192,N_3361);
and U7400 (N_7400,N_3753,N_2816);
nand U7401 (N_7401,N_2916,N_3038);
xnor U7402 (N_7402,N_2669,N_4170);
xnor U7403 (N_7403,N_3283,N_2799);
nand U7404 (N_7404,N_2551,N_4447);
nor U7405 (N_7405,N_3817,N_3025);
xnor U7406 (N_7406,N_3805,N_3038);
nand U7407 (N_7407,N_4091,N_3957);
or U7408 (N_7408,N_4533,N_3812);
nand U7409 (N_7409,N_3428,N_2847);
nor U7410 (N_7410,N_3124,N_3899);
or U7411 (N_7411,N_4877,N_4045);
xor U7412 (N_7412,N_3311,N_4037);
nor U7413 (N_7413,N_2604,N_2819);
and U7414 (N_7414,N_3086,N_3112);
nand U7415 (N_7415,N_2685,N_3515);
or U7416 (N_7416,N_4267,N_3997);
and U7417 (N_7417,N_4988,N_3755);
nand U7418 (N_7418,N_4236,N_3845);
nor U7419 (N_7419,N_4183,N_3968);
nor U7420 (N_7420,N_2836,N_3965);
or U7421 (N_7421,N_4872,N_4639);
or U7422 (N_7422,N_4829,N_4358);
nor U7423 (N_7423,N_3067,N_4170);
nand U7424 (N_7424,N_4570,N_2560);
nor U7425 (N_7425,N_2816,N_4369);
nor U7426 (N_7426,N_4481,N_3264);
xor U7427 (N_7427,N_4269,N_3239);
and U7428 (N_7428,N_4699,N_4004);
and U7429 (N_7429,N_4485,N_4026);
nand U7430 (N_7430,N_4639,N_2650);
xor U7431 (N_7431,N_4050,N_3145);
or U7432 (N_7432,N_4775,N_4633);
or U7433 (N_7433,N_4063,N_4718);
nand U7434 (N_7434,N_3473,N_4432);
xor U7435 (N_7435,N_2608,N_3494);
nor U7436 (N_7436,N_3870,N_4927);
nand U7437 (N_7437,N_4869,N_4191);
and U7438 (N_7438,N_2791,N_3443);
or U7439 (N_7439,N_2857,N_3649);
or U7440 (N_7440,N_3253,N_4127);
nand U7441 (N_7441,N_3492,N_3521);
and U7442 (N_7442,N_4121,N_3598);
nor U7443 (N_7443,N_2738,N_2915);
and U7444 (N_7444,N_4031,N_3945);
or U7445 (N_7445,N_4439,N_3530);
nor U7446 (N_7446,N_2730,N_4444);
or U7447 (N_7447,N_3779,N_4177);
or U7448 (N_7448,N_3994,N_3408);
and U7449 (N_7449,N_4267,N_4008);
or U7450 (N_7450,N_3031,N_4627);
and U7451 (N_7451,N_4688,N_3943);
or U7452 (N_7452,N_4330,N_3533);
nand U7453 (N_7453,N_4803,N_3818);
nor U7454 (N_7454,N_4664,N_4592);
xor U7455 (N_7455,N_3045,N_4947);
and U7456 (N_7456,N_4809,N_2786);
nand U7457 (N_7457,N_3307,N_3381);
or U7458 (N_7458,N_4931,N_3003);
nand U7459 (N_7459,N_3690,N_4960);
xor U7460 (N_7460,N_4264,N_4441);
nand U7461 (N_7461,N_4467,N_3944);
or U7462 (N_7462,N_3434,N_4909);
or U7463 (N_7463,N_2544,N_2623);
xor U7464 (N_7464,N_3468,N_3121);
nor U7465 (N_7465,N_3091,N_2716);
and U7466 (N_7466,N_3507,N_2598);
xnor U7467 (N_7467,N_4378,N_4565);
nor U7468 (N_7468,N_2693,N_3790);
xnor U7469 (N_7469,N_3751,N_3898);
or U7470 (N_7470,N_4211,N_3154);
and U7471 (N_7471,N_4543,N_2774);
or U7472 (N_7472,N_4654,N_4005);
xor U7473 (N_7473,N_3319,N_4057);
and U7474 (N_7474,N_4089,N_3558);
xor U7475 (N_7475,N_3926,N_4165);
nand U7476 (N_7476,N_3156,N_2788);
nand U7477 (N_7477,N_4513,N_4627);
xnor U7478 (N_7478,N_3738,N_3989);
xnor U7479 (N_7479,N_4962,N_2848);
or U7480 (N_7480,N_3280,N_2637);
or U7481 (N_7481,N_4616,N_3019);
nor U7482 (N_7482,N_3330,N_4997);
nor U7483 (N_7483,N_3472,N_3204);
nand U7484 (N_7484,N_3546,N_4080);
and U7485 (N_7485,N_4510,N_4619);
or U7486 (N_7486,N_4784,N_2562);
or U7487 (N_7487,N_4322,N_4541);
nand U7488 (N_7488,N_3334,N_4382);
or U7489 (N_7489,N_3485,N_3800);
or U7490 (N_7490,N_3661,N_3352);
or U7491 (N_7491,N_3140,N_3562);
nand U7492 (N_7492,N_4778,N_3893);
xor U7493 (N_7493,N_2613,N_4026);
or U7494 (N_7494,N_3750,N_4144);
nand U7495 (N_7495,N_2639,N_4101);
nand U7496 (N_7496,N_4901,N_2514);
or U7497 (N_7497,N_4602,N_3999);
or U7498 (N_7498,N_3081,N_3076);
nand U7499 (N_7499,N_4378,N_3251);
nand U7500 (N_7500,N_5290,N_5088);
nor U7501 (N_7501,N_5607,N_6249);
nand U7502 (N_7502,N_7498,N_5740);
nor U7503 (N_7503,N_5315,N_5303);
nand U7504 (N_7504,N_5648,N_6848);
or U7505 (N_7505,N_5757,N_6806);
nor U7506 (N_7506,N_6817,N_5808);
or U7507 (N_7507,N_6576,N_7054);
nand U7508 (N_7508,N_5117,N_6719);
xor U7509 (N_7509,N_7124,N_5908);
and U7510 (N_7510,N_5034,N_6155);
or U7511 (N_7511,N_6051,N_5547);
nor U7512 (N_7512,N_6346,N_6513);
nor U7513 (N_7513,N_5817,N_5717);
and U7514 (N_7514,N_6298,N_5924);
nor U7515 (N_7515,N_6220,N_5076);
xor U7516 (N_7516,N_6038,N_7094);
nor U7517 (N_7517,N_6594,N_7000);
and U7518 (N_7518,N_7217,N_7493);
xor U7519 (N_7519,N_5268,N_5353);
xnor U7520 (N_7520,N_5244,N_5651);
nand U7521 (N_7521,N_5780,N_6482);
nand U7522 (N_7522,N_5529,N_5251);
xor U7523 (N_7523,N_5868,N_7421);
nand U7524 (N_7524,N_6952,N_7106);
or U7525 (N_7525,N_6066,N_6050);
nand U7526 (N_7526,N_7197,N_6932);
nor U7527 (N_7527,N_7039,N_5447);
nand U7528 (N_7528,N_5048,N_6545);
nand U7529 (N_7529,N_6232,N_6444);
and U7530 (N_7530,N_6418,N_6660);
nand U7531 (N_7531,N_5845,N_6803);
and U7532 (N_7532,N_6948,N_7093);
or U7533 (N_7533,N_6369,N_5174);
or U7534 (N_7534,N_6570,N_6309);
xnor U7535 (N_7535,N_7361,N_5570);
nor U7536 (N_7536,N_6668,N_5940);
xor U7537 (N_7537,N_6154,N_5670);
xor U7538 (N_7538,N_5549,N_5140);
nand U7539 (N_7539,N_5974,N_7451);
xor U7540 (N_7540,N_5346,N_7213);
nor U7541 (N_7541,N_5496,N_6588);
nor U7542 (N_7542,N_5618,N_5785);
xor U7543 (N_7543,N_6735,N_5054);
nor U7544 (N_7544,N_7342,N_5952);
or U7545 (N_7545,N_5372,N_6524);
nor U7546 (N_7546,N_6353,N_6006);
xnor U7547 (N_7547,N_5083,N_7363);
nor U7548 (N_7548,N_5595,N_6977);
nor U7549 (N_7549,N_6567,N_6677);
nand U7550 (N_7550,N_5351,N_7476);
or U7551 (N_7551,N_5426,N_5828);
and U7552 (N_7552,N_5402,N_5020);
or U7553 (N_7553,N_6921,N_5914);
or U7554 (N_7554,N_5894,N_5835);
or U7555 (N_7555,N_5374,N_5443);
or U7556 (N_7556,N_5441,N_6207);
nand U7557 (N_7557,N_5359,N_7229);
xor U7558 (N_7558,N_6998,N_6124);
and U7559 (N_7559,N_6111,N_5580);
nand U7560 (N_7560,N_5423,N_7023);
nand U7561 (N_7561,N_7449,N_7326);
xor U7562 (N_7562,N_6800,N_7424);
xnor U7563 (N_7563,N_7276,N_5212);
and U7564 (N_7564,N_6877,N_6486);
and U7565 (N_7565,N_6974,N_5433);
xnor U7566 (N_7566,N_5122,N_7157);
xor U7567 (N_7567,N_5545,N_6151);
nand U7568 (N_7568,N_5225,N_6465);
or U7569 (N_7569,N_6461,N_5142);
nor U7570 (N_7570,N_7154,N_6737);
or U7571 (N_7571,N_7447,N_6655);
nor U7572 (N_7572,N_5532,N_6308);
nor U7573 (N_7573,N_7404,N_6669);
and U7574 (N_7574,N_6022,N_5218);
or U7575 (N_7575,N_6045,N_6264);
xnor U7576 (N_7576,N_5949,N_5900);
nand U7577 (N_7577,N_5652,N_5709);
nand U7578 (N_7578,N_5158,N_5578);
nor U7579 (N_7579,N_5308,N_5234);
and U7580 (N_7580,N_6914,N_6422);
xor U7581 (N_7581,N_5861,N_5653);
nand U7582 (N_7582,N_5171,N_5108);
xor U7583 (N_7583,N_5192,N_6063);
nand U7584 (N_7584,N_5732,N_6724);
nand U7585 (N_7585,N_6879,N_5273);
nor U7586 (N_7586,N_6098,N_6452);
nor U7587 (N_7587,N_5895,N_6603);
nor U7588 (N_7588,N_5756,N_5536);
nand U7589 (N_7589,N_7411,N_6665);
xnor U7590 (N_7590,N_6826,N_6699);
nor U7591 (N_7591,N_6397,N_6640);
xnor U7592 (N_7592,N_6286,N_6752);
nand U7593 (N_7593,N_5472,N_6497);
nor U7594 (N_7594,N_7481,N_6238);
xnor U7595 (N_7595,N_7299,N_5220);
and U7596 (N_7596,N_7012,N_6312);
xor U7597 (N_7597,N_5487,N_6957);
and U7598 (N_7598,N_6454,N_6632);
xnor U7599 (N_7599,N_5797,N_6425);
nor U7600 (N_7600,N_6562,N_7381);
xor U7601 (N_7601,N_7338,N_5502);
or U7602 (N_7602,N_7396,N_7389);
or U7603 (N_7603,N_6233,N_7267);
xor U7604 (N_7604,N_5418,N_6083);
and U7605 (N_7605,N_6389,N_7118);
nand U7606 (N_7606,N_6907,N_5832);
xor U7607 (N_7607,N_5498,N_7475);
xnor U7608 (N_7608,N_7353,N_5465);
nand U7609 (N_7609,N_5405,N_7156);
xnor U7610 (N_7610,N_6873,N_5169);
nand U7611 (N_7611,N_6671,N_7370);
or U7612 (N_7612,N_7444,N_6200);
nor U7613 (N_7613,N_6507,N_6159);
xnor U7614 (N_7614,N_6734,N_5953);
and U7615 (N_7615,N_5456,N_6161);
nor U7616 (N_7616,N_5181,N_5871);
nor U7617 (N_7617,N_6438,N_5593);
xnor U7618 (N_7618,N_7148,N_6287);
and U7619 (N_7619,N_5902,N_5937);
or U7620 (N_7620,N_6673,N_7224);
nor U7621 (N_7621,N_6090,N_6196);
or U7622 (N_7622,N_5379,N_6569);
xor U7623 (N_7623,N_5490,N_6306);
and U7624 (N_7624,N_6980,N_5962);
and U7625 (N_7625,N_6904,N_5544);
and U7626 (N_7626,N_5948,N_7446);
xor U7627 (N_7627,N_5357,N_7251);
or U7628 (N_7628,N_5432,N_5541);
xnor U7629 (N_7629,N_5420,N_6199);
nor U7630 (N_7630,N_5294,N_7019);
and U7631 (N_7631,N_5120,N_5327);
nor U7632 (N_7632,N_5692,N_7105);
xor U7633 (N_7633,N_7349,N_5413);
xor U7634 (N_7634,N_7452,N_5723);
nand U7635 (N_7635,N_6726,N_5104);
nor U7636 (N_7636,N_5912,N_6917);
nor U7637 (N_7637,N_6406,N_5092);
or U7638 (N_7638,N_7335,N_7220);
or U7639 (N_7639,N_6685,N_7170);
nor U7640 (N_7640,N_6981,N_5996);
or U7641 (N_7641,N_5393,N_6221);
nand U7642 (N_7642,N_5086,N_5001);
nand U7643 (N_7643,N_7162,N_6175);
nand U7644 (N_7644,N_5288,N_6197);
and U7645 (N_7645,N_5892,N_5515);
xnor U7646 (N_7646,N_7497,N_6595);
and U7647 (N_7647,N_7115,N_6061);
nand U7648 (N_7648,N_6611,N_5396);
and U7649 (N_7649,N_5950,N_6703);
nand U7650 (N_7650,N_5005,N_5858);
and U7651 (N_7651,N_6709,N_6361);
nand U7652 (N_7652,N_6982,N_5153);
nand U7653 (N_7653,N_7018,N_5622);
nand U7654 (N_7654,N_5792,N_5629);
xnor U7655 (N_7655,N_6700,N_6150);
nor U7656 (N_7656,N_7445,N_6528);
or U7657 (N_7657,N_6635,N_7261);
nand U7658 (N_7658,N_7394,N_6590);
xnor U7659 (N_7659,N_6833,N_7104);
nand U7660 (N_7660,N_6336,N_6598);
nand U7661 (N_7661,N_5317,N_5090);
or U7662 (N_7662,N_5829,N_6008);
and U7663 (N_7663,N_5474,N_5563);
or U7664 (N_7664,N_7400,N_6396);
nand U7665 (N_7665,N_5326,N_6936);
xnor U7666 (N_7666,N_6442,N_7492);
or U7667 (N_7667,N_7319,N_6994);
nor U7668 (N_7668,N_7350,N_6792);
or U7669 (N_7669,N_5781,N_6896);
or U7670 (N_7670,N_5015,N_5056);
and U7671 (N_7671,N_5735,N_6295);
nand U7672 (N_7672,N_6097,N_6906);
nand U7673 (N_7673,N_5210,N_6750);
and U7674 (N_7674,N_5213,N_5237);
nor U7675 (N_7675,N_5719,N_6015);
nand U7676 (N_7676,N_7339,N_5051);
nand U7677 (N_7677,N_5369,N_7056);
or U7678 (N_7678,N_5737,N_5450);
and U7679 (N_7679,N_5554,N_7345);
or U7680 (N_7680,N_5870,N_7264);
nand U7681 (N_7681,N_5577,N_5698);
and U7682 (N_7682,N_5318,N_5833);
nor U7683 (N_7683,N_6368,N_6441);
nand U7684 (N_7684,N_6195,N_5358);
xor U7685 (N_7685,N_7168,N_6972);
nand U7686 (N_7686,N_6717,N_6559);
nand U7687 (N_7687,N_6662,N_6831);
and U7688 (N_7688,N_5846,N_6253);
nor U7689 (N_7689,N_5926,N_6451);
or U7690 (N_7690,N_5149,N_5224);
nand U7691 (N_7691,N_5636,N_6351);
xnor U7692 (N_7692,N_5425,N_5072);
and U7693 (N_7693,N_5451,N_7160);
xor U7694 (N_7694,N_7029,N_5191);
xnor U7695 (N_7695,N_5337,N_6753);
or U7696 (N_7696,N_5795,N_6019);
or U7697 (N_7697,N_5057,N_5036);
xor U7698 (N_7698,N_6518,N_6492);
nand U7699 (N_7699,N_7453,N_6941);
or U7700 (N_7700,N_6202,N_7066);
nor U7701 (N_7701,N_6718,N_6179);
nand U7702 (N_7702,N_6030,N_6321);
or U7703 (N_7703,N_7122,N_5668);
nor U7704 (N_7704,N_6883,N_6416);
nand U7705 (N_7705,N_7373,N_6771);
or U7706 (N_7706,N_6589,N_5066);
nor U7707 (N_7707,N_6341,N_5022);
and U7708 (N_7708,N_6774,N_6934);
and U7709 (N_7709,N_7086,N_5060);
xor U7710 (N_7710,N_6804,N_5935);
and U7711 (N_7711,N_5600,N_5012);
or U7712 (N_7712,N_5582,N_6839);
nand U7713 (N_7713,N_6112,N_5339);
nor U7714 (N_7714,N_5383,N_7020);
and U7715 (N_7715,N_6508,N_6897);
xor U7716 (N_7716,N_5311,N_6781);
or U7717 (N_7717,N_6604,N_6205);
nor U7718 (N_7718,N_6115,N_7006);
or U7719 (N_7719,N_6649,N_6261);
nor U7720 (N_7720,N_6367,N_5528);
xor U7721 (N_7721,N_6095,N_6472);
nor U7722 (N_7722,N_6384,N_5282);
nor U7723 (N_7723,N_5687,N_5062);
nor U7724 (N_7724,N_7418,N_7222);
nand U7725 (N_7725,N_5688,N_7057);
xor U7726 (N_7726,N_7126,N_5306);
or U7727 (N_7727,N_6211,N_6257);
and U7728 (N_7728,N_7485,N_5113);
and U7729 (N_7729,N_5392,N_5127);
nor U7730 (N_7730,N_6775,N_5331);
or U7731 (N_7731,N_5223,N_6946);
and U7732 (N_7732,N_6143,N_5875);
and U7733 (N_7733,N_5074,N_5644);
or U7734 (N_7734,N_5135,N_5242);
xor U7735 (N_7735,N_5973,N_5204);
xor U7736 (N_7736,N_5365,N_5917);
xnor U7737 (N_7737,N_5312,N_5362);
xnor U7738 (N_7738,N_7233,N_7427);
and U7739 (N_7739,N_5232,N_5139);
or U7740 (N_7740,N_6363,N_7185);
and U7741 (N_7741,N_6085,N_6370);
xor U7742 (N_7742,N_6882,N_5931);
nor U7743 (N_7743,N_7190,N_7205);
nand U7744 (N_7744,N_6023,N_5195);
nor U7745 (N_7745,N_6137,N_5998);
nor U7746 (N_7746,N_5475,N_5523);
or U7747 (N_7747,N_7310,N_5459);
xnor U7748 (N_7748,N_7173,N_7042);
nand U7749 (N_7749,N_5274,N_6270);
and U7750 (N_7750,N_5377,N_6653);
and U7751 (N_7751,N_6169,N_6704);
and U7752 (N_7752,N_7180,N_5031);
xor U7753 (N_7753,N_7245,N_7437);
and U7754 (N_7754,N_5132,N_7367);
xor U7755 (N_7755,N_5842,N_5575);
nand U7756 (N_7756,N_5000,N_6987);
and U7757 (N_7757,N_5610,N_7182);
nor U7758 (N_7758,N_5510,N_6905);
xnor U7759 (N_7759,N_5521,N_5412);
nor U7760 (N_7760,N_6012,N_6428);
and U7761 (N_7761,N_6157,N_7322);
xor U7762 (N_7762,N_5626,N_5837);
nand U7763 (N_7763,N_7025,N_7091);
xnor U7764 (N_7764,N_7307,N_7473);
xnor U7765 (N_7765,N_7083,N_6109);
nand U7766 (N_7766,N_6100,N_6072);
or U7767 (N_7767,N_6176,N_6872);
nand U7768 (N_7768,N_6304,N_7030);
and U7769 (N_7769,N_5494,N_6854);
xor U7770 (N_7770,N_6362,N_6477);
or U7771 (N_7771,N_6401,N_6751);
nand U7772 (N_7772,N_6514,N_7199);
nor U7773 (N_7773,N_6612,N_6646);
nand U7774 (N_7774,N_6814,N_7378);
and U7775 (N_7775,N_6229,N_5161);
nor U7776 (N_7776,N_6035,N_7189);
nand U7777 (N_7777,N_5637,N_7323);
nand U7778 (N_7778,N_6509,N_7395);
and U7779 (N_7779,N_5024,N_7358);
nor U7780 (N_7780,N_6104,N_5277);
and U7781 (N_7781,N_6054,N_7232);
xnor U7782 (N_7782,N_5109,N_5363);
and U7783 (N_7783,N_5354,N_6194);
nand U7784 (N_7784,N_5011,N_5107);
or U7785 (N_7785,N_6651,N_6539);
or U7786 (N_7786,N_7332,N_7410);
nand U7787 (N_7787,N_5175,N_6347);
nor U7788 (N_7788,N_5587,N_7316);
or U7789 (N_7789,N_6656,N_5387);
xor U7790 (N_7790,N_5129,N_7055);
or U7791 (N_7791,N_6326,N_7239);
xnor U7792 (N_7792,N_5922,N_5954);
nand U7793 (N_7793,N_5466,N_6754);
and U7794 (N_7794,N_6929,N_5207);
nand U7795 (N_7795,N_7413,N_5635);
xnor U7796 (N_7796,N_7102,N_5517);
and U7797 (N_7797,N_6684,N_5946);
and U7798 (N_7798,N_6376,N_5081);
and U7799 (N_7799,N_5773,N_5576);
nand U7800 (N_7800,N_5979,N_5507);
xnor U7801 (N_7801,N_7372,N_5384);
nand U7802 (N_7802,N_6844,N_5196);
and U7803 (N_7803,N_7419,N_6786);
and U7804 (N_7804,N_6740,N_5550);
xor U7805 (N_7805,N_5253,N_5713);
xor U7806 (N_7806,N_5830,N_5802);
nand U7807 (N_7807,N_6592,N_7070);
and U7808 (N_7808,N_7101,N_6892);
or U7809 (N_7809,N_7169,N_5240);
nor U7810 (N_7810,N_6824,N_7375);
and U7811 (N_7811,N_6573,N_7280);
nor U7812 (N_7812,N_5686,N_6861);
xor U7813 (N_7813,N_6572,N_6899);
nand U7814 (N_7814,N_5604,N_6866);
xnor U7815 (N_7815,N_6556,N_7409);
nor U7816 (N_7816,N_5893,N_5730);
nor U7817 (N_7817,N_7327,N_6440);
and U7818 (N_7818,N_5888,N_5509);
xnor U7819 (N_7819,N_5130,N_7017);
and U7820 (N_7820,N_6144,N_7248);
or U7821 (N_7821,N_5495,N_7163);
nor U7822 (N_7822,N_6760,N_6940);
xnor U7823 (N_7823,N_5873,N_6088);
or U7824 (N_7824,N_5491,N_7405);
or U7825 (N_7825,N_5598,N_7275);
xor U7826 (N_7826,N_7313,N_7430);
and U7827 (N_7827,N_7369,N_5697);
nor U7828 (N_7828,N_6922,N_5907);
nor U7829 (N_7829,N_6092,N_5479);
nand U7830 (N_7830,N_6078,N_5322);
and U7831 (N_7831,N_7121,N_5138);
nand U7832 (N_7832,N_6663,N_6626);
or U7833 (N_7833,N_7416,N_6445);
xnor U7834 (N_7834,N_6617,N_7471);
and U7835 (N_7835,N_7364,N_7348);
or U7836 (N_7836,N_6862,N_6743);
and U7837 (N_7837,N_7406,N_5724);
nor U7838 (N_7838,N_6962,N_5366);
nor U7839 (N_7839,N_6183,N_6639);
nand U7840 (N_7840,N_5275,N_5573);
xor U7841 (N_7841,N_5984,N_6352);
and U7842 (N_7842,N_5766,N_6984);
nand U7843 (N_7843,N_5018,N_7254);
nor U7844 (N_7844,N_6203,N_6496);
nand U7845 (N_7845,N_5506,N_6373);
nand U7846 (N_7846,N_7040,N_7098);
nand U7847 (N_7847,N_6810,N_5304);
xor U7848 (N_7848,N_6447,N_5470);
and U7849 (N_7849,N_6910,N_5033);
nand U7850 (N_7850,N_6003,N_6744);
nor U7851 (N_7851,N_5705,N_6842);
nor U7852 (N_7852,N_6533,N_7371);
nor U7853 (N_7853,N_5305,N_5683);
and U7854 (N_7854,N_7241,N_6519);
xnor U7855 (N_7855,N_5599,N_5546);
nor U7856 (N_7856,N_6170,N_6860);
nand U7857 (N_7857,N_5887,N_6074);
and U7858 (N_7858,N_6620,N_6542);
nor U7859 (N_7859,N_5614,N_7274);
and U7860 (N_7860,N_6535,N_5039);
xor U7861 (N_7861,N_6134,N_6325);
xor U7862 (N_7862,N_5200,N_5767);
xnor U7863 (N_7863,N_7305,N_5776);
and U7864 (N_7864,N_6531,N_5674);
nand U7865 (N_7865,N_7250,N_5044);
or U7866 (N_7866,N_5800,N_5079);
xor U7867 (N_7867,N_6212,N_6033);
nand U7868 (N_7868,N_6385,N_5884);
or U7869 (N_7869,N_7286,N_6727);
and U7870 (N_7870,N_5489,N_6963);
and U7871 (N_7871,N_5816,N_6310);
or U7872 (N_7872,N_7051,N_6628);
nor U7873 (N_7873,N_6344,N_7484);
nand U7874 (N_7874,N_5564,N_6071);
xnor U7875 (N_7875,N_7247,N_7263);
or U7876 (N_7876,N_7103,N_5865);
xnor U7877 (N_7877,N_6087,N_6613);
xnor U7878 (N_7878,N_6606,N_5073);
nand U7879 (N_7879,N_6007,N_7288);
and U7880 (N_7880,N_5178,N_7043);
xor U7881 (N_7881,N_6859,N_5052);
and U7882 (N_7882,N_5748,N_6647);
nand U7883 (N_7883,N_7117,N_5291);
nand U7884 (N_7884,N_7037,N_7044);
and U7885 (N_7885,N_6423,N_5154);
nor U7886 (N_7886,N_7210,N_7318);
xor U7887 (N_7887,N_7393,N_6113);
and U7888 (N_7888,N_7225,N_6667);
xnor U7889 (N_7889,N_5983,N_5002);
or U7890 (N_7890,N_7099,N_7141);
or U7891 (N_7891,N_5819,N_5665);
xnor U7892 (N_7892,N_6431,N_6337);
and U7893 (N_7893,N_5106,N_6721);
and U7894 (N_7894,N_6070,N_5623);
xor U7895 (N_7895,N_5838,N_7278);
xnor U7896 (N_7896,N_6067,N_5565);
nor U7897 (N_7897,N_6123,N_5968);
nand U7898 (N_7898,N_5134,N_6462);
xnor U7899 (N_7899,N_5591,N_6456);
nor U7900 (N_7900,N_6675,N_5221);
nor U7901 (N_7901,N_6210,N_5035);
and U7902 (N_7902,N_6293,N_6457);
and U7903 (N_7903,N_5409,N_7201);
nor U7904 (N_7904,N_6770,N_6748);
and U7905 (N_7905,N_5957,N_6434);
and U7906 (N_7906,N_6827,N_6566);
nand U7907 (N_7907,N_6125,N_5608);
nand U7908 (N_7908,N_6849,N_6165);
xnor U7909 (N_7909,N_5815,N_6268);
nand U7910 (N_7910,N_5347,N_5141);
and U7911 (N_7911,N_6945,N_7420);
nand U7912 (N_7912,N_5089,N_6636);
and U7913 (N_7913,N_7047,N_5631);
nor U7914 (N_7914,N_6674,N_5913);
xnor U7915 (N_7915,N_7314,N_5285);
or U7916 (N_7916,N_6259,N_6291);
xor U7917 (N_7917,N_5116,N_7194);
xor U7918 (N_7918,N_6031,N_7289);
xor U7919 (N_7919,N_5085,N_6690);
nor U7920 (N_7920,N_6029,N_5355);
nand U7921 (N_7921,N_7242,N_6395);
and U7922 (N_7922,N_6329,N_6383);
and U7923 (N_7923,N_6464,N_6117);
nor U7924 (N_7924,N_6918,N_5649);
or U7925 (N_7925,N_7458,N_5016);
or U7926 (N_7926,N_5214,N_7355);
xnor U7927 (N_7927,N_5807,N_5695);
and U7928 (N_7928,N_6392,N_7432);
nand U7929 (N_7929,N_6158,N_6961);
xnor U7930 (N_7930,N_5124,N_6180);
xor U7931 (N_7931,N_6730,N_6439);
or U7932 (N_7932,N_7244,N_5669);
nand U7933 (N_7933,N_6670,N_6487);
and U7934 (N_7934,N_6281,N_5445);
xnor U7935 (N_7935,N_6928,N_6610);
and U7936 (N_7936,N_5524,N_7207);
and U7937 (N_7937,N_7401,N_6412);
xnor U7938 (N_7938,N_7133,N_6358);
and U7939 (N_7939,N_7343,N_6499);
or U7940 (N_7940,N_6271,N_5543);
or U7941 (N_7941,N_6393,N_6342);
nor U7942 (N_7942,N_5457,N_7426);
or U7943 (N_7943,N_6853,N_6887);
or U7944 (N_7944,N_7228,N_5246);
and U7945 (N_7945,N_7320,N_5725);
nor U7946 (N_7946,N_6018,N_7135);
and U7947 (N_7947,N_7137,N_7376);
and U7948 (N_7948,N_5925,N_6933);
and U7949 (N_7949,N_6557,N_6227);
xor U7950 (N_7950,N_5228,N_6537);
xor U7951 (N_7951,N_6517,N_7380);
xnor U7952 (N_7952,N_7067,N_5146);
or U7953 (N_7953,N_7100,N_5026);
nand U7954 (N_7954,N_5676,N_5967);
or U7955 (N_7955,N_6468,N_6919);
and U7956 (N_7956,N_5783,N_6534);
nor U7957 (N_7957,N_5059,N_5400);
xnor U7958 (N_7958,N_6978,N_5985);
xor U7959 (N_7959,N_5332,N_5329);
xor U7960 (N_7960,N_6360,N_5987);
and U7961 (N_7961,N_6511,N_7147);
nand U7962 (N_7962,N_7045,N_7309);
nand U7963 (N_7963,N_5939,N_6729);
nor U7964 (N_7964,N_5170,N_7002);
nand U7965 (N_7965,N_5215,N_6419);
xnor U7966 (N_7966,N_5693,N_6333);
nor U7967 (N_7967,N_6122,N_5818);
nor U7968 (N_7968,N_6413,N_6820);
xor U7969 (N_7969,N_6348,N_6218);
xor U7970 (N_7970,N_5064,N_5438);
nand U7971 (N_7971,N_5839,N_5645);
nand U7972 (N_7972,N_7178,N_5247);
xor U7973 (N_7973,N_7204,N_5508);
or U7974 (N_7974,N_5535,N_6992);
xnor U7975 (N_7975,N_5187,N_7164);
nor U7976 (N_7976,N_6201,N_5114);
nor U7977 (N_7977,N_6224,N_5231);
nor U7978 (N_7978,N_6631,N_6867);
or U7979 (N_7979,N_5157,N_7285);
nor U7980 (N_7980,N_6282,N_7469);
xnor U7981 (N_7981,N_7050,N_5739);
and U7982 (N_7982,N_6789,N_5032);
or U7983 (N_7983,N_7262,N_5264);
nand U7984 (N_7984,N_6579,N_6755);
nor U7985 (N_7985,N_6302,N_6516);
and U7986 (N_7986,N_5639,N_5727);
or U7987 (N_7987,N_5989,N_7028);
nor U7988 (N_7988,N_5848,N_7377);
nand U7989 (N_7989,N_5567,N_7347);
and U7990 (N_7990,N_5981,N_5855);
and U7991 (N_7991,N_5551,N_6583);
nor U7992 (N_7992,N_5663,N_6236);
or U7993 (N_7993,N_6410,N_6317);
xor U7994 (N_7994,N_5620,N_7456);
or U7995 (N_7995,N_6548,N_5970);
and U7996 (N_7996,N_7383,N_5343);
xnor U7997 (N_7997,N_5172,N_5919);
and U7998 (N_7998,N_6911,N_6414);
nor U7999 (N_7999,N_6884,N_5678);
xnor U8000 (N_8000,N_6148,N_6240);
and U8001 (N_8001,N_6262,N_5103);
nor U8002 (N_8002,N_6741,N_6970);
nor U8003 (N_8003,N_6320,N_7079);
nand U8004 (N_8004,N_5988,N_6652);
nor U8005 (N_8005,N_6094,N_7431);
or U8006 (N_8006,N_5881,N_7464);
nand U8007 (N_8007,N_6644,N_5125);
and U8008 (N_8008,N_6616,N_5804);
and U8009 (N_8009,N_7032,N_6068);
nor U8010 (N_8010,N_5841,N_7486);
nand U8011 (N_8011,N_5869,N_5245);
nor U8012 (N_8012,N_6448,N_5722);
nor U8013 (N_8013,N_5473,N_5430);
xor U8014 (N_8014,N_5562,N_7216);
xnor U8015 (N_8015,N_5435,N_6079);
nor U8016 (N_8016,N_6459,N_5289);
nand U8017 (N_8017,N_5042,N_6571);
nor U8018 (N_8018,N_6658,N_7259);
xor U8019 (N_8019,N_7166,N_6601);
or U8020 (N_8020,N_5398,N_6687);
and U8021 (N_8021,N_6185,N_7211);
nor U8022 (N_8022,N_5084,N_5077);
xnor U8023 (N_8023,N_6547,N_6738);
xor U8024 (N_8024,N_7462,N_7113);
and U8025 (N_8025,N_6780,N_6965);
nor U8026 (N_8026,N_7088,N_5606);
nor U8027 (N_8027,N_7330,N_5075);
or U8028 (N_8028,N_6506,N_5386);
and U8029 (N_8029,N_6004,N_6679);
or U8030 (N_8030,N_5186,N_6512);
nand U8031 (N_8031,N_7116,N_6356);
nor U8032 (N_8032,N_5283,N_5879);
nand U8033 (N_8033,N_5316,N_7235);
or U8034 (N_8034,N_5505,N_6455);
xor U8035 (N_8035,N_7120,N_5801);
or U8036 (N_8036,N_5063,N_6565);
and U8037 (N_8037,N_6424,N_7317);
nand U8038 (N_8038,N_7090,N_6664);
nor U8039 (N_8039,N_6335,N_6912);
nand U8040 (N_8040,N_6036,N_7443);
nand U8041 (N_8041,N_7296,N_5778);
nand U8042 (N_8042,N_5381,N_7143);
nand U8043 (N_8043,N_5348,N_5542);
or U8044 (N_8044,N_5690,N_5836);
or U8045 (N_8045,N_5380,N_5266);
xnor U8046 (N_8046,N_6024,N_6648);
nor U8047 (N_8047,N_6235,N_6931);
and U8048 (N_8048,N_6625,N_5779);
and U8049 (N_8049,N_7130,N_6989);
nand U8050 (N_8050,N_6430,N_5341);
or U8051 (N_8051,N_7457,N_7324);
nor U8052 (N_8052,N_6378,N_6387);
and U8053 (N_8053,N_7293,N_6593);
or U8054 (N_8054,N_7408,N_5537);
nand U8055 (N_8055,N_6269,N_6053);
nor U8056 (N_8056,N_5750,N_5611);
nor U8057 (N_8057,N_5731,N_6762);
nand U8058 (N_8058,N_6891,N_6857);
nand U8059 (N_8059,N_5854,N_7391);
and U8060 (N_8060,N_5743,N_6139);
xor U8061 (N_8061,N_7223,N_7321);
nor U8062 (N_8062,N_6327,N_6214);
or U8063 (N_8063,N_5584,N_7459);
nor U8064 (N_8064,N_6162,N_6390);
nand U8065 (N_8065,N_7209,N_6133);
or U8066 (N_8066,N_6947,N_5226);
or U8067 (N_8067,N_6777,N_5501);
and U8068 (N_8068,N_6680,N_5389);
xnor U8069 (N_8069,N_6908,N_7329);
xnor U8070 (N_8070,N_6001,N_6435);
xnor U8071 (N_8071,N_7279,N_6863);
or U8072 (N_8072,N_6756,N_5309);
or U8073 (N_8073,N_6815,N_5333);
nand U8074 (N_8074,N_5934,N_6105);
and U8075 (N_8075,N_5102,N_6836);
xor U8076 (N_8076,N_7052,N_5736);
nor U8077 (N_8077,N_6365,N_5091);
xor U8078 (N_8078,N_5775,N_6119);
or U8079 (N_8079,N_6681,N_5249);
and U8080 (N_8080,N_5219,N_7212);
and U8081 (N_8081,N_5100,N_5301);
and U8082 (N_8082,N_5006,N_7072);
xnor U8083 (N_8083,N_5826,N_6894);
xnor U8084 (N_8084,N_6276,N_6226);
xor U8085 (N_8085,N_7470,N_5199);
or U8086 (N_8086,N_6841,N_6600);
nor U8087 (N_8087,N_5352,N_5552);
or U8088 (N_8088,N_6637,N_7226);
nor U8089 (N_8089,N_5431,N_6044);
xnor U8090 (N_8090,N_6808,N_6252);
and U8091 (N_8091,N_5877,N_6822);
and U8092 (N_8092,N_6340,N_5715);
nand U8093 (N_8093,N_6273,N_6374);
xnor U8094 (N_8094,N_7269,N_5159);
or U8095 (N_8095,N_6234,N_7368);
xnor U8096 (N_8096,N_7461,N_6495);
xor U8097 (N_8097,N_6025,N_6830);
nand U8098 (N_8098,N_7183,N_7328);
and U8099 (N_8099,N_5905,N_6294);
nor U8100 (N_8100,N_6149,N_5193);
nand U8101 (N_8101,N_6446,N_6818);
and U8102 (N_8102,N_6878,N_6091);
and U8103 (N_8103,N_6708,N_6040);
and U8104 (N_8104,N_5596,N_7001);
and U8105 (N_8105,N_7026,N_6417);
xor U8106 (N_8106,N_5173,N_6217);
xor U8107 (N_8107,N_5726,N_5448);
nor U8108 (N_8108,N_6809,N_7027);
xor U8109 (N_8109,N_6114,N_5680);
nand U8110 (N_8110,N_5205,N_5770);
and U8111 (N_8111,N_7294,N_7227);
nand U8112 (N_8112,N_6181,N_6503);
nor U8113 (N_8113,N_7206,N_5977);
nor U8114 (N_8114,N_5370,N_7114);
nor U8115 (N_8115,N_5375,N_6526);
xnor U8116 (N_8116,N_5477,N_5661);
and U8117 (N_8117,N_5444,N_6371);
and U8118 (N_8118,N_5658,N_7301);
and U8119 (N_8119,N_6160,N_7034);
nand U8120 (N_8120,N_5734,N_5112);
and U8121 (N_8121,N_5008,N_6561);
or U8122 (N_8122,N_6108,N_7388);
nor U8123 (N_8123,N_5718,N_7384);
nand U8124 (N_8124,N_6585,N_5202);
or U8125 (N_8125,N_7062,N_6311);
nand U8126 (N_8126,N_5030,N_5694);
and U8127 (N_8127,N_7082,N_5050);
nor U8128 (N_8128,N_5189,N_7312);
nor U8129 (N_8129,N_7298,N_5728);
or U8130 (N_8130,N_5188,N_5302);
nor U8131 (N_8131,N_6243,N_6225);
and U8132 (N_8132,N_5406,N_6856);
nand U8133 (N_8133,N_7127,N_5478);
nor U8134 (N_8134,N_5167,N_6650);
nand U8135 (N_8135,N_5211,N_5558);
nor U8136 (N_8136,N_5632,N_7270);
and U8137 (N_8137,N_6582,N_6676);
xor U8138 (N_8138,N_5930,N_6812);
nand U8139 (N_8139,N_6101,N_6330);
and U8140 (N_8140,N_5455,N_5407);
and U8141 (N_8141,N_6449,N_5896);
nor U8142 (N_8142,N_6301,N_5999);
xnor U8143 (N_8143,N_6868,N_5744);
nor U8144 (N_8144,N_5082,N_5671);
xnor U8145 (N_8145,N_6796,N_5903);
nor U8146 (N_8146,N_5714,N_5638);
and U8147 (N_8147,N_7125,N_5121);
nor U8148 (N_8148,N_6968,N_5373);
nand U8149 (N_8149,N_6504,N_5798);
xnor U8150 (N_8150,N_6136,N_7150);
and U8151 (N_8151,N_7273,N_5045);
and U8152 (N_8152,N_7354,N_5080);
nor U8153 (N_8153,N_6895,N_7177);
and U8154 (N_8154,N_5956,N_6121);
xnor U8155 (N_8155,N_6767,N_5272);
nor U8156 (N_8156,N_6629,N_5229);
nor U8157 (N_8157,N_7334,N_5488);
nand U8158 (N_8158,N_5263,N_5449);
xor U8159 (N_8159,N_6835,N_5704);
or U8160 (N_8160,N_5019,N_6405);
and U8161 (N_8161,N_5061,N_6049);
nor U8162 (N_8162,N_6349,N_6166);
nor U8163 (N_8163,N_6522,N_6386);
nand U8164 (N_8164,N_6081,N_5323);
xor U8165 (N_8165,N_7433,N_5115);
nor U8166 (N_8166,N_6521,N_5556);
and U8167 (N_8167,N_6379,N_5927);
xor U8168 (N_8168,N_5811,N_7290);
xor U8169 (N_8169,N_5874,N_5166);
nand U8170 (N_8170,N_5367,N_6177);
and U8171 (N_8171,N_7240,N_6520);
or U8172 (N_8172,N_6902,N_5824);
or U8173 (N_8173,N_5013,N_6953);
nand U8174 (N_8174,N_6331,N_7089);
xor U8175 (N_8175,N_6782,N_6116);
xor U8176 (N_8176,N_5520,N_6480);
and U8177 (N_8177,N_7340,N_5659);
nand U8178 (N_8178,N_6937,N_5160);
nor U8179 (N_8179,N_5859,N_6705);
or U8180 (N_8180,N_5143,N_7308);
or U8181 (N_8181,N_5217,N_5462);
nor U8182 (N_8182,N_5145,N_7249);
and U8183 (N_8183,N_5793,N_5943);
xnor U8184 (N_8184,N_5437,N_7128);
xor U8185 (N_8185,N_6799,N_7489);
nor U8186 (N_8186,N_6795,N_5738);
or U8187 (N_8187,N_5810,N_6701);
or U8188 (N_8188,N_5960,N_6280);
and U8189 (N_8189,N_5972,N_5571);
nor U8190 (N_8190,N_5321,N_5555);
nor U8191 (N_8191,N_5590,N_5572);
xor U8192 (N_8192,N_5118,N_7035);
and U8193 (N_8193,N_7015,N_5761);
xnor U8194 (N_8194,N_5469,N_6483);
nand U8195 (N_8195,N_5538,N_6925);
nand U8196 (N_8196,N_6107,N_6837);
or U8197 (N_8197,N_6720,N_7144);
or U8198 (N_8198,N_7468,N_5991);
and U8199 (N_8199,N_5483,N_6471);
or U8200 (N_8200,N_6529,N_6283);
or U8201 (N_8201,N_6747,N_5330);
nand U8202 (N_8202,N_6178,N_5882);
or U8203 (N_8203,N_6807,N_6494);
or U8204 (N_8204,N_6265,N_7119);
nand U8205 (N_8205,N_7033,N_5700);
nand U8206 (N_8206,N_6239,N_7390);
or U8207 (N_8207,N_5787,N_5961);
nand U8208 (N_8208,N_7009,N_7078);
and U8209 (N_8209,N_7402,N_5216);
nor U8210 (N_8210,N_5843,N_6855);
nand U8211 (N_8211,N_7188,N_5261);
xor U8212 (N_8212,N_5284,N_5243);
xor U8213 (N_8213,N_7297,N_7193);
nor U8214 (N_8214,N_5643,N_5070);
xnor U8215 (N_8215,N_5920,N_5844);
or U8216 (N_8216,N_7287,N_6924);
xor U8217 (N_8217,N_5650,N_5993);
xor U8218 (N_8218,N_6787,N_5906);
or U8219 (N_8219,N_6059,N_6299);
xnor U8220 (N_8220,N_5360,N_6409);
and U8221 (N_8221,N_6784,N_5630);
nor U8222 (N_8222,N_5548,N_5029);
nor U8223 (N_8223,N_7184,N_6532);
and U8224 (N_8224,N_5069,N_7171);
nand U8225 (N_8225,N_5627,N_5511);
nand U8226 (N_8226,N_5250,N_7474);
or U8227 (N_8227,N_6549,N_6739);
xnor U8228 (N_8228,N_5227,N_7415);
and U8229 (N_8229,N_7454,N_5860);
nand U8230 (N_8230,N_6707,N_7111);
nor U8231 (N_8231,N_6296,N_6219);
or U8232 (N_8232,N_6869,N_6267);
or U8233 (N_8233,N_5982,N_5707);
nand U8234 (N_8234,N_6764,N_6695);
or U8235 (N_8235,N_5759,N_5747);
or U8236 (N_8236,N_6375,N_7038);
xnor U8237 (N_8237,N_6251,N_6791);
and U8238 (N_8238,N_6619,N_6551);
nor U8239 (N_8239,N_6811,N_5238);
or U8240 (N_8240,N_5119,N_6813);
nor U8241 (N_8241,N_6046,N_5641);
nand U8242 (N_8242,N_6502,N_5516);
or U8243 (N_8243,N_7243,N_7136);
nand U8244 (N_8244,N_5752,N_5878);
nor U8245 (N_8245,N_6339,N_6596);
nor U8246 (N_8246,N_5422,N_5853);
or U8247 (N_8247,N_7013,N_6563);
or U8248 (N_8248,N_5471,N_5368);
nor U8249 (N_8249,N_6377,N_7333);
nor U8250 (N_8250,N_6951,N_6716);
nor U8251 (N_8251,N_6076,N_7252);
xnor U8252 (N_8252,N_5612,N_5831);
or U8253 (N_8253,N_7466,N_6303);
nor U8254 (N_8254,N_5666,N_6129);
or U8255 (N_8255,N_6322,N_6850);
and U8256 (N_8256,N_5691,N_6772);
nand U8257 (N_8257,N_6453,N_5821);
xnor U8258 (N_8258,N_6638,N_5568);
and U8259 (N_8259,N_5911,N_6171);
nand U8260 (N_8260,N_6485,N_6042);
and U8261 (N_8261,N_5095,N_5867);
nand U8262 (N_8262,N_5525,N_5856);
nand U8263 (N_8263,N_7386,N_5399);
and U8264 (N_8264,N_5014,N_7112);
and U8265 (N_8265,N_6622,N_5980);
nand U8266 (N_8266,N_6785,N_5677);
nand U8267 (N_8267,N_5165,N_5936);
nor U8268 (N_8268,N_5314,N_6420);
nor U8269 (N_8269,N_5342,N_5148);
or U8270 (N_8270,N_6693,N_7138);
xor U8271 (N_8271,N_7146,N_7208);
xor U8272 (N_8272,N_6725,N_6568);
or U8273 (N_8273,N_6411,N_6880);
nor U8274 (N_8274,N_5128,N_6530);
xor U8275 (N_8275,N_5111,N_5404);
nand U8276 (N_8276,N_5602,N_5794);
and U8277 (N_8277,N_6255,N_6047);
or U8278 (N_8278,N_5850,N_5969);
nor U8279 (N_8279,N_5096,N_7129);
and U8280 (N_8280,N_5763,N_5177);
nand U8281 (N_8281,N_5904,N_5428);
or U8282 (N_8282,N_6942,N_5087);
nand U8283 (N_8283,N_7060,N_7428);
nor U8284 (N_8284,N_5886,N_6927);
or U8285 (N_8285,N_6338,N_5131);
and U8286 (N_8286,N_6900,N_6147);
nand U8287 (N_8287,N_7429,N_6366);
and U8288 (N_8288,N_6591,N_5711);
nor U8289 (N_8289,N_6332,N_6641);
nand U8290 (N_8290,N_7084,N_6256);
nor U8291 (N_8291,N_5769,N_6069);
nand U8292 (N_8292,N_6715,N_6722);
nand U8293 (N_8293,N_5254,N_7292);
and U8294 (N_8294,N_5847,N_7149);
xnor U8295 (N_8295,N_5889,N_5371);
and U8296 (N_8296,N_6958,N_7200);
nand U8297 (N_8297,N_6858,N_6215);
and U8298 (N_8298,N_5446,N_6659);
xnor U8299 (N_8299,N_5270,N_5657);
nor U8300 (N_8300,N_5136,N_5401);
or U8301 (N_8301,N_6909,N_6182);
nand U8302 (N_8302,N_7271,N_6543);
nand U8303 (N_8303,N_6055,N_6969);
nor U8304 (N_8304,N_6976,N_5248);
nand U8305 (N_8305,N_6926,N_5820);
and U8306 (N_8306,N_6759,N_6174);
or U8307 (N_8307,N_5864,N_5163);
nor U8308 (N_8308,N_5439,N_6357);
or U8309 (N_8309,N_6478,N_5286);
nor U8310 (N_8310,N_6450,N_6706);
nor U8311 (N_8311,N_5758,N_5901);
nor U8312 (N_8312,N_7140,N_6840);
nand U8313 (N_8313,N_6761,N_5458);
nand U8314 (N_8314,N_7151,N_6274);
xor U8315 (N_8315,N_6443,N_6578);
xor U8316 (N_8316,N_7365,N_6876);
xor U8317 (N_8317,N_5378,N_5340);
xor U8318 (N_8318,N_6415,N_5672);
and U8319 (N_8319,N_7108,N_5947);
xor U8320 (N_8320,N_6702,N_6564);
nor U8321 (N_8321,N_6614,N_6318);
nand U8322 (N_8322,N_7191,N_5328);
nor U8323 (N_8323,N_7465,N_7494);
nand U8324 (N_8324,N_6246,N_6408);
xor U8325 (N_8325,N_6163,N_6765);
and U8326 (N_8326,N_5975,N_6020);
nand U8327 (N_8327,N_6732,N_6555);
and U8328 (N_8328,N_5746,N_6034);
nor U8329 (N_8329,N_5429,N_6645);
nor U8330 (N_8330,N_7186,N_5771);
and U8331 (N_8331,N_5921,N_5997);
xnor U8332 (N_8332,N_5256,N_5058);
xnor U8333 (N_8333,N_6102,N_7472);
nand U8334 (N_8334,N_5656,N_6797);
or U8335 (N_8335,N_5594,N_7110);
nor U8336 (N_8336,N_5990,N_7007);
nor U8337 (N_8337,N_5176,N_7010);
nand U8338 (N_8338,N_5390,N_6484);
nand U8339 (N_8339,N_6846,N_5588);
nand U8340 (N_8340,N_7016,N_7483);
or U8341 (N_8341,N_6099,N_5279);
nand U8342 (N_8342,N_6580,N_5184);
nor U8343 (N_8343,N_6407,N_5679);
nor U8344 (N_8344,N_6758,N_6481);
or U8345 (N_8345,N_6223,N_6315);
and U8346 (N_8346,N_5126,N_6027);
or U8347 (N_8347,N_6432,N_6017);
xor U8348 (N_8348,N_5995,N_6037);
nor U8349 (N_8349,N_6190,N_6819);
or U8350 (N_8350,N_7360,N_7172);
nor U8351 (N_8351,N_6297,N_6541);
xnor U8352 (N_8352,N_5046,N_5814);
nand U8353 (N_8353,N_5021,N_6307);
or U8354 (N_8354,N_6574,N_7215);
or U8355 (N_8355,N_6285,N_5955);
or U8356 (N_8356,N_6964,N_7266);
or U8357 (N_8357,N_6026,N_7455);
nor U8358 (N_8358,N_5646,N_5361);
or U8359 (N_8359,N_7061,N_6985);
and U8360 (N_8360,N_5932,N_6874);
and U8361 (N_8361,N_5349,N_6713);
and U8362 (N_8362,N_7496,N_7403);
xor U8363 (N_8363,N_5299,N_6893);
or U8364 (N_8364,N_5094,N_6398);
nand U8365 (N_8365,N_7255,N_5897);
xor U8366 (N_8366,N_6275,N_5898);
nor U8367 (N_8367,N_5296,N_7283);
or U8368 (N_8368,N_5492,N_5655);
nor U8369 (N_8369,N_5619,N_6300);
nand U8370 (N_8370,N_7046,N_5464);
or U8371 (N_8371,N_5928,N_5566);
or U8372 (N_8372,N_5105,N_5098);
nor U8373 (N_8373,N_6692,N_6213);
nand U8374 (N_8374,N_6073,N_6802);
xnor U8375 (N_8375,N_6064,N_5929);
and U8376 (N_8376,N_5230,N_7064);
xnor U8377 (N_8377,N_6011,N_5890);
or U8378 (N_8378,N_5963,N_6132);
and U8379 (N_8379,N_6834,N_7253);
xor U8380 (N_8380,N_5786,N_5068);
and U8381 (N_8381,N_7187,N_5442);
or U8382 (N_8382,N_6400,N_7022);
nand U8383 (N_8383,N_5203,N_5667);
and U8384 (N_8384,N_5027,N_5518);
xnor U8385 (N_8385,N_6231,N_7234);
xor U8386 (N_8386,N_6779,N_7085);
or U8387 (N_8387,N_6319,N_5463);
nand U8388 (N_8388,N_6284,N_5603);
xor U8389 (N_8389,N_6277,N_5986);
xor U8390 (N_8390,N_5049,N_7341);
or U8391 (N_8391,N_7387,N_5320);
nor U8392 (N_8392,N_6052,N_7488);
or U8393 (N_8393,N_6474,N_6354);
nor U8394 (N_8394,N_5966,N_5382);
nor U8395 (N_8395,N_5067,N_5239);
xor U8396 (N_8396,N_5287,N_6429);
or U8397 (N_8397,N_5010,N_7434);
nor U8398 (N_8398,N_5880,N_5476);
nor U8399 (N_8399,N_7300,N_5152);
xor U8400 (N_8400,N_6710,N_5156);
nor U8401 (N_8401,N_6935,N_7132);
and U8402 (N_8402,N_6250,N_5742);
or U8403 (N_8403,N_5527,N_5753);
nor U8404 (N_8404,N_7422,N_5689);
xor U8405 (N_8405,N_6798,N_5480);
xor U8406 (N_8406,N_6609,N_6266);
nand U8407 (N_8407,N_5754,N_6768);
or U8408 (N_8408,N_7069,N_5037);
xnor U8409 (N_8409,N_6345,N_6126);
xnor U8410 (N_8410,N_5324,N_7024);
or U8411 (N_8411,N_6248,N_6577);
nand U8412 (N_8412,N_6140,N_6187);
and U8413 (N_8413,N_6954,N_5616);
or U8414 (N_8414,N_6825,N_6686);
nand U8415 (N_8415,N_5197,N_7174);
xor U8416 (N_8416,N_6944,N_7315);
and U8417 (N_8417,N_6145,N_7295);
xor U8418 (N_8418,N_6736,N_7107);
or U8419 (N_8419,N_6131,N_7003);
or U8420 (N_8420,N_6491,N_7436);
or U8421 (N_8421,N_7221,N_7277);
nand U8422 (N_8422,N_6550,N_5038);
nand U8423 (N_8423,N_7303,N_6470);
and U8424 (N_8424,N_7068,N_6314);
or U8425 (N_8425,N_5486,N_6698);
xor U8426 (N_8426,N_6865,N_6821);
xnor U8427 (N_8427,N_5760,N_6463);
or U8428 (N_8428,N_5162,N_7379);
xor U8429 (N_8429,N_5461,N_5512);
and U8430 (N_8430,N_5235,N_7236);
or U8431 (N_8431,N_6164,N_6254);
nor U8432 (N_8432,N_6394,N_5436);
or U8433 (N_8433,N_6916,N_7004);
nand U8434 (N_8434,N_7385,N_7291);
or U8435 (N_8435,N_7071,N_6380);
or U8436 (N_8436,N_5416,N_5345);
nor U8437 (N_8437,N_6028,N_5417);
nor U8438 (N_8438,N_7407,N_7399);
nor U8439 (N_8439,N_6458,N_5621);
or U8440 (N_8440,N_6939,N_6241);
or U8441 (N_8441,N_7477,N_5774);
and U8442 (N_8442,N_5262,N_7282);
nand U8443 (N_8443,N_5712,N_6473);
nand U8444 (N_8444,N_7439,N_6403);
nor U8445 (N_8445,N_5923,N_6643);
xnor U8446 (N_8446,N_6289,N_6082);
nand U8447 (N_8447,N_5703,N_6493);
nor U8448 (N_8448,N_6156,N_5733);
xor U8449 (N_8449,N_5325,N_6075);
and U8450 (N_8450,N_5625,N_5236);
and U8451 (N_8451,N_5183,N_5356);
nor U8452 (N_8452,N_5944,N_7167);
nand U8453 (N_8453,N_6642,N_6152);
or U8454 (N_8454,N_5964,N_7304);
or U8455 (N_8455,N_5403,N_7080);
xnor U8456 (N_8456,N_6237,N_5958);
nand U8457 (N_8457,N_6127,N_6575);
nand U8458 (N_8458,N_7414,N_5526);
nor U8459 (N_8459,N_5681,N_6118);
and U8460 (N_8460,N_5942,N_6845);
and U8461 (N_8461,N_5201,N_7036);
nand U8462 (N_8462,N_5885,N_5751);
or U8463 (N_8463,N_6794,N_6597);
nor U8464 (N_8464,N_7087,N_5706);
xor U8465 (N_8465,N_6621,N_5421);
nor U8466 (N_8466,N_5269,N_6691);
nand U8467 (N_8467,N_6060,N_6956);
xnor U8468 (N_8468,N_6146,N_5796);
xnor U8469 (N_8469,N_5260,N_6847);
and U8470 (N_8470,N_6505,N_5634);
or U8471 (N_8471,N_6168,N_6678);
or U8472 (N_8472,N_5257,N_6885);
xnor U8473 (N_8473,N_5916,N_7161);
and U8474 (N_8474,N_6382,N_5613);
nand U8475 (N_8475,N_5003,N_6120);
or U8476 (N_8476,N_5344,N_7460);
nor U8477 (N_8477,N_5194,N_5994);
nor U8478 (N_8478,N_5190,N_7053);
nand U8479 (N_8479,N_6816,N_6466);
or U8480 (N_8480,N_6404,N_6898);
or U8481 (N_8481,N_6852,N_5685);
or U8482 (N_8482,N_5866,N_6057);
xnor U8483 (N_8483,N_5292,N_7440);
nand U8484 (N_8484,N_7441,N_7256);
and U8485 (N_8485,N_7346,N_6618);
nor U8486 (N_8486,N_7374,N_5721);
or U8487 (N_8487,N_6290,N_6913);
xnor U8488 (N_8488,N_6630,N_5297);
nand U8489 (N_8489,N_7398,N_6623);
and U8490 (N_8490,N_6871,N_5583);
nand U8491 (N_8491,N_6657,N_6584);
and U8492 (N_8492,N_6138,N_5503);
nor U8493 (N_8493,N_6920,N_6581);
or U8494 (N_8494,N_5863,N_5484);
nor U8495 (N_8495,N_7123,N_6666);
nor U8496 (N_8496,N_6776,N_7065);
xor U8497 (N_8497,N_5267,N_5007);
nand U8498 (N_8498,N_5918,N_6490);
nor U8499 (N_8499,N_6399,N_5777);
nand U8500 (N_8500,N_7482,N_6093);
nor U8501 (N_8501,N_6488,N_6959);
or U8502 (N_8502,N_5915,N_7392);
xnor U8503 (N_8503,N_5597,N_6010);
and U8504 (N_8504,N_6607,N_7155);
nand U8505 (N_8505,N_6696,N_6993);
and U8506 (N_8506,N_5300,N_6433);
nor U8507 (N_8507,N_6938,N_6141);
nor U8508 (N_8508,N_5978,N_6950);
or U8509 (N_8509,N_5559,N_7463);
and U8510 (N_8510,N_5255,N_5624);
nor U8511 (N_8511,N_5617,N_6552);
xnor U8512 (N_8512,N_7219,N_5729);
nor U8513 (N_8513,N_5298,N_7442);
and U8514 (N_8514,N_6476,N_5581);
or U8515 (N_8515,N_5702,N_6313);
xnor U8516 (N_8516,N_7356,N_6475);
nor U8517 (N_8517,N_5553,N_7246);
and U8518 (N_8518,N_6694,N_5180);
nand U8519 (N_8519,N_6479,N_5271);
or U8520 (N_8520,N_6381,N_5933);
and U8521 (N_8521,N_5992,N_6184);
nand U8522 (N_8522,N_6634,N_5749);
and U8523 (N_8523,N_6208,N_5971);
nand U8524 (N_8524,N_6783,N_6128);
and U8525 (N_8525,N_5574,N_7479);
nand U8526 (N_8526,N_5813,N_7359);
and U8527 (N_8527,N_6769,N_5540);
or U8528 (N_8528,N_7306,N_6943);
or U8529 (N_8529,N_6080,N_5823);
nand U8530 (N_8530,N_6983,N_6427);
nor U8531 (N_8531,N_5534,N_6500);
nor U8532 (N_8532,N_6013,N_6986);
and U8533 (N_8533,N_6056,N_5976);
xnor U8534 (N_8534,N_5137,N_5799);
and U8535 (N_8535,N_6323,N_5605);
and U8536 (N_8536,N_5338,N_6077);
and U8537 (N_8537,N_5827,N_5410);
or U8538 (N_8538,N_6790,N_7179);
nand U8539 (N_8539,N_6364,N_7005);
nand U8540 (N_8540,N_5640,N_6263);
xnor U8541 (N_8541,N_5682,N_6089);
and U8542 (N_8542,N_5557,N_7218);
nor U8543 (N_8543,N_7139,N_6608);
and U8544 (N_8544,N_6554,N_5852);
xor U8545 (N_8545,N_7257,N_6510);
and U8546 (N_8546,N_6247,N_5664);
xnor U8547 (N_8547,N_6890,N_5209);
nand U8548 (N_8548,N_6106,N_6763);
and U8549 (N_8549,N_5408,N_6209);
xnor U8550 (N_8550,N_5097,N_6173);
nand U8551 (N_8551,N_6216,N_6167);
xnor U8552 (N_8552,N_5293,N_6388);
nor U8553 (N_8553,N_5093,N_6206);
nand U8554 (N_8554,N_5849,N_6540);
xnor U8555 (N_8555,N_6272,N_7336);
xnor U8556 (N_8556,N_7196,N_7351);
nand U8557 (N_8557,N_7272,N_5144);
nor U8558 (N_8558,N_6688,N_6967);
nand U8559 (N_8559,N_6065,N_5499);
xnor U8560 (N_8560,N_5419,N_5805);
nor U8561 (N_8561,N_5350,N_7258);
and U8562 (N_8562,N_7074,N_6191);
or U8563 (N_8563,N_6204,N_5411);
and U8564 (N_8564,N_7325,N_5415);
and U8565 (N_8565,N_5164,N_7281);
and U8566 (N_8566,N_7131,N_6712);
or U8567 (N_8567,N_5601,N_7357);
and U8568 (N_8568,N_5099,N_6469);
xnor U8569 (N_8569,N_6888,N_5909);
nand U8570 (N_8570,N_5385,N_5513);
and U8571 (N_8571,N_6359,N_7435);
nand U8572 (N_8572,N_6605,N_6288);
xnor U8573 (N_8573,N_5589,N_5834);
nor U8574 (N_8574,N_7423,N_7096);
and U8575 (N_8575,N_5806,N_5017);
or U8576 (N_8576,N_6558,N_7049);
or U8577 (N_8577,N_5586,N_6805);
nand U8578 (N_8578,N_6086,N_7480);
nor U8579 (N_8579,N_6553,N_6039);
xor U8580 (N_8580,N_5493,N_7175);
or U8581 (N_8581,N_6870,N_7059);
xor U8582 (N_8582,N_5467,N_6523);
and U8583 (N_8583,N_6437,N_7176);
nand U8584 (N_8584,N_5822,N_5460);
nand U8585 (N_8585,N_6930,N_6096);
nor U8586 (N_8586,N_7014,N_6498);
nor U8587 (N_8587,N_7352,N_6489);
nor U8588 (N_8588,N_7095,N_6189);
or U8589 (N_8589,N_5004,N_5803);
nor U8590 (N_8590,N_6975,N_5123);
nand U8591 (N_8591,N_6142,N_5910);
xor U8592 (N_8592,N_5364,N_7344);
nor U8593 (N_8593,N_6999,N_6258);
nand U8594 (N_8594,N_6279,N_5071);
nand U8595 (N_8595,N_5531,N_6728);
nand U8596 (N_8596,N_6672,N_6766);
nand U8597 (N_8597,N_6372,N_7011);
and U8598 (N_8598,N_6355,N_5397);
or U8599 (N_8599,N_5335,N_7048);
nor U8600 (N_8600,N_7214,N_7142);
xor U8601 (N_8601,N_6005,N_5151);
nor U8602 (N_8602,N_7490,N_6515);
nand U8603 (N_8603,N_7284,N_6749);
nand U8604 (N_8604,N_6683,N_5504);
xor U8605 (N_8605,N_7081,N_5155);
xor U8606 (N_8606,N_5560,N_6501);
nand U8607 (N_8607,N_6426,N_7499);
and U8608 (N_8608,N_5530,N_5514);
xor U8609 (N_8609,N_5009,N_5252);
or U8610 (N_8610,N_7145,N_5041);
and U8611 (N_8611,N_7198,N_7478);
nor U8612 (N_8612,N_7450,N_6714);
nor U8613 (N_8613,N_5522,N_7152);
or U8614 (N_8614,N_6244,N_6742);
xor U8615 (N_8615,N_6014,N_7195);
nand U8616 (N_8616,N_6731,N_5662);
and U8617 (N_8617,N_6536,N_5784);
nand U8618 (N_8618,N_7134,N_5812);
nor U8619 (N_8619,N_6832,N_5208);
xor U8620 (N_8620,N_6654,N_5745);
and U8621 (N_8621,N_5319,N_6000);
nor U8622 (N_8622,N_6793,N_6778);
xnor U8623 (N_8623,N_7260,N_5434);
nor U8624 (N_8624,N_5313,N_5043);
nand U8625 (N_8625,N_6624,N_5394);
nand U8626 (N_8626,N_5395,N_5539);
nand U8627 (N_8627,N_5497,N_6546);
nor U8628 (N_8628,N_7092,N_7268);
nor U8629 (N_8629,N_6062,N_7331);
or U8630 (N_8630,N_6193,N_5628);
nor U8631 (N_8631,N_6633,N_5482);
xor U8632 (N_8632,N_6058,N_6838);
nor U8633 (N_8633,N_7238,N_6402);
or U8634 (N_8634,N_5825,N_6228);
and U8635 (N_8635,N_6278,N_5025);
xnor U8636 (N_8636,N_5684,N_5938);
nand U8637 (N_8637,N_7076,N_6990);
xor U8638 (N_8638,N_6823,N_5768);
and U8639 (N_8639,N_6996,N_5206);
or U8640 (N_8640,N_5533,N_5241);
nor U8641 (N_8641,N_6245,N_5295);
and U8642 (N_8642,N_6222,N_6460);
nand U8643 (N_8643,N_7041,N_7203);
and U8644 (N_8644,N_5592,N_6587);
nand U8645 (N_8645,N_5150,N_5414);
or U8646 (N_8646,N_5182,N_5762);
nand U8647 (N_8647,N_6421,N_6875);
and U8648 (N_8648,N_7153,N_5755);
nand U8649 (N_8649,N_5569,N_6788);
xnor U8650 (N_8650,N_5259,N_6602);
and U8651 (N_8651,N_5047,N_6198);
and U8652 (N_8652,N_7467,N_6110);
nor U8653 (N_8653,N_7073,N_6973);
xor U8654 (N_8654,N_5585,N_6350);
nor U8655 (N_8655,N_5764,N_5633);
xor U8656 (N_8656,N_6316,N_5876);
nor U8657 (N_8657,N_5233,N_5481);
and U8658 (N_8658,N_6544,N_5782);
or U8659 (N_8659,N_5276,N_6084);
and U8660 (N_8660,N_5951,N_7397);
nor U8661 (N_8661,N_5179,N_5790);
xor U8662 (N_8662,N_7109,N_6995);
or U8663 (N_8663,N_6032,N_6851);
nor U8664 (N_8664,N_6016,N_6324);
nor U8665 (N_8665,N_5198,N_7237);
xor U8666 (N_8666,N_5485,N_5965);
nand U8667 (N_8667,N_7031,N_5720);
and U8668 (N_8668,N_7302,N_7058);
or U8669 (N_8669,N_5427,N_7265);
nand U8670 (N_8670,N_6560,N_6723);
xnor U8671 (N_8671,N_6901,N_6343);
and U8672 (N_8672,N_6979,N_5862);
xor U8673 (N_8673,N_7231,N_5579);
nor U8674 (N_8674,N_6773,N_6886);
xnor U8675 (N_8675,N_6697,N_5699);
or U8676 (N_8676,N_6188,N_5615);
xnor U8677 (N_8677,N_5110,N_7021);
or U8678 (N_8678,N_7448,N_6305);
nand U8679 (N_8679,N_5519,N_6889);
and U8680 (N_8680,N_6135,N_5133);
and U8681 (N_8681,N_6903,N_5872);
nand U8682 (N_8682,N_5840,N_6960);
or U8683 (N_8683,N_5899,N_7438);
or U8684 (N_8684,N_6923,N_5883);
or U8685 (N_8685,N_6711,N_6260);
and U8686 (N_8686,N_6009,N_5028);
nand U8687 (N_8687,N_6048,N_7158);
nor U8688 (N_8688,N_5078,N_5101);
nand U8689 (N_8689,N_7495,N_5453);
nand U8690 (N_8690,N_7382,N_5809);
nand U8691 (N_8691,N_7230,N_7202);
and U8692 (N_8692,N_7159,N_6627);
or U8693 (N_8693,N_6328,N_7487);
or U8694 (N_8694,N_6615,N_5647);
or U8695 (N_8695,N_6153,N_5708);
nand U8696 (N_8696,N_5673,N_5185);
xor U8697 (N_8697,N_5851,N_5561);
and U8698 (N_8698,N_6733,N_5452);
or U8699 (N_8699,N_6997,N_6130);
nand U8700 (N_8700,N_5053,N_6757);
xnor U8701 (N_8701,N_5310,N_6971);
nor U8702 (N_8702,N_5660,N_7192);
nand U8703 (N_8703,N_7097,N_5675);
nand U8704 (N_8704,N_6966,N_6843);
or U8705 (N_8705,N_6527,N_6689);
nor U8706 (N_8706,N_6192,N_5765);
and U8707 (N_8707,N_5281,N_5147);
nand U8708 (N_8708,N_7425,N_5701);
nand U8709 (N_8709,N_5716,N_5945);
nor U8710 (N_8710,N_5040,N_5468);
xor U8711 (N_8711,N_5788,N_6746);
nor U8712 (N_8712,N_5391,N_6292);
or U8713 (N_8713,N_6334,N_5222);
xor U8714 (N_8714,N_7337,N_7181);
nor U8715 (N_8715,N_7008,N_5336);
xor U8716 (N_8716,N_7077,N_6991);
or U8717 (N_8717,N_6230,N_5424);
or U8718 (N_8718,N_7417,N_6041);
or U8719 (N_8719,N_5265,N_6586);
or U8720 (N_8720,N_5959,N_5891);
or U8721 (N_8721,N_7075,N_7311);
or U8722 (N_8722,N_7165,N_6829);
and U8723 (N_8723,N_6682,N_6661);
and U8724 (N_8724,N_6988,N_6103);
nand U8725 (N_8725,N_5789,N_6949);
nor U8726 (N_8726,N_5454,N_6002);
or U8727 (N_8727,N_6391,N_6828);
nand U8728 (N_8728,N_6881,N_6186);
nor U8729 (N_8729,N_6525,N_5023);
xnor U8730 (N_8730,N_6864,N_5278);
xor U8731 (N_8731,N_7366,N_5307);
or U8732 (N_8732,N_7362,N_6801);
xor U8733 (N_8733,N_5376,N_6467);
nor U8734 (N_8734,N_6172,N_5500);
xor U8735 (N_8735,N_5941,N_5055);
nor U8736 (N_8736,N_5280,N_5654);
nor U8737 (N_8737,N_5710,N_6436);
xor U8738 (N_8738,N_5772,N_6538);
or U8739 (N_8739,N_5857,N_7412);
nor U8740 (N_8740,N_5440,N_5741);
or U8741 (N_8741,N_5642,N_5791);
and U8742 (N_8742,N_5065,N_5334);
and U8743 (N_8743,N_5609,N_6915);
nand U8744 (N_8744,N_6043,N_6745);
or U8745 (N_8745,N_7063,N_6021);
nor U8746 (N_8746,N_5696,N_7491);
xor U8747 (N_8747,N_6955,N_6242);
nor U8748 (N_8748,N_5168,N_6599);
nand U8749 (N_8749,N_5388,N_5258);
xnor U8750 (N_8750,N_6937,N_6904);
nor U8751 (N_8751,N_6141,N_7405);
nor U8752 (N_8752,N_5199,N_6492);
and U8753 (N_8753,N_6076,N_5527);
nand U8754 (N_8754,N_6803,N_5550);
nand U8755 (N_8755,N_5253,N_6870);
xor U8756 (N_8756,N_6161,N_6932);
and U8757 (N_8757,N_5768,N_6806);
nor U8758 (N_8758,N_5560,N_6006);
and U8759 (N_8759,N_5972,N_7440);
or U8760 (N_8760,N_6193,N_5169);
or U8761 (N_8761,N_7052,N_5954);
or U8762 (N_8762,N_7188,N_6868);
or U8763 (N_8763,N_6782,N_6840);
nor U8764 (N_8764,N_6224,N_5377);
and U8765 (N_8765,N_6275,N_7370);
nand U8766 (N_8766,N_7114,N_6413);
and U8767 (N_8767,N_5810,N_5696);
xnor U8768 (N_8768,N_5735,N_5028);
xnor U8769 (N_8769,N_6759,N_7396);
xor U8770 (N_8770,N_5860,N_6509);
or U8771 (N_8771,N_5149,N_5527);
xnor U8772 (N_8772,N_5249,N_5491);
nor U8773 (N_8773,N_6512,N_6851);
and U8774 (N_8774,N_5674,N_6468);
xor U8775 (N_8775,N_6003,N_7074);
and U8776 (N_8776,N_5767,N_6374);
xor U8777 (N_8777,N_6836,N_6629);
nand U8778 (N_8778,N_7433,N_5956);
nand U8779 (N_8779,N_7192,N_5927);
nand U8780 (N_8780,N_6035,N_5729);
nor U8781 (N_8781,N_5635,N_7417);
nor U8782 (N_8782,N_5541,N_6068);
xor U8783 (N_8783,N_7409,N_5338);
nor U8784 (N_8784,N_7248,N_6070);
and U8785 (N_8785,N_6722,N_7076);
and U8786 (N_8786,N_6072,N_6725);
or U8787 (N_8787,N_6066,N_5790);
and U8788 (N_8788,N_6716,N_5139);
nand U8789 (N_8789,N_6561,N_6589);
nor U8790 (N_8790,N_5035,N_6410);
or U8791 (N_8791,N_6968,N_7272);
nor U8792 (N_8792,N_5292,N_6884);
and U8793 (N_8793,N_6619,N_5813);
nor U8794 (N_8794,N_6337,N_6658);
and U8795 (N_8795,N_7094,N_5524);
xor U8796 (N_8796,N_5053,N_6660);
and U8797 (N_8797,N_5548,N_6994);
nand U8798 (N_8798,N_5050,N_5283);
or U8799 (N_8799,N_5559,N_7478);
and U8800 (N_8800,N_7398,N_5612);
nand U8801 (N_8801,N_7420,N_6172);
xnor U8802 (N_8802,N_6536,N_6026);
or U8803 (N_8803,N_7478,N_7092);
and U8804 (N_8804,N_5064,N_5042);
xor U8805 (N_8805,N_5653,N_5435);
xor U8806 (N_8806,N_6332,N_7347);
nor U8807 (N_8807,N_7346,N_5081);
or U8808 (N_8808,N_5695,N_6222);
xnor U8809 (N_8809,N_7488,N_6851);
nor U8810 (N_8810,N_7355,N_5627);
or U8811 (N_8811,N_5769,N_5112);
and U8812 (N_8812,N_6736,N_6158);
or U8813 (N_8813,N_6830,N_5545);
nand U8814 (N_8814,N_5180,N_7487);
nand U8815 (N_8815,N_6555,N_7064);
nor U8816 (N_8816,N_5534,N_5564);
nor U8817 (N_8817,N_7481,N_7128);
nor U8818 (N_8818,N_7232,N_5619);
nand U8819 (N_8819,N_5202,N_6960);
xnor U8820 (N_8820,N_6367,N_5231);
or U8821 (N_8821,N_7192,N_7313);
or U8822 (N_8822,N_5331,N_5450);
xor U8823 (N_8823,N_6672,N_7373);
nor U8824 (N_8824,N_6407,N_7313);
and U8825 (N_8825,N_5317,N_6175);
and U8826 (N_8826,N_5373,N_5464);
nand U8827 (N_8827,N_5524,N_7277);
nor U8828 (N_8828,N_5737,N_5339);
xor U8829 (N_8829,N_6115,N_6692);
or U8830 (N_8830,N_6704,N_5790);
and U8831 (N_8831,N_5533,N_7414);
and U8832 (N_8832,N_5001,N_6395);
nor U8833 (N_8833,N_6557,N_7167);
nand U8834 (N_8834,N_5487,N_6136);
nor U8835 (N_8835,N_5456,N_5949);
xnor U8836 (N_8836,N_5696,N_6692);
or U8837 (N_8837,N_6890,N_7020);
and U8838 (N_8838,N_6996,N_7060);
nand U8839 (N_8839,N_7252,N_5083);
or U8840 (N_8840,N_6377,N_5346);
or U8841 (N_8841,N_5169,N_6518);
or U8842 (N_8842,N_5356,N_7402);
nor U8843 (N_8843,N_7458,N_5835);
or U8844 (N_8844,N_7059,N_5592);
or U8845 (N_8845,N_6349,N_7464);
xnor U8846 (N_8846,N_7383,N_5582);
or U8847 (N_8847,N_5923,N_5731);
or U8848 (N_8848,N_5452,N_7386);
xor U8849 (N_8849,N_5811,N_5189);
nand U8850 (N_8850,N_7355,N_7277);
or U8851 (N_8851,N_5867,N_6823);
and U8852 (N_8852,N_5457,N_5273);
nor U8853 (N_8853,N_7102,N_5586);
or U8854 (N_8854,N_5733,N_6248);
nand U8855 (N_8855,N_6300,N_5345);
and U8856 (N_8856,N_6267,N_6145);
or U8857 (N_8857,N_7205,N_7252);
and U8858 (N_8858,N_6106,N_5356);
or U8859 (N_8859,N_5313,N_5418);
nand U8860 (N_8860,N_6905,N_6025);
nor U8861 (N_8861,N_6830,N_6417);
nor U8862 (N_8862,N_5689,N_6740);
xnor U8863 (N_8863,N_5197,N_5049);
and U8864 (N_8864,N_6112,N_7226);
and U8865 (N_8865,N_6940,N_6295);
xnor U8866 (N_8866,N_6968,N_5203);
or U8867 (N_8867,N_6445,N_5725);
and U8868 (N_8868,N_6512,N_7470);
or U8869 (N_8869,N_5357,N_5825);
or U8870 (N_8870,N_5266,N_5034);
or U8871 (N_8871,N_6426,N_5467);
nand U8872 (N_8872,N_5678,N_6188);
nand U8873 (N_8873,N_5490,N_5272);
xnor U8874 (N_8874,N_6836,N_5076);
or U8875 (N_8875,N_6180,N_7357);
nor U8876 (N_8876,N_7082,N_7394);
or U8877 (N_8877,N_5270,N_7322);
and U8878 (N_8878,N_6782,N_5990);
nor U8879 (N_8879,N_5327,N_5344);
and U8880 (N_8880,N_5188,N_6763);
or U8881 (N_8881,N_6482,N_5115);
and U8882 (N_8882,N_6724,N_6433);
nor U8883 (N_8883,N_5410,N_5075);
nand U8884 (N_8884,N_6296,N_5159);
or U8885 (N_8885,N_5828,N_6485);
nand U8886 (N_8886,N_6336,N_6981);
xnor U8887 (N_8887,N_5796,N_6790);
xor U8888 (N_8888,N_5155,N_6000);
xnor U8889 (N_8889,N_5181,N_6539);
and U8890 (N_8890,N_7256,N_7350);
xor U8891 (N_8891,N_6573,N_5369);
xor U8892 (N_8892,N_6841,N_5632);
xnor U8893 (N_8893,N_6882,N_5548);
and U8894 (N_8894,N_6233,N_5171);
nor U8895 (N_8895,N_6611,N_5587);
xnor U8896 (N_8896,N_6698,N_6548);
nor U8897 (N_8897,N_6442,N_6120);
nand U8898 (N_8898,N_6475,N_6345);
or U8899 (N_8899,N_5862,N_6452);
nand U8900 (N_8900,N_6880,N_6186);
or U8901 (N_8901,N_5346,N_5972);
nand U8902 (N_8902,N_5646,N_6305);
or U8903 (N_8903,N_5012,N_6564);
and U8904 (N_8904,N_6619,N_5632);
xnor U8905 (N_8905,N_7435,N_6446);
and U8906 (N_8906,N_6494,N_6884);
nor U8907 (N_8907,N_7268,N_6162);
and U8908 (N_8908,N_6455,N_6501);
nor U8909 (N_8909,N_6449,N_6488);
and U8910 (N_8910,N_5718,N_6296);
nand U8911 (N_8911,N_7202,N_7136);
nor U8912 (N_8912,N_6644,N_7107);
and U8913 (N_8913,N_5630,N_5822);
xor U8914 (N_8914,N_5321,N_5487);
and U8915 (N_8915,N_7344,N_6133);
and U8916 (N_8916,N_6188,N_5004);
nor U8917 (N_8917,N_5510,N_6346);
nor U8918 (N_8918,N_7057,N_6773);
or U8919 (N_8919,N_7365,N_6425);
nand U8920 (N_8920,N_6166,N_6422);
and U8921 (N_8921,N_5143,N_5999);
or U8922 (N_8922,N_6730,N_5028);
xor U8923 (N_8923,N_5220,N_6080);
or U8924 (N_8924,N_5343,N_7268);
or U8925 (N_8925,N_7020,N_6953);
or U8926 (N_8926,N_6592,N_5093);
nand U8927 (N_8927,N_5676,N_6519);
nor U8928 (N_8928,N_6642,N_5612);
or U8929 (N_8929,N_6171,N_6095);
nand U8930 (N_8930,N_5254,N_5444);
and U8931 (N_8931,N_5307,N_6852);
and U8932 (N_8932,N_5514,N_5762);
nor U8933 (N_8933,N_7209,N_5594);
nor U8934 (N_8934,N_5084,N_7286);
and U8935 (N_8935,N_5944,N_6799);
nand U8936 (N_8936,N_5751,N_6748);
or U8937 (N_8937,N_7361,N_5010);
nor U8938 (N_8938,N_6587,N_7268);
nand U8939 (N_8939,N_5409,N_5735);
nor U8940 (N_8940,N_6960,N_5317);
and U8941 (N_8941,N_6771,N_5602);
nand U8942 (N_8942,N_5171,N_6388);
and U8943 (N_8943,N_5818,N_5916);
or U8944 (N_8944,N_5506,N_6446);
nand U8945 (N_8945,N_6852,N_6243);
nand U8946 (N_8946,N_7312,N_5512);
or U8947 (N_8947,N_6552,N_6291);
nand U8948 (N_8948,N_6989,N_6300);
nand U8949 (N_8949,N_6913,N_6832);
xnor U8950 (N_8950,N_6659,N_7328);
or U8951 (N_8951,N_6267,N_5943);
nand U8952 (N_8952,N_6639,N_5879);
nand U8953 (N_8953,N_5323,N_6120);
nand U8954 (N_8954,N_7444,N_6004);
or U8955 (N_8955,N_7274,N_5806);
xor U8956 (N_8956,N_6068,N_5288);
nor U8957 (N_8957,N_5743,N_5158);
xor U8958 (N_8958,N_6305,N_6814);
and U8959 (N_8959,N_5799,N_7297);
and U8960 (N_8960,N_7424,N_5341);
and U8961 (N_8961,N_5480,N_5763);
xnor U8962 (N_8962,N_5686,N_5289);
xnor U8963 (N_8963,N_5968,N_5583);
nor U8964 (N_8964,N_5780,N_5025);
nor U8965 (N_8965,N_5351,N_6840);
xnor U8966 (N_8966,N_6897,N_6929);
or U8967 (N_8967,N_7365,N_6085);
or U8968 (N_8968,N_5596,N_5166);
and U8969 (N_8969,N_6648,N_5485);
nor U8970 (N_8970,N_7128,N_5034);
or U8971 (N_8971,N_5482,N_5300);
xnor U8972 (N_8972,N_5050,N_6580);
nor U8973 (N_8973,N_6782,N_6438);
and U8974 (N_8974,N_6454,N_6157);
and U8975 (N_8975,N_6105,N_6635);
nor U8976 (N_8976,N_7133,N_5846);
xor U8977 (N_8977,N_6488,N_5874);
or U8978 (N_8978,N_7304,N_7352);
xnor U8979 (N_8979,N_5002,N_7152);
and U8980 (N_8980,N_5813,N_7415);
xor U8981 (N_8981,N_5627,N_5151);
xnor U8982 (N_8982,N_5974,N_7263);
nand U8983 (N_8983,N_7402,N_6584);
nand U8984 (N_8984,N_6863,N_5834);
xnor U8985 (N_8985,N_6718,N_6223);
and U8986 (N_8986,N_6898,N_6427);
nand U8987 (N_8987,N_6014,N_7455);
or U8988 (N_8988,N_7243,N_5174);
nor U8989 (N_8989,N_7250,N_6023);
xnor U8990 (N_8990,N_5454,N_7004);
xnor U8991 (N_8991,N_7382,N_6864);
nor U8992 (N_8992,N_6561,N_5265);
nor U8993 (N_8993,N_6253,N_6847);
nand U8994 (N_8994,N_6133,N_7308);
xor U8995 (N_8995,N_6711,N_6097);
nand U8996 (N_8996,N_6144,N_6806);
xnor U8997 (N_8997,N_7397,N_5516);
nor U8998 (N_8998,N_5113,N_7462);
nand U8999 (N_8999,N_6679,N_5102);
and U9000 (N_9000,N_6622,N_6517);
and U9001 (N_9001,N_5711,N_6312);
nor U9002 (N_9002,N_5833,N_5997);
nand U9003 (N_9003,N_5622,N_6261);
nor U9004 (N_9004,N_6380,N_5269);
nor U9005 (N_9005,N_5357,N_5826);
xor U9006 (N_9006,N_7494,N_6929);
nand U9007 (N_9007,N_6556,N_6033);
nor U9008 (N_9008,N_5708,N_7397);
or U9009 (N_9009,N_6227,N_6782);
and U9010 (N_9010,N_6439,N_7484);
nor U9011 (N_9011,N_6320,N_6250);
and U9012 (N_9012,N_7195,N_6829);
or U9013 (N_9013,N_5532,N_5605);
or U9014 (N_9014,N_5288,N_7032);
and U9015 (N_9015,N_6071,N_6643);
nand U9016 (N_9016,N_5758,N_5414);
nand U9017 (N_9017,N_7023,N_5781);
xnor U9018 (N_9018,N_7188,N_6445);
nand U9019 (N_9019,N_5951,N_5497);
and U9020 (N_9020,N_7264,N_6514);
or U9021 (N_9021,N_6710,N_5374);
or U9022 (N_9022,N_7080,N_5655);
or U9023 (N_9023,N_5792,N_6072);
and U9024 (N_9024,N_6681,N_5278);
and U9025 (N_9025,N_7226,N_6510);
nor U9026 (N_9026,N_7376,N_5973);
or U9027 (N_9027,N_6943,N_6634);
nor U9028 (N_9028,N_6026,N_5510);
nand U9029 (N_9029,N_7301,N_7446);
or U9030 (N_9030,N_6393,N_6801);
and U9031 (N_9031,N_6841,N_6177);
nor U9032 (N_9032,N_7192,N_7449);
nor U9033 (N_9033,N_5517,N_5671);
or U9034 (N_9034,N_5945,N_7090);
and U9035 (N_9035,N_5186,N_5524);
nor U9036 (N_9036,N_5938,N_6139);
nand U9037 (N_9037,N_6985,N_5386);
or U9038 (N_9038,N_5274,N_6757);
xor U9039 (N_9039,N_6601,N_5301);
and U9040 (N_9040,N_5542,N_5965);
nor U9041 (N_9041,N_5108,N_6210);
or U9042 (N_9042,N_7440,N_6664);
or U9043 (N_9043,N_6933,N_6104);
xor U9044 (N_9044,N_5611,N_6970);
nor U9045 (N_9045,N_7486,N_6801);
nor U9046 (N_9046,N_7300,N_6223);
xnor U9047 (N_9047,N_7197,N_6060);
xor U9048 (N_9048,N_5238,N_7421);
or U9049 (N_9049,N_6266,N_6096);
xor U9050 (N_9050,N_7041,N_5007);
nand U9051 (N_9051,N_6849,N_5676);
xnor U9052 (N_9052,N_5195,N_6698);
nand U9053 (N_9053,N_5706,N_7198);
nand U9054 (N_9054,N_5796,N_5432);
xnor U9055 (N_9055,N_5221,N_7318);
nand U9056 (N_9056,N_5331,N_6480);
nor U9057 (N_9057,N_7098,N_6501);
and U9058 (N_9058,N_6578,N_6399);
nand U9059 (N_9059,N_7343,N_6349);
nor U9060 (N_9060,N_5112,N_6077);
nand U9061 (N_9061,N_5828,N_6271);
or U9062 (N_9062,N_5245,N_5488);
and U9063 (N_9063,N_5904,N_5353);
or U9064 (N_9064,N_7034,N_6865);
and U9065 (N_9065,N_5990,N_5984);
or U9066 (N_9066,N_7214,N_6697);
nand U9067 (N_9067,N_7386,N_5117);
nor U9068 (N_9068,N_5536,N_6208);
nand U9069 (N_9069,N_7038,N_5575);
and U9070 (N_9070,N_7243,N_7317);
nor U9071 (N_9071,N_6010,N_6687);
or U9072 (N_9072,N_7491,N_7495);
or U9073 (N_9073,N_6297,N_6405);
nor U9074 (N_9074,N_5418,N_7273);
and U9075 (N_9075,N_6882,N_6776);
or U9076 (N_9076,N_5480,N_6982);
nand U9077 (N_9077,N_6780,N_5250);
xor U9078 (N_9078,N_6341,N_7132);
xor U9079 (N_9079,N_6302,N_5653);
xnor U9080 (N_9080,N_5237,N_6154);
nand U9081 (N_9081,N_7385,N_6494);
or U9082 (N_9082,N_6924,N_5181);
xor U9083 (N_9083,N_6501,N_5029);
nand U9084 (N_9084,N_6402,N_5464);
nand U9085 (N_9085,N_5590,N_6629);
xnor U9086 (N_9086,N_6589,N_6799);
xor U9087 (N_9087,N_5077,N_6080);
or U9088 (N_9088,N_6001,N_7111);
or U9089 (N_9089,N_6017,N_6507);
xnor U9090 (N_9090,N_7428,N_7244);
or U9091 (N_9091,N_6770,N_6901);
xor U9092 (N_9092,N_6423,N_5758);
and U9093 (N_9093,N_5418,N_7294);
nor U9094 (N_9094,N_5802,N_5820);
and U9095 (N_9095,N_6000,N_6362);
or U9096 (N_9096,N_5411,N_5649);
nor U9097 (N_9097,N_6185,N_6885);
nand U9098 (N_9098,N_6574,N_5764);
nand U9099 (N_9099,N_6073,N_6021);
xnor U9100 (N_9100,N_6924,N_6149);
and U9101 (N_9101,N_6540,N_5978);
nand U9102 (N_9102,N_6501,N_6772);
or U9103 (N_9103,N_7134,N_5496);
nor U9104 (N_9104,N_5059,N_6676);
nor U9105 (N_9105,N_5111,N_6153);
nand U9106 (N_9106,N_5188,N_6489);
nor U9107 (N_9107,N_5922,N_5057);
xor U9108 (N_9108,N_6815,N_5452);
nand U9109 (N_9109,N_5670,N_6232);
nand U9110 (N_9110,N_6404,N_5277);
nor U9111 (N_9111,N_5556,N_6987);
nor U9112 (N_9112,N_6195,N_6350);
nor U9113 (N_9113,N_5385,N_7370);
xor U9114 (N_9114,N_6758,N_6672);
and U9115 (N_9115,N_6869,N_5535);
or U9116 (N_9116,N_5781,N_5615);
and U9117 (N_9117,N_7000,N_7431);
xnor U9118 (N_9118,N_6319,N_5574);
nand U9119 (N_9119,N_6839,N_6876);
nand U9120 (N_9120,N_6670,N_7036);
nand U9121 (N_9121,N_5434,N_6896);
nor U9122 (N_9122,N_5241,N_6312);
nand U9123 (N_9123,N_5796,N_6895);
or U9124 (N_9124,N_7376,N_6648);
nand U9125 (N_9125,N_7306,N_7399);
nand U9126 (N_9126,N_6370,N_6411);
or U9127 (N_9127,N_5212,N_5905);
nand U9128 (N_9128,N_6316,N_6917);
nor U9129 (N_9129,N_6651,N_6043);
xor U9130 (N_9130,N_5391,N_7028);
xnor U9131 (N_9131,N_6081,N_6548);
xor U9132 (N_9132,N_5899,N_6090);
and U9133 (N_9133,N_5748,N_5474);
nor U9134 (N_9134,N_6079,N_7216);
xor U9135 (N_9135,N_5456,N_5977);
or U9136 (N_9136,N_7456,N_6599);
nor U9137 (N_9137,N_5395,N_5574);
nor U9138 (N_9138,N_7072,N_6517);
and U9139 (N_9139,N_5969,N_5897);
nand U9140 (N_9140,N_5059,N_6346);
nand U9141 (N_9141,N_7205,N_5891);
or U9142 (N_9142,N_7415,N_5702);
nor U9143 (N_9143,N_6157,N_6395);
nor U9144 (N_9144,N_6132,N_6366);
or U9145 (N_9145,N_7267,N_6054);
and U9146 (N_9146,N_6591,N_5899);
xor U9147 (N_9147,N_7490,N_7149);
or U9148 (N_9148,N_6742,N_6883);
and U9149 (N_9149,N_6467,N_6954);
nand U9150 (N_9150,N_5779,N_7171);
nand U9151 (N_9151,N_5388,N_6738);
and U9152 (N_9152,N_6810,N_6439);
nand U9153 (N_9153,N_7128,N_6196);
or U9154 (N_9154,N_5689,N_5255);
nand U9155 (N_9155,N_7221,N_5100);
and U9156 (N_9156,N_5758,N_5307);
and U9157 (N_9157,N_6251,N_5921);
nor U9158 (N_9158,N_6353,N_6712);
nor U9159 (N_9159,N_6992,N_6259);
xor U9160 (N_9160,N_7346,N_7264);
nand U9161 (N_9161,N_6740,N_5893);
and U9162 (N_9162,N_7195,N_5248);
nand U9163 (N_9163,N_5290,N_6288);
or U9164 (N_9164,N_6202,N_6112);
nor U9165 (N_9165,N_6415,N_6874);
or U9166 (N_9166,N_6678,N_6476);
xor U9167 (N_9167,N_5306,N_5784);
and U9168 (N_9168,N_6783,N_6552);
nor U9169 (N_9169,N_5419,N_7439);
nor U9170 (N_9170,N_7169,N_6109);
nand U9171 (N_9171,N_5990,N_6386);
or U9172 (N_9172,N_6962,N_5715);
xnor U9173 (N_9173,N_7060,N_6263);
or U9174 (N_9174,N_7038,N_5510);
and U9175 (N_9175,N_6802,N_5973);
xor U9176 (N_9176,N_6953,N_6570);
nand U9177 (N_9177,N_5037,N_5982);
nor U9178 (N_9178,N_5792,N_6939);
xor U9179 (N_9179,N_6990,N_6064);
nand U9180 (N_9180,N_5010,N_6628);
nor U9181 (N_9181,N_7111,N_6587);
xor U9182 (N_9182,N_6646,N_5046);
nand U9183 (N_9183,N_6583,N_6716);
and U9184 (N_9184,N_6664,N_7495);
or U9185 (N_9185,N_5478,N_6435);
or U9186 (N_9186,N_7374,N_7004);
or U9187 (N_9187,N_6394,N_6396);
or U9188 (N_9188,N_6413,N_5012);
nand U9189 (N_9189,N_5198,N_5036);
or U9190 (N_9190,N_6674,N_6446);
nand U9191 (N_9191,N_7208,N_5791);
and U9192 (N_9192,N_6211,N_5914);
xor U9193 (N_9193,N_6567,N_5617);
nand U9194 (N_9194,N_7488,N_6252);
or U9195 (N_9195,N_6551,N_6850);
nor U9196 (N_9196,N_6210,N_7462);
xnor U9197 (N_9197,N_5440,N_7383);
xnor U9198 (N_9198,N_5099,N_7108);
or U9199 (N_9199,N_7269,N_6244);
or U9200 (N_9200,N_7194,N_5049);
xnor U9201 (N_9201,N_6706,N_5193);
nand U9202 (N_9202,N_6374,N_7393);
nand U9203 (N_9203,N_7255,N_6791);
and U9204 (N_9204,N_6187,N_6021);
nor U9205 (N_9205,N_5477,N_7094);
and U9206 (N_9206,N_6342,N_5207);
and U9207 (N_9207,N_7329,N_6564);
and U9208 (N_9208,N_6393,N_6137);
xnor U9209 (N_9209,N_7255,N_6703);
and U9210 (N_9210,N_6321,N_7181);
nor U9211 (N_9211,N_7026,N_7135);
and U9212 (N_9212,N_5767,N_5913);
nand U9213 (N_9213,N_5956,N_5858);
and U9214 (N_9214,N_6245,N_7137);
nand U9215 (N_9215,N_5995,N_5446);
or U9216 (N_9216,N_6861,N_6072);
nand U9217 (N_9217,N_5991,N_7394);
nand U9218 (N_9218,N_7304,N_6863);
or U9219 (N_9219,N_5042,N_5494);
and U9220 (N_9220,N_6452,N_6870);
and U9221 (N_9221,N_6776,N_6089);
xnor U9222 (N_9222,N_7495,N_7251);
and U9223 (N_9223,N_5401,N_5485);
or U9224 (N_9224,N_5216,N_5668);
and U9225 (N_9225,N_5627,N_7034);
and U9226 (N_9226,N_7427,N_5257);
or U9227 (N_9227,N_7413,N_7075);
and U9228 (N_9228,N_5367,N_6111);
nand U9229 (N_9229,N_5194,N_6337);
xor U9230 (N_9230,N_7297,N_6264);
or U9231 (N_9231,N_6763,N_5318);
or U9232 (N_9232,N_6417,N_5707);
and U9233 (N_9233,N_6114,N_6490);
and U9234 (N_9234,N_7103,N_5539);
and U9235 (N_9235,N_6750,N_7399);
nor U9236 (N_9236,N_5619,N_6401);
xor U9237 (N_9237,N_6860,N_6253);
nor U9238 (N_9238,N_5491,N_5766);
or U9239 (N_9239,N_6254,N_6229);
xor U9240 (N_9240,N_7356,N_6583);
nor U9241 (N_9241,N_5987,N_6416);
nand U9242 (N_9242,N_5452,N_5926);
or U9243 (N_9243,N_5304,N_7279);
nand U9244 (N_9244,N_5179,N_6269);
xnor U9245 (N_9245,N_6517,N_5031);
xor U9246 (N_9246,N_7406,N_5863);
or U9247 (N_9247,N_5156,N_7243);
and U9248 (N_9248,N_7044,N_5145);
nand U9249 (N_9249,N_6733,N_6720);
and U9250 (N_9250,N_6152,N_5263);
and U9251 (N_9251,N_5529,N_7405);
or U9252 (N_9252,N_6728,N_6372);
xnor U9253 (N_9253,N_5833,N_5877);
or U9254 (N_9254,N_5239,N_5842);
nand U9255 (N_9255,N_6640,N_7146);
nor U9256 (N_9256,N_5433,N_7240);
and U9257 (N_9257,N_6711,N_6471);
nand U9258 (N_9258,N_6438,N_5062);
xor U9259 (N_9259,N_7192,N_6751);
and U9260 (N_9260,N_6824,N_5705);
or U9261 (N_9261,N_5836,N_6097);
xor U9262 (N_9262,N_6958,N_6708);
nand U9263 (N_9263,N_6939,N_7112);
xor U9264 (N_9264,N_5157,N_5186);
xor U9265 (N_9265,N_6579,N_7045);
nand U9266 (N_9266,N_6901,N_5466);
and U9267 (N_9267,N_6866,N_6507);
nand U9268 (N_9268,N_6712,N_6109);
xnor U9269 (N_9269,N_5240,N_7243);
and U9270 (N_9270,N_7165,N_5499);
and U9271 (N_9271,N_6448,N_7476);
or U9272 (N_9272,N_6154,N_5953);
nor U9273 (N_9273,N_6991,N_5401);
nor U9274 (N_9274,N_6751,N_6739);
and U9275 (N_9275,N_6358,N_6049);
or U9276 (N_9276,N_6596,N_7429);
nor U9277 (N_9277,N_6269,N_5706);
or U9278 (N_9278,N_5000,N_6273);
or U9279 (N_9279,N_5920,N_6541);
nor U9280 (N_9280,N_5005,N_5008);
nor U9281 (N_9281,N_6967,N_5908);
or U9282 (N_9282,N_7199,N_7099);
xor U9283 (N_9283,N_5213,N_6943);
xnor U9284 (N_9284,N_6190,N_7094);
xnor U9285 (N_9285,N_5229,N_7450);
and U9286 (N_9286,N_6044,N_6076);
or U9287 (N_9287,N_7179,N_5960);
or U9288 (N_9288,N_6095,N_7143);
or U9289 (N_9289,N_5444,N_7320);
and U9290 (N_9290,N_6086,N_5313);
xor U9291 (N_9291,N_5477,N_6085);
nand U9292 (N_9292,N_6798,N_6691);
nand U9293 (N_9293,N_5936,N_7481);
or U9294 (N_9294,N_5253,N_6110);
or U9295 (N_9295,N_5090,N_5509);
nor U9296 (N_9296,N_5862,N_6717);
xnor U9297 (N_9297,N_7236,N_5315);
nor U9298 (N_9298,N_5218,N_6227);
xnor U9299 (N_9299,N_5390,N_6881);
nand U9300 (N_9300,N_6081,N_6730);
xnor U9301 (N_9301,N_6708,N_5291);
or U9302 (N_9302,N_6183,N_6480);
xor U9303 (N_9303,N_7311,N_6781);
nand U9304 (N_9304,N_5764,N_7297);
nand U9305 (N_9305,N_5871,N_5364);
nand U9306 (N_9306,N_6761,N_7255);
nor U9307 (N_9307,N_7342,N_5922);
nor U9308 (N_9308,N_5227,N_6467);
and U9309 (N_9309,N_5819,N_5150);
xnor U9310 (N_9310,N_5855,N_6881);
xnor U9311 (N_9311,N_6783,N_5414);
or U9312 (N_9312,N_5048,N_5250);
or U9313 (N_9313,N_7290,N_7315);
and U9314 (N_9314,N_7037,N_6954);
nor U9315 (N_9315,N_6504,N_6426);
and U9316 (N_9316,N_7440,N_6010);
and U9317 (N_9317,N_7238,N_6334);
or U9318 (N_9318,N_6445,N_5160);
and U9319 (N_9319,N_5425,N_5129);
nand U9320 (N_9320,N_6152,N_5958);
or U9321 (N_9321,N_6766,N_5069);
xnor U9322 (N_9322,N_7413,N_6066);
nor U9323 (N_9323,N_6537,N_6094);
nand U9324 (N_9324,N_6244,N_5582);
or U9325 (N_9325,N_5445,N_7320);
and U9326 (N_9326,N_5701,N_5649);
nand U9327 (N_9327,N_5635,N_7019);
and U9328 (N_9328,N_6972,N_5033);
nor U9329 (N_9329,N_5051,N_6236);
xor U9330 (N_9330,N_5342,N_5499);
nor U9331 (N_9331,N_6152,N_5350);
nor U9332 (N_9332,N_6768,N_6443);
nand U9333 (N_9333,N_6759,N_6234);
nor U9334 (N_9334,N_6826,N_5912);
xnor U9335 (N_9335,N_6533,N_5351);
nand U9336 (N_9336,N_7390,N_7255);
nor U9337 (N_9337,N_5339,N_7108);
xor U9338 (N_9338,N_6419,N_5080);
xor U9339 (N_9339,N_6090,N_5991);
xor U9340 (N_9340,N_7442,N_6191);
xor U9341 (N_9341,N_5664,N_5675);
nor U9342 (N_9342,N_6123,N_5557);
nor U9343 (N_9343,N_5511,N_5839);
and U9344 (N_9344,N_6823,N_6770);
nand U9345 (N_9345,N_6253,N_6251);
nand U9346 (N_9346,N_5081,N_6111);
xnor U9347 (N_9347,N_5851,N_5532);
and U9348 (N_9348,N_7042,N_5161);
nor U9349 (N_9349,N_6025,N_5942);
xor U9350 (N_9350,N_6510,N_5867);
xor U9351 (N_9351,N_7460,N_5139);
xor U9352 (N_9352,N_5603,N_6589);
nand U9353 (N_9353,N_5984,N_5437);
or U9354 (N_9354,N_7231,N_5240);
xnor U9355 (N_9355,N_6472,N_6666);
and U9356 (N_9356,N_5578,N_7353);
xor U9357 (N_9357,N_7101,N_6553);
or U9358 (N_9358,N_5379,N_6256);
nor U9359 (N_9359,N_6674,N_6312);
nand U9360 (N_9360,N_7376,N_5617);
nand U9361 (N_9361,N_5663,N_5654);
nor U9362 (N_9362,N_7359,N_6989);
nand U9363 (N_9363,N_6026,N_7428);
xor U9364 (N_9364,N_7165,N_7333);
and U9365 (N_9365,N_6353,N_5982);
or U9366 (N_9366,N_6428,N_5968);
nor U9367 (N_9367,N_6318,N_5436);
nand U9368 (N_9368,N_7392,N_5902);
nand U9369 (N_9369,N_6008,N_5028);
and U9370 (N_9370,N_7386,N_6521);
nor U9371 (N_9371,N_7136,N_5716);
xnor U9372 (N_9372,N_6715,N_7035);
nand U9373 (N_9373,N_6803,N_6783);
nor U9374 (N_9374,N_5360,N_5986);
nand U9375 (N_9375,N_5127,N_7369);
nand U9376 (N_9376,N_6163,N_7488);
nand U9377 (N_9377,N_5219,N_7423);
or U9378 (N_9378,N_7354,N_5085);
nand U9379 (N_9379,N_7310,N_6298);
or U9380 (N_9380,N_6214,N_6377);
nor U9381 (N_9381,N_6656,N_6906);
and U9382 (N_9382,N_7363,N_6302);
nor U9383 (N_9383,N_7419,N_6910);
and U9384 (N_9384,N_6494,N_5854);
nor U9385 (N_9385,N_6318,N_7059);
nor U9386 (N_9386,N_5875,N_5359);
nand U9387 (N_9387,N_6775,N_6442);
nor U9388 (N_9388,N_7183,N_5587);
nand U9389 (N_9389,N_7430,N_5474);
nor U9390 (N_9390,N_5004,N_6882);
nor U9391 (N_9391,N_6275,N_6499);
nand U9392 (N_9392,N_7150,N_5573);
or U9393 (N_9393,N_7091,N_5153);
and U9394 (N_9394,N_5935,N_6673);
nand U9395 (N_9395,N_5076,N_7256);
xnor U9396 (N_9396,N_6676,N_5339);
nor U9397 (N_9397,N_6842,N_5944);
xor U9398 (N_9398,N_5584,N_5136);
nand U9399 (N_9399,N_5104,N_5499);
and U9400 (N_9400,N_5244,N_6508);
or U9401 (N_9401,N_5287,N_5904);
and U9402 (N_9402,N_6622,N_7038);
xor U9403 (N_9403,N_5618,N_5308);
or U9404 (N_9404,N_5100,N_6985);
and U9405 (N_9405,N_6941,N_5584);
xor U9406 (N_9406,N_6693,N_5809);
and U9407 (N_9407,N_5670,N_6393);
and U9408 (N_9408,N_5331,N_6867);
and U9409 (N_9409,N_6327,N_7198);
xnor U9410 (N_9410,N_5316,N_7070);
nor U9411 (N_9411,N_5062,N_7245);
or U9412 (N_9412,N_7046,N_5019);
xor U9413 (N_9413,N_5729,N_6949);
nand U9414 (N_9414,N_6763,N_7464);
nand U9415 (N_9415,N_6765,N_7221);
xor U9416 (N_9416,N_6620,N_5357);
nand U9417 (N_9417,N_6439,N_7454);
nor U9418 (N_9418,N_6501,N_5931);
or U9419 (N_9419,N_7096,N_6813);
nor U9420 (N_9420,N_6878,N_7227);
nor U9421 (N_9421,N_5808,N_6279);
nor U9422 (N_9422,N_6575,N_6061);
and U9423 (N_9423,N_6703,N_7067);
nor U9424 (N_9424,N_5848,N_5787);
nand U9425 (N_9425,N_5867,N_6498);
or U9426 (N_9426,N_6498,N_5259);
nand U9427 (N_9427,N_7400,N_6630);
nor U9428 (N_9428,N_5897,N_5399);
or U9429 (N_9429,N_6717,N_5482);
and U9430 (N_9430,N_6741,N_6527);
nand U9431 (N_9431,N_5122,N_5788);
nor U9432 (N_9432,N_7493,N_5131);
nand U9433 (N_9433,N_5533,N_6578);
or U9434 (N_9434,N_7254,N_7404);
nand U9435 (N_9435,N_7242,N_5316);
and U9436 (N_9436,N_5368,N_5505);
xnor U9437 (N_9437,N_6963,N_7402);
xor U9438 (N_9438,N_5184,N_7208);
or U9439 (N_9439,N_6467,N_6548);
or U9440 (N_9440,N_6318,N_6548);
xnor U9441 (N_9441,N_6498,N_7481);
nand U9442 (N_9442,N_6046,N_6988);
xor U9443 (N_9443,N_6829,N_5708);
xor U9444 (N_9444,N_7387,N_5759);
or U9445 (N_9445,N_5661,N_5328);
nor U9446 (N_9446,N_5203,N_6520);
or U9447 (N_9447,N_6975,N_6176);
nand U9448 (N_9448,N_6018,N_7099);
and U9449 (N_9449,N_6490,N_7042);
nor U9450 (N_9450,N_6519,N_5697);
nand U9451 (N_9451,N_7079,N_5905);
nor U9452 (N_9452,N_6669,N_6211);
nand U9453 (N_9453,N_5449,N_6821);
nand U9454 (N_9454,N_6745,N_6260);
xor U9455 (N_9455,N_7114,N_5203);
xor U9456 (N_9456,N_5250,N_5469);
or U9457 (N_9457,N_6432,N_6509);
nor U9458 (N_9458,N_5939,N_7126);
or U9459 (N_9459,N_7088,N_6915);
nand U9460 (N_9460,N_5349,N_5449);
and U9461 (N_9461,N_5008,N_5527);
and U9462 (N_9462,N_5538,N_6984);
and U9463 (N_9463,N_5084,N_7050);
nand U9464 (N_9464,N_7426,N_7006);
and U9465 (N_9465,N_6430,N_5928);
nor U9466 (N_9466,N_6371,N_7005);
and U9467 (N_9467,N_7260,N_6276);
or U9468 (N_9468,N_5981,N_6036);
xnor U9469 (N_9469,N_7097,N_5197);
and U9470 (N_9470,N_5261,N_6447);
nor U9471 (N_9471,N_6701,N_5490);
and U9472 (N_9472,N_7054,N_5037);
or U9473 (N_9473,N_5917,N_5024);
xor U9474 (N_9474,N_6543,N_6875);
nand U9475 (N_9475,N_5155,N_5379);
and U9476 (N_9476,N_7496,N_5728);
and U9477 (N_9477,N_5401,N_5982);
xor U9478 (N_9478,N_6762,N_5214);
or U9479 (N_9479,N_5878,N_6911);
nand U9480 (N_9480,N_7083,N_6640);
nor U9481 (N_9481,N_7310,N_6222);
nor U9482 (N_9482,N_5765,N_6279);
or U9483 (N_9483,N_7063,N_6614);
nand U9484 (N_9484,N_6920,N_6886);
xnor U9485 (N_9485,N_6842,N_6585);
nor U9486 (N_9486,N_6314,N_6446);
and U9487 (N_9487,N_6357,N_5556);
nand U9488 (N_9488,N_6321,N_7423);
xor U9489 (N_9489,N_5896,N_6331);
and U9490 (N_9490,N_5956,N_6062);
nor U9491 (N_9491,N_6381,N_5929);
and U9492 (N_9492,N_6703,N_6435);
and U9493 (N_9493,N_5064,N_6394);
xor U9494 (N_9494,N_6790,N_6382);
and U9495 (N_9495,N_6273,N_6779);
xor U9496 (N_9496,N_6134,N_6474);
and U9497 (N_9497,N_6074,N_6995);
nor U9498 (N_9498,N_6847,N_7196);
xor U9499 (N_9499,N_7413,N_6389);
xnor U9500 (N_9500,N_7360,N_7290);
nand U9501 (N_9501,N_6862,N_5507);
or U9502 (N_9502,N_5592,N_7457);
nand U9503 (N_9503,N_5262,N_6303);
xnor U9504 (N_9504,N_5904,N_5795);
nor U9505 (N_9505,N_6710,N_7333);
and U9506 (N_9506,N_5606,N_7376);
xnor U9507 (N_9507,N_6781,N_6767);
nor U9508 (N_9508,N_5570,N_5372);
nand U9509 (N_9509,N_5101,N_5448);
or U9510 (N_9510,N_6550,N_7148);
nor U9511 (N_9511,N_6363,N_5052);
nor U9512 (N_9512,N_5426,N_6798);
or U9513 (N_9513,N_5605,N_7213);
nand U9514 (N_9514,N_7124,N_6578);
nor U9515 (N_9515,N_5422,N_6752);
nor U9516 (N_9516,N_6922,N_5844);
or U9517 (N_9517,N_7220,N_5004);
and U9518 (N_9518,N_6454,N_6603);
xor U9519 (N_9519,N_6594,N_6189);
and U9520 (N_9520,N_6151,N_6096);
and U9521 (N_9521,N_5305,N_6728);
or U9522 (N_9522,N_6525,N_7482);
nor U9523 (N_9523,N_5390,N_5113);
or U9524 (N_9524,N_5411,N_7100);
nor U9525 (N_9525,N_7333,N_5335);
nand U9526 (N_9526,N_6730,N_7093);
xor U9527 (N_9527,N_5796,N_6962);
nand U9528 (N_9528,N_7297,N_6282);
or U9529 (N_9529,N_5658,N_6844);
nor U9530 (N_9530,N_6682,N_6314);
and U9531 (N_9531,N_5796,N_6653);
nor U9532 (N_9532,N_6162,N_5703);
nand U9533 (N_9533,N_6468,N_5387);
nand U9534 (N_9534,N_7222,N_7366);
or U9535 (N_9535,N_5411,N_5291);
xor U9536 (N_9536,N_5732,N_6446);
nand U9537 (N_9537,N_6457,N_5655);
or U9538 (N_9538,N_5792,N_7053);
nand U9539 (N_9539,N_6561,N_6842);
and U9540 (N_9540,N_5359,N_5735);
xor U9541 (N_9541,N_6383,N_5038);
or U9542 (N_9542,N_6643,N_5297);
nor U9543 (N_9543,N_5006,N_7088);
nand U9544 (N_9544,N_7081,N_5090);
nand U9545 (N_9545,N_5763,N_5664);
or U9546 (N_9546,N_6569,N_6250);
nand U9547 (N_9547,N_5150,N_6528);
xnor U9548 (N_9548,N_5052,N_6219);
xor U9549 (N_9549,N_6014,N_6938);
xnor U9550 (N_9550,N_5882,N_6098);
and U9551 (N_9551,N_6471,N_5413);
nand U9552 (N_9552,N_5075,N_6277);
nand U9553 (N_9553,N_6185,N_7453);
nor U9554 (N_9554,N_5839,N_5660);
and U9555 (N_9555,N_5542,N_7460);
and U9556 (N_9556,N_5868,N_5007);
or U9557 (N_9557,N_5301,N_7264);
xor U9558 (N_9558,N_5156,N_5110);
and U9559 (N_9559,N_6820,N_6320);
xor U9560 (N_9560,N_6006,N_5274);
xnor U9561 (N_9561,N_6204,N_6790);
nor U9562 (N_9562,N_6630,N_5042);
and U9563 (N_9563,N_5944,N_5763);
or U9564 (N_9564,N_6737,N_5606);
or U9565 (N_9565,N_6463,N_6053);
and U9566 (N_9566,N_6408,N_7402);
or U9567 (N_9567,N_6378,N_6333);
nor U9568 (N_9568,N_6698,N_5284);
nor U9569 (N_9569,N_6036,N_7250);
xnor U9570 (N_9570,N_5002,N_5023);
nand U9571 (N_9571,N_6147,N_5675);
xnor U9572 (N_9572,N_6291,N_6456);
nor U9573 (N_9573,N_5410,N_5800);
or U9574 (N_9574,N_6190,N_6840);
nor U9575 (N_9575,N_6208,N_5106);
and U9576 (N_9576,N_5732,N_5348);
and U9577 (N_9577,N_7143,N_6411);
or U9578 (N_9578,N_6658,N_5626);
xnor U9579 (N_9579,N_7245,N_6795);
and U9580 (N_9580,N_6843,N_6674);
xnor U9581 (N_9581,N_6830,N_5795);
nor U9582 (N_9582,N_6401,N_7283);
or U9583 (N_9583,N_7288,N_5802);
nand U9584 (N_9584,N_7132,N_5486);
xor U9585 (N_9585,N_6408,N_6705);
nand U9586 (N_9586,N_7415,N_7179);
xor U9587 (N_9587,N_7219,N_7231);
and U9588 (N_9588,N_5704,N_5567);
or U9589 (N_9589,N_7368,N_6718);
or U9590 (N_9590,N_6284,N_5066);
and U9591 (N_9591,N_5111,N_6875);
and U9592 (N_9592,N_5214,N_5254);
nor U9593 (N_9593,N_5955,N_5713);
or U9594 (N_9594,N_6639,N_6980);
or U9595 (N_9595,N_5481,N_7445);
or U9596 (N_9596,N_5275,N_6543);
nor U9597 (N_9597,N_5810,N_5793);
or U9598 (N_9598,N_7255,N_5952);
xor U9599 (N_9599,N_5157,N_5682);
nand U9600 (N_9600,N_6424,N_5213);
or U9601 (N_9601,N_5133,N_6663);
or U9602 (N_9602,N_5216,N_6346);
and U9603 (N_9603,N_6412,N_6289);
or U9604 (N_9604,N_6651,N_5843);
or U9605 (N_9605,N_5889,N_6421);
nand U9606 (N_9606,N_7034,N_6554);
xor U9607 (N_9607,N_6612,N_5836);
and U9608 (N_9608,N_5534,N_6071);
nand U9609 (N_9609,N_6411,N_7130);
nand U9610 (N_9610,N_6902,N_5220);
nor U9611 (N_9611,N_5144,N_5030);
or U9612 (N_9612,N_5758,N_5638);
nand U9613 (N_9613,N_6401,N_6793);
nor U9614 (N_9614,N_6487,N_6347);
xor U9615 (N_9615,N_5509,N_5551);
nor U9616 (N_9616,N_5759,N_5948);
nor U9617 (N_9617,N_7041,N_5222);
xor U9618 (N_9618,N_7214,N_5790);
nand U9619 (N_9619,N_5604,N_5206);
or U9620 (N_9620,N_5547,N_5489);
or U9621 (N_9621,N_5793,N_7298);
nor U9622 (N_9622,N_7399,N_5852);
or U9623 (N_9623,N_6297,N_6117);
and U9624 (N_9624,N_5439,N_5603);
or U9625 (N_9625,N_5968,N_6065);
nand U9626 (N_9626,N_7008,N_5106);
or U9627 (N_9627,N_5968,N_6908);
and U9628 (N_9628,N_6709,N_6128);
and U9629 (N_9629,N_5640,N_5336);
nand U9630 (N_9630,N_5587,N_6077);
nand U9631 (N_9631,N_6982,N_6997);
xnor U9632 (N_9632,N_6695,N_7398);
and U9633 (N_9633,N_6043,N_5865);
and U9634 (N_9634,N_7113,N_5180);
or U9635 (N_9635,N_5525,N_6484);
nand U9636 (N_9636,N_6509,N_5012);
or U9637 (N_9637,N_7243,N_7453);
nor U9638 (N_9638,N_5881,N_6987);
nand U9639 (N_9639,N_7316,N_6293);
nor U9640 (N_9640,N_7312,N_5764);
nand U9641 (N_9641,N_7438,N_7020);
nor U9642 (N_9642,N_6470,N_5872);
xnor U9643 (N_9643,N_7275,N_6026);
and U9644 (N_9644,N_6296,N_5179);
nand U9645 (N_9645,N_5867,N_6625);
or U9646 (N_9646,N_7155,N_6554);
xnor U9647 (N_9647,N_6738,N_6966);
xor U9648 (N_9648,N_7324,N_7278);
nor U9649 (N_9649,N_6870,N_6566);
xor U9650 (N_9650,N_5808,N_7306);
xnor U9651 (N_9651,N_6875,N_5846);
and U9652 (N_9652,N_6911,N_5533);
and U9653 (N_9653,N_5674,N_5675);
and U9654 (N_9654,N_5017,N_6368);
and U9655 (N_9655,N_6241,N_5762);
and U9656 (N_9656,N_5565,N_5061);
nand U9657 (N_9657,N_7119,N_5842);
xnor U9658 (N_9658,N_6531,N_6479);
and U9659 (N_9659,N_6679,N_5174);
nand U9660 (N_9660,N_7183,N_7233);
or U9661 (N_9661,N_6453,N_5233);
nor U9662 (N_9662,N_6153,N_7238);
nor U9663 (N_9663,N_6328,N_6932);
nand U9664 (N_9664,N_5357,N_5367);
xor U9665 (N_9665,N_5377,N_6406);
xnor U9666 (N_9666,N_6501,N_6080);
and U9667 (N_9667,N_6554,N_6557);
xnor U9668 (N_9668,N_6848,N_5654);
nor U9669 (N_9669,N_7413,N_5821);
nor U9670 (N_9670,N_6025,N_5696);
and U9671 (N_9671,N_7054,N_7068);
xnor U9672 (N_9672,N_5855,N_5474);
and U9673 (N_9673,N_5841,N_6789);
nor U9674 (N_9674,N_5948,N_6980);
xor U9675 (N_9675,N_7164,N_6140);
xor U9676 (N_9676,N_6470,N_6375);
and U9677 (N_9677,N_5266,N_6401);
or U9678 (N_9678,N_6557,N_6042);
nor U9679 (N_9679,N_6777,N_6748);
xnor U9680 (N_9680,N_6003,N_5338);
or U9681 (N_9681,N_5858,N_7343);
nand U9682 (N_9682,N_5474,N_5381);
nand U9683 (N_9683,N_5630,N_6470);
xor U9684 (N_9684,N_5601,N_5551);
xor U9685 (N_9685,N_5374,N_6059);
nand U9686 (N_9686,N_7147,N_5750);
and U9687 (N_9687,N_7318,N_6980);
or U9688 (N_9688,N_5843,N_5562);
or U9689 (N_9689,N_7402,N_6336);
or U9690 (N_9690,N_6641,N_6639);
xor U9691 (N_9691,N_7160,N_6011);
and U9692 (N_9692,N_7394,N_5060);
xnor U9693 (N_9693,N_5751,N_6418);
nand U9694 (N_9694,N_6482,N_6996);
xor U9695 (N_9695,N_5093,N_6701);
nand U9696 (N_9696,N_6182,N_7252);
xor U9697 (N_9697,N_6001,N_6789);
and U9698 (N_9698,N_5514,N_7157);
nand U9699 (N_9699,N_6492,N_6819);
nand U9700 (N_9700,N_5824,N_7087);
or U9701 (N_9701,N_5051,N_6268);
nand U9702 (N_9702,N_6042,N_6468);
and U9703 (N_9703,N_5259,N_6016);
and U9704 (N_9704,N_7250,N_6675);
or U9705 (N_9705,N_5579,N_5431);
xor U9706 (N_9706,N_5268,N_7090);
and U9707 (N_9707,N_6984,N_5734);
xor U9708 (N_9708,N_5374,N_6072);
nand U9709 (N_9709,N_5857,N_6845);
and U9710 (N_9710,N_7220,N_5068);
xnor U9711 (N_9711,N_5385,N_5649);
and U9712 (N_9712,N_5859,N_5135);
and U9713 (N_9713,N_6900,N_6622);
xnor U9714 (N_9714,N_7242,N_5581);
nand U9715 (N_9715,N_7316,N_5782);
xor U9716 (N_9716,N_5516,N_5650);
or U9717 (N_9717,N_6401,N_7401);
or U9718 (N_9718,N_5487,N_6057);
nand U9719 (N_9719,N_7215,N_6311);
xor U9720 (N_9720,N_6087,N_5872);
xnor U9721 (N_9721,N_5429,N_7245);
xor U9722 (N_9722,N_6818,N_7331);
or U9723 (N_9723,N_5264,N_6420);
nand U9724 (N_9724,N_5694,N_6908);
nand U9725 (N_9725,N_6455,N_5182);
nand U9726 (N_9726,N_6984,N_6878);
nand U9727 (N_9727,N_7308,N_6944);
and U9728 (N_9728,N_6440,N_6221);
nor U9729 (N_9729,N_6348,N_5825);
and U9730 (N_9730,N_6661,N_6743);
xnor U9731 (N_9731,N_6370,N_7270);
and U9732 (N_9732,N_5543,N_5240);
or U9733 (N_9733,N_6713,N_6181);
or U9734 (N_9734,N_6511,N_7301);
nor U9735 (N_9735,N_5017,N_5968);
nand U9736 (N_9736,N_6118,N_5925);
nand U9737 (N_9737,N_6717,N_6796);
xnor U9738 (N_9738,N_5434,N_5932);
or U9739 (N_9739,N_5212,N_5222);
nand U9740 (N_9740,N_6170,N_5849);
or U9741 (N_9741,N_7429,N_5808);
or U9742 (N_9742,N_6514,N_6118);
and U9743 (N_9743,N_5310,N_7024);
and U9744 (N_9744,N_5369,N_6363);
or U9745 (N_9745,N_6293,N_7273);
xnor U9746 (N_9746,N_5005,N_5053);
or U9747 (N_9747,N_5135,N_5895);
or U9748 (N_9748,N_5670,N_6716);
xnor U9749 (N_9749,N_5470,N_5527);
and U9750 (N_9750,N_5971,N_5150);
and U9751 (N_9751,N_5809,N_5899);
and U9752 (N_9752,N_6786,N_5226);
and U9753 (N_9753,N_6337,N_6439);
nor U9754 (N_9754,N_5975,N_6911);
xor U9755 (N_9755,N_5035,N_5338);
nand U9756 (N_9756,N_5856,N_6029);
and U9757 (N_9757,N_5091,N_6197);
and U9758 (N_9758,N_6192,N_5438);
and U9759 (N_9759,N_6467,N_5303);
nand U9760 (N_9760,N_5436,N_6239);
and U9761 (N_9761,N_5895,N_7070);
xor U9762 (N_9762,N_5835,N_7320);
or U9763 (N_9763,N_5002,N_7273);
nand U9764 (N_9764,N_7146,N_6368);
and U9765 (N_9765,N_7014,N_7363);
or U9766 (N_9766,N_6052,N_7364);
or U9767 (N_9767,N_7118,N_7121);
and U9768 (N_9768,N_7392,N_5173);
nand U9769 (N_9769,N_7013,N_6527);
nor U9770 (N_9770,N_6365,N_6740);
xnor U9771 (N_9771,N_7304,N_5487);
nand U9772 (N_9772,N_5464,N_6250);
xnor U9773 (N_9773,N_6087,N_7403);
nor U9774 (N_9774,N_6400,N_6548);
or U9775 (N_9775,N_5239,N_6538);
nor U9776 (N_9776,N_5130,N_6097);
xnor U9777 (N_9777,N_7015,N_7063);
nor U9778 (N_9778,N_7244,N_7208);
or U9779 (N_9779,N_5844,N_7084);
xnor U9780 (N_9780,N_7487,N_7365);
or U9781 (N_9781,N_5337,N_6946);
xnor U9782 (N_9782,N_5593,N_6330);
xnor U9783 (N_9783,N_7384,N_6459);
xor U9784 (N_9784,N_6480,N_7360);
or U9785 (N_9785,N_5890,N_7364);
nand U9786 (N_9786,N_7197,N_5622);
nor U9787 (N_9787,N_6828,N_6465);
xnor U9788 (N_9788,N_6154,N_5957);
or U9789 (N_9789,N_5366,N_5300);
or U9790 (N_9790,N_5576,N_5289);
or U9791 (N_9791,N_5820,N_6610);
or U9792 (N_9792,N_6417,N_5801);
or U9793 (N_9793,N_5963,N_5132);
and U9794 (N_9794,N_6242,N_6855);
nor U9795 (N_9795,N_5886,N_5367);
and U9796 (N_9796,N_6006,N_6383);
xnor U9797 (N_9797,N_5943,N_5362);
and U9798 (N_9798,N_7477,N_6793);
and U9799 (N_9799,N_7474,N_6657);
nand U9800 (N_9800,N_5978,N_5937);
xor U9801 (N_9801,N_6979,N_5083);
nand U9802 (N_9802,N_7412,N_6832);
nand U9803 (N_9803,N_6207,N_5274);
nor U9804 (N_9804,N_5649,N_5258);
nand U9805 (N_9805,N_7427,N_6051);
or U9806 (N_9806,N_5945,N_6971);
nor U9807 (N_9807,N_5054,N_7294);
or U9808 (N_9808,N_7133,N_6798);
nor U9809 (N_9809,N_5786,N_6751);
and U9810 (N_9810,N_5778,N_5913);
xor U9811 (N_9811,N_5524,N_5083);
xnor U9812 (N_9812,N_5483,N_5059);
and U9813 (N_9813,N_5052,N_7460);
and U9814 (N_9814,N_6818,N_5345);
nor U9815 (N_9815,N_6199,N_7424);
nor U9816 (N_9816,N_7039,N_7114);
xnor U9817 (N_9817,N_6960,N_6877);
nor U9818 (N_9818,N_6887,N_6376);
or U9819 (N_9819,N_5702,N_6318);
or U9820 (N_9820,N_5683,N_6947);
nand U9821 (N_9821,N_6342,N_7247);
nand U9822 (N_9822,N_6217,N_5537);
and U9823 (N_9823,N_5396,N_5745);
or U9824 (N_9824,N_6262,N_5376);
xor U9825 (N_9825,N_6526,N_5139);
nand U9826 (N_9826,N_6385,N_6549);
and U9827 (N_9827,N_5559,N_5878);
and U9828 (N_9828,N_5358,N_7377);
xnor U9829 (N_9829,N_6892,N_5942);
and U9830 (N_9830,N_6424,N_5344);
nor U9831 (N_9831,N_5684,N_6954);
nand U9832 (N_9832,N_6308,N_5691);
and U9833 (N_9833,N_6667,N_5017);
xnor U9834 (N_9834,N_6743,N_7150);
and U9835 (N_9835,N_7026,N_6842);
and U9836 (N_9836,N_7332,N_5560);
xor U9837 (N_9837,N_6641,N_6884);
xnor U9838 (N_9838,N_5131,N_6835);
and U9839 (N_9839,N_5585,N_7423);
or U9840 (N_9840,N_5779,N_6636);
and U9841 (N_9841,N_6335,N_6733);
xnor U9842 (N_9842,N_5385,N_6662);
or U9843 (N_9843,N_6143,N_6510);
or U9844 (N_9844,N_6648,N_5474);
and U9845 (N_9845,N_6257,N_6316);
and U9846 (N_9846,N_6844,N_7370);
nand U9847 (N_9847,N_6692,N_5713);
xor U9848 (N_9848,N_5571,N_6673);
nand U9849 (N_9849,N_7374,N_6143);
or U9850 (N_9850,N_6575,N_5712);
and U9851 (N_9851,N_6584,N_7080);
nor U9852 (N_9852,N_5431,N_6575);
and U9853 (N_9853,N_7347,N_7051);
or U9854 (N_9854,N_5295,N_6734);
xnor U9855 (N_9855,N_6179,N_7290);
nand U9856 (N_9856,N_5162,N_7076);
and U9857 (N_9857,N_6801,N_5624);
nor U9858 (N_9858,N_6961,N_5866);
nand U9859 (N_9859,N_6479,N_5094);
or U9860 (N_9860,N_6664,N_5494);
xor U9861 (N_9861,N_5432,N_6394);
and U9862 (N_9862,N_7445,N_5650);
or U9863 (N_9863,N_5191,N_6990);
xor U9864 (N_9864,N_5103,N_5311);
nor U9865 (N_9865,N_5842,N_5799);
and U9866 (N_9866,N_6136,N_6143);
and U9867 (N_9867,N_6733,N_6624);
nor U9868 (N_9868,N_6194,N_7395);
nand U9869 (N_9869,N_5881,N_6739);
nand U9870 (N_9870,N_5464,N_6770);
nor U9871 (N_9871,N_6026,N_5644);
xor U9872 (N_9872,N_6250,N_6969);
xor U9873 (N_9873,N_5122,N_6268);
xnor U9874 (N_9874,N_6693,N_6008);
nor U9875 (N_9875,N_6985,N_6759);
nand U9876 (N_9876,N_6352,N_6870);
nand U9877 (N_9877,N_6391,N_5399);
nor U9878 (N_9878,N_5911,N_5753);
and U9879 (N_9879,N_5711,N_6429);
nand U9880 (N_9880,N_6715,N_5851);
or U9881 (N_9881,N_5349,N_6449);
and U9882 (N_9882,N_7324,N_6543);
nor U9883 (N_9883,N_5877,N_7322);
xnor U9884 (N_9884,N_6239,N_5644);
nand U9885 (N_9885,N_5436,N_5304);
and U9886 (N_9886,N_5868,N_7015);
nor U9887 (N_9887,N_6560,N_7084);
and U9888 (N_9888,N_6979,N_6135);
nor U9889 (N_9889,N_5470,N_6555);
nand U9890 (N_9890,N_5773,N_6103);
nand U9891 (N_9891,N_5610,N_5432);
or U9892 (N_9892,N_6903,N_5463);
nor U9893 (N_9893,N_6936,N_5845);
nor U9894 (N_9894,N_5977,N_6429);
nor U9895 (N_9895,N_6570,N_6492);
nand U9896 (N_9896,N_5512,N_7384);
xnor U9897 (N_9897,N_5123,N_6268);
xnor U9898 (N_9898,N_6522,N_5789);
and U9899 (N_9899,N_5040,N_7437);
or U9900 (N_9900,N_5107,N_7331);
or U9901 (N_9901,N_6638,N_5164);
and U9902 (N_9902,N_5156,N_6687);
xor U9903 (N_9903,N_7003,N_7382);
nor U9904 (N_9904,N_5307,N_6530);
nor U9905 (N_9905,N_6066,N_6676);
and U9906 (N_9906,N_5332,N_6709);
nand U9907 (N_9907,N_5293,N_5079);
and U9908 (N_9908,N_5165,N_6837);
and U9909 (N_9909,N_5274,N_6509);
xor U9910 (N_9910,N_6881,N_5084);
nor U9911 (N_9911,N_5601,N_5502);
nor U9912 (N_9912,N_6326,N_5611);
or U9913 (N_9913,N_7035,N_7057);
nor U9914 (N_9914,N_6698,N_5814);
xor U9915 (N_9915,N_5473,N_6767);
or U9916 (N_9916,N_7299,N_5378);
xor U9917 (N_9917,N_5508,N_7281);
or U9918 (N_9918,N_6278,N_6177);
and U9919 (N_9919,N_7250,N_7444);
and U9920 (N_9920,N_5929,N_5657);
nor U9921 (N_9921,N_5161,N_5460);
nand U9922 (N_9922,N_5769,N_5836);
and U9923 (N_9923,N_6474,N_6635);
xnor U9924 (N_9924,N_7481,N_6532);
or U9925 (N_9925,N_6187,N_7114);
or U9926 (N_9926,N_6603,N_7217);
nor U9927 (N_9927,N_7207,N_7382);
nand U9928 (N_9928,N_6094,N_5074);
and U9929 (N_9929,N_6634,N_6282);
or U9930 (N_9930,N_7156,N_5476);
nand U9931 (N_9931,N_5455,N_5319);
nor U9932 (N_9932,N_5459,N_6557);
or U9933 (N_9933,N_6376,N_6159);
or U9934 (N_9934,N_5524,N_5042);
nand U9935 (N_9935,N_6479,N_7120);
nand U9936 (N_9936,N_5812,N_5646);
xnor U9937 (N_9937,N_6289,N_6151);
or U9938 (N_9938,N_6698,N_5863);
xnor U9939 (N_9939,N_6518,N_6434);
xor U9940 (N_9940,N_7409,N_5358);
xor U9941 (N_9941,N_5033,N_5844);
xnor U9942 (N_9942,N_6346,N_5499);
nand U9943 (N_9943,N_5922,N_5027);
and U9944 (N_9944,N_5604,N_6906);
or U9945 (N_9945,N_5568,N_7353);
and U9946 (N_9946,N_6345,N_5078);
nor U9947 (N_9947,N_7092,N_5540);
or U9948 (N_9948,N_5811,N_5594);
and U9949 (N_9949,N_6094,N_5710);
and U9950 (N_9950,N_7144,N_5597);
or U9951 (N_9951,N_5024,N_5912);
or U9952 (N_9952,N_6003,N_7390);
or U9953 (N_9953,N_5103,N_5962);
xor U9954 (N_9954,N_5044,N_7091);
and U9955 (N_9955,N_7329,N_6344);
nand U9956 (N_9956,N_7380,N_6803);
xor U9957 (N_9957,N_7250,N_6686);
xnor U9958 (N_9958,N_7432,N_6788);
xnor U9959 (N_9959,N_5697,N_6595);
and U9960 (N_9960,N_7036,N_5532);
nor U9961 (N_9961,N_7373,N_6184);
xnor U9962 (N_9962,N_5501,N_5734);
nor U9963 (N_9963,N_7358,N_5911);
nor U9964 (N_9964,N_6007,N_5321);
nand U9965 (N_9965,N_7409,N_5465);
or U9966 (N_9966,N_6418,N_7058);
xor U9967 (N_9967,N_7329,N_5871);
nor U9968 (N_9968,N_5943,N_5307);
xor U9969 (N_9969,N_5609,N_5317);
xnor U9970 (N_9970,N_7152,N_6805);
xor U9971 (N_9971,N_6744,N_7149);
nor U9972 (N_9972,N_6541,N_6725);
xor U9973 (N_9973,N_6931,N_6959);
and U9974 (N_9974,N_7266,N_5876);
nand U9975 (N_9975,N_5682,N_7374);
xnor U9976 (N_9976,N_5923,N_5227);
nand U9977 (N_9977,N_5738,N_6039);
and U9978 (N_9978,N_6321,N_6615);
nor U9979 (N_9979,N_7437,N_6193);
nand U9980 (N_9980,N_7280,N_5651);
xor U9981 (N_9981,N_6723,N_6366);
or U9982 (N_9982,N_5061,N_6870);
nor U9983 (N_9983,N_6564,N_7152);
and U9984 (N_9984,N_6720,N_5260);
nand U9985 (N_9985,N_5191,N_6745);
and U9986 (N_9986,N_5025,N_5690);
and U9987 (N_9987,N_6403,N_6127);
and U9988 (N_9988,N_5033,N_6406);
nand U9989 (N_9989,N_5193,N_5441);
xnor U9990 (N_9990,N_6979,N_5137);
and U9991 (N_9991,N_5375,N_6236);
nor U9992 (N_9992,N_7096,N_5141);
or U9993 (N_9993,N_5866,N_5522);
nand U9994 (N_9994,N_5084,N_7191);
and U9995 (N_9995,N_5506,N_5560);
and U9996 (N_9996,N_6140,N_6347);
nor U9997 (N_9997,N_6683,N_5069);
nor U9998 (N_9998,N_6686,N_6971);
or U9999 (N_9999,N_7433,N_6347);
nand U10000 (N_10000,N_8062,N_8521);
xor U10001 (N_10001,N_9951,N_9457);
nor U10002 (N_10002,N_8622,N_8283);
and U10003 (N_10003,N_8546,N_9008);
or U10004 (N_10004,N_8133,N_7559);
xor U10005 (N_10005,N_7991,N_9865);
xnor U10006 (N_10006,N_8258,N_7858);
nor U10007 (N_10007,N_8468,N_9723);
or U10008 (N_10008,N_7999,N_9000);
xor U10009 (N_10009,N_9855,N_8165);
nand U10010 (N_10010,N_9264,N_9864);
nand U10011 (N_10011,N_8497,N_8120);
or U10012 (N_10012,N_7601,N_9845);
nor U10013 (N_10013,N_9499,N_7655);
and U10014 (N_10014,N_9086,N_8978);
xor U10015 (N_10015,N_9833,N_8585);
nor U10016 (N_10016,N_9069,N_7631);
xor U10017 (N_10017,N_9797,N_8196);
nand U10018 (N_10018,N_9465,N_7543);
nand U10019 (N_10019,N_9458,N_7701);
nand U10020 (N_10020,N_7654,N_9590);
xor U10021 (N_10021,N_8350,N_8892);
nor U10022 (N_10022,N_7956,N_8830);
and U10023 (N_10023,N_7960,N_7607);
nor U10024 (N_10024,N_9419,N_8738);
and U10025 (N_10025,N_8486,N_8436);
xnor U10026 (N_10026,N_9168,N_8739);
and U10027 (N_10027,N_8138,N_9389);
and U10028 (N_10028,N_8243,N_8623);
and U10029 (N_10029,N_8712,N_8379);
or U10030 (N_10030,N_9975,N_7990);
nor U10031 (N_10031,N_9228,N_9853);
and U10032 (N_10032,N_8203,N_9009);
and U10033 (N_10033,N_8643,N_9050);
nor U10034 (N_10034,N_9850,N_8587);
or U10035 (N_10035,N_9130,N_8465);
and U10036 (N_10036,N_8376,N_9564);
xnor U10037 (N_10037,N_7735,N_9369);
and U10038 (N_10038,N_7796,N_9466);
and U10039 (N_10039,N_9659,N_9503);
and U10040 (N_10040,N_9965,N_8837);
xnor U10041 (N_10041,N_8659,N_7888);
or U10042 (N_10042,N_8420,N_7593);
or U10043 (N_10043,N_9212,N_8709);
or U10044 (N_10044,N_9452,N_8921);
nor U10045 (N_10045,N_9891,N_9041);
xor U10046 (N_10046,N_8999,N_8247);
or U10047 (N_10047,N_7859,N_9048);
and U10048 (N_10048,N_9632,N_9644);
nand U10049 (N_10049,N_8224,N_7503);
and U10050 (N_10050,N_9693,N_9029);
xor U10051 (N_10051,N_9910,N_7510);
nand U10052 (N_10052,N_8524,N_9156);
nor U10053 (N_10053,N_8629,N_7520);
or U10054 (N_10054,N_8395,N_9750);
or U10055 (N_10055,N_9587,N_8458);
nor U10056 (N_10056,N_9924,N_8417);
nand U10057 (N_10057,N_7513,N_9570);
nor U10058 (N_10058,N_9770,N_8055);
nor U10059 (N_10059,N_8431,N_9158);
nand U10060 (N_10060,N_8961,N_9201);
nand U10061 (N_10061,N_8366,N_9359);
nand U10062 (N_10062,N_8777,N_9652);
xor U10063 (N_10063,N_8969,N_7538);
nand U10064 (N_10064,N_9640,N_7661);
nor U10065 (N_10065,N_9295,N_7628);
and U10066 (N_10066,N_8344,N_8499);
nand U10067 (N_10067,N_9322,N_8107);
nor U10068 (N_10068,N_7784,N_7569);
or U10069 (N_10069,N_8285,N_9609);
and U10070 (N_10070,N_7689,N_9018);
xor U10071 (N_10071,N_9588,N_8119);
nand U10072 (N_10072,N_8819,N_8783);
and U10073 (N_10073,N_8876,N_9309);
or U10074 (N_10074,N_9710,N_9641);
or U10075 (N_10075,N_9275,N_8040);
nor U10076 (N_10076,N_9353,N_9976);
nor U10077 (N_10077,N_9591,N_8972);
and U10078 (N_10078,N_9516,N_9796);
xnor U10079 (N_10079,N_8687,N_8096);
nand U10080 (N_10080,N_9779,N_7954);
xnor U10081 (N_10081,N_7752,N_9771);
or U10082 (N_10082,N_7723,N_8631);
nand U10083 (N_10083,N_9248,N_9923);
and U10084 (N_10084,N_9550,N_9572);
nor U10085 (N_10085,N_8672,N_7610);
or U10086 (N_10086,N_8759,N_8355);
nand U10087 (N_10087,N_8815,N_7781);
xor U10088 (N_10088,N_8985,N_8901);
xor U10089 (N_10089,N_9935,N_9272);
xor U10090 (N_10090,N_8429,N_9131);
nand U10091 (N_10091,N_8880,N_7973);
nand U10092 (N_10092,N_8520,N_9208);
xnor U10093 (N_10093,N_9594,N_9828);
or U10094 (N_10094,N_9463,N_8028);
nand U10095 (N_10095,N_7774,N_7845);
or U10096 (N_10096,N_9129,N_8085);
xnor U10097 (N_10097,N_9113,N_7736);
xnor U10098 (N_10098,N_9080,N_7816);
and U10099 (N_10099,N_9428,N_9092);
nand U10100 (N_10100,N_8456,N_8691);
xor U10101 (N_10101,N_8769,N_7782);
nor U10102 (N_10102,N_8654,N_8506);
nor U10103 (N_10103,N_9656,N_7545);
nor U10104 (N_10104,N_9585,N_9243);
nand U10105 (N_10105,N_9408,N_9209);
and U10106 (N_10106,N_8141,N_7957);
nor U10107 (N_10107,N_8405,N_9905);
nand U10108 (N_10108,N_8846,N_8128);
nor U10109 (N_10109,N_8515,N_9336);
and U10110 (N_10110,N_9343,N_9645);
nand U10111 (N_10111,N_7721,N_9247);
nor U10112 (N_10112,N_9339,N_9700);
and U10113 (N_10113,N_9973,N_9737);
and U10114 (N_10114,N_9731,N_8638);
nor U10115 (N_10115,N_9945,N_8102);
nor U10116 (N_10116,N_8323,N_8543);
nand U10117 (N_10117,N_9263,N_9062);
and U10118 (N_10118,N_8101,N_9150);
nor U10119 (N_10119,N_7773,N_9616);
nor U10120 (N_10120,N_7617,N_9323);
xor U10121 (N_10121,N_8413,N_9592);
xor U10122 (N_10122,N_8762,N_8162);
or U10123 (N_10123,N_8593,N_9411);
nand U10124 (N_10124,N_9184,N_9692);
or U10125 (N_10125,N_9361,N_9214);
xor U10126 (N_10126,N_8080,N_8232);
nor U10127 (N_10127,N_9227,N_7822);
nor U10128 (N_10128,N_9903,N_7951);
or U10129 (N_10129,N_7547,N_8731);
xor U10130 (N_10130,N_8201,N_7740);
xor U10131 (N_10131,N_8669,N_8216);
or U10132 (N_10132,N_9093,N_7703);
and U10133 (N_10133,N_9374,N_7732);
or U10134 (N_10134,N_8337,N_8866);
xor U10135 (N_10135,N_9380,N_8157);
or U10136 (N_10136,N_8550,N_9174);
or U10137 (N_10137,N_9036,N_9566);
or U10138 (N_10138,N_9812,N_8378);
nor U10139 (N_10139,N_9447,N_9541);
and U10140 (N_10140,N_8888,N_8567);
and U10141 (N_10141,N_9649,N_8195);
nand U10142 (N_10142,N_7779,N_8123);
xor U10143 (N_10143,N_9074,N_8407);
or U10144 (N_10144,N_9991,N_8159);
and U10145 (N_10145,N_9111,N_9904);
xor U10146 (N_10146,N_8733,N_8314);
or U10147 (N_10147,N_9890,N_9674);
nand U10148 (N_10148,N_9962,N_8464);
nor U10149 (N_10149,N_9016,N_8032);
and U10150 (N_10150,N_9509,N_7525);
nor U10151 (N_10151,N_7589,N_9348);
nand U10152 (N_10152,N_9921,N_9291);
nand U10153 (N_10153,N_9027,N_8578);
xor U10154 (N_10154,N_9449,N_8502);
and U10155 (N_10155,N_9416,N_9536);
or U10156 (N_10156,N_8242,N_9267);
or U10157 (N_10157,N_8859,N_7948);
nor U10158 (N_10158,N_7663,N_9147);
and U10159 (N_10159,N_9091,N_8489);
nand U10160 (N_10160,N_8327,N_8516);
or U10161 (N_10161,N_8016,N_9563);
nor U10162 (N_10162,N_9985,N_8217);
and U10163 (N_10163,N_7793,N_7982);
and U10164 (N_10164,N_7687,N_7980);
and U10165 (N_10165,N_8528,N_9047);
or U10166 (N_10166,N_8240,N_8734);
nor U10167 (N_10167,N_8492,N_7965);
xnor U10168 (N_10168,N_8046,N_9250);
xnor U10169 (N_10169,N_9655,N_8112);
xnor U10170 (N_10170,N_7541,N_7931);
or U10171 (N_10171,N_7835,N_7802);
nor U10172 (N_10172,N_7775,N_9998);
nor U10173 (N_10173,N_9537,N_9152);
nand U10174 (N_10174,N_9151,N_8718);
nand U10175 (N_10175,N_8173,N_9835);
nor U10176 (N_10176,N_8656,N_8711);
nor U10177 (N_10177,N_9706,N_8542);
xnor U10178 (N_10178,N_9677,N_8430);
or U10179 (N_10179,N_9341,N_8577);
nand U10180 (N_10180,N_9814,N_7672);
nor U10181 (N_10181,N_9755,N_9884);
xor U10182 (N_10182,N_8403,N_8061);
and U10183 (N_10183,N_7813,N_9347);
and U10184 (N_10184,N_8388,N_8793);
nand U10185 (N_10185,N_8331,N_9546);
nand U10186 (N_10186,N_7800,N_7778);
nand U10187 (N_10187,N_9282,N_7805);
and U10188 (N_10188,N_9846,N_9469);
nand U10189 (N_10189,N_8000,N_9939);
xnor U10190 (N_10190,N_8596,N_8214);
nor U10191 (N_10191,N_7527,N_7578);
and U10192 (N_10192,N_7604,N_9698);
and U10193 (N_10193,N_8938,N_9679);
and U10194 (N_10194,N_9293,N_9171);
or U10195 (N_10195,N_8852,N_7504);
and U10196 (N_10196,N_9090,N_8385);
xor U10197 (N_10197,N_7648,N_8617);
or U10198 (N_10198,N_8661,N_7738);
or U10199 (N_10199,N_8174,N_8570);
nand U10200 (N_10200,N_8955,N_7895);
and U10201 (N_10201,N_9365,N_9799);
xnor U10202 (N_10202,N_8098,N_8618);
or U10203 (N_10203,N_9584,N_7967);
xor U10204 (N_10204,N_8706,N_9787);
and U10205 (N_10205,N_9667,N_8153);
nand U10206 (N_10206,N_8931,N_8073);
and U10207 (N_10207,N_9854,N_7709);
xnor U10208 (N_10208,N_8850,N_8657);
nand U10209 (N_10209,N_9744,N_8988);
and U10210 (N_10210,N_8341,N_9426);
and U10211 (N_10211,N_7814,N_7697);
or U10212 (N_10212,N_9636,N_8775);
nor U10213 (N_10213,N_7587,N_9840);
nor U10214 (N_10214,N_9053,N_9424);
xor U10215 (N_10215,N_8841,N_8911);
or U10216 (N_10216,N_9056,N_9867);
xnor U10217 (N_10217,N_8662,N_9298);
nor U10218 (N_10218,N_9832,N_9709);
xor U10219 (N_10219,N_9699,N_8956);
nor U10220 (N_10220,N_9881,N_7976);
or U10221 (N_10221,N_9598,N_7883);
xor U10222 (N_10222,N_9821,N_9303);
or U10223 (N_10223,N_8150,N_9031);
xnor U10224 (N_10224,N_8071,N_8552);
and U10225 (N_10225,N_7906,N_9626);
nor U10226 (N_10226,N_9034,N_9167);
xor U10227 (N_10227,N_9475,N_9634);
nand U10228 (N_10228,N_9310,N_9072);
xnor U10229 (N_10229,N_8339,N_8668);
nor U10230 (N_10230,N_9540,N_9759);
nand U10231 (N_10231,N_7987,N_9887);
or U10232 (N_10232,N_8462,N_8761);
nand U10233 (N_10233,N_8137,N_9127);
nor U10234 (N_10234,N_9274,N_8472);
xor U10235 (N_10235,N_7627,N_8992);
xnor U10236 (N_10236,N_9751,N_8370);
and U10237 (N_10237,N_9760,N_9245);
xnor U10238 (N_10238,N_8475,N_8386);
or U10239 (N_10239,N_8800,N_9387);
xor U10240 (N_10240,N_8838,N_9862);
or U10241 (N_10241,N_8278,N_7586);
nor U10242 (N_10242,N_9378,N_8716);
nor U10243 (N_10243,N_8504,N_8275);
nor U10244 (N_10244,N_8603,N_7887);
or U10245 (N_10245,N_9547,N_8142);
xnor U10246 (N_10246,N_7584,N_8050);
or U10247 (N_10247,N_9612,N_9173);
nand U10248 (N_10248,N_7935,N_8324);
or U10249 (N_10249,N_7749,N_9415);
xnor U10250 (N_10250,N_8522,N_8879);
and U10251 (N_10251,N_8558,N_8770);
nor U10252 (N_10252,N_9239,N_9085);
xor U10253 (N_10253,N_8758,N_9262);
nor U10254 (N_10254,N_8084,N_8154);
nand U10255 (N_10255,N_7921,N_7850);
or U10256 (N_10256,N_8135,N_8682);
xnor U10257 (N_10257,N_7546,N_7901);
nand U10258 (N_10258,N_8811,N_9077);
and U10259 (N_10259,N_8414,N_7680);
nand U10260 (N_10260,N_8548,N_8151);
nor U10261 (N_10261,N_8963,N_8494);
or U10262 (N_10262,N_8551,N_8074);
nor U10263 (N_10263,N_8373,N_9418);
nand U10264 (N_10264,N_8361,N_9520);
or U10265 (N_10265,N_8658,N_9838);
and U10266 (N_10266,N_9409,N_8438);
nor U10267 (N_10267,N_9648,N_8122);
or U10268 (N_10268,N_9670,N_7675);
and U10269 (N_10269,N_8883,N_9647);
and U10270 (N_10270,N_8336,N_7597);
nand U10271 (N_10271,N_8772,N_8727);
and U10272 (N_10272,N_8227,N_7912);
or U10273 (N_10273,N_8592,N_8047);
and U10274 (N_10274,N_9316,N_8510);
nor U10275 (N_10275,N_8817,N_9108);
xnor U10276 (N_10276,N_9889,N_9581);
nor U10277 (N_10277,N_9763,N_9953);
or U10278 (N_10278,N_8131,N_8997);
nor U10279 (N_10279,N_9933,N_7681);
nand U10280 (N_10280,N_9405,N_8557);
xor U10281 (N_10281,N_7998,N_9492);
nor U10282 (N_10282,N_7539,N_9972);
xor U10283 (N_10283,N_9970,N_8007);
and U10284 (N_10284,N_9314,N_8349);
nor U10285 (N_10285,N_7926,N_7712);
xnor U10286 (N_10286,N_8519,N_7864);
nor U10287 (N_10287,N_9420,N_8724);
or U10288 (N_10288,N_7653,N_8608);
and U10289 (N_10289,N_8559,N_8228);
or U10290 (N_10290,N_8358,N_9715);
and U10291 (N_10291,N_7839,N_9817);
or U10292 (N_10292,N_9721,N_8774);
xnor U10293 (N_10293,N_8375,N_8952);
nand U10294 (N_10294,N_9707,N_9539);
xnor U10295 (N_10295,N_8825,N_9496);
xor U10296 (N_10296,N_8621,N_9868);
nor U10297 (N_10297,N_8418,N_8976);
or U10298 (N_10298,N_9320,N_8936);
or U10299 (N_10299,N_8863,N_8900);
nor U10300 (N_10300,N_8792,N_7571);
xnor U10301 (N_10301,N_8526,N_9913);
xor U10302 (N_10302,N_9193,N_9446);
xor U10303 (N_10303,N_7928,N_9601);
nor U10304 (N_10304,N_7635,N_7599);
and U10305 (N_10305,N_7923,N_9893);
or U10306 (N_10306,N_8615,N_7602);
nor U10307 (N_10307,N_7922,N_8225);
and U10308 (N_10308,N_7910,N_8860);
and U10309 (N_10309,N_8254,N_8649);
and U10310 (N_10310,N_8856,N_8913);
nand U10311 (N_10311,N_7979,N_9164);
nor U10312 (N_10312,N_9617,N_7570);
and U10313 (N_10313,N_8250,N_9067);
xor U10314 (N_10314,N_9522,N_8348);
nand U10315 (N_10315,N_9126,N_9678);
nand U10316 (N_10316,N_8579,N_9392);
xnor U10317 (N_10317,N_7846,N_8894);
and U10318 (N_10318,N_8737,N_9321);
nor U10319 (N_10319,N_8389,N_9882);
nor U10320 (N_10320,N_9103,N_8194);
nor U10321 (N_10321,N_8023,N_9847);
nor U10322 (N_10322,N_8212,N_7620);
nand U10323 (N_10323,N_9631,N_9195);
and U10324 (N_10324,N_8272,N_8234);
xor U10325 (N_10325,N_8459,N_9680);
or U10326 (N_10326,N_9523,N_7757);
or U10327 (N_10327,N_7567,N_9633);
nand U10328 (N_10328,N_9473,N_7772);
or U10329 (N_10329,N_8448,N_9968);
nor U10330 (N_10330,N_8300,N_8466);
and U10331 (N_10331,N_8259,N_8764);
or U10332 (N_10332,N_7684,N_9377);
nor U10333 (N_10333,N_7958,N_7536);
or U10334 (N_10334,N_8732,N_9254);
xor U10335 (N_10335,N_8211,N_8966);
nor U10336 (N_10336,N_8144,N_9725);
nor U10337 (N_10337,N_8208,N_8298);
nor U10338 (N_10338,N_9919,N_8806);
nor U10339 (N_10339,N_7853,N_9338);
nor U10340 (N_10340,N_8589,N_9734);
nand U10341 (N_10341,N_9551,N_9593);
xor U10342 (N_10342,N_9544,N_8090);
nor U10343 (N_10343,N_9906,N_9404);
xor U10344 (N_10344,N_7522,N_9803);
and U10345 (N_10345,N_9914,N_9895);
or U10346 (N_10346,N_8469,N_8789);
nor U10347 (N_10347,N_9824,N_8937);
nor U10348 (N_10348,N_8027,N_8500);
nand U10349 (N_10349,N_9302,N_9289);
or U10350 (N_10350,N_7909,N_9568);
and U10351 (N_10351,N_9046,N_7988);
xnor U10352 (N_10352,N_8357,N_7580);
nor U10353 (N_10353,N_8003,N_8316);
xnor U10354 (N_10354,N_9498,N_9671);
and U10355 (N_10355,N_7529,N_9084);
and U10356 (N_10356,N_8311,N_8518);
nand U10357 (N_10357,N_7564,N_7821);
nand U10358 (N_10358,N_7702,N_9017);
xor U10359 (N_10359,N_8266,N_8313);
nor U10360 (N_10360,N_9186,N_9747);
nor U10361 (N_10361,N_7785,N_7534);
and U10362 (N_10362,N_9181,N_8163);
nor U10363 (N_10363,N_8356,N_9754);
xor U10364 (N_10364,N_9918,N_8257);
xnor U10365 (N_10365,N_8230,N_8176);
nor U10366 (N_10366,N_8571,N_9060);
nand U10367 (N_10367,N_9004,N_9687);
nand U10368 (N_10368,N_9722,N_9764);
or U10369 (N_10369,N_9089,N_7659);
xor U10370 (N_10370,N_7677,N_9055);
xor U10371 (N_10371,N_8594,N_8684);
and U10372 (N_10372,N_9402,N_8008);
and U10373 (N_10373,N_7612,N_9983);
or U10374 (N_10374,N_9682,N_7820);
or U10375 (N_10375,N_9448,N_9507);
xor U10376 (N_10376,N_9542,N_9495);
nor U10377 (N_10377,N_7843,N_9524);
and U10378 (N_10378,N_8322,N_9619);
nand U10379 (N_10379,N_9159,N_8487);
or U10380 (N_10380,N_8083,N_9144);
or U10381 (N_10381,N_8219,N_9468);
xnor U10382 (N_10382,N_8501,N_8610);
and U10383 (N_10383,N_7986,N_9015);
or U10384 (N_10384,N_7652,N_7933);
xor U10385 (N_10385,N_7598,N_9800);
and U10386 (N_10386,N_7575,N_9500);
xor U10387 (N_10387,N_9717,N_7632);
nor U10388 (N_10388,N_9413,N_9255);
or U10389 (N_10389,N_7947,N_9638);
and U10390 (N_10390,N_9329,N_9197);
and U10391 (N_10391,N_9765,N_9746);
or U10392 (N_10392,N_9326,N_8069);
and U10393 (N_10393,N_8044,N_9714);
or U10394 (N_10394,N_7940,N_9741);
or U10395 (N_10395,N_9476,N_9608);
nor U10396 (N_10396,N_9234,N_8663);
and U10397 (N_10397,N_8103,N_8580);
or U10398 (N_10398,N_8523,N_9519);
xnor U10399 (N_10399,N_8480,N_8872);
and U10400 (N_10400,N_9940,N_8493);
nor U10401 (N_10401,N_7566,N_9372);
or U10402 (N_10402,N_7556,N_8435);
nand U10403 (N_10403,N_9531,N_8155);
or U10404 (N_10404,N_9400,N_9830);
nor U10405 (N_10405,N_8803,N_8694);
and U10406 (N_10406,N_9020,N_9664);
xor U10407 (N_10407,N_8508,N_7505);
and U10408 (N_10408,N_7968,N_7874);
nor U10409 (N_10409,N_9001,N_7907);
nand U10410 (N_10410,N_8199,N_9161);
nand U10411 (N_10411,N_7949,N_9102);
or U10412 (N_10412,N_9061,N_9773);
and U10413 (N_10413,N_7501,N_9916);
or U10414 (N_10414,N_9777,N_8929);
or U10415 (N_10415,N_7695,N_8118);
nor U10416 (N_10416,N_8517,N_9752);
nor U10417 (N_10417,N_7729,N_7885);
and U10418 (N_10418,N_8625,N_9058);
xor U10419 (N_10419,N_7758,N_8152);
nor U10420 (N_10420,N_9101,N_9534);
and U10421 (N_10421,N_7915,N_9858);
nand U10422 (N_10422,N_7561,N_9358);
and U10423 (N_10423,N_8039,N_8511);
and U10424 (N_10424,N_9560,N_8399);
xnor U10425 (N_10425,N_8757,N_8095);
nand U10426 (N_10426,N_8941,N_8626);
xnor U10427 (N_10427,N_8893,N_9256);
and U10428 (N_10428,N_8873,N_9530);
and U10429 (N_10429,N_9440,N_8875);
xor U10430 (N_10430,N_7838,N_9283);
nor U10431 (N_10431,N_9467,N_9988);
or U10432 (N_10432,N_9624,N_8235);
and U10433 (N_10433,N_8916,N_9444);
xor U10434 (N_10434,N_8532,N_7902);
nor U10435 (N_10435,N_8576,N_8400);
xor U10436 (N_10436,N_7603,N_7867);
xnor U10437 (N_10437,N_9815,N_9567);
or U10438 (N_10438,N_8994,N_8384);
xnor U10439 (N_10439,N_9872,N_8460);
nor U10440 (N_10440,N_7876,N_8364);
nor U10441 (N_10441,N_7699,N_7582);
xor U10442 (N_10442,N_8612,N_8467);
or U10443 (N_10443,N_7667,N_8710);
or U10444 (N_10444,N_9486,N_8114);
xor U10445 (N_10445,N_9116,N_8392);
nand U10446 (N_10446,N_8943,N_8110);
nand U10447 (N_10447,N_7879,N_9877);
and U10448 (N_10448,N_9296,N_7719);
and U10449 (N_10449,N_9816,N_9225);
and U10450 (N_10450,N_9573,N_9139);
or U10451 (N_10451,N_8882,N_9650);
and U10452 (N_10452,N_9820,N_7725);
xor U10453 (N_10453,N_7553,N_7548);
xnor U10454 (N_10454,N_9928,N_7975);
nor U10455 (N_10455,N_8168,N_7996);
and U10456 (N_10456,N_9176,N_9947);
nor U10457 (N_10457,N_9253,N_7953);
nand U10458 (N_10458,N_9204,N_8108);
nor U10459 (N_10459,N_9182,N_8642);
or U10460 (N_10460,N_9927,N_8443);
nor U10461 (N_10461,N_8012,N_7894);
nand U10462 (N_10462,N_9472,N_8804);
xnor U10463 (N_10463,N_8805,N_8918);
nor U10464 (N_10464,N_9860,N_9528);
and U10465 (N_10465,N_9287,N_8671);
nand U10466 (N_10466,N_9386,N_7830);
and U10467 (N_10467,N_7756,N_9070);
or U10468 (N_10468,N_9346,N_8041);
nor U10469 (N_10469,N_7583,N_7925);
or U10470 (N_10470,N_7896,N_9460);
nor U10471 (N_10471,N_9284,N_8908);
nor U10472 (N_10472,N_7669,N_9148);
and U10473 (N_10473,N_9484,N_8425);
nor U10474 (N_10474,N_8049,N_8799);
nand U10475 (N_10475,N_9271,N_8832);
or U10476 (N_10476,N_8390,N_8834);
and U10477 (N_10477,N_9880,N_8575);
nor U10478 (N_10478,N_9571,N_8091);
xor U10479 (N_10479,N_7765,N_9911);
xnor U10480 (N_10480,N_8320,N_8268);
and U10481 (N_10481,N_8333,N_8784);
xor U10482 (N_10482,N_8426,N_8717);
or U10483 (N_10483,N_8088,N_8263);
and U10484 (N_10484,N_7633,N_9595);
or U10485 (N_10485,N_9954,N_9857);
and U10486 (N_10486,N_9974,N_8409);
xor U10487 (N_10487,N_9602,N_9574);
or U10488 (N_10488,N_9257,N_8043);
nor U10489 (N_10489,N_9097,N_8685);
xnor U10490 (N_10490,N_8175,N_8686);
and U10491 (N_10491,N_8001,N_8676);
nor U10492 (N_10492,N_8309,N_7962);
or U10493 (N_10493,N_8801,N_7606);
nor U10494 (N_10494,N_7831,N_9280);
nor U10495 (N_10495,N_8476,N_8845);
or U10496 (N_10496,N_7562,N_9175);
xor U10497 (N_10497,N_9705,N_7777);
and U10498 (N_10498,N_7834,N_8035);
and U10499 (N_10499,N_8011,N_8124);
xor U10500 (N_10500,N_8248,N_8981);
xor U10501 (N_10501,N_9926,N_8197);
and U10502 (N_10502,N_8267,N_9745);
xnor U10503 (N_10503,N_8813,N_9170);
nand U10504 (N_10504,N_8530,N_8944);
or U10505 (N_10505,N_9125,N_7673);
and U10506 (N_10506,N_7969,N_9642);
xor U10507 (N_10507,N_7787,N_9900);
or U10508 (N_10508,N_9733,N_7881);
and U10509 (N_10509,N_9695,N_9431);
nand U10510 (N_10510,N_8332,N_9512);
nand U10511 (N_10511,N_7718,N_8149);
and U10512 (N_10512,N_9549,N_8996);
nand U10513 (N_10513,N_7727,N_8289);
nor U10514 (N_10514,N_8393,N_9436);
nand U10515 (N_10515,N_8346,N_9166);
nor U10516 (N_10516,N_8787,N_8351);
xnor U10517 (N_10517,N_9966,N_8321);
nand U10518 (N_10518,N_9909,N_9217);
or U10519 (N_10519,N_8072,N_9340);
or U10520 (N_10520,N_9580,N_7944);
nand U10521 (N_10521,N_9313,N_7827);
nor U10522 (N_10522,N_9774,N_7824);
or U10523 (N_10523,N_9822,N_9100);
xnor U10524 (N_10524,N_9653,N_8296);
and U10525 (N_10525,N_9141,N_9133);
nor U10526 (N_10526,N_9081,N_7739);
xor U10527 (N_10527,N_9871,N_8261);
or U10528 (N_10528,N_9727,N_9666);
nor U10529 (N_10529,N_7741,N_9479);
xor U10530 (N_10530,N_9719,N_7993);
or U10531 (N_10531,N_9260,N_7857);
nor U10532 (N_10532,N_8536,N_7528);
or U10533 (N_10533,N_8613,N_9545);
nand U10534 (N_10534,N_8920,N_9044);
nor U10535 (N_10535,N_8369,N_8984);
xnor U10536 (N_10536,N_7786,N_9605);
nand U10537 (N_10537,N_9930,N_9805);
or U10538 (N_10538,N_9117,N_9761);
or U10539 (N_10539,N_7861,N_9482);
nand U10540 (N_10540,N_8531,N_8054);
nor U10541 (N_10541,N_8848,N_9012);
and U10542 (N_10542,N_8697,N_8485);
xor U10543 (N_10543,N_8954,N_9767);
and U10544 (N_10544,N_9007,N_9478);
xnor U10545 (N_10545,N_9456,N_8291);
nand U10546 (N_10546,N_7856,N_7704);
nand U10547 (N_10547,N_7966,N_9963);
or U10548 (N_10548,N_7705,N_7748);
nand U10549 (N_10549,N_7776,N_7507);
and U10550 (N_10550,N_8304,N_9399);
or U10551 (N_10551,N_9888,N_8134);
nand U10552 (N_10552,N_9236,N_9997);
nor U10553 (N_10553,N_8914,N_8223);
and U10554 (N_10554,N_9562,N_7688);
nor U10555 (N_10555,N_7666,N_8946);
and U10556 (N_10556,N_8514,N_9979);
or U10557 (N_10557,N_7970,N_7558);
and U10558 (N_10558,N_8253,N_8878);
xor U10559 (N_10559,N_8262,N_9397);
xnor U10560 (N_10560,N_7789,N_9357);
and U10561 (N_10561,N_7823,N_8802);
and U10562 (N_10562,N_9596,N_9376);
or U10563 (N_10563,N_8974,N_9912);
nor U10564 (N_10564,N_9268,N_9439);
xor U10565 (N_10565,N_8719,N_7849);
and U10566 (N_10566,N_8810,N_7530);
nand U10567 (N_10567,N_9501,N_8870);
nor U10568 (N_10568,N_8708,N_9690);
nor U10569 (N_10569,N_9354,N_9780);
nor U10570 (N_10570,N_8473,N_8447);
and U10571 (N_10571,N_8912,N_9736);
nand U10572 (N_10572,N_8288,N_9504);
or U10573 (N_10573,N_8231,N_8563);
nor U10574 (N_10574,N_9952,N_7509);
or U10575 (N_10575,N_9639,N_7691);
or U10576 (N_10576,N_9224,N_8750);
and U10577 (N_10577,N_9829,N_7851);
xor U10578 (N_10578,N_7611,N_9417);
and U10579 (N_10579,N_8844,N_9388);
xor U10580 (N_10580,N_9730,N_8455);
nor U10581 (N_10581,N_9791,N_9334);
nor U10582 (N_10582,N_8013,N_7812);
and U10583 (N_10583,N_7518,N_8639);
and U10584 (N_10584,N_7780,N_8689);
or U10585 (N_10585,N_9371,N_9600);
nor U10586 (N_10586,N_9230,N_9223);
nor U10587 (N_10587,N_7646,N_9785);
and U10588 (N_10588,N_7515,N_7616);
nand U10589 (N_10589,N_9265,N_8640);
nor U10590 (N_10590,N_8190,N_8675);
xnor U10591 (N_10591,N_8015,N_8308);
nand U10592 (N_10592,N_8359,N_8868);
nand U10593 (N_10593,N_9095,N_8645);
or U10594 (N_10594,N_9367,N_7994);
or U10595 (N_10595,N_8187,N_8544);
and U10596 (N_10596,N_7581,N_7595);
xnor U10597 (N_10597,N_8269,N_9775);
xor U10598 (N_10598,N_9989,N_8495);
nor U10599 (N_10599,N_7639,N_8714);
nand U10600 (N_10600,N_9898,N_9781);
nor U10601 (N_10601,N_8633,N_8360);
or U10602 (N_10602,N_8591,N_8780);
or U10603 (N_10603,N_9792,N_8301);
nand U10604 (N_10604,N_7523,N_8186);
nor U10605 (N_10605,N_9211,N_8045);
nand U10606 (N_10606,N_9481,N_9035);
and U10607 (N_10607,N_8564,N_9277);
and U10608 (N_10608,N_7594,N_8886);
nand U10609 (N_10609,N_9238,N_8983);
and U10610 (N_10610,N_7640,N_9586);
xor U10611 (N_10611,N_8068,N_8965);
or U10612 (N_10612,N_9307,N_8881);
xor U10613 (N_10613,N_7526,N_7624);
xnor U10614 (N_10614,N_9879,N_7565);
or U10615 (N_10615,N_8644,N_8290);
nand U10616 (N_10616,N_9140,N_8094);
nand U10617 (N_10617,N_9143,N_9464);
nor U10618 (N_10618,N_9668,N_8809);
xnor U10619 (N_10619,N_8767,N_8446);
xor U10620 (N_10620,N_9177,N_8627);
nand U10621 (N_10621,N_9646,N_8527);
nand U10622 (N_10622,N_9603,N_8652);
nor U10623 (N_10623,N_9178,N_9163);
or U10624 (N_10624,N_9735,N_9704);
nand U10625 (N_10625,N_8857,N_9215);
and U10626 (N_10626,N_7854,N_9762);
nand U10627 (N_10627,N_8949,N_8451);
nand U10628 (N_10628,N_9042,N_8816);
xnor U10629 (N_10629,N_8693,N_7792);
xnor U10630 (N_10630,N_8220,N_8056);
nor U10631 (N_10631,N_9237,N_8555);
xor U10632 (N_10632,N_9681,N_9697);
or U10633 (N_10633,N_8024,N_9028);
nand U10634 (N_10634,N_8265,N_8445);
xnor U10635 (N_10635,N_7555,N_9366);
nand U10636 (N_10636,N_8745,N_7614);
nor U10637 (N_10637,N_8971,N_8031);
xor U10638 (N_10638,N_8125,N_7521);
nand U10639 (N_10639,N_9949,N_7657);
nand U10640 (N_10640,N_9393,N_9453);
xor U10641 (N_10641,N_9381,N_9794);
or U10642 (N_10642,N_8547,N_8057);
nand U10643 (N_10643,N_8950,N_8701);
or U10644 (N_10644,N_8287,N_8415);
or U10645 (N_10645,N_9010,N_7934);
xor U10646 (N_10646,N_9390,N_8534);
nor U10647 (N_10647,N_7615,N_8034);
or U10648 (N_10648,N_9818,N_8922);
or U10649 (N_10649,N_9929,N_9720);
or U10650 (N_10650,N_9724,N_8233);
and U10651 (N_10651,N_7516,N_8670);
nand U10652 (N_10652,N_8885,N_7563);
nor U10653 (N_10653,N_9806,N_7918);
nand U10654 (N_10654,N_9967,N_8746);
or U10655 (N_10655,N_9360,N_7724);
or U10656 (N_10656,N_8160,N_8509);
xor U10657 (N_10657,N_9957,N_8822);
nand U10658 (N_10658,N_8897,N_8334);
nor U10659 (N_10659,N_9703,N_7726);
and U10660 (N_10660,N_8067,N_8730);
nand U10661 (N_10661,N_8840,N_9491);
xnor U10662 (N_10662,N_8089,N_9969);
xnor U10663 (N_10663,N_9876,N_9434);
nor U10664 (N_10664,N_8121,N_8616);
nor U10665 (N_10665,N_8006,N_8010);
and U10666 (N_10666,N_9210,N_8206);
nand U10667 (N_10667,N_8947,N_9308);
and U10668 (N_10668,N_7744,N_8241);
and U10669 (N_10669,N_8791,N_7942);
xnor U10670 (N_10670,N_9474,N_8855);
nand U10671 (N_10671,N_9827,N_8172);
nor U10672 (N_10672,N_9269,N_9852);
and U10673 (N_10673,N_8319,N_8973);
or U10674 (N_10674,N_7502,N_9937);
nand U10675 (N_10675,N_8692,N_7517);
nand U10676 (N_10676,N_8239,N_8678);
nand U10677 (N_10677,N_9057,N_7806);
nor U10678 (N_10678,N_8363,N_8345);
and U10679 (N_10679,N_7638,N_8236);
or U10680 (N_10680,N_9192,N_8765);
or U10681 (N_10681,N_8092,N_8421);
nor U10682 (N_10682,N_9789,N_7917);
and U10683 (N_10683,N_9637,N_7985);
nand U10684 (N_10684,N_7764,N_9425);
xor U10685 (N_10685,N_7730,N_8680);
nor U10686 (N_10686,N_9943,N_7535);
and U10687 (N_10687,N_9105,N_9863);
nand U10688 (N_10688,N_7574,N_8401);
and U10689 (N_10689,N_8541,N_8058);
xnor U10690 (N_10690,N_9673,N_9716);
or U10691 (N_10691,N_8915,N_9024);
nand U10692 (N_10692,N_8909,N_8115);
nor U10693 (N_10693,N_9013,N_7692);
nand U10694 (N_10694,N_7750,N_9987);
or U10695 (N_10695,N_7643,N_7936);
xnor U10696 (N_10696,N_8038,N_8484);
nor U10697 (N_10697,N_8720,N_8722);
nor U10698 (N_10698,N_8847,N_9944);
and U10699 (N_10699,N_8178,N_9960);
xnor U10700 (N_10700,N_7880,N_8540);
or U10701 (N_10701,N_8729,N_8778);
or U10702 (N_10702,N_9356,N_7621);
xor U10703 (N_10703,N_9599,N_8797);
and U10704 (N_10704,N_9373,N_9096);
or U10705 (N_10705,N_9043,N_9836);
nor U10706 (N_10706,N_9980,N_7745);
or U10707 (N_10707,N_7608,N_8060);
nand U10708 (N_10708,N_9442,N_9153);
or U10709 (N_10709,N_8831,N_8398);
xor U10710 (N_10710,N_7848,N_8889);
xor U10711 (N_10711,N_8771,N_9757);
and U10712 (N_10712,N_7919,N_8702);
xnor U10713 (N_10713,N_9790,N_9485);
nor U10714 (N_10714,N_8681,N_8752);
or U10715 (N_10715,N_8198,N_9123);
xnor U10716 (N_10716,N_9157,N_8650);
xnor U10717 (N_10717,N_8244,N_9273);
nor U10718 (N_10718,N_8158,N_7506);
or U10719 (N_10719,N_8926,N_9662);
xor U10720 (N_10720,N_9902,N_7540);
or U10721 (N_10721,N_8136,N_8326);
xor U10722 (N_10722,N_7696,N_8939);
nand U10723 (N_10723,N_9742,N_8814);
nand U10724 (N_10724,N_7656,N_7671);
and U10725 (N_10725,N_8440,N_9749);
nand U10726 (N_10726,N_8294,N_9433);
and U10727 (N_10727,N_9819,N_8812);
or U10728 (N_10728,N_8582,N_8651);
nand U10729 (N_10729,N_8664,N_9142);
nand U10730 (N_10730,N_7841,N_9410);
nor U10731 (N_10731,N_7807,N_7929);
or U10732 (N_10732,N_9083,N_9992);
or U10733 (N_10733,N_8191,N_9455);
nor U10734 (N_10734,N_8820,N_7770);
or U10735 (N_10735,N_9990,N_9187);
and U10736 (N_10736,N_8581,N_8823);
and U10737 (N_10737,N_8507,N_8340);
and U10738 (N_10738,N_9235,N_9450);
and U10739 (N_10739,N_7891,N_8100);
nor U10740 (N_10740,N_8679,N_9708);
or U10741 (N_10741,N_8858,N_7716);
or U10742 (N_10742,N_9565,N_8673);
nor U10743 (N_10743,N_8279,N_9219);
and U10744 (N_10744,N_9702,N_8167);
xor U10745 (N_10745,N_9146,N_8751);
nor U10746 (N_10746,N_8574,N_9038);
and U10747 (N_10747,N_7664,N_8910);
nor U10748 (N_10748,N_9231,N_7600);
and U10749 (N_10749,N_8932,N_8183);
and U10750 (N_10750,N_9834,N_7573);
or U10751 (N_10751,N_7768,N_8595);
and U10752 (N_10752,N_9849,N_9578);
or U10753 (N_10753,N_8599,N_8461);
or U10754 (N_10754,N_8590,N_9993);
or U10755 (N_10755,N_9607,N_8782);
nand U10756 (N_10756,N_8307,N_8807);
nor U10757 (N_10757,N_8960,N_7751);
nand U10758 (N_10758,N_9555,N_7592);
nor U10759 (N_10759,N_8884,N_8365);
or U10760 (N_10760,N_8632,N_9300);
nand U10761 (N_10761,N_9206,N_9040);
and U10762 (N_10762,N_9285,N_9134);
nand U10763 (N_10763,N_9786,N_8735);
nor U10764 (N_10764,N_8568,N_8014);
and U10765 (N_10765,N_9885,N_9629);
xor U10766 (N_10766,N_8556,N_9241);
or U10767 (N_10767,N_9961,N_9489);
nor U10768 (N_10768,N_8018,N_9931);
nor U10769 (N_10769,N_9892,N_7678);
nor U10770 (N_10770,N_9432,N_7647);
and U10771 (N_10771,N_9807,N_8896);
nand U10772 (N_10772,N_8525,N_9191);
and U10773 (N_10773,N_9527,N_9301);
nor U10774 (N_10774,N_9497,N_9202);
xnor U10775 (N_10775,N_7971,N_8786);
or U10776 (N_10776,N_8412,N_9559);
nor U10777 (N_10777,N_9620,N_9597);
xnor U10778 (N_10778,N_8410,N_9866);
and U10779 (N_10779,N_8433,N_9441);
or U10780 (N_10780,N_9946,N_8372);
nand U10781 (N_10781,N_9207,N_9330);
nor U10782 (N_10782,N_8990,N_9270);
or U10783 (N_10783,N_8048,N_9063);
nor U10784 (N_10784,N_8628,N_9793);
nor U10785 (N_10785,N_9213,N_8002);
nand U10786 (N_10786,N_9136,N_9842);
or U10787 (N_10787,N_9621,N_8276);
or U10788 (N_10788,N_8925,N_9874);
xnor U10789 (N_10789,N_9327,N_7537);
and U10790 (N_10790,N_8200,N_9396);
or U10791 (N_10791,N_9643,N_9030);
or U10792 (N_10792,N_9319,N_9222);
xor U10793 (N_10793,N_8747,N_9242);
or U10794 (N_10794,N_8260,N_7755);
and U10795 (N_10795,N_7722,N_7679);
xnor U10796 (N_10796,N_8026,N_9623);
nor U10797 (N_10797,N_7710,N_7791);
and U10798 (N_10798,N_9922,N_7715);
or U10799 (N_10799,N_9312,N_8086);
and U10800 (N_10800,N_8665,N_9753);
and U10801 (N_10801,N_8829,N_7662);
nand U10802 (N_10802,N_9611,N_7872);
and U10803 (N_10803,N_8968,N_8713);
xnor U10804 (N_10804,N_8980,N_9011);
or U10805 (N_10805,N_8688,N_8005);
nor U10806 (N_10806,N_9493,N_8601);
xnor U10807 (N_10807,N_8827,N_8169);
xor U10808 (N_10808,N_7508,N_8042);
or U10809 (N_10809,N_8207,N_9613);
or U10810 (N_10810,N_8808,N_8953);
xor U10811 (N_10811,N_8958,N_9932);
xor U10812 (N_10812,N_7809,N_9233);
and U10813 (N_10813,N_7803,N_9506);
and U10814 (N_10814,N_9878,N_9886);
xnor U10815 (N_10815,N_9487,N_9363);
and U10816 (N_10816,N_9627,N_9065);
or U10817 (N_10817,N_8967,N_8143);
nand U10818 (N_10818,N_8328,N_8053);
nor U10819 (N_10819,N_8419,N_7868);
and U10820 (N_10820,N_8907,N_8940);
or U10821 (N_10821,N_9869,N_8744);
nor U10822 (N_10822,N_9897,N_8471);
nor U10823 (N_10823,N_8677,N_9772);
xor U10824 (N_10824,N_9982,N_9756);
nand U10825 (N_10825,N_8093,N_7690);
or U10826 (N_10826,N_8624,N_9115);
and U10827 (N_10827,N_9407,N_8021);
nor U10828 (N_10828,N_8779,N_8019);
nand U10829 (N_10829,N_8353,N_9610);
xnor U10830 (N_10830,N_8229,N_8871);
xor U10831 (N_10831,N_8063,N_7808);
and U10832 (N_10832,N_9732,N_7889);
and U10833 (N_10833,N_9335,N_8842);
and U10834 (N_10834,N_7837,N_9826);
nand U10835 (N_10835,N_9379,N_7683);
nand U10836 (N_10836,N_7898,N_8648);
xor U10837 (N_10837,N_9414,N_7618);
xor U10838 (N_10838,N_7625,N_9286);
or U10839 (N_10839,N_9875,N_8218);
nor U10840 (N_10840,N_8317,N_8371);
nor U10841 (N_10841,N_8634,N_9936);
nand U10842 (N_10842,N_9899,N_8902);
and U10843 (N_10843,N_7763,N_8660);
xnor U10844 (N_10844,N_7795,N_9345);
nor U10845 (N_10845,N_7810,N_9614);
or U10846 (N_10846,N_8302,N_9955);
or U10847 (N_10847,N_8606,N_8970);
and U10848 (N_10848,N_7650,N_7514);
nand U10849 (N_10849,N_7961,N_8315);
nor U10850 (N_10850,N_9669,N_8156);
and U10851 (N_10851,N_9778,N_8743);
and U10852 (N_10852,N_8106,N_8853);
and U10853 (N_10853,N_8835,N_9145);
and U10854 (N_10854,N_8064,N_9576);
nor U10855 (N_10855,N_9279,N_9856);
and U10856 (N_10856,N_7899,N_7544);
xor U10857 (N_10857,N_9554,N_9331);
or U10858 (N_10858,N_8930,N_9368);
nor U10859 (N_10859,N_9200,N_8277);
xor U10860 (N_10860,N_7676,N_7630);
xor U10861 (N_10861,N_7645,N_8394);
and U10862 (N_10862,N_7769,N_9451);
nand U10863 (N_10863,N_9615,N_8204);
nor U10864 (N_10864,N_8698,N_8188);
nand U10865 (N_10865,N_9232,N_9606);
xor U10866 (N_10866,N_8437,N_9934);
and U10867 (N_10867,N_8998,N_8202);
xnor U10868 (N_10868,N_9124,N_9977);
or U10869 (N_10869,N_8274,N_7819);
nand U10870 (N_10870,N_9811,N_8766);
nor U10871 (N_10871,N_7707,N_8620);
nand U10872 (N_10872,N_8139,N_9691);
or U10873 (N_10873,N_8303,N_7882);
and U10874 (N_10874,N_9385,N_7875);
nor U10875 (N_10875,N_9342,N_8740);
xor U10876 (N_10876,N_9094,N_9844);
xor U10877 (N_10877,N_9438,N_9383);
xor U10878 (N_10878,N_8736,N_9005);
and U10879 (N_10879,N_8699,N_9552);
xor U10880 (N_10880,N_9128,N_7927);
and U10881 (N_10881,N_8256,N_9938);
or U10882 (N_10882,N_9579,N_7869);
nand U10883 (N_10883,N_9768,N_8411);
and U10884 (N_10884,N_7870,N_9251);
xnor U10885 (N_10885,N_9663,N_9684);
xor U10886 (N_10886,N_9006,N_8600);
nor U10887 (N_10887,N_9324,N_9494);
nor U10888 (N_10888,N_7963,N_7766);
nand U10889 (N_10889,N_9461,N_9683);
and U10890 (N_10890,N_8111,N_9395);
and U10891 (N_10891,N_9651,N_9873);
or U10892 (N_10892,N_8904,N_9686);
xnor U10893 (N_10893,N_7576,N_9517);
xor U10894 (N_10894,N_8674,N_9654);
nand U10895 (N_10895,N_8029,N_9813);
xnor U10896 (N_10896,N_9630,N_8991);
nand U10897 (N_10897,N_8513,N_8444);
or U10898 (N_10898,N_7660,N_9196);
nand U10899 (N_10899,N_7908,N_9412);
nor U10900 (N_10900,N_7930,N_8306);
nand U10901 (N_10901,N_9801,N_9798);
or U10902 (N_10902,N_8776,N_9883);
nor U10903 (N_10903,N_7833,N_9317);
xnor U10904 (N_10904,N_8635,N_8760);
xnor U10905 (N_10905,N_8756,N_9318);
nor U10906 (N_10906,N_8252,N_8935);
nand U10907 (N_10907,N_7577,N_8826);
xor U10908 (N_10908,N_8281,N_9221);
and U10909 (N_10909,N_7711,N_8295);
nand U10910 (N_10910,N_7568,N_8117);
xor U10911 (N_10911,N_8849,N_7743);
xor U10912 (N_10912,N_8488,N_8449);
or U10913 (N_10913,N_9526,N_8052);
xor U10914 (N_10914,N_7801,N_8905);
nand U10915 (N_10915,N_8075,N_8382);
or U10916 (N_10916,N_8491,N_7759);
nor U10917 (N_10917,N_7694,N_8919);
or U10918 (N_10918,N_8982,N_7613);
xor U10919 (N_10919,N_9299,N_9557);
nor U10920 (N_10920,N_7911,N_8077);
nand U10921 (N_10921,N_8066,N_8836);
or U10922 (N_10922,N_8667,N_9430);
xor U10923 (N_10923,N_9344,N_7533);
nor U10924 (N_10924,N_9259,N_7978);
xor U10925 (N_10925,N_8051,N_7767);
or U10926 (N_10926,N_7890,N_7840);
and U10927 (N_10927,N_8193,N_8641);
xor U10928 (N_10928,N_8942,N_9518);
nor U10929 (N_10929,N_8923,N_8185);
nor U10930 (N_10930,N_9118,N_9713);
and U10931 (N_10931,N_8478,N_8795);
nor U10932 (N_10932,N_8293,N_9216);
nand U10933 (N_10933,N_9401,N_9783);
nand U10934 (N_10934,N_9471,N_8569);
nand U10935 (N_10935,N_9548,N_9406);
xnor U10936 (N_10936,N_8821,N_7609);
xnor U10937 (N_10937,N_9978,N_8347);
nand U10938 (N_10938,N_8383,N_8282);
or U10939 (N_10939,N_9421,N_8647);
xor U10940 (N_10940,N_9635,N_9054);
nand U10941 (N_10941,N_8387,N_8362);
or U10942 (N_10942,N_9942,N_9026);
xor U10943 (N_10943,N_8636,N_7591);
or U10944 (N_10944,N_9477,N_7892);
xnor U10945 (N_10945,N_9252,N_8690);
nor U10946 (N_10946,N_9025,N_8605);
or U10947 (N_10947,N_7642,N_9459);
and U10948 (N_10948,N_9538,N_8022);
nor U10949 (N_10949,N_7815,N_8964);
nand U10950 (N_10950,N_9205,N_8145);
nor U10951 (N_10951,N_7714,N_9795);
xor U10952 (N_10952,N_9726,N_8877);
and U10953 (N_10953,N_9311,N_9454);
nor U10954 (N_10954,N_9132,N_9870);
xnor U10955 (N_10955,N_8742,N_9831);
or U10956 (N_10956,N_7878,N_9740);
and U10957 (N_10957,N_8402,N_7873);
nand U10958 (N_10958,N_8105,N_9194);
nor U10959 (N_10959,N_7720,N_9604);
and U10960 (N_10960,N_8251,N_8538);
and U10961 (N_10961,N_8354,N_9694);
nand U10962 (N_10962,N_8588,N_7531);
xor U10963 (N_10963,N_7579,N_9297);
xnor U10964 (N_10964,N_8989,N_9333);
nand U10965 (N_10965,N_7984,N_8025);
nand U10966 (N_10966,N_8132,N_9160);
xor U10967 (N_10967,N_8004,N_8442);
nor U10968 (N_10968,N_8927,N_9370);
nand U10969 (N_10969,N_7619,N_7826);
or U10970 (N_10970,N_9337,N_8423);
or U10971 (N_10971,N_9362,N_7992);
nor U10972 (N_10972,N_9782,N_9351);
and U10973 (N_10973,N_8479,N_9021);
and U10974 (N_10974,N_8009,N_7728);
nor U10975 (N_10975,N_7596,N_8696);
and U10976 (N_10976,N_7877,N_7836);
or U10977 (N_10977,N_9110,N_9515);
nor U10978 (N_10978,N_9185,N_9290);
and U10979 (N_10979,N_8377,N_9525);
xnor U10980 (N_10980,N_9003,N_8284);
xor U10981 (N_10981,N_9022,N_9808);
or U10982 (N_10982,N_7914,N_7955);
nor U10983 (N_10983,N_8583,N_9508);
nor U10984 (N_10984,N_8245,N_8246);
or U10985 (N_10985,N_9658,N_9106);
nor U10986 (N_10986,N_8338,N_9825);
nand U10987 (N_10987,N_8368,N_8427);
and U10988 (N_10988,N_8367,N_8033);
nor U10989 (N_10989,N_9188,N_9138);
nor U10990 (N_10990,N_9244,N_7941);
nor U10991 (N_10991,N_7964,N_9437);
nor U10992 (N_10992,N_9051,N_9529);
xnor U10993 (N_10993,N_9082,N_9422);
and U10994 (N_10994,N_8539,N_8164);
nor U10995 (N_10995,N_7818,N_9622);
nand U10996 (N_10996,N_9901,N_9240);
xor U10997 (N_10997,N_9908,N_8422);
nand U10998 (N_10998,N_7959,N_7983);
xnor U10999 (N_10999,N_8979,N_7524);
xnor U11000 (N_11000,N_8097,N_8104);
and U11001 (N_11001,N_8503,N_8554);
xnor U11002 (N_11002,N_9514,N_8147);
and U11003 (N_11003,N_7871,N_7798);
xor U11004 (N_11004,N_8951,N_8993);
nor U11005 (N_11005,N_8434,N_9033);
or U11006 (N_11006,N_9350,N_9014);
nand U11007 (N_11007,N_7811,N_7626);
or U11008 (N_11008,N_8391,N_8130);
or U11009 (N_11009,N_7788,N_9964);
nand U11010 (N_11010,N_7897,N_7674);
nand U11011 (N_11011,N_9470,N_8975);
xor U11012 (N_11012,N_8934,N_8987);
xor U11013 (N_11013,N_8609,N_9510);
or U11014 (N_11014,N_8796,N_7670);
and U11015 (N_11015,N_9660,N_8604);
and U11016 (N_11016,N_8381,N_9304);
nor U11017 (N_11017,N_8899,N_9848);
and U11018 (N_11018,N_9075,N_8828);
nor U11019 (N_11019,N_9037,N_9558);
and U11020 (N_11020,N_9994,N_8210);
nand U11021 (N_11021,N_9073,N_9718);
nand U11022 (N_11022,N_7588,N_8129);
or U11023 (N_11023,N_9220,N_7731);
and U11024 (N_11024,N_8505,N_7644);
or U11025 (N_11025,N_8030,N_9278);
xnor U11026 (N_11026,N_9098,N_7742);
or U11027 (N_11027,N_9743,N_9332);
nand U11028 (N_11028,N_9375,N_9533);
or U11029 (N_11029,N_9583,N_8703);
or U11030 (N_11030,N_9249,N_9229);
xnor U11031 (N_11031,N_8725,N_9305);
nand U11032 (N_11032,N_7651,N_7753);
and U11033 (N_11033,N_9521,N_9701);
xnor U11034 (N_11034,N_7952,N_9099);
xor U11035 (N_11035,N_8237,N_9788);
or U11036 (N_11036,N_9068,N_9738);
or U11037 (N_11037,N_8790,N_9915);
nand U11038 (N_11038,N_8335,N_8781);
or U11039 (N_11039,N_8177,N_9577);
or U11040 (N_11040,N_9996,N_7761);
xnor U11041 (N_11041,N_8614,N_7733);
and U11042 (N_11042,N_9758,N_8653);
and U11043 (N_11043,N_8127,N_8749);
xor U11044 (N_11044,N_8305,N_7665);
xnor U11045 (N_11045,N_9079,N_8655);
and U11046 (N_11046,N_8463,N_9784);
nand U11047 (N_11047,N_9306,N_7997);
nor U11048 (N_11048,N_7771,N_8226);
nand U11049 (N_11049,N_8598,N_8310);
nor U11050 (N_11050,N_9618,N_9261);
xnor U11051 (N_11051,N_9019,N_8561);
xor U11052 (N_11052,N_8406,N_8535);
xnor U11053 (N_11053,N_7797,N_8318);
nand U11054 (N_11054,N_7995,N_8962);
nor U11055 (N_11055,N_7939,N_8182);
xnor U11056 (N_11056,N_9582,N_7855);
nor U11057 (N_11057,N_8213,N_9950);
nor U11058 (N_11058,N_7734,N_8428);
nor U11059 (N_11059,N_9711,N_8113);
nor U11060 (N_11060,N_8325,N_9023);
xnor U11061 (N_11061,N_7981,N_9907);
xnor U11062 (N_11062,N_8148,N_7832);
xnor U11063 (N_11063,N_9959,N_8948);
xor U11064 (N_11064,N_7825,N_7737);
and U11065 (N_11065,N_8404,N_8562);
or U11066 (N_11066,N_8454,N_8903);
nand U11067 (N_11067,N_8728,N_7629);
nand U11068 (N_11068,N_8768,N_9190);
and U11069 (N_11069,N_8146,N_7549);
nor U11070 (N_11070,N_9505,N_9689);
or U11071 (N_11071,N_9948,N_8566);
and U11072 (N_11072,N_9059,N_9294);
nand U11073 (N_11073,N_8330,N_8439);
xnor U11074 (N_11074,N_7886,N_7828);
nand U11075 (N_11075,N_8529,N_9039);
or U11076 (N_11076,N_8895,N_9513);
or U11077 (N_11077,N_8861,N_9382);
and U11078 (N_11078,N_7542,N_9535);
or U11079 (N_11079,N_7685,N_9920);
nand U11080 (N_11080,N_7989,N_9104);
nor U11081 (N_11081,N_7866,N_9064);
or U11082 (N_11082,N_8959,N_7817);
and U11083 (N_11083,N_8481,N_7698);
nor U11084 (N_11084,N_9569,N_9122);
nor U11085 (N_11085,N_8721,N_8611);
xnor U11086 (N_11086,N_7937,N_7790);
nor U11087 (N_11087,N_9052,N_9198);
or U11088 (N_11088,N_7700,N_8065);
xor U11089 (N_11089,N_9589,N_9384);
nor U11090 (N_11090,N_8891,N_7590);
xor U11091 (N_11091,N_7794,N_8788);
or U11092 (N_11092,N_7649,N_9149);
nand U11093 (N_11093,N_7946,N_9403);
xnor U11094 (N_11094,N_8079,N_8352);
or U11095 (N_11095,N_8082,N_9328);
and U11096 (N_11096,N_9266,N_9199);
and U11097 (N_11097,N_8264,N_7686);
and U11098 (N_11098,N_8560,N_8565);
nand U11099 (N_11099,N_9002,N_8470);
nor U11100 (N_11100,N_9841,N_8700);
or U11101 (N_11101,N_9218,N_8755);
and U11102 (N_11102,N_7511,N_8630);
xnor U11103 (N_11103,N_9045,N_8457);
and U11104 (N_11104,N_8584,N_7829);
and U11105 (N_11105,N_8887,N_8715);
and U11106 (N_11106,N_7550,N_9203);
nor U11107 (N_11107,N_8537,N_8059);
and U11108 (N_11108,N_7903,N_8161);
nand U11109 (N_11109,N_8189,N_8180);
nor U11110 (N_11110,N_8477,N_8070);
or U11111 (N_11111,N_7658,N_9435);
and U11112 (N_11112,N_8833,N_8553);
xnor U11113 (N_11113,N_9180,N_9676);
nand U11114 (N_11114,N_8773,N_9179);
or U11115 (N_11115,N_9398,N_9352);
or U11116 (N_11116,N_8851,N_7532);
nand U11117 (N_11117,N_7972,N_7844);
xor U11118 (N_11118,N_8977,N_9971);
or U11119 (N_11119,N_9391,N_7862);
and U11120 (N_11120,N_9675,N_9917);
xor U11121 (N_11121,N_9804,N_8184);
and U11122 (N_11122,N_8273,N_8753);
nand U11123 (N_11123,N_9189,N_8824);
nand U11124 (N_11124,N_7977,N_8986);
nand U11125 (N_11125,N_9999,N_8474);
nand U11126 (N_11126,N_9986,N_9511);
nor U11127 (N_11127,N_8441,N_9502);
nor U11128 (N_11128,N_8099,N_8865);
nand U11129 (N_11129,N_8898,N_9837);
or U11130 (N_11130,N_7713,N_8343);
xor U11131 (N_11131,N_8222,N_8205);
nor U11132 (N_11132,N_7634,N_8933);
nand U11133 (N_11133,N_7519,N_7920);
and U11134 (N_11134,N_9155,N_9315);
and U11135 (N_11135,N_7924,N_8249);
and U11136 (N_11136,N_8255,N_7938);
or U11137 (N_11137,N_7904,N_7762);
nand U11138 (N_11138,N_9748,N_9532);
nor U11139 (N_11139,N_9488,N_8704);
and U11140 (N_11140,N_7950,N_9628);
and U11141 (N_11141,N_9958,N_8748);
or U11142 (N_11142,N_7900,N_7860);
xnor U11143 (N_11143,N_7865,N_8695);
xnor U11144 (N_11144,N_9258,N_8839);
or U11145 (N_11145,N_9066,N_7974);
nor U11146 (N_11146,N_8864,N_8726);
nor U11147 (N_11147,N_9112,N_8549);
nand U11148 (N_11148,N_9809,N_9276);
xor U11149 (N_11149,N_8867,N_8496);
nand U11150 (N_11150,N_7641,N_8181);
and U11151 (N_11151,N_7500,N_8637);
nand U11152 (N_11152,N_8299,N_9107);
nor U11153 (N_11153,N_8928,N_9292);
and U11154 (N_11154,N_8741,N_7552);
or U11155 (N_11155,N_8572,N_8924);
and U11156 (N_11156,N_8607,N_9728);
xor U11157 (N_11157,N_9561,N_7905);
nand U11158 (N_11158,N_8297,N_8906);
nand U11159 (N_11159,N_9665,N_9109);
and U11160 (N_11160,N_8483,N_7708);
and U11161 (N_11161,N_8862,N_9325);
or U11162 (N_11162,N_7913,N_8945);
nand U11163 (N_11163,N_7622,N_9137);
and U11164 (N_11164,N_8452,N_7637);
xnor U11165 (N_11165,N_9165,N_8116);
and U11166 (N_11166,N_9851,N_8170);
or U11167 (N_11167,N_8854,N_8020);
and U11168 (N_11168,N_7754,N_7557);
xor U11169 (N_11169,N_9739,N_9364);
nor U11170 (N_11170,N_8646,N_7893);
xnor U11171 (N_11171,N_9995,N_8271);
and U11172 (N_11172,N_9894,N_8416);
or U11173 (N_11173,N_9859,N_9553);
xnor U11174 (N_11174,N_8081,N_7623);
nor U11175 (N_11175,N_8221,N_9823);
or U11176 (N_11176,N_8707,N_9810);
and U11177 (N_11177,N_9078,N_9226);
nand U11178 (N_11178,N_8017,N_7760);
nand U11179 (N_11179,N_7717,N_9429);
and U11180 (N_11180,N_8798,N_9423);
and U11181 (N_11181,N_9729,N_8037);
xor U11182 (N_11182,N_9712,N_9657);
and U11183 (N_11183,N_9556,N_7847);
xnor U11184 (N_11184,N_8342,N_7668);
and U11185 (N_11185,N_9246,N_8533);
and U11186 (N_11186,N_9925,N_7932);
and U11187 (N_11187,N_9769,N_9288);
nor U11188 (N_11188,N_8215,N_9076);
xor U11189 (N_11189,N_8723,N_9861);
nand U11190 (N_11190,N_9087,N_7945);
nand U11191 (N_11191,N_9154,N_9049);
nor U11192 (N_11192,N_8763,N_8209);
or U11193 (N_11193,N_8597,N_9941);
nand U11194 (N_11194,N_7799,N_7706);
nor U11195 (N_11195,N_8586,N_8076);
nand U11196 (N_11196,N_8794,N_9984);
nand U11197 (N_11197,N_9071,N_8036);
nor U11198 (N_11198,N_8573,N_9672);
or U11199 (N_11199,N_9427,N_9120);
and U11200 (N_11200,N_9121,N_8329);
and U11201 (N_11201,N_7943,N_9896);
xnor U11202 (N_11202,N_8424,N_8380);
nand U11203 (N_11203,N_7512,N_7585);
nor U11204 (N_11204,N_9114,N_9543);
nor U11205 (N_11205,N_8498,N_7804);
and U11206 (N_11206,N_7747,N_8818);
and U11207 (N_11207,N_9088,N_7560);
nor U11208 (N_11208,N_8109,N_8192);
or U11209 (N_11209,N_7572,N_8087);
nor U11210 (N_11210,N_8619,N_9688);
xnor U11211 (N_11211,N_8666,N_7636);
and U11212 (N_11212,N_9776,N_9480);
nor U11213 (N_11213,N_8890,N_8602);
nor U11214 (N_11214,N_9135,N_9169);
or U11215 (N_11215,N_8171,N_7746);
nor U11216 (N_11216,N_8490,N_9172);
nand U11217 (N_11217,N_9981,N_8238);
xor U11218 (N_11218,N_8396,N_8995);
nor U11219 (N_11219,N_9162,N_9355);
or U11220 (N_11220,N_9462,N_9349);
or U11221 (N_11221,N_8179,N_7783);
nor U11222 (N_11222,N_8408,N_7916);
or U11223 (N_11223,N_8374,N_8785);
nor U11224 (N_11224,N_8270,N_7842);
and U11225 (N_11225,N_9839,N_8754);
xor U11226 (N_11226,N_8292,N_8432);
nand U11227 (N_11227,N_8453,N_9443);
or U11228 (N_11228,N_9625,N_9956);
or U11229 (N_11229,N_8280,N_9575);
or U11230 (N_11230,N_8705,N_9032);
and U11231 (N_11231,N_8512,N_9445);
nand U11232 (N_11232,N_9281,N_8312);
xnor U11233 (N_11233,N_9843,N_8078);
nor U11234 (N_11234,N_9802,N_7884);
nand U11235 (N_11235,N_8545,N_7693);
nor U11236 (N_11236,N_8286,N_8397);
nor U11237 (N_11237,N_8140,N_8683);
nand U11238 (N_11238,N_8843,N_9483);
nand U11239 (N_11239,N_8869,N_8126);
nor U11240 (N_11240,N_8917,N_8957);
or U11241 (N_11241,N_7551,N_8166);
and U11242 (N_11242,N_9661,N_9119);
nand U11243 (N_11243,N_9490,N_7554);
or U11244 (N_11244,N_8874,N_7682);
nor U11245 (N_11245,N_8450,N_9696);
and U11246 (N_11246,N_9183,N_8482);
nor U11247 (N_11247,N_7605,N_9394);
or U11248 (N_11248,N_7863,N_7852);
xor U11249 (N_11249,N_9685,N_9766);
and U11250 (N_11250,N_8660,N_7733);
nor U11251 (N_11251,N_7514,N_8267);
or U11252 (N_11252,N_9560,N_9245);
nand U11253 (N_11253,N_9115,N_7876);
nor U11254 (N_11254,N_9739,N_8488);
and U11255 (N_11255,N_7546,N_7549);
nand U11256 (N_11256,N_7738,N_9632);
nand U11257 (N_11257,N_7677,N_8716);
nor U11258 (N_11258,N_9549,N_8895);
nor U11259 (N_11259,N_8389,N_9849);
nor U11260 (N_11260,N_9325,N_9352);
and U11261 (N_11261,N_7551,N_8623);
nor U11262 (N_11262,N_8935,N_9264);
or U11263 (N_11263,N_9706,N_9787);
and U11264 (N_11264,N_9818,N_8732);
and U11265 (N_11265,N_8002,N_7534);
xnor U11266 (N_11266,N_8796,N_9389);
xnor U11267 (N_11267,N_7918,N_7684);
xnor U11268 (N_11268,N_9638,N_7924);
and U11269 (N_11269,N_7919,N_8682);
xor U11270 (N_11270,N_9730,N_8024);
or U11271 (N_11271,N_9162,N_7981);
nand U11272 (N_11272,N_8544,N_9035);
or U11273 (N_11273,N_8276,N_9167);
or U11274 (N_11274,N_9279,N_9182);
xor U11275 (N_11275,N_8470,N_8861);
and U11276 (N_11276,N_8072,N_7970);
nand U11277 (N_11277,N_9102,N_8509);
and U11278 (N_11278,N_8348,N_9168);
or U11279 (N_11279,N_8111,N_7697);
or U11280 (N_11280,N_8778,N_9594);
xnor U11281 (N_11281,N_8832,N_9198);
xnor U11282 (N_11282,N_9924,N_8521);
nand U11283 (N_11283,N_8973,N_9617);
or U11284 (N_11284,N_8030,N_8010);
and U11285 (N_11285,N_8820,N_9314);
and U11286 (N_11286,N_7748,N_9375);
or U11287 (N_11287,N_8241,N_7588);
nor U11288 (N_11288,N_7941,N_7783);
and U11289 (N_11289,N_7887,N_8876);
nor U11290 (N_11290,N_8656,N_8503);
nand U11291 (N_11291,N_7554,N_9651);
or U11292 (N_11292,N_9895,N_9715);
or U11293 (N_11293,N_7548,N_9264);
and U11294 (N_11294,N_9028,N_9959);
xor U11295 (N_11295,N_9148,N_8072);
nor U11296 (N_11296,N_8669,N_7961);
and U11297 (N_11297,N_8442,N_7669);
and U11298 (N_11298,N_8289,N_8893);
and U11299 (N_11299,N_9866,N_7814);
xor U11300 (N_11300,N_9503,N_9428);
nor U11301 (N_11301,N_9139,N_9944);
and U11302 (N_11302,N_9847,N_8563);
nor U11303 (N_11303,N_8865,N_9361);
and U11304 (N_11304,N_8174,N_8811);
and U11305 (N_11305,N_9838,N_7710);
xor U11306 (N_11306,N_9460,N_8114);
xnor U11307 (N_11307,N_8372,N_9792);
nor U11308 (N_11308,N_8739,N_8676);
nand U11309 (N_11309,N_8660,N_9128);
nand U11310 (N_11310,N_9554,N_7942);
or U11311 (N_11311,N_9586,N_9313);
xor U11312 (N_11312,N_8236,N_8772);
or U11313 (N_11313,N_8019,N_8816);
nor U11314 (N_11314,N_7514,N_7518);
and U11315 (N_11315,N_7652,N_9245);
nand U11316 (N_11316,N_9891,N_8076);
xnor U11317 (N_11317,N_9689,N_9961);
xnor U11318 (N_11318,N_8126,N_7960);
xor U11319 (N_11319,N_9499,N_9000);
xnor U11320 (N_11320,N_9814,N_7894);
and U11321 (N_11321,N_9430,N_8238);
nor U11322 (N_11322,N_9355,N_9202);
and U11323 (N_11323,N_8178,N_9021);
xnor U11324 (N_11324,N_9927,N_8312);
xnor U11325 (N_11325,N_9545,N_8707);
nand U11326 (N_11326,N_7647,N_9062);
or U11327 (N_11327,N_9781,N_7923);
nor U11328 (N_11328,N_9350,N_9483);
nor U11329 (N_11329,N_8612,N_8464);
nand U11330 (N_11330,N_7733,N_8092);
and U11331 (N_11331,N_8855,N_7581);
and U11332 (N_11332,N_9979,N_8320);
nor U11333 (N_11333,N_8088,N_7545);
and U11334 (N_11334,N_7554,N_8024);
and U11335 (N_11335,N_9448,N_8115);
and U11336 (N_11336,N_7736,N_8663);
nor U11337 (N_11337,N_8702,N_8283);
nor U11338 (N_11338,N_7966,N_9423);
and U11339 (N_11339,N_7605,N_9922);
or U11340 (N_11340,N_9451,N_9061);
or U11341 (N_11341,N_9538,N_8225);
nand U11342 (N_11342,N_9357,N_7969);
or U11343 (N_11343,N_8624,N_9962);
or U11344 (N_11344,N_7938,N_7527);
and U11345 (N_11345,N_9120,N_8898);
nand U11346 (N_11346,N_9618,N_9125);
xnor U11347 (N_11347,N_8181,N_7756);
nand U11348 (N_11348,N_8968,N_8906);
or U11349 (N_11349,N_8344,N_9905);
and U11350 (N_11350,N_8570,N_8238);
nor U11351 (N_11351,N_9151,N_9923);
and U11352 (N_11352,N_9472,N_7647);
and U11353 (N_11353,N_7648,N_9371);
or U11354 (N_11354,N_7810,N_7657);
and U11355 (N_11355,N_7571,N_9224);
nand U11356 (N_11356,N_7729,N_7959);
nor U11357 (N_11357,N_8945,N_9685);
and U11358 (N_11358,N_9860,N_9742);
or U11359 (N_11359,N_8649,N_7646);
and U11360 (N_11360,N_8029,N_9523);
or U11361 (N_11361,N_7544,N_7750);
nand U11362 (N_11362,N_7565,N_7886);
nor U11363 (N_11363,N_9430,N_9038);
nor U11364 (N_11364,N_8815,N_9576);
xor U11365 (N_11365,N_8979,N_7739);
xor U11366 (N_11366,N_9779,N_9091);
or U11367 (N_11367,N_8903,N_9736);
nand U11368 (N_11368,N_7531,N_9390);
nor U11369 (N_11369,N_7654,N_8928);
nor U11370 (N_11370,N_9630,N_8103);
xnor U11371 (N_11371,N_9199,N_8599);
nand U11372 (N_11372,N_7707,N_7615);
nor U11373 (N_11373,N_9134,N_8775);
nor U11374 (N_11374,N_8245,N_9429);
or U11375 (N_11375,N_9495,N_8873);
and U11376 (N_11376,N_8106,N_9789);
nand U11377 (N_11377,N_8089,N_8449);
or U11378 (N_11378,N_9344,N_7745);
nand U11379 (N_11379,N_8449,N_9837);
and U11380 (N_11380,N_7817,N_7760);
nor U11381 (N_11381,N_7640,N_7708);
nand U11382 (N_11382,N_9147,N_9199);
xor U11383 (N_11383,N_9917,N_9321);
xor U11384 (N_11384,N_8747,N_7849);
and U11385 (N_11385,N_9657,N_8632);
nor U11386 (N_11386,N_9968,N_8797);
nor U11387 (N_11387,N_8849,N_8243);
xnor U11388 (N_11388,N_7706,N_9704);
nor U11389 (N_11389,N_9552,N_9571);
and U11390 (N_11390,N_8757,N_8585);
or U11391 (N_11391,N_8457,N_9644);
or U11392 (N_11392,N_8089,N_8727);
nor U11393 (N_11393,N_9307,N_7969);
or U11394 (N_11394,N_9974,N_8428);
nand U11395 (N_11395,N_7626,N_9897);
nor U11396 (N_11396,N_8713,N_9896);
and U11397 (N_11397,N_9468,N_8304);
and U11398 (N_11398,N_8174,N_9009);
xor U11399 (N_11399,N_7848,N_8193);
or U11400 (N_11400,N_8412,N_9634);
and U11401 (N_11401,N_9651,N_9246);
and U11402 (N_11402,N_7721,N_9440);
xor U11403 (N_11403,N_9531,N_8480);
xor U11404 (N_11404,N_8992,N_8917);
or U11405 (N_11405,N_7833,N_8073);
nor U11406 (N_11406,N_8967,N_8122);
or U11407 (N_11407,N_9682,N_8259);
nand U11408 (N_11408,N_9616,N_9145);
or U11409 (N_11409,N_9209,N_8092);
xnor U11410 (N_11410,N_8384,N_9075);
nand U11411 (N_11411,N_9088,N_8074);
nor U11412 (N_11412,N_8029,N_8635);
or U11413 (N_11413,N_8443,N_8410);
and U11414 (N_11414,N_9308,N_8887);
xnor U11415 (N_11415,N_7580,N_8624);
or U11416 (N_11416,N_9548,N_8530);
or U11417 (N_11417,N_8367,N_9232);
or U11418 (N_11418,N_9821,N_9214);
or U11419 (N_11419,N_7999,N_8182);
nor U11420 (N_11420,N_8724,N_9479);
or U11421 (N_11421,N_8577,N_7976);
and U11422 (N_11422,N_8050,N_7914);
nor U11423 (N_11423,N_9760,N_8846);
xor U11424 (N_11424,N_8578,N_8110);
or U11425 (N_11425,N_9485,N_9208);
nor U11426 (N_11426,N_8988,N_9117);
nand U11427 (N_11427,N_8556,N_7969);
nor U11428 (N_11428,N_8797,N_9293);
xnor U11429 (N_11429,N_7977,N_9602);
nand U11430 (N_11430,N_9933,N_9898);
nor U11431 (N_11431,N_8110,N_8140);
nand U11432 (N_11432,N_8718,N_9255);
or U11433 (N_11433,N_9131,N_7854);
xnor U11434 (N_11434,N_8438,N_9307);
nor U11435 (N_11435,N_9314,N_7581);
nor U11436 (N_11436,N_8989,N_9422);
nand U11437 (N_11437,N_9773,N_7910);
and U11438 (N_11438,N_9620,N_8230);
nor U11439 (N_11439,N_9902,N_8176);
or U11440 (N_11440,N_9264,N_9403);
or U11441 (N_11441,N_8770,N_7554);
xnor U11442 (N_11442,N_8308,N_8870);
and U11443 (N_11443,N_8545,N_7593);
or U11444 (N_11444,N_9214,N_9869);
xor U11445 (N_11445,N_9868,N_9791);
nand U11446 (N_11446,N_8156,N_8754);
nand U11447 (N_11447,N_7578,N_9810);
xnor U11448 (N_11448,N_9822,N_8208);
nand U11449 (N_11449,N_8895,N_9953);
nand U11450 (N_11450,N_9117,N_7707);
nand U11451 (N_11451,N_8201,N_9489);
nand U11452 (N_11452,N_9229,N_7629);
nor U11453 (N_11453,N_8477,N_9742);
nand U11454 (N_11454,N_9747,N_9140);
and U11455 (N_11455,N_8655,N_7560);
and U11456 (N_11456,N_7735,N_8015);
nor U11457 (N_11457,N_8034,N_8797);
xnor U11458 (N_11458,N_8306,N_8180);
nor U11459 (N_11459,N_7795,N_9246);
nor U11460 (N_11460,N_9183,N_7555);
nor U11461 (N_11461,N_9134,N_8765);
xor U11462 (N_11462,N_8652,N_8881);
nand U11463 (N_11463,N_7795,N_8355);
nand U11464 (N_11464,N_9823,N_9332);
nand U11465 (N_11465,N_9159,N_8920);
nor U11466 (N_11466,N_9479,N_9711);
nor U11467 (N_11467,N_8802,N_9225);
nor U11468 (N_11468,N_9106,N_8782);
nand U11469 (N_11469,N_7549,N_9243);
xor U11470 (N_11470,N_7638,N_9500);
nand U11471 (N_11471,N_9323,N_8382);
xnor U11472 (N_11472,N_8008,N_7840);
nor U11473 (N_11473,N_8238,N_8185);
xor U11474 (N_11474,N_8283,N_8350);
xnor U11475 (N_11475,N_9923,N_9801);
nand U11476 (N_11476,N_8222,N_9453);
nand U11477 (N_11477,N_9844,N_9829);
nand U11478 (N_11478,N_8039,N_9841);
xnor U11479 (N_11479,N_8295,N_9430);
xnor U11480 (N_11480,N_8345,N_8836);
or U11481 (N_11481,N_8164,N_7655);
or U11482 (N_11482,N_9216,N_8389);
nor U11483 (N_11483,N_9512,N_7848);
xnor U11484 (N_11484,N_8368,N_9257);
nand U11485 (N_11485,N_9588,N_8831);
and U11486 (N_11486,N_7590,N_9332);
nor U11487 (N_11487,N_7836,N_8121);
or U11488 (N_11488,N_9000,N_8770);
and U11489 (N_11489,N_9496,N_8675);
nor U11490 (N_11490,N_7694,N_9241);
xnor U11491 (N_11491,N_9094,N_9948);
nand U11492 (N_11492,N_8571,N_9324);
nand U11493 (N_11493,N_8974,N_9515);
nand U11494 (N_11494,N_8797,N_8227);
xnor U11495 (N_11495,N_8742,N_9451);
xnor U11496 (N_11496,N_8298,N_8440);
or U11497 (N_11497,N_7855,N_9747);
and U11498 (N_11498,N_8048,N_7730);
nand U11499 (N_11499,N_7559,N_8304);
nand U11500 (N_11500,N_9535,N_7814);
nand U11501 (N_11501,N_7529,N_9974);
and U11502 (N_11502,N_7613,N_9714);
nor U11503 (N_11503,N_9719,N_8129);
xnor U11504 (N_11504,N_7969,N_9059);
or U11505 (N_11505,N_8557,N_8843);
nor U11506 (N_11506,N_9446,N_9101);
nor U11507 (N_11507,N_8270,N_9930);
or U11508 (N_11508,N_8756,N_7873);
or U11509 (N_11509,N_9239,N_8712);
and U11510 (N_11510,N_7542,N_8229);
nor U11511 (N_11511,N_8141,N_9247);
or U11512 (N_11512,N_7996,N_7905);
xor U11513 (N_11513,N_8678,N_8153);
xnor U11514 (N_11514,N_9532,N_7669);
xnor U11515 (N_11515,N_8773,N_8799);
and U11516 (N_11516,N_8943,N_9891);
and U11517 (N_11517,N_7999,N_9050);
and U11518 (N_11518,N_8417,N_8150);
and U11519 (N_11519,N_8332,N_7909);
nand U11520 (N_11520,N_9974,N_8866);
nor U11521 (N_11521,N_8504,N_7520);
xor U11522 (N_11522,N_7760,N_8270);
xor U11523 (N_11523,N_8087,N_8717);
or U11524 (N_11524,N_9069,N_8222);
nor U11525 (N_11525,N_8853,N_7965);
nor U11526 (N_11526,N_7547,N_9519);
and U11527 (N_11527,N_8986,N_9855);
nand U11528 (N_11528,N_7613,N_7504);
nand U11529 (N_11529,N_7508,N_8222);
nor U11530 (N_11530,N_9742,N_7611);
nor U11531 (N_11531,N_8096,N_9378);
and U11532 (N_11532,N_9687,N_9727);
nand U11533 (N_11533,N_9433,N_9718);
or U11534 (N_11534,N_8853,N_9559);
nand U11535 (N_11535,N_8081,N_8020);
nor U11536 (N_11536,N_7640,N_8790);
nand U11537 (N_11537,N_7761,N_8325);
nand U11538 (N_11538,N_9150,N_8986);
nor U11539 (N_11539,N_7597,N_8254);
and U11540 (N_11540,N_7698,N_9434);
xnor U11541 (N_11541,N_8835,N_8382);
nor U11542 (N_11542,N_9321,N_8158);
xor U11543 (N_11543,N_9904,N_9516);
and U11544 (N_11544,N_8356,N_9799);
nor U11545 (N_11545,N_9719,N_8631);
nand U11546 (N_11546,N_9842,N_9229);
or U11547 (N_11547,N_9258,N_8808);
xnor U11548 (N_11548,N_9323,N_9809);
nor U11549 (N_11549,N_8345,N_9387);
xnor U11550 (N_11550,N_8079,N_8757);
or U11551 (N_11551,N_9184,N_7640);
or U11552 (N_11552,N_9668,N_9916);
and U11553 (N_11553,N_8020,N_9954);
nand U11554 (N_11554,N_8564,N_8128);
xor U11555 (N_11555,N_8205,N_8624);
nor U11556 (N_11556,N_8796,N_9395);
nor U11557 (N_11557,N_7993,N_7678);
xnor U11558 (N_11558,N_8066,N_8779);
nor U11559 (N_11559,N_7633,N_7860);
nand U11560 (N_11560,N_9875,N_8557);
and U11561 (N_11561,N_9092,N_9355);
nor U11562 (N_11562,N_9198,N_8287);
or U11563 (N_11563,N_8808,N_7987);
nor U11564 (N_11564,N_9199,N_7593);
nor U11565 (N_11565,N_8950,N_9863);
nand U11566 (N_11566,N_7920,N_8308);
nor U11567 (N_11567,N_9872,N_8473);
nor U11568 (N_11568,N_7934,N_7803);
nor U11569 (N_11569,N_9765,N_7712);
nor U11570 (N_11570,N_8170,N_7810);
and U11571 (N_11571,N_8213,N_7580);
nor U11572 (N_11572,N_8260,N_9666);
and U11573 (N_11573,N_8112,N_7549);
xor U11574 (N_11574,N_8454,N_8715);
and U11575 (N_11575,N_7680,N_9611);
nor U11576 (N_11576,N_7592,N_9655);
nand U11577 (N_11577,N_8500,N_8846);
or U11578 (N_11578,N_8018,N_8353);
nand U11579 (N_11579,N_9427,N_9621);
or U11580 (N_11580,N_9591,N_8639);
and U11581 (N_11581,N_9598,N_9888);
nor U11582 (N_11582,N_9732,N_9718);
xnor U11583 (N_11583,N_7572,N_9307);
xor U11584 (N_11584,N_8925,N_7805);
or U11585 (N_11585,N_9454,N_9041);
xnor U11586 (N_11586,N_9192,N_9552);
xor U11587 (N_11587,N_8642,N_9846);
or U11588 (N_11588,N_7916,N_7709);
or U11589 (N_11589,N_9262,N_9312);
nand U11590 (N_11590,N_7938,N_7705);
or U11591 (N_11591,N_8045,N_9412);
xnor U11592 (N_11592,N_7821,N_8403);
xnor U11593 (N_11593,N_9999,N_8258);
xor U11594 (N_11594,N_9731,N_8473);
xnor U11595 (N_11595,N_8673,N_7921);
or U11596 (N_11596,N_9295,N_8192);
and U11597 (N_11597,N_8169,N_9713);
nor U11598 (N_11598,N_8523,N_9366);
nor U11599 (N_11599,N_9504,N_9124);
nand U11600 (N_11600,N_9586,N_8861);
xnor U11601 (N_11601,N_7751,N_9701);
nand U11602 (N_11602,N_7639,N_8012);
or U11603 (N_11603,N_9976,N_8774);
xnor U11604 (N_11604,N_8037,N_9626);
and U11605 (N_11605,N_9799,N_8629);
and U11606 (N_11606,N_9401,N_9683);
nand U11607 (N_11607,N_9464,N_9472);
or U11608 (N_11608,N_8706,N_9733);
or U11609 (N_11609,N_7886,N_8586);
nor U11610 (N_11610,N_8178,N_8289);
nor U11611 (N_11611,N_8382,N_9352);
xor U11612 (N_11612,N_9836,N_8835);
xor U11613 (N_11613,N_8895,N_8936);
nand U11614 (N_11614,N_9900,N_8364);
xor U11615 (N_11615,N_9654,N_8092);
and U11616 (N_11616,N_9207,N_9245);
or U11617 (N_11617,N_8093,N_8214);
and U11618 (N_11618,N_8851,N_7682);
nand U11619 (N_11619,N_9400,N_9287);
nor U11620 (N_11620,N_9048,N_8132);
xnor U11621 (N_11621,N_9061,N_9482);
or U11622 (N_11622,N_9385,N_9261);
and U11623 (N_11623,N_9817,N_8222);
nand U11624 (N_11624,N_8660,N_8986);
nor U11625 (N_11625,N_9374,N_8155);
nor U11626 (N_11626,N_7845,N_8757);
or U11627 (N_11627,N_9029,N_8343);
and U11628 (N_11628,N_8192,N_7789);
or U11629 (N_11629,N_7668,N_7804);
xnor U11630 (N_11630,N_9544,N_9598);
xnor U11631 (N_11631,N_8984,N_8468);
or U11632 (N_11632,N_9290,N_8979);
or U11633 (N_11633,N_9063,N_9379);
nor U11634 (N_11634,N_9526,N_8641);
nor U11635 (N_11635,N_8942,N_9923);
or U11636 (N_11636,N_9837,N_7976);
xor U11637 (N_11637,N_8943,N_8488);
and U11638 (N_11638,N_9718,N_8264);
xor U11639 (N_11639,N_9531,N_7745);
or U11640 (N_11640,N_9578,N_9503);
nand U11641 (N_11641,N_8921,N_8826);
xor U11642 (N_11642,N_7912,N_8328);
xnor U11643 (N_11643,N_7617,N_7896);
nand U11644 (N_11644,N_8156,N_7667);
xnor U11645 (N_11645,N_8391,N_9299);
nand U11646 (N_11646,N_8678,N_8277);
and U11647 (N_11647,N_9755,N_7584);
or U11648 (N_11648,N_9564,N_7557);
nor U11649 (N_11649,N_9058,N_8347);
and U11650 (N_11650,N_9531,N_9540);
or U11651 (N_11651,N_9548,N_9961);
xnor U11652 (N_11652,N_9966,N_7614);
and U11653 (N_11653,N_8020,N_7512);
nor U11654 (N_11654,N_7986,N_9379);
nand U11655 (N_11655,N_7521,N_9058);
xnor U11656 (N_11656,N_8058,N_7820);
nand U11657 (N_11657,N_7747,N_8865);
xnor U11658 (N_11658,N_9045,N_8742);
and U11659 (N_11659,N_7884,N_7893);
nor U11660 (N_11660,N_8427,N_8762);
xor U11661 (N_11661,N_9117,N_7927);
nor U11662 (N_11662,N_8384,N_9334);
nand U11663 (N_11663,N_9437,N_8833);
nor U11664 (N_11664,N_9848,N_8151);
nor U11665 (N_11665,N_9527,N_8978);
nor U11666 (N_11666,N_8142,N_8812);
xor U11667 (N_11667,N_7758,N_9098);
and U11668 (N_11668,N_9929,N_7773);
nor U11669 (N_11669,N_8836,N_8154);
nand U11670 (N_11670,N_8051,N_9363);
nand U11671 (N_11671,N_9043,N_9362);
nand U11672 (N_11672,N_9617,N_7791);
nor U11673 (N_11673,N_8423,N_9401);
and U11674 (N_11674,N_8587,N_8988);
or U11675 (N_11675,N_7618,N_7692);
xnor U11676 (N_11676,N_7986,N_9795);
nor U11677 (N_11677,N_8951,N_9070);
xor U11678 (N_11678,N_8896,N_8894);
nand U11679 (N_11679,N_7804,N_7654);
or U11680 (N_11680,N_9437,N_9352);
and U11681 (N_11681,N_8816,N_9982);
nand U11682 (N_11682,N_8605,N_9627);
xor U11683 (N_11683,N_7505,N_7912);
or U11684 (N_11684,N_9830,N_7706);
nand U11685 (N_11685,N_9489,N_8289);
nand U11686 (N_11686,N_8612,N_9072);
or U11687 (N_11687,N_7529,N_8235);
and U11688 (N_11688,N_9984,N_7669);
and U11689 (N_11689,N_9444,N_8692);
and U11690 (N_11690,N_9477,N_8491);
xor U11691 (N_11691,N_9774,N_9337);
and U11692 (N_11692,N_8651,N_9883);
nand U11693 (N_11693,N_8064,N_9592);
nor U11694 (N_11694,N_9659,N_9153);
xor U11695 (N_11695,N_7888,N_9971);
and U11696 (N_11696,N_9184,N_8151);
nor U11697 (N_11697,N_9979,N_9319);
nor U11698 (N_11698,N_9067,N_8109);
xnor U11699 (N_11699,N_8229,N_7625);
or U11700 (N_11700,N_9351,N_9018);
xnor U11701 (N_11701,N_7987,N_9397);
or U11702 (N_11702,N_7805,N_7849);
or U11703 (N_11703,N_9019,N_8687);
and U11704 (N_11704,N_9064,N_9192);
nand U11705 (N_11705,N_8835,N_9529);
nor U11706 (N_11706,N_9035,N_7699);
nor U11707 (N_11707,N_9159,N_9101);
nand U11708 (N_11708,N_8519,N_9762);
or U11709 (N_11709,N_8389,N_9540);
nand U11710 (N_11710,N_9332,N_7617);
xnor U11711 (N_11711,N_9885,N_9600);
and U11712 (N_11712,N_8702,N_9544);
or U11713 (N_11713,N_9909,N_8219);
xor U11714 (N_11714,N_9322,N_9365);
xor U11715 (N_11715,N_9009,N_7988);
xnor U11716 (N_11716,N_9859,N_7710);
nor U11717 (N_11717,N_8437,N_8985);
or U11718 (N_11718,N_7567,N_8601);
or U11719 (N_11719,N_8541,N_9814);
or U11720 (N_11720,N_8490,N_8009);
and U11721 (N_11721,N_7825,N_8315);
or U11722 (N_11722,N_7795,N_7953);
and U11723 (N_11723,N_7860,N_8113);
xnor U11724 (N_11724,N_9451,N_9490);
and U11725 (N_11725,N_7898,N_9046);
nand U11726 (N_11726,N_7693,N_8696);
or U11727 (N_11727,N_9783,N_7600);
nor U11728 (N_11728,N_9181,N_9628);
and U11729 (N_11729,N_9417,N_9685);
nand U11730 (N_11730,N_9951,N_8812);
nor U11731 (N_11731,N_9152,N_9950);
xnor U11732 (N_11732,N_8480,N_9387);
nand U11733 (N_11733,N_8302,N_8623);
or U11734 (N_11734,N_9810,N_7924);
and U11735 (N_11735,N_8285,N_8282);
nor U11736 (N_11736,N_8906,N_9505);
xor U11737 (N_11737,N_9446,N_8635);
or U11738 (N_11738,N_8351,N_7565);
xnor U11739 (N_11739,N_9207,N_8151);
xor U11740 (N_11740,N_9332,N_8693);
nand U11741 (N_11741,N_8970,N_8651);
xor U11742 (N_11742,N_9256,N_9937);
nor U11743 (N_11743,N_8684,N_8896);
nor U11744 (N_11744,N_9479,N_9248);
nand U11745 (N_11745,N_9039,N_7734);
xor U11746 (N_11746,N_8377,N_9999);
xor U11747 (N_11747,N_8753,N_7543);
nand U11748 (N_11748,N_7965,N_7931);
xnor U11749 (N_11749,N_8661,N_8279);
and U11750 (N_11750,N_9647,N_8020);
nand U11751 (N_11751,N_9962,N_8801);
nor U11752 (N_11752,N_8296,N_8391);
or U11753 (N_11753,N_9999,N_7540);
nand U11754 (N_11754,N_9221,N_8337);
nand U11755 (N_11755,N_9866,N_9077);
xor U11756 (N_11756,N_8874,N_9967);
nor U11757 (N_11757,N_8961,N_8766);
nor U11758 (N_11758,N_7774,N_7889);
and U11759 (N_11759,N_8060,N_8789);
and U11760 (N_11760,N_7674,N_7959);
nor U11761 (N_11761,N_7908,N_8026);
xor U11762 (N_11762,N_7923,N_7924);
xnor U11763 (N_11763,N_9976,N_7658);
xor U11764 (N_11764,N_9042,N_8998);
or U11765 (N_11765,N_7563,N_8673);
xor U11766 (N_11766,N_9096,N_8162);
xnor U11767 (N_11767,N_8485,N_9511);
xnor U11768 (N_11768,N_7534,N_8514);
and U11769 (N_11769,N_8908,N_7863);
or U11770 (N_11770,N_7990,N_8534);
nand U11771 (N_11771,N_9050,N_8270);
and U11772 (N_11772,N_9999,N_7708);
and U11773 (N_11773,N_8757,N_7747);
nor U11774 (N_11774,N_7945,N_7654);
xnor U11775 (N_11775,N_7889,N_9017);
xnor U11776 (N_11776,N_9281,N_9637);
xor U11777 (N_11777,N_9984,N_9550);
and U11778 (N_11778,N_9460,N_7969);
nor U11779 (N_11779,N_7671,N_8860);
nand U11780 (N_11780,N_8555,N_8610);
xor U11781 (N_11781,N_9489,N_7847);
and U11782 (N_11782,N_9882,N_7870);
xnor U11783 (N_11783,N_7984,N_7998);
nand U11784 (N_11784,N_8139,N_9513);
or U11785 (N_11785,N_9817,N_8288);
and U11786 (N_11786,N_8036,N_7868);
xor U11787 (N_11787,N_7706,N_9241);
xnor U11788 (N_11788,N_8670,N_8455);
nor U11789 (N_11789,N_9669,N_8138);
xor U11790 (N_11790,N_9170,N_8020);
xnor U11791 (N_11791,N_9666,N_9028);
nor U11792 (N_11792,N_9535,N_7671);
and U11793 (N_11793,N_7800,N_8361);
nand U11794 (N_11794,N_9887,N_9804);
xnor U11795 (N_11795,N_7619,N_9034);
or U11796 (N_11796,N_9315,N_8654);
or U11797 (N_11797,N_9961,N_8996);
or U11798 (N_11798,N_8576,N_8300);
nand U11799 (N_11799,N_9008,N_9901);
and U11800 (N_11800,N_9874,N_9924);
xnor U11801 (N_11801,N_8726,N_8225);
and U11802 (N_11802,N_8888,N_9687);
or U11803 (N_11803,N_9925,N_8315);
or U11804 (N_11804,N_7891,N_9399);
and U11805 (N_11805,N_7867,N_8964);
and U11806 (N_11806,N_9327,N_8888);
nor U11807 (N_11807,N_7660,N_8526);
xor U11808 (N_11808,N_8583,N_8115);
nor U11809 (N_11809,N_7549,N_7554);
or U11810 (N_11810,N_9767,N_7547);
nand U11811 (N_11811,N_9239,N_7677);
xnor U11812 (N_11812,N_9151,N_8062);
nor U11813 (N_11813,N_8684,N_8846);
nor U11814 (N_11814,N_8948,N_8483);
and U11815 (N_11815,N_9715,N_7558);
and U11816 (N_11816,N_9320,N_8238);
or U11817 (N_11817,N_9048,N_8126);
and U11818 (N_11818,N_9798,N_9840);
or U11819 (N_11819,N_7542,N_7555);
nor U11820 (N_11820,N_8029,N_8964);
xnor U11821 (N_11821,N_9900,N_9311);
nor U11822 (N_11822,N_8611,N_8352);
or U11823 (N_11823,N_9258,N_7981);
xor U11824 (N_11824,N_7733,N_9070);
or U11825 (N_11825,N_8748,N_9168);
nand U11826 (N_11826,N_9204,N_7653);
xnor U11827 (N_11827,N_8054,N_8445);
or U11828 (N_11828,N_9141,N_9352);
nor U11829 (N_11829,N_7850,N_8214);
and U11830 (N_11830,N_8606,N_9275);
nand U11831 (N_11831,N_9793,N_9151);
and U11832 (N_11832,N_7554,N_8977);
or U11833 (N_11833,N_7551,N_8627);
nor U11834 (N_11834,N_8266,N_9946);
xor U11835 (N_11835,N_7950,N_7927);
and U11836 (N_11836,N_8193,N_8586);
and U11837 (N_11837,N_8602,N_9477);
xor U11838 (N_11838,N_8104,N_9582);
or U11839 (N_11839,N_7875,N_9039);
xnor U11840 (N_11840,N_8856,N_8905);
xnor U11841 (N_11841,N_8436,N_8128);
nor U11842 (N_11842,N_9296,N_8409);
nand U11843 (N_11843,N_7934,N_9912);
and U11844 (N_11844,N_8821,N_9266);
nor U11845 (N_11845,N_7581,N_7883);
and U11846 (N_11846,N_9526,N_9428);
and U11847 (N_11847,N_9247,N_8856);
nand U11848 (N_11848,N_8171,N_8027);
nand U11849 (N_11849,N_9340,N_7692);
nand U11850 (N_11850,N_9005,N_8559);
and U11851 (N_11851,N_9676,N_9030);
or U11852 (N_11852,N_8552,N_8746);
nor U11853 (N_11853,N_7866,N_9775);
xor U11854 (N_11854,N_9123,N_8627);
nor U11855 (N_11855,N_8936,N_7917);
or U11856 (N_11856,N_9055,N_8358);
or U11857 (N_11857,N_8446,N_9790);
nor U11858 (N_11858,N_8283,N_8761);
xnor U11859 (N_11859,N_7992,N_8285);
and U11860 (N_11860,N_9592,N_9780);
nor U11861 (N_11861,N_9179,N_8435);
or U11862 (N_11862,N_9402,N_7689);
nor U11863 (N_11863,N_7695,N_8069);
and U11864 (N_11864,N_8760,N_8590);
or U11865 (N_11865,N_9262,N_8236);
or U11866 (N_11866,N_9804,N_8063);
nand U11867 (N_11867,N_7533,N_8399);
nor U11868 (N_11868,N_9528,N_9834);
nor U11869 (N_11869,N_8445,N_9706);
nor U11870 (N_11870,N_9283,N_9287);
nand U11871 (N_11871,N_7812,N_7627);
nor U11872 (N_11872,N_8609,N_9706);
and U11873 (N_11873,N_8969,N_9483);
nor U11874 (N_11874,N_8018,N_8267);
or U11875 (N_11875,N_9152,N_7828);
or U11876 (N_11876,N_8715,N_7979);
or U11877 (N_11877,N_8130,N_9985);
nor U11878 (N_11878,N_8713,N_9346);
xor U11879 (N_11879,N_8646,N_9776);
or U11880 (N_11880,N_9572,N_9763);
nand U11881 (N_11881,N_8048,N_8675);
or U11882 (N_11882,N_9524,N_9893);
nor U11883 (N_11883,N_9858,N_9859);
nor U11884 (N_11884,N_7586,N_7812);
xnor U11885 (N_11885,N_8389,N_7628);
or U11886 (N_11886,N_9719,N_9402);
and U11887 (N_11887,N_8353,N_7529);
nor U11888 (N_11888,N_8591,N_8617);
nor U11889 (N_11889,N_8815,N_9470);
or U11890 (N_11890,N_7686,N_8357);
or U11891 (N_11891,N_9323,N_8480);
nand U11892 (N_11892,N_9578,N_7661);
xor U11893 (N_11893,N_8441,N_8836);
or U11894 (N_11894,N_8887,N_8291);
nor U11895 (N_11895,N_8791,N_9069);
or U11896 (N_11896,N_9646,N_8414);
nand U11897 (N_11897,N_8746,N_9311);
nand U11898 (N_11898,N_9839,N_9745);
xor U11899 (N_11899,N_8173,N_8772);
nand U11900 (N_11900,N_8175,N_8497);
or U11901 (N_11901,N_8361,N_8651);
and U11902 (N_11902,N_8629,N_8768);
nor U11903 (N_11903,N_8477,N_9375);
nor U11904 (N_11904,N_8199,N_9427);
or U11905 (N_11905,N_9607,N_7558);
or U11906 (N_11906,N_9319,N_9244);
nor U11907 (N_11907,N_9880,N_7503);
xor U11908 (N_11908,N_8400,N_8999);
nor U11909 (N_11909,N_8526,N_7942);
nand U11910 (N_11910,N_8307,N_9595);
and U11911 (N_11911,N_9891,N_9734);
nor U11912 (N_11912,N_8234,N_7719);
nor U11913 (N_11913,N_9113,N_9911);
nand U11914 (N_11914,N_9122,N_8869);
nand U11915 (N_11915,N_8611,N_9396);
nand U11916 (N_11916,N_9368,N_8924);
xor U11917 (N_11917,N_7745,N_9662);
or U11918 (N_11918,N_7826,N_8783);
and U11919 (N_11919,N_9682,N_8951);
or U11920 (N_11920,N_9848,N_7949);
nor U11921 (N_11921,N_8120,N_8539);
nor U11922 (N_11922,N_8546,N_7728);
nand U11923 (N_11923,N_8112,N_9456);
xnor U11924 (N_11924,N_7788,N_8224);
xnor U11925 (N_11925,N_9440,N_9364);
xor U11926 (N_11926,N_7648,N_7524);
xnor U11927 (N_11927,N_8923,N_8437);
xor U11928 (N_11928,N_7789,N_8477);
or U11929 (N_11929,N_8529,N_8979);
and U11930 (N_11930,N_9186,N_8498);
and U11931 (N_11931,N_8359,N_9195);
nand U11932 (N_11932,N_8619,N_8809);
nor U11933 (N_11933,N_8626,N_8222);
xor U11934 (N_11934,N_9449,N_9626);
and U11935 (N_11935,N_7812,N_7564);
nor U11936 (N_11936,N_9804,N_9864);
and U11937 (N_11937,N_8176,N_9559);
xor U11938 (N_11938,N_8088,N_9662);
nor U11939 (N_11939,N_9053,N_9042);
or U11940 (N_11940,N_9275,N_8063);
xnor U11941 (N_11941,N_9430,N_9254);
nand U11942 (N_11942,N_7630,N_7507);
nand U11943 (N_11943,N_7901,N_8588);
and U11944 (N_11944,N_8163,N_8809);
and U11945 (N_11945,N_9415,N_9953);
xor U11946 (N_11946,N_8695,N_9701);
nand U11947 (N_11947,N_8861,N_7521);
nor U11948 (N_11948,N_8001,N_8983);
nor U11949 (N_11949,N_8407,N_8415);
or U11950 (N_11950,N_9510,N_8207);
nand U11951 (N_11951,N_8726,N_7596);
or U11952 (N_11952,N_8584,N_8953);
and U11953 (N_11953,N_8037,N_7758);
or U11954 (N_11954,N_8814,N_8691);
xnor U11955 (N_11955,N_7719,N_7865);
nand U11956 (N_11956,N_9746,N_8564);
xnor U11957 (N_11957,N_8190,N_8469);
and U11958 (N_11958,N_8996,N_7975);
or U11959 (N_11959,N_8137,N_9457);
xor U11960 (N_11960,N_9510,N_8345);
nor U11961 (N_11961,N_8080,N_9073);
nand U11962 (N_11962,N_9487,N_8353);
nand U11963 (N_11963,N_9080,N_9708);
xor U11964 (N_11964,N_7754,N_9561);
xor U11965 (N_11965,N_7923,N_8410);
nand U11966 (N_11966,N_7553,N_9773);
nand U11967 (N_11967,N_9225,N_8634);
xor U11968 (N_11968,N_7717,N_8521);
xnor U11969 (N_11969,N_9417,N_8567);
and U11970 (N_11970,N_8598,N_8055);
or U11971 (N_11971,N_8289,N_7735);
nand U11972 (N_11972,N_9334,N_9242);
and U11973 (N_11973,N_9809,N_8695);
nor U11974 (N_11974,N_8719,N_8802);
xnor U11975 (N_11975,N_9931,N_8998);
and U11976 (N_11976,N_7885,N_9161);
and U11977 (N_11977,N_9526,N_8379);
and U11978 (N_11978,N_8245,N_7679);
nand U11979 (N_11979,N_7696,N_8060);
and U11980 (N_11980,N_9172,N_8225);
xnor U11981 (N_11981,N_8392,N_8633);
nand U11982 (N_11982,N_8126,N_8200);
and U11983 (N_11983,N_9030,N_8997);
and U11984 (N_11984,N_9466,N_8229);
nand U11985 (N_11985,N_9367,N_8965);
nand U11986 (N_11986,N_9027,N_7906);
and U11987 (N_11987,N_9591,N_9143);
nor U11988 (N_11988,N_8093,N_8000);
nor U11989 (N_11989,N_8302,N_7952);
and U11990 (N_11990,N_8181,N_7967);
nor U11991 (N_11991,N_8595,N_9654);
xnor U11992 (N_11992,N_9773,N_9078);
nand U11993 (N_11993,N_9639,N_9249);
nand U11994 (N_11994,N_9983,N_8804);
nor U11995 (N_11995,N_7972,N_8096);
or U11996 (N_11996,N_9569,N_8221);
xnor U11997 (N_11997,N_8526,N_7535);
nand U11998 (N_11998,N_7880,N_7727);
xor U11999 (N_11999,N_7661,N_9836);
and U12000 (N_12000,N_7882,N_9367);
xnor U12001 (N_12001,N_8798,N_8537);
nor U12002 (N_12002,N_8176,N_9615);
or U12003 (N_12003,N_8652,N_8091);
nand U12004 (N_12004,N_9626,N_9874);
xor U12005 (N_12005,N_8069,N_9662);
nand U12006 (N_12006,N_9608,N_9884);
or U12007 (N_12007,N_8801,N_7867);
nand U12008 (N_12008,N_9557,N_8942);
nand U12009 (N_12009,N_8804,N_9741);
and U12010 (N_12010,N_9443,N_9881);
and U12011 (N_12011,N_9728,N_8080);
nor U12012 (N_12012,N_8892,N_9012);
nor U12013 (N_12013,N_8513,N_9517);
and U12014 (N_12014,N_9568,N_8397);
or U12015 (N_12015,N_8139,N_9701);
or U12016 (N_12016,N_8923,N_9389);
or U12017 (N_12017,N_8761,N_8789);
and U12018 (N_12018,N_7857,N_7758);
nand U12019 (N_12019,N_7722,N_9888);
xor U12020 (N_12020,N_7836,N_8484);
xnor U12021 (N_12021,N_8193,N_8210);
xnor U12022 (N_12022,N_7784,N_9745);
nand U12023 (N_12023,N_8140,N_8161);
or U12024 (N_12024,N_9953,N_8257);
nand U12025 (N_12025,N_9423,N_9980);
nor U12026 (N_12026,N_7806,N_9847);
xnor U12027 (N_12027,N_7753,N_9337);
and U12028 (N_12028,N_8870,N_9894);
nand U12029 (N_12029,N_9336,N_8315);
xnor U12030 (N_12030,N_8606,N_9353);
and U12031 (N_12031,N_9242,N_9508);
or U12032 (N_12032,N_9328,N_9755);
nand U12033 (N_12033,N_8648,N_8340);
and U12034 (N_12034,N_9572,N_8252);
xor U12035 (N_12035,N_9790,N_8714);
nand U12036 (N_12036,N_9986,N_9452);
nand U12037 (N_12037,N_8078,N_9646);
xor U12038 (N_12038,N_9687,N_9269);
and U12039 (N_12039,N_9695,N_8073);
and U12040 (N_12040,N_8739,N_8820);
or U12041 (N_12041,N_8709,N_9010);
or U12042 (N_12042,N_9477,N_9051);
nand U12043 (N_12043,N_9487,N_9861);
or U12044 (N_12044,N_9826,N_9675);
or U12045 (N_12045,N_9784,N_9920);
xor U12046 (N_12046,N_7576,N_7601);
xor U12047 (N_12047,N_8676,N_9196);
and U12048 (N_12048,N_7825,N_9018);
nor U12049 (N_12049,N_8617,N_9717);
and U12050 (N_12050,N_9392,N_8783);
and U12051 (N_12051,N_9723,N_8144);
xor U12052 (N_12052,N_9921,N_9995);
xnor U12053 (N_12053,N_9238,N_7975);
nand U12054 (N_12054,N_8800,N_9771);
xnor U12055 (N_12055,N_9968,N_9701);
and U12056 (N_12056,N_9248,N_8436);
nor U12057 (N_12057,N_8708,N_9174);
nand U12058 (N_12058,N_7965,N_9802);
xnor U12059 (N_12059,N_9484,N_7521);
nor U12060 (N_12060,N_7841,N_8380);
or U12061 (N_12061,N_9394,N_8814);
nand U12062 (N_12062,N_9264,N_9709);
nor U12063 (N_12063,N_7937,N_8908);
and U12064 (N_12064,N_9593,N_9705);
or U12065 (N_12065,N_9383,N_9834);
nand U12066 (N_12066,N_8493,N_9766);
and U12067 (N_12067,N_8932,N_8601);
and U12068 (N_12068,N_7684,N_8451);
nand U12069 (N_12069,N_8694,N_9716);
nor U12070 (N_12070,N_9836,N_8359);
and U12071 (N_12071,N_8668,N_7600);
xnor U12072 (N_12072,N_9334,N_7909);
and U12073 (N_12073,N_9920,N_8097);
and U12074 (N_12074,N_8400,N_7706);
or U12075 (N_12075,N_9372,N_8397);
and U12076 (N_12076,N_9822,N_8795);
nand U12077 (N_12077,N_9156,N_9808);
nor U12078 (N_12078,N_9176,N_9152);
nor U12079 (N_12079,N_9731,N_7622);
and U12080 (N_12080,N_9800,N_9393);
nand U12081 (N_12081,N_9368,N_7845);
nor U12082 (N_12082,N_9467,N_8628);
nor U12083 (N_12083,N_8835,N_8060);
or U12084 (N_12084,N_8798,N_8052);
xnor U12085 (N_12085,N_8954,N_9094);
or U12086 (N_12086,N_8442,N_9382);
nor U12087 (N_12087,N_8380,N_8670);
nor U12088 (N_12088,N_8375,N_7914);
nor U12089 (N_12089,N_9584,N_9999);
xnor U12090 (N_12090,N_9657,N_8759);
nand U12091 (N_12091,N_7871,N_9835);
nor U12092 (N_12092,N_8653,N_7858);
and U12093 (N_12093,N_8664,N_9556);
nor U12094 (N_12094,N_7738,N_8514);
and U12095 (N_12095,N_9214,N_7579);
or U12096 (N_12096,N_8957,N_7848);
nor U12097 (N_12097,N_8600,N_9180);
nand U12098 (N_12098,N_9576,N_9532);
nor U12099 (N_12099,N_9121,N_9393);
or U12100 (N_12100,N_9612,N_7518);
nand U12101 (N_12101,N_8309,N_8257);
xor U12102 (N_12102,N_9653,N_7689);
and U12103 (N_12103,N_7596,N_7535);
nor U12104 (N_12104,N_9002,N_7851);
xor U12105 (N_12105,N_8044,N_7814);
xnor U12106 (N_12106,N_9477,N_8314);
nand U12107 (N_12107,N_9757,N_8503);
and U12108 (N_12108,N_9014,N_8277);
or U12109 (N_12109,N_9296,N_9798);
nor U12110 (N_12110,N_9327,N_8129);
or U12111 (N_12111,N_8385,N_9359);
nand U12112 (N_12112,N_7541,N_7980);
and U12113 (N_12113,N_9830,N_8128);
nor U12114 (N_12114,N_7911,N_8522);
xor U12115 (N_12115,N_7789,N_9732);
nand U12116 (N_12116,N_8170,N_8367);
or U12117 (N_12117,N_8966,N_9976);
xnor U12118 (N_12118,N_7535,N_9397);
and U12119 (N_12119,N_8233,N_8380);
xor U12120 (N_12120,N_8593,N_9844);
nor U12121 (N_12121,N_8516,N_9156);
nor U12122 (N_12122,N_8574,N_9881);
nor U12123 (N_12123,N_9588,N_8628);
and U12124 (N_12124,N_9690,N_8811);
and U12125 (N_12125,N_8920,N_8855);
and U12126 (N_12126,N_7883,N_8780);
nor U12127 (N_12127,N_9336,N_8294);
nor U12128 (N_12128,N_9280,N_8417);
or U12129 (N_12129,N_9868,N_9354);
nor U12130 (N_12130,N_8257,N_7884);
xor U12131 (N_12131,N_9485,N_8664);
nor U12132 (N_12132,N_9560,N_9409);
xor U12133 (N_12133,N_9338,N_8026);
nor U12134 (N_12134,N_9659,N_8952);
nor U12135 (N_12135,N_9944,N_9433);
nor U12136 (N_12136,N_8053,N_7957);
nor U12137 (N_12137,N_8309,N_8382);
or U12138 (N_12138,N_7876,N_8127);
or U12139 (N_12139,N_8760,N_8840);
and U12140 (N_12140,N_8919,N_8957);
and U12141 (N_12141,N_9874,N_8485);
and U12142 (N_12142,N_9082,N_7534);
and U12143 (N_12143,N_7910,N_9898);
nand U12144 (N_12144,N_7552,N_7798);
and U12145 (N_12145,N_8560,N_7980);
or U12146 (N_12146,N_8016,N_7652);
xor U12147 (N_12147,N_9585,N_9177);
or U12148 (N_12148,N_7650,N_7988);
nand U12149 (N_12149,N_8251,N_9058);
nor U12150 (N_12150,N_8506,N_7503);
and U12151 (N_12151,N_7629,N_9276);
nor U12152 (N_12152,N_7999,N_8909);
or U12153 (N_12153,N_8097,N_8860);
and U12154 (N_12154,N_8446,N_9414);
xor U12155 (N_12155,N_9995,N_8805);
nor U12156 (N_12156,N_9077,N_9059);
or U12157 (N_12157,N_8579,N_9592);
and U12158 (N_12158,N_7881,N_8161);
and U12159 (N_12159,N_8069,N_8353);
nor U12160 (N_12160,N_8745,N_8069);
and U12161 (N_12161,N_8955,N_7502);
nand U12162 (N_12162,N_7970,N_9867);
nor U12163 (N_12163,N_8266,N_7567);
nand U12164 (N_12164,N_7901,N_9896);
or U12165 (N_12165,N_9239,N_7943);
and U12166 (N_12166,N_8200,N_9094);
or U12167 (N_12167,N_8048,N_7933);
and U12168 (N_12168,N_8703,N_8767);
or U12169 (N_12169,N_8771,N_8661);
and U12170 (N_12170,N_8972,N_8174);
or U12171 (N_12171,N_8728,N_8304);
nand U12172 (N_12172,N_9121,N_8117);
and U12173 (N_12173,N_7510,N_9788);
or U12174 (N_12174,N_8880,N_8114);
or U12175 (N_12175,N_9606,N_9683);
or U12176 (N_12176,N_7857,N_7739);
and U12177 (N_12177,N_8704,N_9757);
and U12178 (N_12178,N_8868,N_7502);
nand U12179 (N_12179,N_8367,N_8971);
nor U12180 (N_12180,N_7929,N_7757);
or U12181 (N_12181,N_8731,N_8106);
xnor U12182 (N_12182,N_8485,N_7870);
xnor U12183 (N_12183,N_9318,N_9710);
and U12184 (N_12184,N_9713,N_9683);
nand U12185 (N_12185,N_9026,N_9688);
or U12186 (N_12186,N_7787,N_8786);
and U12187 (N_12187,N_7828,N_8210);
nand U12188 (N_12188,N_8334,N_7796);
xor U12189 (N_12189,N_8849,N_9698);
nand U12190 (N_12190,N_8093,N_8354);
nand U12191 (N_12191,N_7935,N_9346);
nand U12192 (N_12192,N_9762,N_7780);
nor U12193 (N_12193,N_9767,N_8228);
xor U12194 (N_12194,N_8314,N_8493);
or U12195 (N_12195,N_7535,N_8552);
and U12196 (N_12196,N_7712,N_8718);
and U12197 (N_12197,N_9395,N_9740);
or U12198 (N_12198,N_8267,N_9331);
and U12199 (N_12199,N_9331,N_9896);
xor U12200 (N_12200,N_9620,N_8905);
and U12201 (N_12201,N_9307,N_7797);
xnor U12202 (N_12202,N_9757,N_8287);
or U12203 (N_12203,N_7574,N_8416);
nor U12204 (N_12204,N_9145,N_8047);
or U12205 (N_12205,N_8107,N_9179);
nor U12206 (N_12206,N_9765,N_9576);
nand U12207 (N_12207,N_7961,N_8980);
xnor U12208 (N_12208,N_9787,N_9431);
or U12209 (N_12209,N_8313,N_9444);
or U12210 (N_12210,N_7838,N_8482);
and U12211 (N_12211,N_9558,N_8245);
and U12212 (N_12212,N_7631,N_7991);
nand U12213 (N_12213,N_9987,N_7702);
nand U12214 (N_12214,N_8920,N_9038);
or U12215 (N_12215,N_9199,N_9859);
or U12216 (N_12216,N_9817,N_8441);
xnor U12217 (N_12217,N_9566,N_7760);
nand U12218 (N_12218,N_7954,N_9242);
nor U12219 (N_12219,N_9517,N_9408);
nand U12220 (N_12220,N_8684,N_8169);
nand U12221 (N_12221,N_8068,N_8995);
nor U12222 (N_12222,N_9042,N_8213);
nor U12223 (N_12223,N_8727,N_8580);
or U12224 (N_12224,N_8681,N_9231);
nand U12225 (N_12225,N_9110,N_9510);
or U12226 (N_12226,N_8948,N_9781);
and U12227 (N_12227,N_8038,N_7733);
or U12228 (N_12228,N_7742,N_7962);
nor U12229 (N_12229,N_9708,N_7790);
nand U12230 (N_12230,N_7627,N_9853);
xnor U12231 (N_12231,N_8246,N_8673);
or U12232 (N_12232,N_8247,N_9982);
or U12233 (N_12233,N_9610,N_7869);
and U12234 (N_12234,N_8415,N_9700);
or U12235 (N_12235,N_9053,N_8002);
nand U12236 (N_12236,N_9875,N_8169);
xnor U12237 (N_12237,N_9920,N_8884);
xnor U12238 (N_12238,N_7755,N_8452);
and U12239 (N_12239,N_9894,N_9063);
nor U12240 (N_12240,N_8831,N_9185);
xor U12241 (N_12241,N_8118,N_9843);
nor U12242 (N_12242,N_9970,N_8500);
or U12243 (N_12243,N_8296,N_8895);
nand U12244 (N_12244,N_9391,N_8523);
or U12245 (N_12245,N_7566,N_9922);
or U12246 (N_12246,N_9039,N_9802);
xnor U12247 (N_12247,N_9284,N_9797);
nand U12248 (N_12248,N_8756,N_8222);
and U12249 (N_12249,N_8330,N_8106);
nand U12250 (N_12250,N_9855,N_8250);
and U12251 (N_12251,N_9979,N_8634);
xnor U12252 (N_12252,N_8462,N_8458);
or U12253 (N_12253,N_8958,N_7635);
nand U12254 (N_12254,N_8189,N_7534);
or U12255 (N_12255,N_8335,N_7553);
or U12256 (N_12256,N_7839,N_9912);
and U12257 (N_12257,N_8685,N_7741);
nor U12258 (N_12258,N_8106,N_9907);
or U12259 (N_12259,N_7645,N_9349);
and U12260 (N_12260,N_8986,N_9613);
and U12261 (N_12261,N_7973,N_9996);
nand U12262 (N_12262,N_8538,N_7970);
xnor U12263 (N_12263,N_7930,N_8235);
nor U12264 (N_12264,N_7713,N_9122);
nand U12265 (N_12265,N_8126,N_9295);
xor U12266 (N_12266,N_8280,N_9956);
nand U12267 (N_12267,N_7939,N_8481);
or U12268 (N_12268,N_9672,N_7515);
nor U12269 (N_12269,N_8673,N_9566);
nor U12270 (N_12270,N_9368,N_9277);
and U12271 (N_12271,N_7759,N_7674);
xor U12272 (N_12272,N_8213,N_8160);
or U12273 (N_12273,N_8275,N_9022);
and U12274 (N_12274,N_7614,N_7735);
xnor U12275 (N_12275,N_9313,N_9267);
nand U12276 (N_12276,N_8368,N_9662);
nor U12277 (N_12277,N_8535,N_9832);
nand U12278 (N_12278,N_9599,N_9025);
and U12279 (N_12279,N_9743,N_8741);
nand U12280 (N_12280,N_9287,N_9694);
or U12281 (N_12281,N_8699,N_8797);
or U12282 (N_12282,N_9634,N_8515);
and U12283 (N_12283,N_8622,N_7575);
or U12284 (N_12284,N_9923,N_9252);
xnor U12285 (N_12285,N_9120,N_9873);
nand U12286 (N_12286,N_9364,N_9168);
nor U12287 (N_12287,N_8072,N_9856);
nand U12288 (N_12288,N_9014,N_8330);
nor U12289 (N_12289,N_9193,N_9709);
and U12290 (N_12290,N_8807,N_8484);
nand U12291 (N_12291,N_8956,N_8621);
nand U12292 (N_12292,N_9591,N_8005);
nor U12293 (N_12293,N_9690,N_8956);
and U12294 (N_12294,N_8850,N_8751);
xnor U12295 (N_12295,N_9153,N_8146);
nand U12296 (N_12296,N_8423,N_9380);
and U12297 (N_12297,N_8791,N_8473);
and U12298 (N_12298,N_8906,N_7917);
or U12299 (N_12299,N_7866,N_8315);
nor U12300 (N_12300,N_7926,N_8675);
nand U12301 (N_12301,N_8829,N_9836);
or U12302 (N_12302,N_9404,N_8618);
nand U12303 (N_12303,N_8610,N_9526);
nand U12304 (N_12304,N_9937,N_8021);
and U12305 (N_12305,N_8486,N_9326);
nor U12306 (N_12306,N_7537,N_8439);
and U12307 (N_12307,N_9940,N_9369);
nor U12308 (N_12308,N_9288,N_9421);
nand U12309 (N_12309,N_7776,N_8577);
nand U12310 (N_12310,N_8972,N_9692);
nand U12311 (N_12311,N_8851,N_9411);
xor U12312 (N_12312,N_8566,N_7593);
xor U12313 (N_12313,N_9586,N_9398);
and U12314 (N_12314,N_7596,N_9748);
nor U12315 (N_12315,N_7546,N_8953);
nor U12316 (N_12316,N_9040,N_9489);
nand U12317 (N_12317,N_8298,N_7578);
nand U12318 (N_12318,N_9447,N_8385);
and U12319 (N_12319,N_7503,N_8819);
or U12320 (N_12320,N_8742,N_9906);
nor U12321 (N_12321,N_7746,N_8678);
or U12322 (N_12322,N_9971,N_9126);
and U12323 (N_12323,N_9654,N_9760);
nor U12324 (N_12324,N_9641,N_8620);
nor U12325 (N_12325,N_9186,N_8732);
nand U12326 (N_12326,N_7560,N_8909);
or U12327 (N_12327,N_8279,N_7606);
nor U12328 (N_12328,N_7982,N_8366);
or U12329 (N_12329,N_8193,N_9176);
and U12330 (N_12330,N_7611,N_7957);
nand U12331 (N_12331,N_8023,N_9457);
and U12332 (N_12332,N_7853,N_9701);
nor U12333 (N_12333,N_9686,N_7890);
nand U12334 (N_12334,N_8964,N_8663);
nand U12335 (N_12335,N_8610,N_8803);
nor U12336 (N_12336,N_7551,N_7614);
or U12337 (N_12337,N_9744,N_8557);
nand U12338 (N_12338,N_8690,N_8065);
nand U12339 (N_12339,N_8144,N_7842);
nor U12340 (N_12340,N_9349,N_7915);
or U12341 (N_12341,N_9852,N_9765);
or U12342 (N_12342,N_7580,N_8196);
and U12343 (N_12343,N_7868,N_9978);
and U12344 (N_12344,N_9435,N_8268);
and U12345 (N_12345,N_8343,N_8356);
or U12346 (N_12346,N_7717,N_9042);
xor U12347 (N_12347,N_7627,N_9812);
nand U12348 (N_12348,N_8742,N_9511);
nor U12349 (N_12349,N_7946,N_8954);
nor U12350 (N_12350,N_8418,N_7584);
nor U12351 (N_12351,N_8346,N_9612);
or U12352 (N_12352,N_8296,N_7915);
xnor U12353 (N_12353,N_8489,N_9940);
xor U12354 (N_12354,N_9058,N_7766);
nand U12355 (N_12355,N_9492,N_9812);
xnor U12356 (N_12356,N_8343,N_7718);
nand U12357 (N_12357,N_8914,N_9530);
nor U12358 (N_12358,N_9886,N_9450);
or U12359 (N_12359,N_9399,N_8185);
or U12360 (N_12360,N_7603,N_8240);
nand U12361 (N_12361,N_8126,N_9676);
nand U12362 (N_12362,N_9543,N_8294);
nand U12363 (N_12363,N_8177,N_9744);
and U12364 (N_12364,N_8513,N_9273);
nand U12365 (N_12365,N_8551,N_9441);
xor U12366 (N_12366,N_9110,N_7699);
or U12367 (N_12367,N_8389,N_8742);
and U12368 (N_12368,N_8985,N_8474);
nor U12369 (N_12369,N_9754,N_7789);
or U12370 (N_12370,N_9234,N_8183);
nand U12371 (N_12371,N_9301,N_9019);
or U12372 (N_12372,N_8501,N_9502);
nand U12373 (N_12373,N_8371,N_8134);
or U12374 (N_12374,N_9474,N_8610);
nor U12375 (N_12375,N_8025,N_8028);
or U12376 (N_12376,N_9667,N_8436);
xnor U12377 (N_12377,N_8194,N_9596);
or U12378 (N_12378,N_8075,N_9364);
nand U12379 (N_12379,N_8852,N_9795);
xnor U12380 (N_12380,N_8459,N_8217);
and U12381 (N_12381,N_8423,N_9141);
xnor U12382 (N_12382,N_9088,N_7803);
nand U12383 (N_12383,N_8160,N_9487);
nand U12384 (N_12384,N_9575,N_9398);
xor U12385 (N_12385,N_9445,N_9081);
xor U12386 (N_12386,N_8962,N_9568);
xor U12387 (N_12387,N_9503,N_9194);
and U12388 (N_12388,N_8546,N_9139);
nor U12389 (N_12389,N_9871,N_7655);
xor U12390 (N_12390,N_9131,N_9476);
nor U12391 (N_12391,N_7681,N_9562);
nand U12392 (N_12392,N_9909,N_9662);
and U12393 (N_12393,N_7924,N_9674);
xnor U12394 (N_12394,N_8359,N_7534);
or U12395 (N_12395,N_9492,N_8625);
nor U12396 (N_12396,N_8474,N_8439);
xnor U12397 (N_12397,N_9469,N_8033);
nor U12398 (N_12398,N_8326,N_9266);
nand U12399 (N_12399,N_8109,N_7657);
nor U12400 (N_12400,N_8150,N_9402);
or U12401 (N_12401,N_9923,N_8184);
xnor U12402 (N_12402,N_9187,N_9394);
and U12403 (N_12403,N_9759,N_8305);
nand U12404 (N_12404,N_9139,N_9599);
nand U12405 (N_12405,N_7590,N_9743);
nor U12406 (N_12406,N_9495,N_9071);
nand U12407 (N_12407,N_8570,N_7765);
or U12408 (N_12408,N_7615,N_8948);
nand U12409 (N_12409,N_9171,N_8936);
xor U12410 (N_12410,N_9045,N_9427);
xnor U12411 (N_12411,N_7993,N_9226);
and U12412 (N_12412,N_9573,N_8162);
nor U12413 (N_12413,N_8751,N_8599);
and U12414 (N_12414,N_7686,N_9300);
or U12415 (N_12415,N_8864,N_8432);
xnor U12416 (N_12416,N_7964,N_8581);
xnor U12417 (N_12417,N_7965,N_9599);
nor U12418 (N_12418,N_8450,N_8055);
nor U12419 (N_12419,N_9670,N_8280);
and U12420 (N_12420,N_9444,N_7692);
nor U12421 (N_12421,N_7691,N_7636);
nand U12422 (N_12422,N_8802,N_9870);
or U12423 (N_12423,N_9567,N_8541);
or U12424 (N_12424,N_7670,N_8830);
xnor U12425 (N_12425,N_8612,N_8528);
nand U12426 (N_12426,N_8259,N_9385);
nor U12427 (N_12427,N_9897,N_9111);
or U12428 (N_12428,N_8620,N_8169);
nand U12429 (N_12429,N_7967,N_9287);
nor U12430 (N_12430,N_8184,N_9033);
nand U12431 (N_12431,N_8738,N_9247);
and U12432 (N_12432,N_8758,N_8402);
and U12433 (N_12433,N_9792,N_8385);
nand U12434 (N_12434,N_9742,N_8811);
nand U12435 (N_12435,N_9933,N_8943);
xnor U12436 (N_12436,N_9954,N_9408);
or U12437 (N_12437,N_9035,N_9182);
and U12438 (N_12438,N_8862,N_9871);
and U12439 (N_12439,N_8590,N_9455);
xnor U12440 (N_12440,N_9900,N_9099);
nor U12441 (N_12441,N_8269,N_9301);
xnor U12442 (N_12442,N_7684,N_7872);
xnor U12443 (N_12443,N_7620,N_9624);
and U12444 (N_12444,N_9596,N_9445);
and U12445 (N_12445,N_7962,N_8308);
nor U12446 (N_12446,N_8309,N_9405);
nor U12447 (N_12447,N_9341,N_8474);
and U12448 (N_12448,N_8467,N_9465);
and U12449 (N_12449,N_9087,N_8394);
and U12450 (N_12450,N_8704,N_8205);
xnor U12451 (N_12451,N_7666,N_8432);
nand U12452 (N_12452,N_7767,N_9323);
or U12453 (N_12453,N_8379,N_9715);
or U12454 (N_12454,N_8879,N_7914);
and U12455 (N_12455,N_7995,N_9192);
xnor U12456 (N_12456,N_9389,N_9191);
nor U12457 (N_12457,N_7844,N_8602);
and U12458 (N_12458,N_8442,N_9687);
nand U12459 (N_12459,N_9055,N_8265);
or U12460 (N_12460,N_7739,N_9704);
or U12461 (N_12461,N_8347,N_7797);
xor U12462 (N_12462,N_9467,N_9616);
nor U12463 (N_12463,N_8971,N_8417);
or U12464 (N_12464,N_9881,N_9474);
and U12465 (N_12465,N_9038,N_9805);
or U12466 (N_12466,N_9948,N_8460);
or U12467 (N_12467,N_8191,N_8832);
nor U12468 (N_12468,N_7503,N_8159);
nor U12469 (N_12469,N_9815,N_9630);
nor U12470 (N_12470,N_8027,N_7678);
and U12471 (N_12471,N_9431,N_9163);
nor U12472 (N_12472,N_9575,N_9131);
and U12473 (N_12473,N_9565,N_9454);
nand U12474 (N_12474,N_8930,N_7663);
or U12475 (N_12475,N_9558,N_8171);
nor U12476 (N_12476,N_9402,N_8425);
nand U12477 (N_12477,N_8828,N_8383);
and U12478 (N_12478,N_9904,N_8737);
or U12479 (N_12479,N_9372,N_9166);
nor U12480 (N_12480,N_9661,N_9337);
nor U12481 (N_12481,N_8514,N_8484);
xor U12482 (N_12482,N_8086,N_9555);
nand U12483 (N_12483,N_9487,N_7653);
nand U12484 (N_12484,N_8385,N_9044);
xor U12485 (N_12485,N_7839,N_9770);
nor U12486 (N_12486,N_8942,N_9738);
and U12487 (N_12487,N_9744,N_7976);
xnor U12488 (N_12488,N_7542,N_8314);
nor U12489 (N_12489,N_9692,N_9557);
nand U12490 (N_12490,N_9554,N_9996);
xor U12491 (N_12491,N_9042,N_9056);
xnor U12492 (N_12492,N_7700,N_9574);
or U12493 (N_12493,N_8611,N_8847);
xor U12494 (N_12494,N_8523,N_8812);
xor U12495 (N_12495,N_8949,N_9153);
nor U12496 (N_12496,N_8936,N_8952);
xor U12497 (N_12497,N_8891,N_8454);
and U12498 (N_12498,N_9617,N_9687);
nor U12499 (N_12499,N_9124,N_8968);
nand U12500 (N_12500,N_11613,N_11487);
and U12501 (N_12501,N_10476,N_10047);
nor U12502 (N_12502,N_10541,N_10084);
and U12503 (N_12503,N_10037,N_11037);
and U12504 (N_12504,N_11745,N_10546);
or U12505 (N_12505,N_10358,N_12385);
xor U12506 (N_12506,N_10866,N_10748);
xnor U12507 (N_12507,N_10421,N_10780);
nand U12508 (N_12508,N_10096,N_10225);
nor U12509 (N_12509,N_10255,N_10584);
or U12510 (N_12510,N_11220,N_10191);
or U12511 (N_12511,N_12197,N_12348);
nand U12512 (N_12512,N_12148,N_12196);
nor U12513 (N_12513,N_10134,N_10574);
xor U12514 (N_12514,N_11917,N_11579);
and U12515 (N_12515,N_10439,N_10272);
and U12516 (N_12516,N_12422,N_11863);
nand U12517 (N_12517,N_12330,N_11359);
nand U12518 (N_12518,N_12134,N_10199);
or U12519 (N_12519,N_11654,N_10766);
and U12520 (N_12520,N_10934,N_10465);
nand U12521 (N_12521,N_10107,N_10741);
and U12522 (N_12522,N_11635,N_12103);
nor U12523 (N_12523,N_10553,N_10326);
and U12524 (N_12524,N_10391,N_11480);
xnor U12525 (N_12525,N_10052,N_12432);
nand U12526 (N_12526,N_11248,N_12256);
nand U12527 (N_12527,N_10538,N_11665);
nand U12528 (N_12528,N_11615,N_12358);
or U12529 (N_12529,N_11755,N_10186);
nand U12530 (N_12530,N_12277,N_10880);
xnor U12531 (N_12531,N_10147,N_10341);
xnor U12532 (N_12532,N_11992,N_11216);
or U12533 (N_12533,N_12396,N_10455);
nand U12534 (N_12534,N_10607,N_11908);
nor U12535 (N_12535,N_11943,N_10148);
xor U12536 (N_12536,N_10166,N_11746);
or U12537 (N_12537,N_11846,N_10975);
nor U12538 (N_12538,N_12125,N_11573);
nand U12539 (N_12539,N_11965,N_11970);
nand U12540 (N_12540,N_11675,N_10536);
nor U12541 (N_12541,N_10757,N_10935);
nor U12542 (N_12542,N_12364,N_10280);
or U12543 (N_12543,N_12313,N_10818);
xnor U12544 (N_12544,N_10817,N_10789);
and U12545 (N_12545,N_10240,N_11454);
or U12546 (N_12546,N_11088,N_10742);
and U12547 (N_12547,N_11121,N_11731);
nand U12548 (N_12548,N_11137,N_10839);
nand U12549 (N_12549,N_11086,N_11477);
nor U12550 (N_12550,N_11204,N_10704);
xnor U12551 (N_12551,N_10020,N_11829);
and U12552 (N_12552,N_11488,N_11663);
nand U12553 (N_12553,N_12319,N_11483);
nor U12554 (N_12554,N_10198,N_11647);
xor U12555 (N_12555,N_11624,N_10259);
and U12556 (N_12556,N_10964,N_11592);
or U12557 (N_12557,N_10786,N_12462);
nor U12558 (N_12558,N_11369,N_11447);
nor U12559 (N_12559,N_10236,N_10159);
nand U12560 (N_12560,N_11641,N_11761);
and U12561 (N_12561,N_11340,N_10699);
nand U12562 (N_12562,N_11017,N_10746);
xor U12563 (N_12563,N_11571,N_12060);
nor U12564 (N_12564,N_12048,N_11307);
nor U12565 (N_12565,N_11680,N_10090);
and U12566 (N_12566,N_10970,N_10739);
xnor U12567 (N_12567,N_12494,N_11628);
or U12568 (N_12568,N_12051,N_11182);
or U12569 (N_12569,N_10908,N_10302);
or U12570 (N_12570,N_11678,N_10734);
nor U12571 (N_12571,N_11486,N_11691);
or U12572 (N_12572,N_11374,N_11033);
xnor U12573 (N_12573,N_11219,N_10078);
and U12574 (N_12574,N_11365,N_12447);
nor U12575 (N_12575,N_12219,N_11253);
and U12576 (N_12576,N_10851,N_11223);
nor U12577 (N_12577,N_11566,N_11558);
xor U12578 (N_12578,N_11695,N_10565);
nand U12579 (N_12579,N_11116,N_12244);
nand U12580 (N_12580,N_10383,N_12053);
nand U12581 (N_12581,N_11740,N_12220);
xor U12582 (N_12582,N_11267,N_10234);
nor U12583 (N_12583,N_10070,N_11156);
nand U12584 (N_12584,N_12231,N_11881);
nand U12585 (N_12585,N_11031,N_11354);
nand U12586 (N_12586,N_12440,N_10622);
nor U12587 (N_12587,N_10625,N_11660);
nand U12588 (N_12588,N_12332,N_11471);
nand U12589 (N_12589,N_12105,N_11021);
or U12590 (N_12590,N_11569,N_12362);
and U12591 (N_12591,N_12002,N_10406);
nor U12592 (N_12592,N_12423,N_10129);
and U12593 (N_12593,N_11949,N_12446);
or U12594 (N_12594,N_11437,N_11952);
nand U12595 (N_12595,N_12482,N_12207);
nor U12596 (N_12596,N_11744,N_10710);
nor U12597 (N_12597,N_11562,N_11495);
nor U12598 (N_12598,N_12107,N_10106);
or U12599 (N_12599,N_10137,N_11777);
nand U12600 (N_12600,N_10123,N_12007);
nor U12601 (N_12601,N_10130,N_11318);
nor U12602 (N_12602,N_12340,N_10893);
nor U12603 (N_12603,N_10629,N_10097);
and U12604 (N_12604,N_11371,N_11742);
xor U12605 (N_12605,N_11986,N_12088);
xor U12606 (N_12606,N_12185,N_11699);
nand U12607 (N_12607,N_11728,N_11105);
xnor U12608 (N_12608,N_11854,N_10680);
nor U12609 (N_12609,N_11705,N_12343);
and U12610 (N_12610,N_11865,N_11337);
xor U12611 (N_12611,N_10454,N_11030);
xor U12612 (N_12612,N_11463,N_12056);
or U12613 (N_12613,N_10450,N_10400);
xnor U12614 (N_12614,N_11738,N_10953);
and U12615 (N_12615,N_12229,N_12467);
nor U12616 (N_12616,N_12089,N_12283);
nand U12617 (N_12617,N_11589,N_11912);
nand U12618 (N_12618,N_12085,N_11423);
or U12619 (N_12619,N_10585,N_11672);
or U12620 (N_12620,N_10060,N_10904);
or U12621 (N_12621,N_12486,N_11529);
and U12622 (N_12622,N_10493,N_12307);
and U12623 (N_12623,N_11377,N_10505);
or U12624 (N_12624,N_10411,N_10842);
nand U12625 (N_12625,N_10478,N_12435);
xnor U12626 (N_12626,N_10924,N_10248);
nand U12627 (N_12627,N_10775,N_11370);
and U12628 (N_12628,N_12475,N_10928);
xnor U12629 (N_12629,N_10164,N_11472);
xnor U12630 (N_12630,N_11298,N_10260);
nand U12631 (N_12631,N_12427,N_10050);
xor U12632 (N_12632,N_10188,N_11417);
xnor U12633 (N_12633,N_11736,N_11181);
and U12634 (N_12634,N_11297,N_11656);
xnor U12635 (N_12635,N_11481,N_11536);
nor U12636 (N_12636,N_10435,N_10937);
xnor U12637 (N_12637,N_12291,N_11773);
nand U12638 (N_12638,N_11963,N_10885);
and U12639 (N_12639,N_10049,N_12328);
nor U12640 (N_12640,N_12442,N_10602);
and U12641 (N_12641,N_10868,N_10600);
and U12642 (N_12642,N_11788,N_10808);
xor U12643 (N_12643,N_11391,N_11585);
or U12644 (N_12644,N_12320,N_12287);
nor U12645 (N_12645,N_10556,N_11351);
xor U12646 (N_12646,N_11467,N_10557);
nor U12647 (N_12647,N_11428,N_11382);
nor U12648 (N_12648,N_12177,N_11389);
xor U12649 (N_12649,N_10224,N_11543);
nor U12650 (N_12650,N_12428,N_11978);
nor U12651 (N_12651,N_10561,N_12111);
and U12652 (N_12652,N_12096,N_12221);
xor U12653 (N_12653,N_12081,N_11385);
nand U12654 (N_12654,N_10495,N_10196);
or U12655 (N_12655,N_10811,N_12157);
nor U12656 (N_12656,N_11233,N_10879);
nor U12657 (N_12657,N_12294,N_10145);
nand U12658 (N_12658,N_11140,N_11063);
xor U12659 (N_12659,N_11144,N_11878);
or U12660 (N_12660,N_11452,N_12175);
xnor U12661 (N_12661,N_11496,N_10061);
and U12662 (N_12662,N_11449,N_10407);
and U12663 (N_12663,N_11927,N_10008);
xor U12664 (N_12664,N_10163,N_10282);
xor U12665 (N_12665,N_10350,N_11526);
xor U12666 (N_12666,N_10017,N_10544);
xnor U12667 (N_12667,N_10484,N_12210);
nand U12668 (N_12668,N_11299,N_10679);
nand U12669 (N_12669,N_10362,N_11619);
nor U12670 (N_12670,N_12415,N_10591);
nor U12671 (N_12671,N_10183,N_11443);
nor U12672 (N_12672,N_10001,N_10870);
or U12673 (N_12673,N_11859,N_11826);
and U12674 (N_12674,N_11556,N_11231);
nor U12675 (N_12675,N_10313,N_10416);
or U12676 (N_12676,N_12091,N_10921);
xor U12677 (N_12677,N_10192,N_11876);
xor U12678 (N_12678,N_11520,N_12267);
nand U12679 (N_12679,N_10686,N_11686);
nand U12680 (N_12680,N_10624,N_11780);
and U12681 (N_12681,N_10731,N_10687);
nand U12682 (N_12682,N_11545,N_10216);
and U12683 (N_12683,N_12444,N_11507);
or U12684 (N_12684,N_10551,N_10628);
nor U12685 (N_12685,N_12372,N_11157);
nand U12686 (N_12686,N_11247,N_12420);
nand U12687 (N_12687,N_10357,N_11008);
and U12688 (N_12688,N_10141,N_11727);
and U12689 (N_12689,N_10048,N_11919);
or U12690 (N_12690,N_10366,N_12086);
xnor U12691 (N_12691,N_12241,N_11112);
xor U12692 (N_12692,N_10906,N_11295);
or U12693 (N_12693,N_10267,N_10284);
nor U12694 (N_12694,N_10896,N_11333);
nor U12695 (N_12695,N_11711,N_10000);
nand U12696 (N_12696,N_10269,N_10728);
or U12697 (N_12697,N_11990,N_10511);
and U12698 (N_12698,N_10709,N_10103);
and U12699 (N_12699,N_10570,N_11578);
nor U12700 (N_12700,N_10719,N_10480);
xnor U12701 (N_12701,N_11850,N_10499);
nand U12702 (N_12702,N_10669,N_11929);
or U12703 (N_12703,N_11830,N_12174);
nor U12704 (N_12704,N_10278,N_12335);
or U12705 (N_12705,N_10841,N_10189);
nand U12706 (N_12706,N_11768,N_10014);
or U12707 (N_12707,N_11099,N_12414);
xor U12708 (N_12708,N_10913,N_10577);
and U12709 (N_12709,N_10694,N_11683);
and U12710 (N_12710,N_12128,N_12416);
nor U12711 (N_12711,N_11089,N_11835);
xor U12712 (N_12712,N_11807,N_12278);
nor U12713 (N_12713,N_10412,N_11421);
xor U12714 (N_12714,N_11210,N_11614);
nand U12715 (N_12715,N_11873,N_10243);
nor U12716 (N_12716,N_11870,N_12226);
and U12717 (N_12717,N_10562,N_10093);
nor U12718 (N_12718,N_10079,N_11776);
nand U12719 (N_12719,N_10946,N_11898);
nor U12720 (N_12720,N_11276,N_12303);
nor U12721 (N_12721,N_10251,N_10344);
nor U12722 (N_12722,N_11796,N_12084);
xnor U12723 (N_12723,N_12457,N_11015);
or U12724 (N_12724,N_11726,N_11268);
nand U12725 (N_12725,N_10333,N_11386);
and U12726 (N_12726,N_11858,N_12190);
or U12727 (N_12727,N_11714,N_12222);
xnor U12728 (N_12728,N_10816,N_10005);
nor U12729 (N_12729,N_11430,N_10914);
or U12730 (N_12730,N_10316,N_11152);
xor U12731 (N_12731,N_11759,N_11213);
xor U12732 (N_12732,N_10498,N_11587);
nor U12733 (N_12733,N_11574,N_12458);
nor U12734 (N_12734,N_11074,N_12251);
xnor U12735 (N_12735,N_11117,N_12351);
nor U12736 (N_12736,N_12421,N_12160);
nand U12737 (N_12737,N_10778,N_12201);
nor U12738 (N_12738,N_11747,N_11521);
xnor U12739 (N_12739,N_10559,N_11294);
nor U12740 (N_12740,N_11228,N_12264);
nand U12741 (N_12741,N_11819,N_11923);
and U12742 (N_12742,N_11100,N_12299);
nor U12743 (N_12743,N_11277,N_10170);
nand U12744 (N_12744,N_10526,N_12382);
xnor U12745 (N_12745,N_11668,N_11674);
and U12746 (N_12746,N_11713,N_10449);
nor U12747 (N_12747,N_11518,N_12489);
nor U12748 (N_12748,N_11468,N_12285);
and U12749 (N_12749,N_11143,N_12314);
or U12750 (N_12750,N_10174,N_12132);
and U12751 (N_12751,N_11888,N_11261);
xnor U12752 (N_12752,N_11363,N_10457);
and U12753 (N_12753,N_10675,N_10098);
nand U12754 (N_12754,N_10609,N_11304);
xor U12755 (N_12755,N_11644,N_10788);
xnor U12756 (N_12756,N_12472,N_10900);
nand U12757 (N_12757,N_11630,N_10395);
nand U12758 (N_12758,N_12225,N_11597);
nand U12759 (N_12759,N_11110,N_11851);
xnor U12760 (N_12760,N_10214,N_11075);
xnor U12761 (N_12761,N_10140,N_12247);
or U12762 (N_12762,N_10616,N_10382);
nand U12763 (N_12763,N_11384,N_11190);
or U12764 (N_12764,N_10122,N_10066);
or U12765 (N_12765,N_10714,N_10545);
or U12766 (N_12766,N_10530,N_11230);
or U12767 (N_12767,N_12217,N_11073);
nand U12768 (N_12768,N_11909,N_12498);
and U12769 (N_12769,N_10614,N_11046);
nor U12770 (N_12770,N_10925,N_10678);
xor U12771 (N_12771,N_12471,N_12437);
nand U12772 (N_12772,N_10723,N_10144);
or U12773 (N_12773,N_10238,N_11650);
nand U12774 (N_12774,N_11308,N_10510);
xnor U12775 (N_12775,N_11448,N_12377);
xnor U12776 (N_12776,N_11300,N_10007);
nor U12777 (N_12777,N_11476,N_10340);
nor U12778 (N_12778,N_10294,N_11042);
xor U12779 (N_12779,N_10652,N_11249);
xor U12780 (N_12780,N_11921,N_10581);
nand U12781 (N_12781,N_11195,N_10810);
nor U12782 (N_12782,N_11489,N_11062);
xnor U12783 (N_12783,N_11779,N_11406);
xor U12784 (N_12784,N_12391,N_11080);
and U12785 (N_12785,N_11244,N_11887);
xnor U12786 (N_12786,N_10524,N_11122);
and U12787 (N_12787,N_10104,N_11013);
and U12788 (N_12788,N_12071,N_10286);
and U12789 (N_12789,N_12109,N_12337);
nand U12790 (N_12790,N_10402,N_12191);
nor U12791 (N_12791,N_11068,N_10749);
and U12792 (N_12792,N_11131,N_12090);
xnor U12793 (N_12793,N_10620,N_11425);
nand U12794 (N_12794,N_11024,N_11688);
xnor U12795 (N_12795,N_10506,N_11200);
nor U12796 (N_12796,N_10279,N_10057);
or U12797 (N_12797,N_10051,N_11994);
nor U12798 (N_12798,N_10427,N_11607);
and U12799 (N_12799,N_10094,N_11314);
nand U12800 (N_12800,N_11372,N_12139);
and U12801 (N_12801,N_10100,N_10590);
or U12802 (N_12802,N_11458,N_10024);
nand U12803 (N_12803,N_10138,N_11439);
and U12804 (N_12804,N_10301,N_10884);
or U12805 (N_12805,N_11052,N_10025);
and U12806 (N_12806,N_12376,N_11262);
or U12807 (N_12807,N_12024,N_11344);
xor U12808 (N_12808,N_12245,N_10401);
nand U12809 (N_12809,N_12099,N_11186);
nand U12810 (N_12810,N_12413,N_11153);
nor U12811 (N_12811,N_10273,N_12055);
nor U12812 (N_12812,N_11381,N_11014);
and U12813 (N_12813,N_10772,N_11453);
and U12814 (N_12814,N_11517,N_10167);
xnor U12815 (N_12815,N_11828,N_10998);
xor U12816 (N_12816,N_10660,N_10515);
nor U12817 (N_12817,N_10359,N_12082);
and U12818 (N_12818,N_10887,N_10783);
and U12819 (N_12819,N_12126,N_10462);
nand U12820 (N_12820,N_12115,N_11225);
nand U12821 (N_12821,N_11178,N_11580);
xnor U12822 (N_12822,N_10330,N_11135);
xor U12823 (N_12823,N_11633,N_11217);
xnor U12824 (N_12824,N_11968,N_12490);
nor U12825 (N_12825,N_12270,N_11154);
xor U12826 (N_12826,N_10448,N_11810);
and U12827 (N_12827,N_12466,N_12401);
xnor U12828 (N_12828,N_10262,N_11065);
and U12829 (N_12829,N_11836,N_11816);
nor U12830 (N_12830,N_11706,N_11938);
nand U12831 (N_12831,N_11955,N_12434);
xnor U12832 (N_12832,N_10488,N_11281);
and U12833 (N_12833,N_10006,N_11632);
or U12834 (N_12834,N_12030,N_11111);
nand U12835 (N_12835,N_11698,N_12093);
or U12836 (N_12836,N_10555,N_11685);
nand U12837 (N_12837,N_10927,N_10054);
nand U12838 (N_12838,N_11682,N_11595);
and U12839 (N_12839,N_11050,N_10867);
nor U12840 (N_12840,N_10873,N_11191);
nand U12841 (N_12841,N_10994,N_11269);
nand U12842 (N_12842,N_10434,N_11162);
or U12843 (N_12843,N_11522,N_10899);
nor U12844 (N_12844,N_10012,N_12312);
nor U12845 (N_12845,N_10663,N_11842);
xor U12846 (N_12846,N_11882,N_10954);
xor U12847 (N_12847,N_11911,N_11331);
xnor U12848 (N_12848,N_10764,N_11513);
nor U12849 (N_12849,N_10860,N_10840);
nand U12850 (N_12850,N_10745,N_10948);
or U12851 (N_12851,N_11862,N_10863);
and U12852 (N_12852,N_11786,N_12315);
and U12853 (N_12853,N_12306,N_10485);
or U12854 (N_12854,N_12187,N_11918);
nand U12855 (N_12855,N_10275,N_12483);
xor U12856 (N_12856,N_10959,N_11266);
or U12857 (N_12857,N_12321,N_11885);
nand U12858 (N_12858,N_12189,N_10833);
nor U12859 (N_12859,N_11038,N_10339);
nand U12860 (N_12860,N_10227,N_10747);
and U12861 (N_12861,N_11018,N_12150);
and U12862 (N_12862,N_10056,N_11469);
nand U12863 (N_12863,N_10437,N_11916);
or U12864 (N_12864,N_10328,N_11960);
or U12865 (N_12865,N_10794,N_10389);
xnor U12866 (N_12866,N_11681,N_12037);
and U12867 (N_12867,N_11928,N_11551);
nor U12868 (N_12868,N_12159,N_10299);
xor U12869 (N_12869,N_10689,N_11944);
and U12870 (N_12870,N_10185,N_10666);
nand U12871 (N_12871,N_12459,N_10509);
nand U12872 (N_12872,N_11168,N_10667);
or U12873 (N_12873,N_11765,N_11808);
nand U12874 (N_12874,N_10676,N_11067);
or U12875 (N_12875,N_10417,N_12014);
nor U12876 (N_12876,N_10608,N_12106);
nand U12877 (N_12877,N_12327,N_10315);
nand U12878 (N_12878,N_12246,N_10968);
and U12879 (N_12879,N_12393,N_10949);
and U12880 (N_12880,N_10826,N_10931);
xnor U12881 (N_12881,N_11546,N_11948);
and U12882 (N_12882,N_10086,N_10977);
nand U12883 (N_12883,N_11723,N_11240);
nor U12884 (N_12884,N_11679,N_10119);
xnor U12885 (N_12885,N_11342,N_11833);
nor U12886 (N_12886,N_12417,N_12145);
nor U12887 (N_12887,N_11202,N_11523);
nand U12888 (N_12888,N_10367,N_12443);
xor U12889 (N_12889,N_10518,N_10635);
or U12890 (N_12890,N_11227,N_11673);
nand U12891 (N_12891,N_11733,N_10612);
nand U12892 (N_12892,N_11565,N_10408);
nor U12893 (N_12893,N_10035,N_10324);
nand U12894 (N_12894,N_10712,N_10211);
or U12895 (N_12895,N_12322,N_10642);
or U12896 (N_12896,N_10685,N_12478);
nand U12897 (N_12897,N_11512,N_10588);
nand U12898 (N_12898,N_12117,N_10398);
nor U12899 (N_12899,N_11766,N_12405);
nor U12900 (N_12900,N_10309,N_12381);
nor U12901 (N_12901,N_11514,N_12023);
nor U12902 (N_12902,N_10662,N_10763);
xor U12903 (N_12903,N_10563,N_11016);
or U12904 (N_12904,N_10149,N_10318);
or U12905 (N_12905,N_11756,N_11598);
or U12906 (N_12906,N_10319,N_11964);
and U12907 (N_12907,N_10997,N_11362);
nand U12908 (N_12908,N_11877,N_11504);
xnor U12909 (N_12909,N_12133,N_11288);
nand U12910 (N_12910,N_12326,N_10752);
xnor U12911 (N_12911,N_10882,N_11940);
or U12912 (N_12912,N_11555,N_10529);
and U12913 (N_12913,N_10071,N_12269);
and U12914 (N_12914,N_10296,N_10158);
nand U12915 (N_12915,N_12176,N_11023);
or U12916 (N_12916,N_11236,N_10569);
or U12917 (N_12917,N_11827,N_12250);
and U12918 (N_12918,N_10869,N_10467);
and U12919 (N_12919,N_10632,N_11383);
and U12920 (N_12920,N_10753,N_12006);
xor U12921 (N_12921,N_12110,N_10823);
xor U12922 (N_12922,N_11567,N_11801);
or U12923 (N_12923,N_11412,N_10907);
and U12924 (N_12924,N_11102,N_12238);
and U12925 (N_12925,N_11606,N_11302);
nand U12926 (N_12926,N_10289,N_10571);
nand U12927 (N_12927,N_10649,N_11222);
nor U12928 (N_12928,N_10168,N_11638);
and U12929 (N_12929,N_12078,N_10597);
and U12930 (N_12930,N_10990,N_10938);
or U12931 (N_12931,N_12281,N_11956);
nor U12932 (N_12932,N_10985,N_10876);
nor U12933 (N_12933,N_12412,N_10637);
nand U12934 (N_12934,N_10472,N_11915);
or U12935 (N_12935,N_11857,N_11081);
nor U12936 (N_12936,N_10356,N_11404);
or U12937 (N_12937,N_12441,N_11159);
or U12938 (N_12938,N_10456,N_12480);
nor U12939 (N_12939,N_12016,N_11811);
and U12940 (N_12940,N_11474,N_10743);
and U12941 (N_12941,N_11519,N_10068);
xor U12942 (N_12942,N_10564,N_10724);
xnor U12943 (N_12943,N_10598,N_11799);
nor U12944 (N_12944,N_10777,N_11749);
or U12945 (N_12945,N_10043,N_12469);
xnor U12946 (N_12946,N_12384,N_11951);
nand U12947 (N_12947,N_11677,N_10983);
nor U12948 (N_12948,N_11303,N_10305);
or U12949 (N_12949,N_11588,N_11239);
or U12950 (N_12950,N_10253,N_11957);
and U12951 (N_12951,N_10349,N_11378);
nor U12952 (N_12952,N_12453,N_10862);
and U12953 (N_12953,N_12212,N_10836);
and U12954 (N_12954,N_10072,N_10871);
xnor U12955 (N_12955,N_12274,N_10226);
nand U12956 (N_12956,N_12325,N_11265);
nor U12957 (N_12957,N_10257,N_10800);
nand U12958 (N_12958,N_10706,N_10926);
and U12959 (N_12959,N_11712,N_11534);
nand U12960 (N_12960,N_11586,N_12476);
and U12961 (N_12961,N_10410,N_10082);
xnor U12962 (N_12962,N_11954,N_10396);
xor U12963 (N_12963,N_11690,N_11500);
nor U12964 (N_12964,N_10814,N_12034);
nor U12965 (N_12965,N_11648,N_11662);
nor U12966 (N_12966,N_11831,N_12293);
xnor U12967 (N_12967,N_11490,N_12266);
and U12968 (N_12968,N_10821,N_12079);
nor U12969 (N_12969,N_10321,N_10418);
nand U12970 (N_12970,N_11338,N_12012);
nand U12971 (N_12971,N_12013,N_12272);
nand U12972 (N_12972,N_10837,N_10827);
and U12973 (N_12973,N_11169,N_11456);
and U12974 (N_12974,N_10604,N_11118);
nand U12975 (N_12975,N_12027,N_12033);
xor U12976 (N_12976,N_11871,N_11703);
xnor U12977 (N_12977,N_10322,N_10774);
xnor U12978 (N_12978,N_11506,N_10105);
or U12979 (N_12979,N_11446,N_11245);
xor U12980 (N_12980,N_11492,N_11041);
nand U12981 (N_12981,N_11405,N_10522);
nor U12982 (N_12982,N_12067,N_11361);
nor U12983 (N_12983,N_11572,N_11339);
nand U12984 (N_12984,N_10508,N_12404);
or U12985 (N_12985,N_11791,N_12204);
nand U12986 (N_12986,N_11892,N_11762);
nor U12987 (N_12987,N_10930,N_11064);
xor U12988 (N_12988,N_11364,N_11130);
nor U12989 (N_12989,N_10481,N_12025);
xor U12990 (N_12990,N_10342,N_10424);
or U12991 (N_12991,N_10233,N_10756);
and U12992 (N_12992,N_10220,N_12049);
and U12993 (N_12993,N_11621,N_11947);
or U12994 (N_12994,N_10258,N_12263);
or U12995 (N_12995,N_11590,N_12010);
nand U12996 (N_12996,N_11634,N_11394);
nand U12997 (N_12997,N_10327,N_11601);
or U12998 (N_12998,N_10630,N_12346);
and U12999 (N_12999,N_11557,N_10092);
xor U13000 (N_13000,N_11287,N_11465);
xnor U13001 (N_13001,N_12248,N_12112);
or U13002 (N_13002,N_12387,N_11473);
nand U13003 (N_13003,N_11760,N_11860);
nor U13004 (N_13004,N_10067,N_10965);
nand U13005 (N_13005,N_10787,N_12101);
nor U13006 (N_13006,N_12029,N_11005);
nand U13007 (N_13007,N_10791,N_11974);
xor U13008 (N_13008,N_10219,N_11839);
and U13009 (N_13009,N_11272,N_11198);
and U13010 (N_13010,N_11925,N_10594);
or U13011 (N_13011,N_10673,N_10102);
nand U13012 (N_13012,N_10539,N_10343);
nor U13013 (N_13013,N_10956,N_10650);
xor U13014 (N_13014,N_10263,N_11187);
nand U13015 (N_13015,N_10125,N_10374);
nand U13016 (N_13016,N_10197,N_10194);
nand U13017 (N_13017,N_12257,N_12156);
or U13018 (N_13018,N_11150,N_11540);
or U13019 (N_13019,N_11501,N_10618);
nor U13020 (N_13020,N_11785,N_11460);
and U13021 (N_13021,N_10773,N_11750);
or U13022 (N_13022,N_12309,N_10807);
or U13023 (N_13023,N_10202,N_11071);
nand U13024 (N_13024,N_11098,N_11470);
or U13025 (N_13025,N_11258,N_12410);
or U13026 (N_13026,N_10041,N_12230);
nor U13027 (N_13027,N_10180,N_10247);
nand U13028 (N_13028,N_10601,N_10824);
or U13029 (N_13029,N_12301,N_10592);
or U13030 (N_13030,N_11864,N_10468);
xnor U13031 (N_13031,N_10274,N_11893);
nor U13032 (N_13032,N_11667,N_10187);
or U13033 (N_13033,N_12203,N_10781);
xnor U13034 (N_13034,N_12211,N_12041);
and U13035 (N_13035,N_12279,N_12436);
nand U13036 (N_13036,N_11532,N_11241);
and U13037 (N_13037,N_10804,N_12493);
nand U13038 (N_13038,N_12454,N_11719);
nor U13039 (N_13039,N_12038,N_12066);
nor U13040 (N_13040,N_11164,N_12073);
nor U13041 (N_13041,N_10973,N_12242);
or U13042 (N_13042,N_11855,N_11511);
or U13043 (N_13043,N_10626,N_12198);
nor U13044 (N_13044,N_12465,N_11790);
or U13045 (N_13045,N_10423,N_11356);
xor U13046 (N_13046,N_10769,N_11352);
xor U13047 (N_13047,N_10979,N_10392);
xnor U13048 (N_13048,N_11988,N_11834);
nor U13049 (N_13049,N_11379,N_12186);
nor U13050 (N_13050,N_11348,N_11172);
nand U13051 (N_13051,N_11704,N_10390);
nand U13052 (N_13052,N_11524,N_12292);
and U13053 (N_13053,N_10252,N_10702);
nor U13054 (N_13054,N_10475,N_11375);
nor U13055 (N_13055,N_10815,N_11966);
xor U13056 (N_13056,N_12429,N_12040);
and U13057 (N_13057,N_11914,N_11962);
nor U13058 (N_13058,N_10135,N_12044);
nor U13059 (N_13059,N_12094,N_10665);
or U13060 (N_13060,N_12365,N_11895);
nor U13061 (N_13061,N_10266,N_11026);
nand U13062 (N_13062,N_11399,N_11946);
or U13063 (N_13063,N_11547,N_10157);
nand U13064 (N_13064,N_11044,N_11051);
and U13065 (N_13065,N_10737,N_11193);
nor U13066 (N_13066,N_11637,N_11004);
or U13067 (N_13067,N_11411,N_10636);
or U13068 (N_13068,N_11285,N_10380);
and U13069 (N_13069,N_12171,N_12324);
nor U13070 (N_13070,N_12182,N_10184);
nor U13071 (N_13071,N_11935,N_11196);
and U13072 (N_13072,N_12298,N_12140);
nand U13073 (N_13073,N_11321,N_10785);
xor U13074 (N_13074,N_11737,N_10169);
or U13075 (N_13075,N_11035,N_11097);
xnor U13076 (N_13076,N_10910,N_11279);
xor U13077 (N_13077,N_10765,N_11120);
xor U13078 (N_13078,N_10044,N_11967);
xnor U13079 (N_13079,N_12181,N_12121);
and U13080 (N_13080,N_12026,N_10120);
xnor U13081 (N_13081,N_12172,N_10021);
or U13082 (N_13082,N_11060,N_10492);
and U13083 (N_13083,N_12092,N_10451);
or U13084 (N_13084,N_12481,N_10543);
and U13085 (N_13085,N_11320,N_10645);
nand U13086 (N_13086,N_10182,N_12149);
and U13087 (N_13087,N_12046,N_11392);
xnor U13088 (N_13088,N_10069,N_12380);
and U13089 (N_13089,N_12152,N_10771);
nor U13090 (N_13090,N_12202,N_11076);
or U13091 (N_13091,N_11684,N_11748);
nor U13092 (N_13092,N_10820,N_10311);
nand U13093 (N_13093,N_12288,N_11027);
nand U13094 (N_13094,N_10915,N_11502);
and U13095 (N_13095,N_11402,N_10801);
xnor U13096 (N_13096,N_12487,N_11145);
or U13097 (N_13097,N_11350,N_12297);
and U13098 (N_13098,N_10363,N_11129);
nand U13099 (N_13099,N_10809,N_11128);
nand U13100 (N_13100,N_12379,N_12032);
or U13101 (N_13101,N_11692,N_10063);
xor U13102 (N_13102,N_11257,N_10354);
and U13103 (N_13103,N_12147,N_11313);
nand U13104 (N_13104,N_11427,N_11069);
or U13105 (N_13105,N_10671,N_12122);
nor U13106 (N_13106,N_10372,N_12456);
nand U13107 (N_13107,N_11082,N_10320);
nand U13108 (N_13108,N_10894,N_10034);
or U13109 (N_13109,N_10428,N_10982);
xor U13110 (N_13110,N_10916,N_11782);
nor U13111 (N_13111,N_10890,N_12399);
or U13112 (N_13112,N_10993,N_11701);
xnor U13113 (N_13113,N_10829,N_11188);
or U13114 (N_13114,N_10798,N_10429);
and U13115 (N_13115,N_12461,N_10782);
xnor U13116 (N_13116,N_10974,N_11772);
and U13117 (N_13117,N_10955,N_11366);
nor U13118 (N_13118,N_10325,N_11256);
nor U13119 (N_13119,N_11757,N_10576);
xnor U13120 (N_13120,N_11920,N_12261);
and U13121 (N_13121,N_11867,N_11904);
nand U13122 (N_13122,N_12057,N_12375);
xnor U13123 (N_13123,N_10348,N_11401);
or U13124 (N_13124,N_10381,N_10674);
nor U13125 (N_13125,N_11937,N_10115);
xor U13126 (N_13126,N_10466,N_11158);
nor U13127 (N_13127,N_12496,N_11900);
xnor U13128 (N_13128,N_11327,N_11505);
and U13129 (N_13129,N_10483,N_12463);
nand U13130 (N_13130,N_11409,N_11301);
and U13131 (N_13131,N_10287,N_12015);
xnor U13132 (N_13132,N_11019,N_11194);
nor U13133 (N_13133,N_10696,N_11848);
nand U13134 (N_13134,N_10797,N_10958);
nand U13135 (N_13135,N_11687,N_11720);
and U13136 (N_13136,N_10203,N_10083);
nor U13137 (N_13137,N_10615,N_10572);
xor U13138 (N_13138,N_11197,N_12276);
xor U13139 (N_13139,N_10175,N_12050);
or U13140 (N_13140,N_12497,N_10204);
xnor U13141 (N_13141,N_11028,N_11292);
or U13142 (N_13142,N_10101,N_11141);
or U13143 (N_13143,N_10761,N_11326);
and U13144 (N_13144,N_11090,N_10770);
nand U13145 (N_13145,N_11455,N_11436);
or U13146 (N_13146,N_11432,N_10889);
and U13147 (N_13147,N_12195,N_11175);
nand U13148 (N_13148,N_12113,N_12495);
nand U13149 (N_13149,N_10834,N_11959);
nor U13150 (N_13150,N_12237,N_11508);
nor U13151 (N_13151,N_10075,N_10235);
nand U13152 (N_13152,N_10293,N_10245);
xnor U13153 (N_13153,N_11189,N_11840);
xnor U13154 (N_13154,N_11218,N_10845);
nor U13155 (N_13155,N_11419,N_12223);
or U13156 (N_13156,N_10981,N_11767);
and U13157 (N_13157,N_11996,N_11347);
nor U13158 (N_13158,N_11397,N_10528);
nand U13159 (N_13159,N_11003,N_12061);
and U13160 (N_13160,N_11653,N_10422);
xnor U13161 (N_13161,N_12452,N_10205);
and U13162 (N_13162,N_12083,N_10828);
or U13163 (N_13163,N_11484,N_11626);
or U13164 (N_13164,N_10643,N_10853);
or U13165 (N_13165,N_11091,N_10672);
xor U13166 (N_13166,N_11124,N_10099);
nand U13167 (N_13167,N_11445,N_10623);
nor U13168 (N_13168,N_11771,N_10393);
and U13169 (N_13169,N_10943,N_10795);
xnor U13170 (N_13170,N_10019,N_10110);
nor U13171 (N_13171,N_12339,N_11570);
and U13172 (N_13172,N_10911,N_11984);
xnor U13173 (N_13173,N_11146,N_11510);
nand U13174 (N_13174,N_11132,N_12116);
nand U13175 (N_13175,N_12043,N_10659);
xnor U13176 (N_13176,N_11612,N_11408);
nand U13177 (N_13177,N_11328,N_10221);
or U13178 (N_13178,N_11527,N_10668);
xnor U13179 (N_13179,N_10496,N_10088);
xnor U13180 (N_13180,N_12333,N_10897);
nor U13181 (N_13181,N_10246,N_10690);
or U13182 (N_13182,N_12477,N_12445);
xor U13183 (N_13183,N_12076,N_11694);
nor U13184 (N_13184,N_10856,N_10038);
and U13185 (N_13185,N_12154,N_12499);
and U13186 (N_13186,N_12068,N_11661);
xor U13187 (N_13187,N_10514,N_11079);
nand U13188 (N_13188,N_10270,N_11553);
nor U13189 (N_13189,N_12304,N_10314);
nor U13190 (N_13190,N_11537,N_12227);
nand U13191 (N_13191,N_10947,N_12123);
xnor U13192 (N_13192,N_10160,N_12252);
or U13193 (N_13193,N_11642,N_11092);
nor U13194 (N_13194,N_11903,N_11910);
xor U13195 (N_13195,N_10684,N_10352);
or U13196 (N_13196,N_11906,N_11853);
nand U13197 (N_13197,N_11815,N_11787);
xnor U13198 (N_13198,N_10939,N_10718);
or U13199 (N_13199,N_11113,N_11400);
nand U13200 (N_13200,N_12350,N_10989);
nor U13201 (N_13201,N_10903,N_12361);
or U13202 (N_13202,N_10420,N_10713);
nor U13203 (N_13203,N_10015,N_11336);
xnor U13204 (N_13204,N_10368,N_10504);
and U13205 (N_13205,N_10888,N_11055);
or U13206 (N_13206,N_11497,N_10586);
xor U13207 (N_13207,N_11999,N_11306);
and U13208 (N_13208,N_11861,N_11594);
nor U13209 (N_13209,N_12450,N_10936);
or U13210 (N_13210,N_12100,N_10790);
xnor U13211 (N_13211,N_12273,N_12419);
or U13212 (N_13212,N_12161,N_10444);
nor U13213 (N_13213,N_10074,N_11376);
nor U13214 (N_13214,N_10688,N_10846);
and U13215 (N_13215,N_11979,N_11096);
and U13216 (N_13216,N_11142,N_12017);
nand U13217 (N_13217,N_10447,N_11725);
xor U13218 (N_13218,N_10150,N_11010);
nand U13219 (N_13219,N_12193,N_10986);
or U13220 (N_13220,N_10587,N_11373);
xnor U13221 (N_13221,N_10707,N_10336);
nor U13222 (N_13222,N_11319,N_10653);
and U13223 (N_13223,N_11732,N_10469);
nor U13224 (N_13224,N_10634,N_10089);
or U13225 (N_13225,N_11869,N_11897);
xnor U13226 (N_13226,N_10857,N_10045);
or U13227 (N_13227,N_11094,N_11413);
xnor U13228 (N_13228,N_10497,N_12383);
nand U13229 (N_13229,N_11972,N_11913);
nand U13230 (N_13230,N_10874,N_10568);
xnor U13231 (N_13231,N_11709,N_10479);
xor U13232 (N_13232,N_10657,N_10369);
xor U13233 (N_13233,N_11973,N_11464);
nand U13234 (N_13234,N_10039,N_11568);
xnor U13235 (N_13235,N_11657,N_10230);
nand U13236 (N_13236,N_11237,N_12228);
xnor U13237 (N_13237,N_11208,N_11316);
nor U13238 (N_13238,N_10292,N_11211);
xor U13239 (N_13239,N_10875,N_11907);
or U13240 (N_13240,N_11971,N_11891);
or U13241 (N_13241,N_11783,N_10131);
nand U13242 (N_13242,N_10346,N_10805);
nor U13243 (N_13243,N_10691,N_11533);
and U13244 (N_13244,N_12430,N_12000);
or U13245 (N_13245,N_10835,N_10819);
and U13246 (N_13246,N_10040,N_10201);
nor U13247 (N_13247,N_10533,N_12433);
and U13248 (N_13248,N_11611,N_11671);
xor U13249 (N_13249,N_11410,N_10579);
nand U13250 (N_13250,N_11289,N_10283);
nand U13251 (N_13251,N_11104,N_10881);
xor U13252 (N_13252,N_12102,N_11173);
and U13253 (N_13253,N_10384,N_10337);
and U13254 (N_13254,N_10682,N_11093);
nor U13255 (N_13255,N_12114,N_11420);
xor U13256 (N_13256,N_10295,N_10222);
xor U13257 (N_13257,N_11866,N_10338);
or U13258 (N_13258,N_12289,N_10987);
nor U13259 (N_13259,N_10854,N_12199);
xor U13260 (N_13260,N_11651,N_11775);
nand U13261 (N_13261,N_11631,N_11958);
nor U13262 (N_13262,N_12035,N_10213);
or U13263 (N_13263,N_10064,N_12143);
nand U13264 (N_13264,N_10995,N_11623);
nand U13265 (N_13265,N_11056,N_12005);
and U13266 (N_13266,N_11491,N_11280);
or U13267 (N_13267,N_11147,N_11002);
xnor U13268 (N_13268,N_10441,N_10619);
nor U13269 (N_13269,N_10961,N_10831);
and U13270 (N_13270,N_10729,N_11604);
or U13271 (N_13271,N_10861,N_12260);
nand U13272 (N_13272,N_10443,N_11323);
and U13273 (N_13273,N_11134,N_10080);
nand U13274 (N_13274,N_11345,N_10371);
and U13275 (N_13275,N_11942,N_12426);
nand U13276 (N_13276,N_10901,N_10976);
or U13277 (N_13277,N_11541,N_11753);
and U13278 (N_13278,N_11479,N_12259);
nand U13279 (N_13279,N_10580,N_12371);
nand U13280 (N_13280,N_10277,N_11133);
and U13281 (N_13281,N_10517,N_10055);
nand U13282 (N_13282,N_10419,N_10026);
or U13283 (N_13283,N_11426,N_10285);
nand U13284 (N_13284,N_11561,N_12208);
nand U13285 (N_13285,N_11416,N_12151);
or U13286 (N_13286,N_12265,N_11812);
nand U13287 (N_13287,N_10030,N_11538);
nand U13288 (N_13288,N_11263,N_10918);
nand U13289 (N_13289,N_11563,N_10172);
nor U13290 (N_13290,N_11123,N_11707);
nand U13291 (N_13291,N_10963,N_12438);
and U13292 (N_13292,N_11933,N_10631);
or U13293 (N_13293,N_12200,N_11264);
nor U13294 (N_13294,N_10606,N_10784);
nor U13295 (N_13295,N_11360,N_12439);
and U13296 (N_13296,N_11794,N_10722);
and U13297 (N_13297,N_10859,N_12047);
or U13298 (N_13298,N_10980,N_11856);
nor U13299 (N_13299,N_10596,N_12234);
and U13300 (N_13300,N_12268,N_11270);
or U13301 (N_13301,N_11544,N_12164);
nor U13302 (N_13302,N_10849,N_11503);
xnor U13303 (N_13303,N_10117,N_11346);
or U13304 (N_13304,N_10754,N_11291);
or U13305 (N_13305,N_10218,N_10291);
and U13306 (N_13306,N_11185,N_11357);
nand U13307 (N_13307,N_10502,N_10345);
nor U13308 (N_13308,N_10452,N_10109);
xnor U13309 (N_13309,N_10459,N_11599);
nand U13310 (N_13310,N_11161,N_10178);
xor U13311 (N_13311,N_10118,N_11192);
and U13312 (N_13312,N_12008,N_12402);
and U13313 (N_13313,N_12310,N_10877);
xnor U13314 (N_13314,N_10241,N_10647);
or U13315 (N_13315,N_11975,N_10507);
and U13316 (N_13316,N_12070,N_11059);
xnor U13317 (N_13317,N_12386,N_10377);
nand U13318 (N_13318,N_12136,N_12407);
nor U13319 (N_13319,N_11620,N_12243);
xnor U13320 (N_13320,N_11125,N_10491);
xor U13321 (N_13321,N_11778,N_12464);
nand U13322 (N_13322,N_11459,N_11462);
nor U13323 (N_13323,N_10513,N_10486);
nor U13324 (N_13324,N_12170,N_10059);
nor U13325 (N_13325,N_11214,N_12474);
and U13326 (N_13326,N_11012,N_10290);
nand U13327 (N_13327,N_11792,N_12468);
and U13328 (N_13328,N_11845,N_11822);
nand U13329 (N_13329,N_10641,N_11250);
nor U13330 (N_13330,N_10654,N_11981);
and U13331 (N_13331,N_10951,N_11229);
nor U13332 (N_13332,N_10822,N_10540);
or U13333 (N_13333,N_10085,N_10992);
nor U13334 (N_13334,N_11058,N_11066);
and U13335 (N_13335,N_12323,N_11243);
and U13336 (N_13336,N_11552,N_11034);
xnor U13337 (N_13337,N_12236,N_10112);
xnor U13338 (N_13338,N_10477,N_11640);
and U13339 (N_13339,N_11708,N_11325);
nor U13340 (N_13340,N_11542,N_12166);
xnor U13341 (N_13341,N_11431,N_10500);
xor U13342 (N_13342,N_11509,N_10531);
nand U13343 (N_13343,N_10193,N_11006);
xor U13344 (N_13344,N_11025,N_12233);
nor U13345 (N_13345,N_10512,N_11109);
nand U13346 (N_13346,N_12129,N_10844);
or U13347 (N_13347,N_11255,N_11151);
and U13348 (N_13348,N_10969,N_10171);
or U13349 (N_13349,N_11166,N_11057);
nand U13350 (N_13350,N_10229,N_11054);
and U13351 (N_13351,N_11539,N_11224);
or U13352 (N_13352,N_10409,N_10173);
and U13353 (N_13353,N_10076,N_10898);
xor U13354 (N_13354,N_11355,N_12137);
and U13355 (N_13355,N_10683,N_11206);
nor U13356 (N_13356,N_10593,N_12300);
or U13357 (N_13357,N_10121,N_10058);
and U13358 (N_13358,N_10825,N_11393);
or U13359 (N_13359,N_12180,N_12357);
and U13360 (N_13360,N_10523,N_11179);
or U13361 (N_13361,N_12188,N_12173);
nor U13362 (N_13362,N_10029,N_10433);
and U13363 (N_13363,N_10658,N_11883);
and U13364 (N_13364,N_11724,N_12394);
nand U13365 (N_13365,N_12165,N_10611);
nor U13366 (N_13366,N_12028,N_12296);
nand U13367 (N_13367,N_11741,N_12213);
or U13368 (N_13368,N_12425,N_10310);
and U13369 (N_13369,N_11924,N_10864);
nand U13370 (N_13370,N_10440,N_12080);
nand U13371 (N_13371,N_10489,N_11837);
xnor U13372 (N_13372,N_11482,N_10206);
nor U13373 (N_13373,N_11645,N_10603);
nor U13374 (N_13374,N_12131,N_11078);
or U13375 (N_13375,N_11926,N_10376);
or U13376 (N_13376,N_11061,N_11781);
nor U13377 (N_13377,N_12138,N_11330);
and U13378 (N_13378,N_10132,N_10031);
nand U13379 (N_13379,N_11009,N_10331);
or U13380 (N_13380,N_11106,N_10482);
or U13381 (N_13381,N_11315,N_10733);
and U13382 (N_13382,N_10087,N_11387);
or U13383 (N_13383,N_12488,N_11203);
xor U13384 (N_13384,N_11485,N_10028);
nor U13385 (N_13385,N_11278,N_10566);
and U13386 (N_13386,N_10463,N_12215);
xor U13387 (N_13387,N_10902,N_11309);
nand U13388 (N_13388,N_10207,N_10432);
nor U13389 (N_13389,N_12018,N_11886);
and U13390 (N_13390,N_11717,N_10548);
nand U13391 (N_13391,N_11843,N_12052);
nor U13392 (N_13392,N_11138,N_11183);
or U13393 (N_13393,N_11583,N_11581);
nand U13394 (N_13394,N_10490,N_10334);
and U13395 (N_13395,N_11126,N_10720);
nor U13396 (N_13396,N_10375,N_10200);
or U13397 (N_13397,N_12075,N_10032);
and U13398 (N_13398,N_12262,N_10776);
or U13399 (N_13399,N_11390,N_12003);
xor U13400 (N_13400,N_12409,N_10053);
nand U13401 (N_13401,N_11659,N_12206);
nand U13402 (N_13402,N_11077,N_11011);
or U13403 (N_13403,N_10143,N_11721);
nor U13404 (N_13404,N_10139,N_12308);
and U13405 (N_13405,N_10848,N_10516);
and U13406 (N_13406,N_12119,N_11872);
or U13407 (N_13407,N_10397,N_10062);
and U13408 (N_13408,N_10971,N_10655);
xor U13409 (N_13409,N_11273,N_11548);
nand U13410 (N_13410,N_10458,N_12194);
nand U13411 (N_13411,N_11901,N_10646);
nor U13412 (N_13412,N_10046,N_10677);
nand U13413 (N_13413,N_12183,N_11424);
and U13414 (N_13414,N_11395,N_10223);
xnor U13415 (N_13415,N_10966,N_11655);
or U13416 (N_13416,N_11989,N_10960);
or U13417 (N_13417,N_11311,N_10697);
xor U13418 (N_13418,N_12098,N_10036);
xnor U13419 (N_13419,N_11305,N_10312);
nor U13420 (N_13420,N_11841,N_11433);
or U13421 (N_13421,N_11969,N_11875);
xor U13422 (N_13422,N_12097,N_12280);
nand U13423 (N_13423,N_10304,N_11184);
nor U13424 (N_13424,N_12009,N_11442);
or U13425 (N_13425,N_12485,N_11160);
or U13426 (N_13426,N_12039,N_12368);
nand U13427 (N_13427,N_10471,N_11032);
and U13428 (N_13428,N_12059,N_12130);
xnor U13429 (N_13429,N_11498,N_11976);
xnor U13430 (N_13430,N_11201,N_11629);
or U13431 (N_13431,N_11450,N_11422);
xnor U13432 (N_13432,N_11095,N_11283);
and U13433 (N_13433,N_12366,N_12178);
nand U13434 (N_13434,N_10700,N_10547);
nand U13435 (N_13435,N_10250,N_10942);
and U13436 (N_13436,N_10560,N_12124);
nor U13437 (N_13437,N_11879,N_10307);
xor U13438 (N_13438,N_10405,N_10360);
xor U13439 (N_13439,N_10519,N_11139);
nor U13440 (N_13440,N_10212,N_11722);
nand U13441 (N_13441,N_10308,N_11136);
nor U13442 (N_13442,N_10351,N_10288);
nand U13443 (N_13443,N_11931,N_11809);
xnor U13444 (N_13444,N_10181,N_12249);
nand U13445 (N_13445,N_10883,N_10276);
nor U13446 (N_13446,N_11209,N_12127);
or U13447 (N_13447,N_10162,N_11652);
nor U13448 (N_13448,N_12072,N_10850);
and U13449 (N_13449,N_12155,N_10177);
nor U13450 (N_13450,N_10128,N_11029);
and U13451 (N_13451,N_12162,N_11494);
and U13452 (N_13452,N_11444,N_11751);
or U13453 (N_13453,N_11324,N_12403);
nand U13454 (N_13454,N_10779,N_12232);
and U13455 (N_13455,N_12011,N_11884);
and U13456 (N_13456,N_10004,N_11535);
nor U13457 (N_13457,N_10578,N_10190);
xnor U13458 (N_13458,N_10751,N_12374);
nand U13459 (N_13459,N_12054,N_11380);
nor U13460 (N_13460,N_12318,N_10487);
or U13461 (N_13461,N_10306,N_10582);
nand U13462 (N_13462,N_11290,N_10740);
and U13463 (N_13463,N_11212,N_10126);
xor U13464 (N_13464,N_10767,N_12214);
xor U13465 (N_13465,N_12065,N_11739);
xor U13466 (N_13466,N_11457,N_12253);
or U13467 (N_13467,N_11602,N_12218);
nor U13468 (N_13468,N_11286,N_10535);
or U13469 (N_13469,N_11403,N_11242);
and U13470 (N_13470,N_10146,N_10249);
or U13471 (N_13471,N_11932,N_11894);
or U13472 (N_13472,N_11368,N_11103);
nand U13473 (N_13473,N_10865,N_10403);
nand U13474 (N_13474,N_11438,N_10165);
nor U13475 (N_13475,N_11849,N_10210);
nand U13476 (N_13476,N_11155,N_10151);
or U13477 (N_13477,N_12334,N_11922);
nor U13478 (N_13478,N_11950,N_10847);
nor U13479 (N_13479,N_12022,N_12311);
or U13480 (N_13480,N_10520,N_11575);
xnor U13481 (N_13481,N_12369,N_11070);
xnor U13482 (N_13482,N_10638,N_11817);
nor U13483 (N_13483,N_11774,N_12144);
and U13484 (N_13484,N_10988,N_11669);
and U13485 (N_13485,N_10727,N_10473);
and U13486 (N_13486,N_10575,N_12063);
xor U13487 (N_13487,N_10744,N_10011);
or U13488 (N_13488,N_11813,N_12036);
or U13489 (N_13489,N_10648,N_10365);
nand U13490 (N_13490,N_10081,N_11689);
and U13491 (N_13491,N_12135,N_12255);
or U13492 (N_13492,N_11149,N_10027);
nor U13493 (N_13493,N_12373,N_10022);
or U13494 (N_13494,N_11554,N_12209);
nand U13495 (N_13495,N_10018,N_10176);
and U13496 (N_13496,N_12449,N_11022);
or U13497 (N_13497,N_10991,N_12354);
and U13498 (N_13498,N_11844,N_10735);
nor U13499 (N_13499,N_10161,N_10549);
xor U13500 (N_13500,N_10681,N_11639);
and U13501 (N_13501,N_11047,N_11702);
and U13502 (N_13502,N_11007,N_11693);
nand U13503 (N_13503,N_10978,N_10999);
nand U13504 (N_13504,N_10812,N_11603);
xnor U13505 (N_13505,N_12336,N_10335);
nand U13506 (N_13506,N_10373,N_11199);
nor U13507 (N_13507,N_10525,N_11176);
and U13508 (N_13508,N_10256,N_12077);
nor U13509 (N_13509,N_10445,N_11758);
xor U13510 (N_13510,N_11939,N_10550);
and U13511 (N_13511,N_10156,N_11789);
and U13512 (N_13512,N_11605,N_10425);
and U13513 (N_13513,N_11234,N_11127);
and U13514 (N_13514,N_11797,N_11997);
nor U13515 (N_13515,N_11429,N_10399);
nor U13516 (N_13516,N_11770,N_10133);
nor U13517 (N_13517,N_11254,N_11735);
xor U13518 (N_13518,N_11226,N_12389);
nand U13519 (N_13519,N_11205,N_11743);
nand U13520 (N_13520,N_11564,N_10661);
and U13521 (N_13521,N_12347,N_10919);
or U13522 (N_13522,N_11805,N_12295);
and U13523 (N_13523,N_12120,N_10558);
nand U13524 (N_13524,N_11284,N_11530);
xor U13525 (N_13525,N_11930,N_12395);
xor U13526 (N_13526,N_12169,N_11716);
or U13527 (N_13527,N_11730,N_11880);
nor U13528 (N_13528,N_11610,N_10347);
xnor U13529 (N_13529,N_10379,N_12341);
nand U13530 (N_13530,N_11823,N_12146);
nand U13531 (N_13531,N_10627,N_11591);
and U13532 (N_13532,N_11821,N_11418);
nand U13533 (N_13533,N_11165,N_11609);
nand U13534 (N_13534,N_10599,N_10802);
nor U13535 (N_13535,N_12342,N_12491);
or U13536 (N_13536,N_10474,N_10917);
nand U13537 (N_13537,N_12360,N_10153);
xor U13538 (N_13538,N_10656,N_10532);
or U13539 (N_13539,N_11550,N_10361);
and U13540 (N_13540,N_10537,N_12271);
nor U13541 (N_13541,N_11329,N_12359);
nand U13542 (N_13542,N_11806,N_11259);
nand U13543 (N_13543,N_10716,N_11310);
xor U13544 (N_13544,N_10127,N_10009);
and U13545 (N_13545,N_11646,N_12069);
xor U13546 (N_13546,N_10114,N_11045);
xnor U13547 (N_13547,N_10695,N_10759);
nand U13548 (N_13548,N_12020,N_11953);
xnor U13549 (N_13549,N_10715,N_10261);
and U13550 (N_13550,N_11322,N_11838);
xnor U13551 (N_13551,N_11043,N_10179);
nand U13552 (N_13552,N_12331,N_11804);
xnor U13553 (N_13553,N_10542,N_11293);
nand U13554 (N_13554,N_12424,N_11119);
nor U13555 (N_13555,N_10353,N_11396);
nand U13556 (N_13556,N_10941,N_10464);
or U13557 (N_13557,N_11048,N_12397);
xor U13558 (N_13558,N_10111,N_12344);
xnor U13559 (N_13559,N_12224,N_11697);
xor U13560 (N_13560,N_11358,N_10378);
and U13561 (N_13561,N_10832,N_12282);
and U13562 (N_13562,N_10155,N_10813);
or U13563 (N_13563,N_10793,N_12286);
nand U13564 (N_13564,N_11961,N_11083);
and U13565 (N_13565,N_10268,N_11221);
nand U13566 (N_13566,N_11945,N_11666);
nor U13567 (N_13567,N_12431,N_11617);
or U13568 (N_13568,N_10501,N_10527);
nor U13569 (N_13569,N_10228,N_12275);
nor U13570 (N_13570,N_11874,N_12338);
nand U13571 (N_13571,N_10154,N_11341);
or U13572 (N_13572,N_12470,N_10639);
and U13573 (N_13573,N_10152,N_10552);
nor U13574 (N_13574,N_10962,N_12418);
nand U13575 (N_13575,N_11349,N_10933);
xor U13576 (N_13576,N_10923,N_10705);
and U13577 (N_13577,N_11718,N_10388);
nand U13578 (N_13578,N_12353,N_11108);
nor U13579 (N_13579,N_11941,N_10414);
or U13580 (N_13580,N_10217,N_10920);
and U13581 (N_13581,N_10426,N_11072);
xor U13582 (N_13582,N_10944,N_11896);
and U13583 (N_13583,N_10438,N_12317);
nand U13584 (N_13584,N_11084,N_10878);
xnor U13585 (N_13585,N_12479,N_10693);
nand U13586 (N_13586,N_10905,N_12258);
or U13587 (N_13587,N_10317,N_11670);
or U13588 (N_13588,N_11754,N_10461);
xnor U13589 (N_13589,N_11824,N_11260);
xnor U13590 (N_13590,N_10095,N_11991);
or U13591 (N_13591,N_12400,N_10843);
or U13592 (N_13592,N_11171,N_10755);
and U13593 (N_13593,N_10431,N_11414);
xor U13594 (N_13594,N_10701,N_11715);
xor U13595 (N_13595,N_12064,N_12158);
or U13596 (N_13596,N_10265,N_10470);
xor U13597 (N_13597,N_11235,N_12345);
nor U13598 (N_13598,N_10300,N_10413);
or U13599 (N_13599,N_11802,N_11115);
and U13600 (N_13600,N_12142,N_10387);
nor U13601 (N_13601,N_11818,N_12473);
xor U13602 (N_13602,N_11275,N_12087);
nor U13603 (N_13603,N_11852,N_12104);
nor U13604 (N_13604,N_10303,N_11317);
nor U13605 (N_13605,N_10952,N_10792);
nand U13606 (N_13606,N_11982,N_11734);
xnor U13607 (N_13607,N_12392,N_12021);
nor U13608 (N_13608,N_12254,N_11312);
or U13609 (N_13609,N_12302,N_10010);
and U13610 (N_13610,N_10922,N_12305);
or U13611 (N_13611,N_10692,N_10237);
and U13612 (N_13612,N_11576,N_11478);
nor U13613 (N_13613,N_11868,N_11899);
nand U13614 (N_13614,N_10023,N_10730);
nand U13615 (N_13615,N_10909,N_10838);
xor U13616 (N_13616,N_11890,N_10891);
or U13617 (N_13617,N_11475,N_10886);
or U13618 (N_13618,N_11085,N_11232);
nor U13619 (N_13619,N_12378,N_10726);
nand U13620 (N_13620,N_12141,N_11549);
and U13621 (N_13621,N_11434,N_11001);
and U13622 (N_13622,N_11367,N_11252);
and U13623 (N_13623,N_11847,N_10803);
nand U13624 (N_13624,N_10073,N_10996);
xnor U13625 (N_13625,N_10239,N_12167);
or U13626 (N_13626,N_10003,N_10945);
nor U13627 (N_13627,N_10698,N_11049);
and U13628 (N_13628,N_10385,N_11101);
and U13629 (N_13629,N_12398,N_11516);
nor U13630 (N_13630,N_10940,N_10573);
nand U13631 (N_13631,N_12492,N_11388);
nor U13632 (N_13632,N_11700,N_11784);
nor U13633 (N_13633,N_10855,N_11087);
or U13634 (N_13634,N_12058,N_11451);
nand U13635 (N_13635,N_11608,N_10567);
nor U13636 (N_13636,N_11795,N_12095);
and U13637 (N_13637,N_12451,N_10605);
nand U13638 (N_13638,N_11461,N_11577);
or U13639 (N_13639,N_10370,N_12042);
or U13640 (N_13640,N_11902,N_10329);
or U13641 (N_13641,N_11763,N_11889);
nor U13642 (N_13642,N_10950,N_11167);
and U13643 (N_13643,N_10215,N_11625);
and U13644 (N_13644,N_10583,N_12460);
nand U13645 (N_13645,N_10892,N_10297);
xnor U13646 (N_13646,N_11998,N_12216);
nor U13647 (N_13647,N_10033,N_11798);
xor U13648 (N_13648,N_12019,N_12004);
xor U13649 (N_13649,N_10670,N_11415);
or U13650 (N_13650,N_12179,N_10589);
nor U13651 (N_13651,N_10610,N_11710);
xor U13652 (N_13652,N_12411,N_10394);
xnor U13653 (N_13653,N_11676,N_10016);
nand U13654 (N_13654,N_11177,N_10972);
nand U13655 (N_13655,N_10453,N_10065);
or U13656 (N_13656,N_12367,N_10760);
or U13657 (N_13657,N_10332,N_10703);
and U13658 (N_13658,N_11039,N_12355);
nand U13659 (N_13659,N_11398,N_10929);
nand U13660 (N_13660,N_11934,N_11180);
xor U13661 (N_13661,N_12388,N_11803);
or U13662 (N_13662,N_12192,N_11246);
or U13663 (N_13663,N_10762,N_12408);
nor U13664 (N_13664,N_10002,N_11525);
xnor U13665 (N_13665,N_10750,N_10858);
or U13666 (N_13666,N_11752,N_11040);
nand U13667 (N_13667,N_12001,N_11238);
and U13668 (N_13668,N_12329,N_10430);
and U13669 (N_13669,N_12074,N_11985);
nor U13670 (N_13670,N_11560,N_11441);
or U13671 (N_13671,N_10932,N_10124);
xor U13672 (N_13672,N_10796,N_11020);
or U13673 (N_13673,N_10613,N_11769);
and U13674 (N_13674,N_10617,N_11170);
or U13675 (N_13675,N_12118,N_12062);
xnor U13676 (N_13676,N_10799,N_11649);
xnor U13677 (N_13677,N_11053,N_10644);
nand U13678 (N_13678,N_10091,N_10651);
and U13679 (N_13679,N_12031,N_10758);
and U13680 (N_13680,N_11148,N_12316);
or U13681 (N_13681,N_12235,N_10554);
nand U13682 (N_13682,N_11832,N_11905);
nor U13683 (N_13683,N_12363,N_11296);
nand U13684 (N_13684,N_12356,N_10254);
and U13685 (N_13685,N_12168,N_10415);
or U13686 (N_13686,N_10142,N_11658);
nand U13687 (N_13687,N_11036,N_10446);
nor U13688 (N_13688,N_11793,N_11000);
xor U13689 (N_13689,N_10209,N_11596);
xnor U13690 (N_13690,N_10116,N_11643);
nor U13691 (N_13691,N_10806,N_11800);
xnor U13692 (N_13692,N_12448,N_10732);
and U13693 (N_13693,N_10323,N_10721);
nand U13694 (N_13694,N_11251,N_12205);
or U13695 (N_13695,N_11493,N_10355);
nand U13696 (N_13696,N_11215,N_10113);
or U13697 (N_13697,N_11174,N_10830);
or U13698 (N_13698,N_10231,N_11343);
nand U13699 (N_13699,N_10494,N_10264);
or U13700 (N_13700,N_11466,N_10436);
or U13701 (N_13701,N_10852,N_11274);
nor U13702 (N_13702,N_11499,N_12390);
nor U13703 (N_13703,N_11814,N_10364);
xor U13704 (N_13704,N_11114,N_11334);
and U13705 (N_13705,N_12406,N_11993);
and U13706 (N_13706,N_10195,N_10711);
and U13707 (N_13707,N_10534,N_11616);
or U13708 (N_13708,N_10717,N_12352);
and U13709 (N_13709,N_12370,N_11627);
or U13710 (N_13710,N_11980,N_12153);
nand U13711 (N_13711,N_10621,N_10208);
or U13712 (N_13712,N_11282,N_11618);
or U13713 (N_13713,N_11559,N_10708);
and U13714 (N_13714,N_11983,N_11528);
xnor U13715 (N_13715,N_10872,N_10442);
and U13716 (N_13716,N_11936,N_12290);
or U13717 (N_13717,N_11531,N_11107);
nor U13718 (N_13718,N_10967,N_10895);
and U13719 (N_13719,N_10404,N_10281);
and U13720 (N_13720,N_11593,N_11729);
and U13721 (N_13721,N_11353,N_10957);
nor U13722 (N_13722,N_11163,N_11995);
nor U13723 (N_13723,N_11407,N_11764);
nand U13724 (N_13724,N_12239,N_11600);
or U13725 (N_13725,N_11515,N_11207);
and U13726 (N_13726,N_11582,N_11440);
nor U13727 (N_13727,N_10503,N_10738);
and U13728 (N_13728,N_10108,N_12349);
nand U13729 (N_13729,N_10242,N_12045);
or U13730 (N_13730,N_10460,N_12484);
or U13731 (N_13731,N_10736,N_12455);
nor U13732 (N_13732,N_10640,N_10984);
and U13733 (N_13733,N_10298,N_11271);
nand U13734 (N_13734,N_10768,N_11435);
nor U13735 (N_13735,N_11977,N_11696);
nor U13736 (N_13736,N_10595,N_10271);
nand U13737 (N_13737,N_11825,N_10912);
and U13738 (N_13738,N_12163,N_10386);
and U13739 (N_13739,N_12108,N_10042);
or U13740 (N_13740,N_10232,N_10521);
or U13741 (N_13741,N_12184,N_12284);
and U13742 (N_13742,N_11664,N_11820);
xnor U13743 (N_13743,N_12240,N_10013);
or U13744 (N_13744,N_11332,N_11584);
and U13745 (N_13745,N_11987,N_11636);
nand U13746 (N_13746,N_10136,N_10664);
nor U13747 (N_13747,N_10725,N_11335);
xnor U13748 (N_13748,N_11622,N_10633);
and U13749 (N_13749,N_10077,N_10244);
xor U13750 (N_13750,N_11363,N_12192);
xor U13751 (N_13751,N_12284,N_12439);
or U13752 (N_13752,N_10383,N_12287);
nand U13753 (N_13753,N_10647,N_11052);
and U13754 (N_13754,N_11219,N_10904);
nor U13755 (N_13755,N_11975,N_10174);
or U13756 (N_13756,N_11341,N_10505);
and U13757 (N_13757,N_10765,N_11042);
and U13758 (N_13758,N_11973,N_10751);
xnor U13759 (N_13759,N_11857,N_11059);
nand U13760 (N_13760,N_11900,N_12194);
or U13761 (N_13761,N_10351,N_11570);
and U13762 (N_13762,N_10813,N_10996);
xnor U13763 (N_13763,N_11361,N_12456);
nor U13764 (N_13764,N_10852,N_10500);
nand U13765 (N_13765,N_10340,N_10154);
xor U13766 (N_13766,N_11169,N_10565);
xnor U13767 (N_13767,N_11381,N_11793);
nand U13768 (N_13768,N_11360,N_10000);
or U13769 (N_13769,N_10960,N_11916);
nand U13770 (N_13770,N_11684,N_10261);
and U13771 (N_13771,N_11059,N_10717);
xor U13772 (N_13772,N_12318,N_11350);
nor U13773 (N_13773,N_11571,N_10083);
nor U13774 (N_13774,N_10600,N_12417);
nor U13775 (N_13775,N_11381,N_10382);
and U13776 (N_13776,N_12241,N_11419);
xnor U13777 (N_13777,N_11616,N_10626);
and U13778 (N_13778,N_10531,N_10362);
and U13779 (N_13779,N_11853,N_10798);
and U13780 (N_13780,N_11091,N_10062);
nand U13781 (N_13781,N_11626,N_10621);
xor U13782 (N_13782,N_12404,N_11194);
or U13783 (N_13783,N_12271,N_11693);
and U13784 (N_13784,N_10210,N_12064);
and U13785 (N_13785,N_10350,N_12204);
or U13786 (N_13786,N_10829,N_10968);
or U13787 (N_13787,N_10276,N_12212);
nand U13788 (N_13788,N_11747,N_10980);
and U13789 (N_13789,N_10336,N_10873);
and U13790 (N_13790,N_12202,N_10006);
xnor U13791 (N_13791,N_11551,N_10233);
nor U13792 (N_13792,N_12174,N_12027);
or U13793 (N_13793,N_12076,N_12342);
or U13794 (N_13794,N_10769,N_11568);
nor U13795 (N_13795,N_10216,N_11209);
or U13796 (N_13796,N_11402,N_12018);
xor U13797 (N_13797,N_10192,N_10955);
and U13798 (N_13798,N_11888,N_12293);
and U13799 (N_13799,N_11119,N_12336);
nand U13800 (N_13800,N_12328,N_12319);
nor U13801 (N_13801,N_10920,N_10471);
and U13802 (N_13802,N_10208,N_10817);
and U13803 (N_13803,N_11014,N_12121);
nand U13804 (N_13804,N_12392,N_12251);
nand U13805 (N_13805,N_12089,N_10944);
or U13806 (N_13806,N_10784,N_10768);
nor U13807 (N_13807,N_10327,N_11174);
nor U13808 (N_13808,N_11985,N_10112);
or U13809 (N_13809,N_12369,N_11410);
and U13810 (N_13810,N_12456,N_10109);
nor U13811 (N_13811,N_11399,N_11992);
nand U13812 (N_13812,N_12329,N_10247);
and U13813 (N_13813,N_11175,N_10046);
xor U13814 (N_13814,N_12278,N_11892);
and U13815 (N_13815,N_10846,N_11585);
nand U13816 (N_13816,N_11582,N_10773);
and U13817 (N_13817,N_12291,N_10928);
nor U13818 (N_13818,N_11819,N_10198);
or U13819 (N_13819,N_12414,N_11139);
and U13820 (N_13820,N_12383,N_10869);
nor U13821 (N_13821,N_11203,N_10885);
and U13822 (N_13822,N_10116,N_12003);
xor U13823 (N_13823,N_10341,N_10139);
or U13824 (N_13824,N_11086,N_11667);
nor U13825 (N_13825,N_10745,N_11887);
xnor U13826 (N_13826,N_10732,N_12488);
and U13827 (N_13827,N_11004,N_11176);
xnor U13828 (N_13828,N_12053,N_10130);
xnor U13829 (N_13829,N_10142,N_11645);
nand U13830 (N_13830,N_12044,N_11453);
nand U13831 (N_13831,N_10667,N_10705);
xor U13832 (N_13832,N_11065,N_11093);
nand U13833 (N_13833,N_10403,N_11419);
nor U13834 (N_13834,N_11479,N_12281);
xnor U13835 (N_13835,N_10604,N_11816);
xor U13836 (N_13836,N_10634,N_12442);
nand U13837 (N_13837,N_10937,N_12042);
and U13838 (N_13838,N_10375,N_10476);
nor U13839 (N_13839,N_11187,N_10193);
and U13840 (N_13840,N_11870,N_12128);
xnor U13841 (N_13841,N_10391,N_12489);
nand U13842 (N_13842,N_11852,N_11024);
nor U13843 (N_13843,N_12205,N_11064);
and U13844 (N_13844,N_10571,N_11899);
or U13845 (N_13845,N_10544,N_12265);
nand U13846 (N_13846,N_11202,N_11925);
xor U13847 (N_13847,N_11212,N_10184);
and U13848 (N_13848,N_10994,N_10728);
nand U13849 (N_13849,N_10522,N_11389);
nand U13850 (N_13850,N_11197,N_11319);
and U13851 (N_13851,N_11378,N_11781);
and U13852 (N_13852,N_11321,N_11922);
and U13853 (N_13853,N_10648,N_12127);
xor U13854 (N_13854,N_11060,N_11842);
nor U13855 (N_13855,N_12458,N_10872);
and U13856 (N_13856,N_12485,N_11168);
nor U13857 (N_13857,N_11330,N_11590);
and U13858 (N_13858,N_10064,N_11134);
or U13859 (N_13859,N_10276,N_10508);
or U13860 (N_13860,N_10950,N_10796);
and U13861 (N_13861,N_10141,N_11679);
or U13862 (N_13862,N_11296,N_11243);
or U13863 (N_13863,N_10217,N_10819);
or U13864 (N_13864,N_11679,N_11991);
nor U13865 (N_13865,N_10213,N_10851);
and U13866 (N_13866,N_12119,N_10023);
or U13867 (N_13867,N_11656,N_11112);
xnor U13868 (N_13868,N_11864,N_10770);
nand U13869 (N_13869,N_11677,N_10606);
xor U13870 (N_13870,N_12291,N_11759);
nand U13871 (N_13871,N_10116,N_10513);
nor U13872 (N_13872,N_11275,N_10060);
nand U13873 (N_13873,N_10901,N_11380);
nor U13874 (N_13874,N_11700,N_10589);
and U13875 (N_13875,N_10103,N_12376);
or U13876 (N_13876,N_10456,N_11059);
nor U13877 (N_13877,N_10681,N_11718);
xor U13878 (N_13878,N_12368,N_12431);
nand U13879 (N_13879,N_12019,N_11914);
xor U13880 (N_13880,N_10977,N_10684);
xnor U13881 (N_13881,N_12259,N_11807);
and U13882 (N_13882,N_10720,N_12142);
xnor U13883 (N_13883,N_12006,N_11671);
and U13884 (N_13884,N_10181,N_11688);
and U13885 (N_13885,N_10159,N_10891);
or U13886 (N_13886,N_11422,N_10338);
nor U13887 (N_13887,N_11752,N_11781);
or U13888 (N_13888,N_11046,N_11510);
or U13889 (N_13889,N_11727,N_11417);
nand U13890 (N_13890,N_11000,N_11449);
or U13891 (N_13891,N_11552,N_10503);
and U13892 (N_13892,N_10210,N_11571);
and U13893 (N_13893,N_10541,N_11893);
xor U13894 (N_13894,N_10987,N_10249);
xor U13895 (N_13895,N_11973,N_11235);
xor U13896 (N_13896,N_12460,N_11715);
nand U13897 (N_13897,N_10402,N_11099);
nor U13898 (N_13898,N_10518,N_11279);
or U13899 (N_13899,N_10257,N_10271);
nand U13900 (N_13900,N_10188,N_10486);
xor U13901 (N_13901,N_11256,N_10354);
and U13902 (N_13902,N_10144,N_12026);
or U13903 (N_13903,N_11243,N_12151);
or U13904 (N_13904,N_10165,N_11797);
and U13905 (N_13905,N_10069,N_10836);
or U13906 (N_13906,N_10582,N_12465);
nand U13907 (N_13907,N_11242,N_10317);
and U13908 (N_13908,N_11759,N_11987);
xnor U13909 (N_13909,N_10220,N_10772);
nand U13910 (N_13910,N_12115,N_10026);
or U13911 (N_13911,N_11502,N_12165);
or U13912 (N_13912,N_11519,N_12353);
or U13913 (N_13913,N_10370,N_12363);
nand U13914 (N_13914,N_12361,N_11572);
and U13915 (N_13915,N_10659,N_11346);
and U13916 (N_13916,N_10923,N_11107);
nand U13917 (N_13917,N_12390,N_10431);
or U13918 (N_13918,N_11315,N_10403);
and U13919 (N_13919,N_10417,N_11716);
or U13920 (N_13920,N_12000,N_10751);
xor U13921 (N_13921,N_11011,N_10631);
nor U13922 (N_13922,N_11306,N_12045);
xor U13923 (N_13923,N_11953,N_12239);
xor U13924 (N_13924,N_12131,N_10004);
or U13925 (N_13925,N_12115,N_12227);
nand U13926 (N_13926,N_10857,N_10213);
nand U13927 (N_13927,N_10692,N_10365);
nor U13928 (N_13928,N_11187,N_10890);
xor U13929 (N_13929,N_10122,N_10503);
xnor U13930 (N_13930,N_11473,N_11819);
xnor U13931 (N_13931,N_11448,N_10384);
nand U13932 (N_13932,N_11890,N_10737);
xnor U13933 (N_13933,N_11054,N_10330);
and U13934 (N_13934,N_12112,N_11062);
and U13935 (N_13935,N_11381,N_10289);
xor U13936 (N_13936,N_10430,N_12271);
and U13937 (N_13937,N_11485,N_10595);
xnor U13938 (N_13938,N_12280,N_11285);
or U13939 (N_13939,N_10825,N_11102);
or U13940 (N_13940,N_10467,N_12175);
nor U13941 (N_13941,N_10850,N_10114);
nand U13942 (N_13942,N_11465,N_11743);
xnor U13943 (N_13943,N_11855,N_11655);
nand U13944 (N_13944,N_11228,N_10756);
and U13945 (N_13945,N_12433,N_10696);
and U13946 (N_13946,N_12127,N_11773);
nor U13947 (N_13947,N_11904,N_11741);
xor U13948 (N_13948,N_10472,N_11487);
nand U13949 (N_13949,N_12325,N_11079);
xor U13950 (N_13950,N_10436,N_10468);
or U13951 (N_13951,N_12363,N_11935);
xor U13952 (N_13952,N_11349,N_11180);
nor U13953 (N_13953,N_11406,N_10914);
xnor U13954 (N_13954,N_12416,N_10362);
nand U13955 (N_13955,N_10947,N_10570);
and U13956 (N_13956,N_11381,N_11519);
or U13957 (N_13957,N_11496,N_11352);
nor U13958 (N_13958,N_11639,N_10341);
nor U13959 (N_13959,N_12204,N_11880);
nor U13960 (N_13960,N_12419,N_10400);
or U13961 (N_13961,N_10913,N_11131);
or U13962 (N_13962,N_11627,N_12084);
and U13963 (N_13963,N_10198,N_10142);
nand U13964 (N_13964,N_11914,N_12242);
nor U13965 (N_13965,N_10772,N_11776);
nand U13966 (N_13966,N_12132,N_10027);
xor U13967 (N_13967,N_11248,N_12183);
nand U13968 (N_13968,N_11722,N_11343);
xnor U13969 (N_13969,N_10881,N_12106);
xor U13970 (N_13970,N_11014,N_10770);
nand U13971 (N_13971,N_12210,N_11699);
and U13972 (N_13972,N_10935,N_11817);
nor U13973 (N_13973,N_10994,N_12063);
and U13974 (N_13974,N_11467,N_10397);
and U13975 (N_13975,N_11027,N_10100);
nand U13976 (N_13976,N_11210,N_10150);
or U13977 (N_13977,N_11570,N_11023);
xor U13978 (N_13978,N_11915,N_10140);
xnor U13979 (N_13979,N_11622,N_11926);
nor U13980 (N_13980,N_11293,N_10784);
nand U13981 (N_13981,N_10664,N_12261);
xor U13982 (N_13982,N_11490,N_10500);
xnor U13983 (N_13983,N_11480,N_10013);
xnor U13984 (N_13984,N_10337,N_11479);
nand U13985 (N_13985,N_10333,N_11058);
or U13986 (N_13986,N_11685,N_11531);
and U13987 (N_13987,N_11101,N_10618);
xnor U13988 (N_13988,N_11945,N_11949);
nand U13989 (N_13989,N_12408,N_11658);
and U13990 (N_13990,N_12079,N_11514);
or U13991 (N_13991,N_10429,N_10056);
or U13992 (N_13992,N_11753,N_11592);
or U13993 (N_13993,N_12158,N_10993);
xor U13994 (N_13994,N_12127,N_12294);
or U13995 (N_13995,N_10764,N_10129);
xor U13996 (N_13996,N_11752,N_11233);
nand U13997 (N_13997,N_10051,N_11265);
nand U13998 (N_13998,N_11290,N_12473);
and U13999 (N_13999,N_11938,N_12246);
xnor U14000 (N_14000,N_10140,N_12219);
nor U14001 (N_14001,N_10731,N_10373);
or U14002 (N_14002,N_12124,N_12333);
xor U14003 (N_14003,N_12496,N_11359);
or U14004 (N_14004,N_11909,N_10256);
or U14005 (N_14005,N_12310,N_10685);
nor U14006 (N_14006,N_10467,N_11993);
or U14007 (N_14007,N_11002,N_12063);
and U14008 (N_14008,N_11747,N_10723);
and U14009 (N_14009,N_11283,N_11074);
xnor U14010 (N_14010,N_12157,N_10410);
xor U14011 (N_14011,N_10072,N_10461);
xnor U14012 (N_14012,N_11003,N_11250);
nand U14013 (N_14013,N_10388,N_11235);
or U14014 (N_14014,N_11064,N_11955);
xnor U14015 (N_14015,N_12191,N_11182);
nor U14016 (N_14016,N_10054,N_10417);
or U14017 (N_14017,N_12204,N_11719);
nor U14018 (N_14018,N_11546,N_10294);
and U14019 (N_14019,N_11775,N_11838);
or U14020 (N_14020,N_12017,N_11315);
and U14021 (N_14021,N_10228,N_12183);
or U14022 (N_14022,N_10139,N_10612);
and U14023 (N_14023,N_11405,N_10174);
xnor U14024 (N_14024,N_11493,N_10653);
or U14025 (N_14025,N_10602,N_11894);
xnor U14026 (N_14026,N_11339,N_11089);
xnor U14027 (N_14027,N_12413,N_10279);
or U14028 (N_14028,N_11572,N_10931);
xor U14029 (N_14029,N_10454,N_11730);
and U14030 (N_14030,N_11799,N_11838);
nand U14031 (N_14031,N_11562,N_10890);
xnor U14032 (N_14032,N_10061,N_11198);
and U14033 (N_14033,N_12379,N_11889);
and U14034 (N_14034,N_11759,N_11829);
nor U14035 (N_14035,N_11582,N_11080);
xnor U14036 (N_14036,N_12460,N_11552);
nor U14037 (N_14037,N_10335,N_11136);
xnor U14038 (N_14038,N_11621,N_12100);
or U14039 (N_14039,N_11527,N_10735);
nor U14040 (N_14040,N_10336,N_11702);
xor U14041 (N_14041,N_12285,N_11278);
and U14042 (N_14042,N_11148,N_10986);
nor U14043 (N_14043,N_10696,N_10846);
or U14044 (N_14044,N_10135,N_11354);
nor U14045 (N_14045,N_10235,N_10597);
nor U14046 (N_14046,N_12112,N_11059);
nor U14047 (N_14047,N_10125,N_11227);
and U14048 (N_14048,N_12123,N_11733);
xnor U14049 (N_14049,N_10602,N_11178);
nor U14050 (N_14050,N_10817,N_10382);
and U14051 (N_14051,N_10539,N_10671);
nor U14052 (N_14052,N_10228,N_10561);
and U14053 (N_14053,N_12036,N_10315);
and U14054 (N_14054,N_10638,N_10957);
xor U14055 (N_14055,N_10964,N_10555);
nor U14056 (N_14056,N_12194,N_10985);
and U14057 (N_14057,N_11681,N_10201);
or U14058 (N_14058,N_11755,N_12406);
and U14059 (N_14059,N_11339,N_10638);
and U14060 (N_14060,N_12271,N_10082);
nor U14061 (N_14061,N_12126,N_10301);
xnor U14062 (N_14062,N_12023,N_10329);
xor U14063 (N_14063,N_10145,N_12277);
nand U14064 (N_14064,N_11247,N_11056);
nor U14065 (N_14065,N_12299,N_11618);
or U14066 (N_14066,N_11244,N_10381);
xnor U14067 (N_14067,N_12013,N_10144);
and U14068 (N_14068,N_10759,N_11979);
or U14069 (N_14069,N_11886,N_11428);
and U14070 (N_14070,N_10473,N_10472);
and U14071 (N_14071,N_11350,N_10153);
or U14072 (N_14072,N_10810,N_10760);
and U14073 (N_14073,N_11736,N_10356);
and U14074 (N_14074,N_11607,N_12234);
nor U14075 (N_14075,N_12055,N_11410);
xor U14076 (N_14076,N_11307,N_11522);
nor U14077 (N_14077,N_12288,N_10498);
nand U14078 (N_14078,N_12128,N_10989);
xnor U14079 (N_14079,N_11218,N_10761);
and U14080 (N_14080,N_11910,N_10884);
and U14081 (N_14081,N_10353,N_11329);
nor U14082 (N_14082,N_11148,N_11552);
and U14083 (N_14083,N_12163,N_11792);
or U14084 (N_14084,N_11586,N_11715);
or U14085 (N_14085,N_11626,N_10994);
and U14086 (N_14086,N_10453,N_10625);
or U14087 (N_14087,N_10621,N_10366);
xor U14088 (N_14088,N_10226,N_10635);
nor U14089 (N_14089,N_11531,N_11548);
nor U14090 (N_14090,N_10072,N_11678);
nor U14091 (N_14091,N_11555,N_10119);
and U14092 (N_14092,N_10707,N_12281);
xnor U14093 (N_14093,N_12368,N_10137);
or U14094 (N_14094,N_12104,N_11069);
nand U14095 (N_14095,N_11049,N_11404);
and U14096 (N_14096,N_10393,N_12396);
and U14097 (N_14097,N_10577,N_10508);
and U14098 (N_14098,N_10757,N_11401);
or U14099 (N_14099,N_11538,N_10702);
and U14100 (N_14100,N_12361,N_10237);
nand U14101 (N_14101,N_11526,N_11490);
or U14102 (N_14102,N_11079,N_11200);
nor U14103 (N_14103,N_10039,N_11078);
and U14104 (N_14104,N_11371,N_12289);
nor U14105 (N_14105,N_11872,N_10801);
xnor U14106 (N_14106,N_11403,N_10732);
and U14107 (N_14107,N_12335,N_11583);
nand U14108 (N_14108,N_11059,N_10856);
or U14109 (N_14109,N_11891,N_12096);
xor U14110 (N_14110,N_11383,N_10068);
and U14111 (N_14111,N_11934,N_11053);
nor U14112 (N_14112,N_10656,N_11616);
and U14113 (N_14113,N_10215,N_11940);
nand U14114 (N_14114,N_12476,N_10106);
and U14115 (N_14115,N_10663,N_11908);
xnor U14116 (N_14116,N_11163,N_11058);
or U14117 (N_14117,N_12202,N_11208);
or U14118 (N_14118,N_12341,N_10931);
nand U14119 (N_14119,N_11497,N_10827);
nand U14120 (N_14120,N_11796,N_10153);
or U14121 (N_14121,N_11201,N_11809);
nor U14122 (N_14122,N_11794,N_11909);
xnor U14123 (N_14123,N_10084,N_10244);
nand U14124 (N_14124,N_10630,N_10309);
nand U14125 (N_14125,N_10332,N_10009);
or U14126 (N_14126,N_12015,N_11007);
nand U14127 (N_14127,N_10473,N_10927);
or U14128 (N_14128,N_10325,N_12223);
nand U14129 (N_14129,N_10076,N_11628);
nand U14130 (N_14130,N_11641,N_11698);
nor U14131 (N_14131,N_10847,N_12458);
and U14132 (N_14132,N_10568,N_10945);
and U14133 (N_14133,N_12099,N_11296);
and U14134 (N_14134,N_11839,N_11412);
and U14135 (N_14135,N_11433,N_10422);
nor U14136 (N_14136,N_11118,N_11017);
nor U14137 (N_14137,N_10041,N_10543);
nor U14138 (N_14138,N_11486,N_10878);
and U14139 (N_14139,N_10757,N_12292);
nor U14140 (N_14140,N_10733,N_10755);
xor U14141 (N_14141,N_11677,N_12263);
nand U14142 (N_14142,N_11314,N_10012);
and U14143 (N_14143,N_10147,N_10493);
nor U14144 (N_14144,N_10613,N_11081);
and U14145 (N_14145,N_11106,N_11574);
or U14146 (N_14146,N_12421,N_11995);
and U14147 (N_14147,N_11375,N_10636);
xor U14148 (N_14148,N_10435,N_11154);
or U14149 (N_14149,N_10854,N_11960);
and U14150 (N_14150,N_10475,N_11356);
or U14151 (N_14151,N_10460,N_11143);
nor U14152 (N_14152,N_12116,N_10157);
xor U14153 (N_14153,N_11763,N_11528);
nor U14154 (N_14154,N_11939,N_11166);
nand U14155 (N_14155,N_11799,N_12290);
xor U14156 (N_14156,N_11262,N_10532);
nor U14157 (N_14157,N_11941,N_11933);
nor U14158 (N_14158,N_10298,N_10167);
nand U14159 (N_14159,N_12269,N_11901);
xor U14160 (N_14160,N_10172,N_10513);
nor U14161 (N_14161,N_10608,N_11303);
nor U14162 (N_14162,N_12302,N_10374);
nand U14163 (N_14163,N_10820,N_11676);
or U14164 (N_14164,N_10048,N_12316);
or U14165 (N_14165,N_12294,N_11923);
or U14166 (N_14166,N_11946,N_11890);
or U14167 (N_14167,N_10600,N_11548);
xnor U14168 (N_14168,N_12167,N_10080);
xor U14169 (N_14169,N_11043,N_10426);
xor U14170 (N_14170,N_11655,N_10983);
xor U14171 (N_14171,N_10693,N_11529);
nor U14172 (N_14172,N_11747,N_11300);
nand U14173 (N_14173,N_10642,N_10379);
nand U14174 (N_14174,N_11366,N_11782);
xnor U14175 (N_14175,N_12186,N_11433);
and U14176 (N_14176,N_11119,N_11314);
and U14177 (N_14177,N_10779,N_10587);
and U14178 (N_14178,N_12067,N_12085);
xnor U14179 (N_14179,N_10049,N_12490);
nand U14180 (N_14180,N_10724,N_10362);
and U14181 (N_14181,N_10252,N_11090);
or U14182 (N_14182,N_10532,N_12361);
nand U14183 (N_14183,N_11389,N_11807);
nor U14184 (N_14184,N_11641,N_11640);
and U14185 (N_14185,N_10100,N_10495);
nor U14186 (N_14186,N_12488,N_10695);
or U14187 (N_14187,N_10093,N_12383);
or U14188 (N_14188,N_10861,N_11001);
and U14189 (N_14189,N_10468,N_11023);
nor U14190 (N_14190,N_10395,N_12484);
or U14191 (N_14191,N_11454,N_12295);
xor U14192 (N_14192,N_11852,N_10497);
nand U14193 (N_14193,N_11772,N_11513);
xor U14194 (N_14194,N_10708,N_11675);
nand U14195 (N_14195,N_11276,N_10064);
nand U14196 (N_14196,N_12088,N_11631);
nand U14197 (N_14197,N_10309,N_12340);
nor U14198 (N_14198,N_11148,N_12031);
or U14199 (N_14199,N_11224,N_10455);
nor U14200 (N_14200,N_11385,N_12321);
nand U14201 (N_14201,N_11849,N_10446);
xnor U14202 (N_14202,N_10640,N_11225);
nand U14203 (N_14203,N_11112,N_11093);
or U14204 (N_14204,N_12335,N_10470);
nand U14205 (N_14205,N_10476,N_12065);
or U14206 (N_14206,N_10924,N_10682);
nand U14207 (N_14207,N_10974,N_10128);
or U14208 (N_14208,N_12267,N_11755);
xnor U14209 (N_14209,N_11661,N_11049);
and U14210 (N_14210,N_10739,N_12340);
nand U14211 (N_14211,N_11774,N_10296);
nand U14212 (N_14212,N_11761,N_11490);
xnor U14213 (N_14213,N_10790,N_12455);
or U14214 (N_14214,N_10044,N_11560);
nor U14215 (N_14215,N_12175,N_11292);
nor U14216 (N_14216,N_12298,N_10940);
nand U14217 (N_14217,N_12479,N_11238);
or U14218 (N_14218,N_10629,N_11332);
or U14219 (N_14219,N_10077,N_10234);
or U14220 (N_14220,N_11256,N_12035);
and U14221 (N_14221,N_11755,N_10960);
nand U14222 (N_14222,N_11796,N_11134);
nor U14223 (N_14223,N_10429,N_11296);
nor U14224 (N_14224,N_10076,N_11293);
nor U14225 (N_14225,N_10752,N_12259);
or U14226 (N_14226,N_10510,N_10015);
and U14227 (N_14227,N_11200,N_11301);
nand U14228 (N_14228,N_10565,N_11856);
nand U14229 (N_14229,N_11648,N_12166);
nand U14230 (N_14230,N_11582,N_12443);
xnor U14231 (N_14231,N_12407,N_11495);
nand U14232 (N_14232,N_12360,N_10855);
xor U14233 (N_14233,N_12167,N_10044);
nor U14234 (N_14234,N_12289,N_10711);
xnor U14235 (N_14235,N_10368,N_11068);
xnor U14236 (N_14236,N_11416,N_10036);
and U14237 (N_14237,N_10218,N_12224);
and U14238 (N_14238,N_10725,N_10431);
or U14239 (N_14239,N_10420,N_10030);
or U14240 (N_14240,N_11597,N_11795);
nand U14241 (N_14241,N_11365,N_10976);
or U14242 (N_14242,N_11258,N_10614);
or U14243 (N_14243,N_11082,N_10477);
xnor U14244 (N_14244,N_11514,N_12174);
nor U14245 (N_14245,N_10719,N_12228);
nor U14246 (N_14246,N_11250,N_12294);
nor U14247 (N_14247,N_11987,N_11533);
and U14248 (N_14248,N_11193,N_11751);
nor U14249 (N_14249,N_12486,N_10472);
nand U14250 (N_14250,N_10212,N_11691);
xor U14251 (N_14251,N_11154,N_10770);
nand U14252 (N_14252,N_10539,N_10058);
or U14253 (N_14253,N_10241,N_10586);
xor U14254 (N_14254,N_12109,N_11547);
nand U14255 (N_14255,N_11094,N_11241);
nand U14256 (N_14256,N_11511,N_10596);
nand U14257 (N_14257,N_11715,N_10464);
xnor U14258 (N_14258,N_11290,N_11116);
nor U14259 (N_14259,N_12171,N_12087);
or U14260 (N_14260,N_10463,N_11114);
nor U14261 (N_14261,N_10694,N_11093);
xor U14262 (N_14262,N_12221,N_10764);
and U14263 (N_14263,N_11397,N_11969);
or U14264 (N_14264,N_10283,N_10638);
nor U14265 (N_14265,N_12320,N_10404);
or U14266 (N_14266,N_10268,N_11809);
and U14267 (N_14267,N_10894,N_10650);
and U14268 (N_14268,N_10826,N_11675);
nand U14269 (N_14269,N_10844,N_11154);
nand U14270 (N_14270,N_12400,N_10871);
nor U14271 (N_14271,N_10116,N_10257);
and U14272 (N_14272,N_11431,N_11973);
and U14273 (N_14273,N_11103,N_10219);
nor U14274 (N_14274,N_10427,N_11272);
or U14275 (N_14275,N_11973,N_12045);
nand U14276 (N_14276,N_11270,N_10313);
xnor U14277 (N_14277,N_12124,N_11722);
nor U14278 (N_14278,N_10550,N_10884);
and U14279 (N_14279,N_10014,N_10618);
and U14280 (N_14280,N_11022,N_11286);
nor U14281 (N_14281,N_12494,N_11147);
or U14282 (N_14282,N_11851,N_11723);
and U14283 (N_14283,N_11753,N_10466);
and U14284 (N_14284,N_10932,N_11730);
nor U14285 (N_14285,N_10854,N_10267);
nand U14286 (N_14286,N_12185,N_10529);
xnor U14287 (N_14287,N_10931,N_11876);
nor U14288 (N_14288,N_12113,N_12206);
nand U14289 (N_14289,N_11573,N_12098);
nand U14290 (N_14290,N_10927,N_11672);
xnor U14291 (N_14291,N_11953,N_12150);
nand U14292 (N_14292,N_10127,N_11719);
xor U14293 (N_14293,N_10120,N_10205);
and U14294 (N_14294,N_10224,N_10787);
and U14295 (N_14295,N_12113,N_11071);
nand U14296 (N_14296,N_12285,N_12455);
nor U14297 (N_14297,N_10413,N_10582);
nor U14298 (N_14298,N_10080,N_10186);
or U14299 (N_14299,N_10057,N_11664);
and U14300 (N_14300,N_10479,N_12265);
xnor U14301 (N_14301,N_12413,N_12431);
or U14302 (N_14302,N_11466,N_11288);
nand U14303 (N_14303,N_10473,N_10748);
nand U14304 (N_14304,N_11075,N_10719);
xor U14305 (N_14305,N_10121,N_12235);
nor U14306 (N_14306,N_12084,N_12189);
nand U14307 (N_14307,N_12174,N_11649);
xor U14308 (N_14308,N_11115,N_12067);
or U14309 (N_14309,N_12107,N_11856);
and U14310 (N_14310,N_10842,N_11790);
and U14311 (N_14311,N_12396,N_10646);
xnor U14312 (N_14312,N_12401,N_12450);
nor U14313 (N_14313,N_10091,N_11404);
xnor U14314 (N_14314,N_12046,N_10058);
nand U14315 (N_14315,N_11964,N_12037);
or U14316 (N_14316,N_12141,N_12284);
nand U14317 (N_14317,N_10388,N_12011);
nor U14318 (N_14318,N_12184,N_10220);
or U14319 (N_14319,N_12401,N_10900);
or U14320 (N_14320,N_11770,N_10911);
nor U14321 (N_14321,N_10553,N_12383);
nor U14322 (N_14322,N_10551,N_10073);
nand U14323 (N_14323,N_10277,N_11905);
nand U14324 (N_14324,N_10674,N_11815);
xnor U14325 (N_14325,N_12032,N_10431);
or U14326 (N_14326,N_12017,N_11657);
nand U14327 (N_14327,N_11107,N_10742);
xor U14328 (N_14328,N_11666,N_10285);
or U14329 (N_14329,N_10013,N_10180);
nand U14330 (N_14330,N_10188,N_11277);
and U14331 (N_14331,N_11517,N_11095);
or U14332 (N_14332,N_10250,N_11348);
nor U14333 (N_14333,N_10193,N_12270);
or U14334 (N_14334,N_10136,N_11250);
xnor U14335 (N_14335,N_12197,N_10674);
and U14336 (N_14336,N_10358,N_11725);
or U14337 (N_14337,N_11108,N_10978);
nand U14338 (N_14338,N_10431,N_11691);
and U14339 (N_14339,N_10291,N_11655);
nand U14340 (N_14340,N_10349,N_11215);
nor U14341 (N_14341,N_10649,N_12192);
or U14342 (N_14342,N_12225,N_11216);
or U14343 (N_14343,N_10490,N_10815);
and U14344 (N_14344,N_12440,N_10619);
nor U14345 (N_14345,N_10757,N_10548);
nand U14346 (N_14346,N_10480,N_11877);
xnor U14347 (N_14347,N_11723,N_11399);
nor U14348 (N_14348,N_11688,N_11525);
xor U14349 (N_14349,N_10367,N_11059);
nand U14350 (N_14350,N_10858,N_12382);
or U14351 (N_14351,N_11485,N_11009);
nand U14352 (N_14352,N_12223,N_11832);
nor U14353 (N_14353,N_10361,N_10733);
xnor U14354 (N_14354,N_10485,N_10745);
nand U14355 (N_14355,N_11636,N_10310);
or U14356 (N_14356,N_12275,N_11077);
xnor U14357 (N_14357,N_10895,N_11637);
nor U14358 (N_14358,N_11621,N_12286);
nand U14359 (N_14359,N_11237,N_10288);
or U14360 (N_14360,N_12119,N_11588);
xnor U14361 (N_14361,N_11699,N_12112);
nand U14362 (N_14362,N_11978,N_11951);
or U14363 (N_14363,N_12139,N_10245);
xnor U14364 (N_14364,N_11363,N_11153);
nand U14365 (N_14365,N_11501,N_10993);
xnor U14366 (N_14366,N_10072,N_12089);
or U14367 (N_14367,N_11455,N_11921);
xor U14368 (N_14368,N_12366,N_11316);
and U14369 (N_14369,N_12321,N_10873);
xnor U14370 (N_14370,N_11816,N_10937);
nor U14371 (N_14371,N_12346,N_11290);
and U14372 (N_14372,N_10939,N_11121);
or U14373 (N_14373,N_10867,N_11692);
or U14374 (N_14374,N_10694,N_10546);
nor U14375 (N_14375,N_10830,N_12181);
nand U14376 (N_14376,N_11411,N_12056);
or U14377 (N_14377,N_12199,N_11779);
xnor U14378 (N_14378,N_12488,N_10687);
or U14379 (N_14379,N_10191,N_11504);
nor U14380 (N_14380,N_11521,N_10149);
xor U14381 (N_14381,N_10897,N_10914);
nand U14382 (N_14382,N_10221,N_10900);
nand U14383 (N_14383,N_11631,N_10437);
nand U14384 (N_14384,N_11186,N_11746);
or U14385 (N_14385,N_11509,N_11783);
and U14386 (N_14386,N_12095,N_11713);
and U14387 (N_14387,N_10715,N_10390);
nand U14388 (N_14388,N_11881,N_11836);
nor U14389 (N_14389,N_12092,N_10120);
nand U14390 (N_14390,N_11574,N_10416);
and U14391 (N_14391,N_11153,N_12327);
xor U14392 (N_14392,N_11436,N_11110);
nand U14393 (N_14393,N_12394,N_10799);
xor U14394 (N_14394,N_11305,N_11380);
and U14395 (N_14395,N_12396,N_11105);
nor U14396 (N_14396,N_12339,N_10878);
and U14397 (N_14397,N_11206,N_10227);
nor U14398 (N_14398,N_12450,N_11185);
xnor U14399 (N_14399,N_11318,N_11683);
or U14400 (N_14400,N_10744,N_11913);
or U14401 (N_14401,N_10443,N_10165);
and U14402 (N_14402,N_11718,N_10019);
nor U14403 (N_14403,N_10419,N_10610);
and U14404 (N_14404,N_10569,N_11569);
or U14405 (N_14405,N_12365,N_10554);
or U14406 (N_14406,N_10379,N_10988);
nor U14407 (N_14407,N_11168,N_10444);
xor U14408 (N_14408,N_11781,N_10369);
nand U14409 (N_14409,N_10019,N_11171);
xor U14410 (N_14410,N_10858,N_11286);
nand U14411 (N_14411,N_10302,N_11688);
nor U14412 (N_14412,N_12100,N_10859);
and U14413 (N_14413,N_10008,N_11749);
nand U14414 (N_14414,N_10812,N_11562);
or U14415 (N_14415,N_11671,N_11559);
nand U14416 (N_14416,N_10620,N_12242);
or U14417 (N_14417,N_12308,N_10901);
xor U14418 (N_14418,N_11902,N_10245);
and U14419 (N_14419,N_11042,N_12135);
xnor U14420 (N_14420,N_11805,N_12326);
and U14421 (N_14421,N_12240,N_11054);
nand U14422 (N_14422,N_11329,N_11880);
xnor U14423 (N_14423,N_10955,N_11929);
and U14424 (N_14424,N_11662,N_11749);
nor U14425 (N_14425,N_10963,N_11092);
and U14426 (N_14426,N_11905,N_12474);
or U14427 (N_14427,N_10488,N_10027);
or U14428 (N_14428,N_11303,N_11399);
and U14429 (N_14429,N_12173,N_10436);
nor U14430 (N_14430,N_11073,N_11266);
or U14431 (N_14431,N_12231,N_10058);
or U14432 (N_14432,N_10176,N_12449);
nor U14433 (N_14433,N_10776,N_12176);
nand U14434 (N_14434,N_10099,N_12047);
nand U14435 (N_14435,N_12277,N_10813);
nor U14436 (N_14436,N_11019,N_11912);
and U14437 (N_14437,N_12165,N_10746);
nor U14438 (N_14438,N_12479,N_11155);
nor U14439 (N_14439,N_10440,N_12157);
and U14440 (N_14440,N_12405,N_11313);
nand U14441 (N_14441,N_12365,N_12247);
nor U14442 (N_14442,N_10555,N_12385);
nand U14443 (N_14443,N_11772,N_11844);
xor U14444 (N_14444,N_11935,N_11529);
nor U14445 (N_14445,N_10676,N_11143);
nand U14446 (N_14446,N_10258,N_10807);
xor U14447 (N_14447,N_10238,N_11969);
and U14448 (N_14448,N_11062,N_10259);
nor U14449 (N_14449,N_11391,N_12282);
and U14450 (N_14450,N_11752,N_11134);
and U14451 (N_14451,N_10024,N_11603);
xnor U14452 (N_14452,N_10576,N_11736);
nand U14453 (N_14453,N_10921,N_11076);
nand U14454 (N_14454,N_12392,N_12029);
nand U14455 (N_14455,N_12323,N_10452);
nor U14456 (N_14456,N_11562,N_10767);
nor U14457 (N_14457,N_11033,N_12409);
nand U14458 (N_14458,N_11445,N_11572);
nand U14459 (N_14459,N_11811,N_12004);
xnor U14460 (N_14460,N_12446,N_12486);
or U14461 (N_14461,N_11442,N_12102);
nand U14462 (N_14462,N_11578,N_12293);
or U14463 (N_14463,N_12368,N_12497);
nand U14464 (N_14464,N_12392,N_12254);
and U14465 (N_14465,N_11243,N_11367);
and U14466 (N_14466,N_11588,N_11705);
nor U14467 (N_14467,N_10168,N_11566);
nand U14468 (N_14468,N_11687,N_10331);
and U14469 (N_14469,N_11316,N_10063);
nand U14470 (N_14470,N_11922,N_12497);
or U14471 (N_14471,N_11459,N_10477);
and U14472 (N_14472,N_10344,N_11153);
nor U14473 (N_14473,N_11967,N_10962);
nor U14474 (N_14474,N_11276,N_11934);
and U14475 (N_14475,N_10578,N_10081);
nand U14476 (N_14476,N_10392,N_11333);
and U14477 (N_14477,N_11031,N_11755);
or U14478 (N_14478,N_12229,N_10138);
or U14479 (N_14479,N_12200,N_11816);
or U14480 (N_14480,N_11634,N_10653);
xor U14481 (N_14481,N_11145,N_10312);
nor U14482 (N_14482,N_10907,N_11483);
and U14483 (N_14483,N_12104,N_10553);
or U14484 (N_14484,N_12059,N_12263);
nor U14485 (N_14485,N_11451,N_12281);
and U14486 (N_14486,N_11490,N_11165);
nand U14487 (N_14487,N_10131,N_10240);
or U14488 (N_14488,N_12479,N_11961);
nand U14489 (N_14489,N_12361,N_10637);
and U14490 (N_14490,N_10408,N_10474);
nand U14491 (N_14491,N_10966,N_11177);
and U14492 (N_14492,N_10373,N_10603);
nor U14493 (N_14493,N_12405,N_11264);
nand U14494 (N_14494,N_12285,N_11347);
and U14495 (N_14495,N_10333,N_10220);
or U14496 (N_14496,N_10723,N_10955);
nand U14497 (N_14497,N_11499,N_12263);
and U14498 (N_14498,N_12362,N_11468);
xnor U14499 (N_14499,N_10654,N_10631);
xor U14500 (N_14500,N_10336,N_10924);
and U14501 (N_14501,N_10104,N_12234);
and U14502 (N_14502,N_11274,N_10144);
xnor U14503 (N_14503,N_10507,N_12470);
and U14504 (N_14504,N_10406,N_11815);
or U14505 (N_14505,N_11777,N_11699);
nor U14506 (N_14506,N_12013,N_11356);
nor U14507 (N_14507,N_10922,N_11234);
nand U14508 (N_14508,N_10728,N_12482);
nor U14509 (N_14509,N_10135,N_11423);
nor U14510 (N_14510,N_11844,N_10754);
and U14511 (N_14511,N_10914,N_12363);
nor U14512 (N_14512,N_11615,N_11725);
or U14513 (N_14513,N_10433,N_10270);
nand U14514 (N_14514,N_12113,N_12466);
xnor U14515 (N_14515,N_11942,N_11482);
nand U14516 (N_14516,N_10156,N_11824);
or U14517 (N_14517,N_11095,N_10190);
and U14518 (N_14518,N_10632,N_11919);
xnor U14519 (N_14519,N_11996,N_11881);
and U14520 (N_14520,N_10751,N_11219);
or U14521 (N_14521,N_11261,N_11712);
or U14522 (N_14522,N_11512,N_10482);
or U14523 (N_14523,N_11753,N_10438);
and U14524 (N_14524,N_12220,N_11196);
or U14525 (N_14525,N_11288,N_10639);
nor U14526 (N_14526,N_12254,N_11281);
nand U14527 (N_14527,N_12427,N_11938);
xnor U14528 (N_14528,N_10775,N_12101);
nor U14529 (N_14529,N_12374,N_12172);
and U14530 (N_14530,N_11907,N_12251);
or U14531 (N_14531,N_11321,N_11996);
or U14532 (N_14532,N_10721,N_10943);
nor U14533 (N_14533,N_10281,N_11555);
and U14534 (N_14534,N_11574,N_11873);
nand U14535 (N_14535,N_11408,N_11410);
and U14536 (N_14536,N_11143,N_11874);
xnor U14537 (N_14537,N_12308,N_11026);
nor U14538 (N_14538,N_11750,N_10729);
or U14539 (N_14539,N_10894,N_10295);
xnor U14540 (N_14540,N_10038,N_11795);
nor U14541 (N_14541,N_10594,N_11259);
or U14542 (N_14542,N_11198,N_11638);
nand U14543 (N_14543,N_11951,N_12095);
nand U14544 (N_14544,N_10570,N_10745);
or U14545 (N_14545,N_10395,N_10608);
nand U14546 (N_14546,N_10443,N_11021);
nand U14547 (N_14547,N_11400,N_10773);
xnor U14548 (N_14548,N_12403,N_11565);
xnor U14549 (N_14549,N_12406,N_11824);
nand U14550 (N_14550,N_12025,N_12207);
and U14551 (N_14551,N_11326,N_11167);
nor U14552 (N_14552,N_10761,N_11211);
xnor U14553 (N_14553,N_11971,N_12254);
or U14554 (N_14554,N_11825,N_10881);
and U14555 (N_14555,N_11102,N_11825);
nand U14556 (N_14556,N_12364,N_10615);
or U14557 (N_14557,N_12127,N_11087);
xnor U14558 (N_14558,N_11407,N_10260);
nand U14559 (N_14559,N_12145,N_10841);
nor U14560 (N_14560,N_11024,N_10194);
xor U14561 (N_14561,N_11865,N_10565);
and U14562 (N_14562,N_11867,N_11272);
nand U14563 (N_14563,N_11753,N_10205);
nor U14564 (N_14564,N_12450,N_11760);
nor U14565 (N_14565,N_11643,N_10989);
xor U14566 (N_14566,N_12164,N_10078);
nand U14567 (N_14567,N_11763,N_12287);
nor U14568 (N_14568,N_10621,N_11703);
and U14569 (N_14569,N_11131,N_10402);
or U14570 (N_14570,N_10656,N_10778);
nor U14571 (N_14571,N_12472,N_10069);
nand U14572 (N_14572,N_11083,N_10036);
nor U14573 (N_14573,N_10961,N_11192);
xnor U14574 (N_14574,N_11650,N_10473);
nor U14575 (N_14575,N_12196,N_12165);
nor U14576 (N_14576,N_11396,N_11664);
or U14577 (N_14577,N_12094,N_12243);
nand U14578 (N_14578,N_11995,N_10289);
or U14579 (N_14579,N_11437,N_12005);
xor U14580 (N_14580,N_10691,N_11003);
or U14581 (N_14581,N_12157,N_12399);
nand U14582 (N_14582,N_11962,N_11588);
nand U14583 (N_14583,N_12257,N_11803);
and U14584 (N_14584,N_11187,N_10483);
xor U14585 (N_14585,N_11417,N_10283);
or U14586 (N_14586,N_10121,N_10622);
nor U14587 (N_14587,N_10186,N_11133);
xor U14588 (N_14588,N_12098,N_12399);
and U14589 (N_14589,N_12281,N_12156);
or U14590 (N_14590,N_10369,N_10700);
or U14591 (N_14591,N_12446,N_10333);
xor U14592 (N_14592,N_11291,N_12104);
and U14593 (N_14593,N_10311,N_10184);
nand U14594 (N_14594,N_10135,N_11920);
xnor U14595 (N_14595,N_10839,N_11345);
nor U14596 (N_14596,N_11442,N_10156);
and U14597 (N_14597,N_11143,N_11095);
nor U14598 (N_14598,N_10421,N_11919);
nor U14599 (N_14599,N_11323,N_10174);
nand U14600 (N_14600,N_10826,N_10441);
and U14601 (N_14601,N_12011,N_11705);
nor U14602 (N_14602,N_10249,N_11737);
xor U14603 (N_14603,N_12277,N_10207);
nand U14604 (N_14604,N_12047,N_11913);
nand U14605 (N_14605,N_10622,N_11207);
or U14606 (N_14606,N_10130,N_10429);
and U14607 (N_14607,N_10713,N_10158);
and U14608 (N_14608,N_12119,N_11212);
or U14609 (N_14609,N_10482,N_11290);
nand U14610 (N_14610,N_12387,N_11406);
nor U14611 (N_14611,N_11878,N_10768);
nor U14612 (N_14612,N_10014,N_12211);
nor U14613 (N_14613,N_10845,N_11997);
or U14614 (N_14614,N_11280,N_12217);
and U14615 (N_14615,N_10690,N_11358);
nor U14616 (N_14616,N_11411,N_10894);
and U14617 (N_14617,N_11690,N_11470);
or U14618 (N_14618,N_12381,N_10396);
and U14619 (N_14619,N_10780,N_10963);
xnor U14620 (N_14620,N_11784,N_10581);
and U14621 (N_14621,N_11695,N_11497);
and U14622 (N_14622,N_12263,N_11310);
nor U14623 (N_14623,N_10357,N_12188);
and U14624 (N_14624,N_12308,N_11915);
and U14625 (N_14625,N_11381,N_11707);
xor U14626 (N_14626,N_11735,N_12221);
xor U14627 (N_14627,N_11269,N_12162);
xnor U14628 (N_14628,N_11016,N_12289);
and U14629 (N_14629,N_12238,N_11823);
xnor U14630 (N_14630,N_12108,N_12223);
nand U14631 (N_14631,N_11610,N_11579);
or U14632 (N_14632,N_10706,N_11084);
or U14633 (N_14633,N_12415,N_12305);
and U14634 (N_14634,N_10369,N_11824);
or U14635 (N_14635,N_11983,N_12123);
or U14636 (N_14636,N_10683,N_10550);
nand U14637 (N_14637,N_10307,N_12355);
nor U14638 (N_14638,N_12301,N_10147);
nand U14639 (N_14639,N_11194,N_10919);
nand U14640 (N_14640,N_10462,N_11864);
xor U14641 (N_14641,N_12419,N_12142);
xor U14642 (N_14642,N_11232,N_12209);
or U14643 (N_14643,N_10727,N_10607);
nand U14644 (N_14644,N_10719,N_11752);
and U14645 (N_14645,N_12328,N_12423);
xnor U14646 (N_14646,N_10268,N_11470);
xor U14647 (N_14647,N_10814,N_12285);
xor U14648 (N_14648,N_11991,N_12064);
or U14649 (N_14649,N_12035,N_11842);
nand U14650 (N_14650,N_10738,N_10977);
and U14651 (N_14651,N_10418,N_11120);
xor U14652 (N_14652,N_11241,N_12043);
xor U14653 (N_14653,N_12043,N_10509);
or U14654 (N_14654,N_11710,N_12412);
xnor U14655 (N_14655,N_10974,N_11470);
or U14656 (N_14656,N_12471,N_11032);
nor U14657 (N_14657,N_11494,N_11591);
nand U14658 (N_14658,N_12081,N_10555);
xnor U14659 (N_14659,N_12126,N_12466);
nor U14660 (N_14660,N_10681,N_10283);
xor U14661 (N_14661,N_10590,N_10485);
nand U14662 (N_14662,N_10089,N_10607);
nand U14663 (N_14663,N_11865,N_10143);
nor U14664 (N_14664,N_10665,N_10447);
and U14665 (N_14665,N_10216,N_10236);
or U14666 (N_14666,N_11678,N_11858);
or U14667 (N_14667,N_10192,N_11950);
and U14668 (N_14668,N_12094,N_11101);
and U14669 (N_14669,N_12331,N_12403);
nor U14670 (N_14670,N_11505,N_11045);
and U14671 (N_14671,N_12186,N_11695);
xor U14672 (N_14672,N_11060,N_10524);
and U14673 (N_14673,N_10967,N_10697);
or U14674 (N_14674,N_10597,N_11378);
nand U14675 (N_14675,N_10818,N_11974);
and U14676 (N_14676,N_10750,N_11248);
nor U14677 (N_14677,N_11166,N_11053);
nor U14678 (N_14678,N_12399,N_11891);
or U14679 (N_14679,N_11259,N_12216);
nor U14680 (N_14680,N_11937,N_12184);
xnor U14681 (N_14681,N_11598,N_10364);
nor U14682 (N_14682,N_10304,N_11125);
nor U14683 (N_14683,N_10554,N_10912);
xnor U14684 (N_14684,N_10951,N_12028);
xnor U14685 (N_14685,N_11177,N_10786);
xor U14686 (N_14686,N_12040,N_11570);
or U14687 (N_14687,N_10299,N_10989);
xor U14688 (N_14688,N_10036,N_10944);
nor U14689 (N_14689,N_11377,N_10640);
and U14690 (N_14690,N_12019,N_11350);
and U14691 (N_14691,N_11767,N_10679);
xnor U14692 (N_14692,N_11373,N_11677);
and U14693 (N_14693,N_10024,N_12229);
and U14694 (N_14694,N_11416,N_11154);
nor U14695 (N_14695,N_12246,N_11369);
nand U14696 (N_14696,N_12482,N_11481);
or U14697 (N_14697,N_12276,N_11240);
nor U14698 (N_14698,N_10698,N_12464);
or U14699 (N_14699,N_10389,N_11753);
nor U14700 (N_14700,N_11436,N_12441);
nand U14701 (N_14701,N_10307,N_11643);
nor U14702 (N_14702,N_12455,N_12292);
nand U14703 (N_14703,N_12401,N_10210);
or U14704 (N_14704,N_10472,N_12473);
xor U14705 (N_14705,N_12462,N_11874);
or U14706 (N_14706,N_12163,N_11888);
nand U14707 (N_14707,N_11011,N_12379);
nand U14708 (N_14708,N_10744,N_10142);
or U14709 (N_14709,N_10100,N_10202);
nor U14710 (N_14710,N_11155,N_11596);
nand U14711 (N_14711,N_10003,N_11651);
or U14712 (N_14712,N_11333,N_11846);
nor U14713 (N_14713,N_10244,N_10387);
xor U14714 (N_14714,N_11862,N_12184);
xor U14715 (N_14715,N_10425,N_10296);
or U14716 (N_14716,N_10329,N_11519);
xor U14717 (N_14717,N_11180,N_10789);
or U14718 (N_14718,N_11412,N_12059);
nand U14719 (N_14719,N_11855,N_12273);
nand U14720 (N_14720,N_10601,N_11875);
or U14721 (N_14721,N_10138,N_11229);
and U14722 (N_14722,N_10716,N_11673);
nand U14723 (N_14723,N_12322,N_11026);
nand U14724 (N_14724,N_11812,N_11457);
and U14725 (N_14725,N_12438,N_10216);
nand U14726 (N_14726,N_10076,N_10149);
xor U14727 (N_14727,N_11247,N_10209);
and U14728 (N_14728,N_11453,N_11030);
and U14729 (N_14729,N_11779,N_10244);
xor U14730 (N_14730,N_11227,N_10826);
nand U14731 (N_14731,N_10508,N_11545);
nand U14732 (N_14732,N_12409,N_11564);
or U14733 (N_14733,N_11930,N_10265);
or U14734 (N_14734,N_10561,N_12100);
nor U14735 (N_14735,N_10862,N_12055);
xor U14736 (N_14736,N_11140,N_10917);
nor U14737 (N_14737,N_10671,N_12235);
or U14738 (N_14738,N_12051,N_10580);
xnor U14739 (N_14739,N_11567,N_11251);
xor U14740 (N_14740,N_12451,N_10272);
nor U14741 (N_14741,N_12410,N_11774);
and U14742 (N_14742,N_12277,N_11571);
nor U14743 (N_14743,N_11530,N_10514);
xnor U14744 (N_14744,N_11135,N_10100);
and U14745 (N_14745,N_11986,N_11479);
xor U14746 (N_14746,N_11423,N_10476);
nor U14747 (N_14747,N_11380,N_11716);
nor U14748 (N_14748,N_12309,N_12414);
and U14749 (N_14749,N_12479,N_11936);
and U14750 (N_14750,N_11339,N_11229);
xnor U14751 (N_14751,N_11428,N_10082);
and U14752 (N_14752,N_12108,N_12499);
or U14753 (N_14753,N_12298,N_11158);
nand U14754 (N_14754,N_11470,N_11686);
xnor U14755 (N_14755,N_11780,N_10364);
xor U14756 (N_14756,N_11734,N_10702);
xor U14757 (N_14757,N_10410,N_12077);
and U14758 (N_14758,N_10388,N_10115);
nor U14759 (N_14759,N_10875,N_10578);
or U14760 (N_14760,N_11400,N_10025);
and U14761 (N_14761,N_10453,N_11536);
or U14762 (N_14762,N_10655,N_10337);
nand U14763 (N_14763,N_11939,N_12496);
nand U14764 (N_14764,N_11932,N_10704);
xnor U14765 (N_14765,N_10180,N_10364);
or U14766 (N_14766,N_11825,N_11488);
xor U14767 (N_14767,N_12398,N_10662);
or U14768 (N_14768,N_10411,N_11461);
xor U14769 (N_14769,N_10140,N_10428);
and U14770 (N_14770,N_12066,N_12048);
nor U14771 (N_14771,N_10180,N_11630);
or U14772 (N_14772,N_11845,N_12125);
and U14773 (N_14773,N_10763,N_10169);
or U14774 (N_14774,N_11185,N_10519);
xor U14775 (N_14775,N_10434,N_12057);
or U14776 (N_14776,N_10117,N_11975);
nor U14777 (N_14777,N_12492,N_11423);
nor U14778 (N_14778,N_12405,N_11940);
xor U14779 (N_14779,N_11065,N_11491);
nand U14780 (N_14780,N_10158,N_12205);
and U14781 (N_14781,N_11292,N_12220);
or U14782 (N_14782,N_10110,N_11231);
or U14783 (N_14783,N_11831,N_10737);
or U14784 (N_14784,N_12396,N_10337);
or U14785 (N_14785,N_10552,N_10975);
and U14786 (N_14786,N_10656,N_12445);
nand U14787 (N_14787,N_12199,N_11466);
xor U14788 (N_14788,N_12384,N_12337);
xnor U14789 (N_14789,N_12187,N_11529);
xor U14790 (N_14790,N_10409,N_11029);
and U14791 (N_14791,N_10495,N_12483);
nand U14792 (N_14792,N_10808,N_10511);
nor U14793 (N_14793,N_11402,N_10348);
and U14794 (N_14794,N_10202,N_10183);
or U14795 (N_14795,N_11228,N_10827);
and U14796 (N_14796,N_11747,N_11772);
and U14797 (N_14797,N_10884,N_11906);
or U14798 (N_14798,N_10188,N_10972);
or U14799 (N_14799,N_11926,N_11959);
and U14800 (N_14800,N_12192,N_10555);
xor U14801 (N_14801,N_12206,N_10558);
xnor U14802 (N_14802,N_10190,N_10265);
nor U14803 (N_14803,N_10609,N_11876);
and U14804 (N_14804,N_11436,N_10536);
and U14805 (N_14805,N_10398,N_10236);
nor U14806 (N_14806,N_11360,N_10909);
or U14807 (N_14807,N_10848,N_12043);
and U14808 (N_14808,N_11222,N_12098);
or U14809 (N_14809,N_10753,N_10188);
or U14810 (N_14810,N_12112,N_11747);
nand U14811 (N_14811,N_12030,N_10320);
xor U14812 (N_14812,N_10233,N_10662);
or U14813 (N_14813,N_12279,N_10597);
or U14814 (N_14814,N_10107,N_11604);
nor U14815 (N_14815,N_10901,N_11853);
nor U14816 (N_14816,N_10515,N_10716);
or U14817 (N_14817,N_11188,N_12198);
xor U14818 (N_14818,N_10851,N_10698);
xor U14819 (N_14819,N_10100,N_10016);
xor U14820 (N_14820,N_11145,N_11614);
and U14821 (N_14821,N_11691,N_11533);
and U14822 (N_14822,N_10943,N_11143);
and U14823 (N_14823,N_11086,N_10203);
or U14824 (N_14824,N_11055,N_11077);
nand U14825 (N_14825,N_11923,N_10237);
nand U14826 (N_14826,N_11082,N_10406);
and U14827 (N_14827,N_10078,N_11258);
and U14828 (N_14828,N_12480,N_11304);
or U14829 (N_14829,N_11169,N_11715);
or U14830 (N_14830,N_11267,N_10796);
and U14831 (N_14831,N_11514,N_10571);
nand U14832 (N_14832,N_10746,N_12439);
nor U14833 (N_14833,N_11529,N_10351);
or U14834 (N_14834,N_10272,N_10770);
and U14835 (N_14835,N_11883,N_10773);
nor U14836 (N_14836,N_11177,N_10948);
nand U14837 (N_14837,N_10751,N_11557);
or U14838 (N_14838,N_10604,N_11776);
or U14839 (N_14839,N_11155,N_11743);
nor U14840 (N_14840,N_10980,N_11365);
nor U14841 (N_14841,N_11194,N_11347);
or U14842 (N_14842,N_11198,N_10753);
nor U14843 (N_14843,N_11861,N_11630);
xnor U14844 (N_14844,N_11646,N_12317);
or U14845 (N_14845,N_11532,N_10258);
xnor U14846 (N_14846,N_11473,N_12116);
or U14847 (N_14847,N_12218,N_10410);
nand U14848 (N_14848,N_12110,N_11531);
nand U14849 (N_14849,N_11200,N_10709);
or U14850 (N_14850,N_11722,N_10352);
xnor U14851 (N_14851,N_12115,N_10477);
nand U14852 (N_14852,N_10081,N_10402);
xor U14853 (N_14853,N_11673,N_11607);
nand U14854 (N_14854,N_10651,N_11918);
nor U14855 (N_14855,N_11703,N_11432);
or U14856 (N_14856,N_10948,N_12017);
nand U14857 (N_14857,N_10909,N_11167);
and U14858 (N_14858,N_11935,N_11849);
xnor U14859 (N_14859,N_11157,N_12348);
nand U14860 (N_14860,N_10701,N_11814);
nand U14861 (N_14861,N_11715,N_12085);
and U14862 (N_14862,N_11679,N_11835);
xnor U14863 (N_14863,N_12467,N_11068);
nor U14864 (N_14864,N_10809,N_11390);
and U14865 (N_14865,N_11153,N_10590);
and U14866 (N_14866,N_11277,N_10102);
or U14867 (N_14867,N_10410,N_11120);
or U14868 (N_14868,N_10089,N_11805);
xnor U14869 (N_14869,N_10081,N_10555);
nor U14870 (N_14870,N_11314,N_10253);
and U14871 (N_14871,N_12235,N_11410);
or U14872 (N_14872,N_10578,N_10639);
or U14873 (N_14873,N_11112,N_10531);
nand U14874 (N_14874,N_10307,N_11864);
or U14875 (N_14875,N_10385,N_11649);
and U14876 (N_14876,N_10325,N_11711);
nand U14877 (N_14877,N_11167,N_10178);
nand U14878 (N_14878,N_12271,N_12366);
nand U14879 (N_14879,N_10429,N_12135);
nor U14880 (N_14880,N_10679,N_10781);
and U14881 (N_14881,N_11368,N_10977);
nand U14882 (N_14882,N_11516,N_11991);
or U14883 (N_14883,N_10435,N_10458);
nand U14884 (N_14884,N_10823,N_10070);
nor U14885 (N_14885,N_10212,N_11241);
nor U14886 (N_14886,N_10532,N_10945);
or U14887 (N_14887,N_11690,N_10337);
xnor U14888 (N_14888,N_11163,N_10954);
xnor U14889 (N_14889,N_10215,N_10758);
or U14890 (N_14890,N_10124,N_11371);
nor U14891 (N_14891,N_12155,N_11419);
or U14892 (N_14892,N_11544,N_10931);
nor U14893 (N_14893,N_10719,N_11947);
and U14894 (N_14894,N_10388,N_12356);
xor U14895 (N_14895,N_10825,N_10094);
nand U14896 (N_14896,N_11349,N_11426);
xnor U14897 (N_14897,N_10560,N_11869);
and U14898 (N_14898,N_11779,N_10276);
nor U14899 (N_14899,N_12416,N_10718);
and U14900 (N_14900,N_12328,N_10234);
nand U14901 (N_14901,N_10878,N_10251);
or U14902 (N_14902,N_10595,N_11261);
or U14903 (N_14903,N_12196,N_10532);
nand U14904 (N_14904,N_12059,N_10185);
xor U14905 (N_14905,N_10424,N_11958);
nand U14906 (N_14906,N_11715,N_10555);
and U14907 (N_14907,N_11845,N_11875);
or U14908 (N_14908,N_11715,N_12372);
xnor U14909 (N_14909,N_11812,N_12069);
or U14910 (N_14910,N_11474,N_11167);
or U14911 (N_14911,N_10305,N_10879);
xor U14912 (N_14912,N_10198,N_12365);
or U14913 (N_14913,N_10398,N_10067);
or U14914 (N_14914,N_11347,N_11153);
nor U14915 (N_14915,N_12259,N_11344);
or U14916 (N_14916,N_11978,N_11552);
or U14917 (N_14917,N_10871,N_10120);
and U14918 (N_14918,N_10566,N_10662);
xnor U14919 (N_14919,N_12308,N_11365);
or U14920 (N_14920,N_10054,N_12149);
nand U14921 (N_14921,N_10674,N_12021);
nand U14922 (N_14922,N_10930,N_11080);
nand U14923 (N_14923,N_11981,N_11510);
and U14924 (N_14924,N_10829,N_11476);
nor U14925 (N_14925,N_10649,N_10973);
and U14926 (N_14926,N_10318,N_10359);
and U14927 (N_14927,N_10193,N_10120);
nand U14928 (N_14928,N_11243,N_11128);
xor U14929 (N_14929,N_10265,N_10244);
and U14930 (N_14930,N_11789,N_11140);
nand U14931 (N_14931,N_11522,N_11083);
or U14932 (N_14932,N_11234,N_12195);
or U14933 (N_14933,N_11503,N_12091);
nor U14934 (N_14934,N_12278,N_10015);
or U14935 (N_14935,N_11010,N_12489);
or U14936 (N_14936,N_12420,N_11038);
or U14937 (N_14937,N_10666,N_10283);
nor U14938 (N_14938,N_12356,N_12489);
xnor U14939 (N_14939,N_12409,N_11038);
xor U14940 (N_14940,N_11239,N_10371);
xor U14941 (N_14941,N_11839,N_12295);
nor U14942 (N_14942,N_11463,N_12350);
and U14943 (N_14943,N_11326,N_11804);
and U14944 (N_14944,N_11134,N_11196);
or U14945 (N_14945,N_10609,N_12085);
nand U14946 (N_14946,N_12155,N_11351);
nand U14947 (N_14947,N_11822,N_12078);
nand U14948 (N_14948,N_12160,N_11091);
nand U14949 (N_14949,N_11554,N_11957);
or U14950 (N_14950,N_12318,N_11479);
nand U14951 (N_14951,N_10289,N_10232);
or U14952 (N_14952,N_10650,N_12185);
or U14953 (N_14953,N_11065,N_11229);
and U14954 (N_14954,N_10584,N_11363);
nor U14955 (N_14955,N_10146,N_11430);
nand U14956 (N_14956,N_12060,N_11455);
nor U14957 (N_14957,N_10977,N_10372);
nand U14958 (N_14958,N_11760,N_12392);
or U14959 (N_14959,N_10145,N_10590);
nand U14960 (N_14960,N_11425,N_11750);
xnor U14961 (N_14961,N_10206,N_11591);
or U14962 (N_14962,N_11529,N_10183);
xnor U14963 (N_14963,N_10668,N_11218);
xor U14964 (N_14964,N_11835,N_11564);
and U14965 (N_14965,N_11825,N_10624);
xnor U14966 (N_14966,N_11156,N_12323);
xor U14967 (N_14967,N_12226,N_10772);
xnor U14968 (N_14968,N_10040,N_11968);
xnor U14969 (N_14969,N_10689,N_10680);
or U14970 (N_14970,N_10106,N_12179);
xnor U14971 (N_14971,N_10091,N_12265);
or U14972 (N_14972,N_10528,N_12022);
nor U14973 (N_14973,N_11157,N_10218);
xnor U14974 (N_14974,N_10216,N_10791);
or U14975 (N_14975,N_10006,N_11452);
and U14976 (N_14976,N_10623,N_12136);
nand U14977 (N_14977,N_10399,N_12382);
nand U14978 (N_14978,N_10237,N_10716);
xor U14979 (N_14979,N_11218,N_10677);
nand U14980 (N_14980,N_12398,N_11263);
and U14981 (N_14981,N_11523,N_10298);
or U14982 (N_14982,N_10920,N_10925);
nor U14983 (N_14983,N_12381,N_11810);
xor U14984 (N_14984,N_10438,N_11507);
or U14985 (N_14985,N_11936,N_10555);
or U14986 (N_14986,N_10104,N_11347);
and U14987 (N_14987,N_11669,N_12112);
nor U14988 (N_14988,N_11742,N_10633);
xor U14989 (N_14989,N_11702,N_12040);
xnor U14990 (N_14990,N_12365,N_12024);
nor U14991 (N_14991,N_11769,N_11351);
and U14992 (N_14992,N_10792,N_11820);
nor U14993 (N_14993,N_10763,N_12141);
nand U14994 (N_14994,N_12269,N_10063);
or U14995 (N_14995,N_10328,N_10487);
nand U14996 (N_14996,N_11696,N_10331);
or U14997 (N_14997,N_12233,N_11501);
xor U14998 (N_14998,N_12393,N_11331);
and U14999 (N_14999,N_11068,N_10905);
nand U15000 (N_15000,N_14267,N_12531);
nor U15001 (N_15001,N_12610,N_13068);
or U15002 (N_15002,N_13573,N_13272);
nand U15003 (N_15003,N_12590,N_14503);
nand U15004 (N_15004,N_14942,N_13689);
nor U15005 (N_15005,N_14715,N_13442);
nor U15006 (N_15006,N_14001,N_14656);
xor U15007 (N_15007,N_14180,N_14821);
and U15008 (N_15008,N_13301,N_14875);
and U15009 (N_15009,N_12803,N_12672);
and U15010 (N_15010,N_12928,N_13993);
or U15011 (N_15011,N_13174,N_14599);
or U15012 (N_15012,N_13487,N_13679);
xor U15013 (N_15013,N_13878,N_13186);
xnor U15014 (N_15014,N_14673,N_13447);
and U15015 (N_15015,N_13118,N_13499);
nor U15016 (N_15016,N_14049,N_13371);
nor U15017 (N_15017,N_14570,N_14008);
and U15018 (N_15018,N_12796,N_14865);
or U15019 (N_15019,N_13514,N_14392);
xor U15020 (N_15020,N_12683,N_12638);
nand U15021 (N_15021,N_13526,N_13386);
nand U15022 (N_15022,N_12527,N_13937);
and U15023 (N_15023,N_13469,N_12876);
nor U15024 (N_15024,N_14544,N_12771);
xnor U15025 (N_15025,N_14457,N_12757);
and U15026 (N_15026,N_14595,N_14591);
nor U15027 (N_15027,N_12680,N_13010);
or U15028 (N_15028,N_14533,N_14375);
nor U15029 (N_15029,N_12572,N_14402);
nand U15030 (N_15030,N_14859,N_13042);
nor U15031 (N_15031,N_13777,N_13388);
or U15032 (N_15032,N_13567,N_13095);
and U15033 (N_15033,N_13012,N_12563);
xnor U15034 (N_15034,N_14224,N_13971);
nand U15035 (N_15035,N_14824,N_14210);
xor U15036 (N_15036,N_13646,N_13458);
xnor U15037 (N_15037,N_14346,N_12510);
and U15038 (N_15038,N_13998,N_14858);
or U15039 (N_15039,N_14361,N_14214);
nor U15040 (N_15040,N_13819,N_13846);
and U15041 (N_15041,N_14442,N_12724);
nor U15042 (N_15042,N_14809,N_12877);
and U15043 (N_15043,N_14028,N_14076);
and U15044 (N_15044,N_13451,N_12750);
nor U15045 (N_15045,N_13252,N_14275);
nand U15046 (N_15046,N_13733,N_13184);
or U15047 (N_15047,N_14571,N_14886);
nand U15048 (N_15048,N_13420,N_13064);
xnor U15049 (N_15049,N_14371,N_14054);
xor U15050 (N_15050,N_12935,N_13385);
nand U15051 (N_15051,N_14469,N_12565);
nor U15052 (N_15052,N_13531,N_12788);
or U15053 (N_15053,N_13670,N_14631);
nor U15054 (N_15054,N_13961,N_13464);
nor U15055 (N_15055,N_13204,N_13340);
and U15056 (N_15056,N_13255,N_14430);
xnor U15057 (N_15057,N_14157,N_14789);
and U15058 (N_15058,N_13857,N_13744);
or U15059 (N_15059,N_14385,N_12653);
and U15060 (N_15060,N_13545,N_14063);
and U15061 (N_15061,N_12785,N_13604);
nand U15062 (N_15062,N_12577,N_13112);
nor U15063 (N_15063,N_13591,N_14056);
or U15064 (N_15064,N_12846,N_13434);
xnor U15065 (N_15065,N_12606,N_12743);
xnor U15066 (N_15066,N_12548,N_12944);
nand U15067 (N_15067,N_14542,N_13401);
nor U15068 (N_15068,N_12635,N_14717);
nand U15069 (N_15069,N_13889,N_13157);
nand U15070 (N_15070,N_14272,N_13962);
nand U15071 (N_15071,N_13579,N_12979);
xor U15072 (N_15072,N_13077,N_14616);
nor U15073 (N_15073,N_14070,N_12773);
nand U15074 (N_15074,N_14409,N_14983);
or U15075 (N_15075,N_13953,N_14448);
nand U15076 (N_15076,N_14101,N_13087);
and U15077 (N_15077,N_14728,N_14651);
and U15078 (N_15078,N_14421,N_14030);
and U15079 (N_15079,N_12582,N_13779);
nand U15080 (N_15080,N_13368,N_12669);
nor U15081 (N_15081,N_14990,N_13078);
and U15082 (N_15082,N_14319,N_14085);
nor U15083 (N_15083,N_14559,N_13872);
xnor U15084 (N_15084,N_12860,N_14829);
and U15085 (N_15085,N_14832,N_13043);
or U15086 (N_15086,N_13022,N_12916);
or U15087 (N_15087,N_14225,N_12865);
nor U15088 (N_15088,N_14221,N_14065);
or U15089 (N_15089,N_14936,N_14863);
xor U15090 (N_15090,N_14802,N_13577);
or U15091 (N_15091,N_14033,N_13675);
and U15092 (N_15092,N_13182,N_14188);
or U15093 (N_15093,N_14439,N_13045);
and U15094 (N_15094,N_14572,N_14680);
nor U15095 (N_15095,N_13466,N_13952);
nor U15096 (N_15096,N_13822,N_12908);
nand U15097 (N_15097,N_14201,N_13349);
or U15098 (N_15098,N_14851,N_14138);
xnor U15099 (N_15099,N_14646,N_14771);
and U15100 (N_15100,N_14709,N_14742);
xnor U15101 (N_15101,N_12856,N_13904);
nor U15102 (N_15102,N_14499,N_13132);
xor U15103 (N_15103,N_13774,N_13807);
xnor U15104 (N_15104,N_14429,N_14973);
nor U15105 (N_15105,N_13212,N_12904);
or U15106 (N_15106,N_13922,N_14252);
nor U15107 (N_15107,N_14686,N_13741);
and U15108 (N_15108,N_12782,N_12601);
nor U15109 (N_15109,N_14949,N_14736);
and U15110 (N_15110,N_13334,N_13437);
nor U15111 (N_15111,N_12681,N_14089);
xnor U15112 (N_15112,N_14426,N_13826);
and U15113 (N_15113,N_14432,N_14543);
nor U15114 (N_15114,N_13601,N_13175);
xnor U15115 (N_15115,N_14060,N_14038);
nor U15116 (N_15116,N_14286,N_13919);
xnor U15117 (N_15117,N_14075,N_14337);
nand U15118 (N_15118,N_13335,N_14333);
nand U15119 (N_15119,N_14348,N_12991);
and U15120 (N_15120,N_13151,N_13938);
nand U15121 (N_15121,N_13202,N_14116);
xnor U15122 (N_15122,N_12661,N_12640);
xor U15123 (N_15123,N_14769,N_13685);
and U15124 (N_15124,N_14250,N_14372);
nor U15125 (N_15125,N_13185,N_14383);
or U15126 (N_15126,N_14080,N_12535);
or U15127 (N_15127,N_14172,N_14557);
nor U15128 (N_15128,N_14605,N_12826);
nor U15129 (N_15129,N_14522,N_13605);
nor U15130 (N_15130,N_13377,N_13793);
nand U15131 (N_15131,N_13425,N_12686);
xnor U15132 (N_15132,N_14545,N_13477);
nand U15133 (N_15133,N_13413,N_13153);
or U15134 (N_15134,N_14512,N_14561);
xor U15135 (N_15135,N_14611,N_14549);
nand U15136 (N_15136,N_13897,N_13711);
or U15137 (N_15137,N_13622,N_13109);
or U15138 (N_15138,N_12814,N_12626);
nor U15139 (N_15139,N_14456,N_12684);
and U15140 (N_15140,N_13221,N_13483);
nand U15141 (N_15141,N_13480,N_12732);
xor U15142 (N_15142,N_14305,N_12566);
and U15143 (N_15143,N_14240,N_13626);
or U15144 (N_15144,N_12585,N_13900);
nor U15145 (N_15145,N_14123,N_13438);
nor U15146 (N_15146,N_14168,N_12975);
nor U15147 (N_15147,N_14885,N_13122);
nor U15148 (N_15148,N_13417,N_13721);
or U15149 (N_15149,N_12618,N_13885);
xor U15150 (N_15150,N_13170,N_14810);
or U15151 (N_15151,N_14438,N_13770);
nor U15152 (N_15152,N_13419,N_14854);
nor U15153 (N_15153,N_12532,N_13674);
xnor U15154 (N_15154,N_14282,N_12940);
or U15155 (N_15155,N_14694,N_14342);
nand U15156 (N_15156,N_14470,N_12967);
xor U15157 (N_15157,N_13942,N_14704);
or U15158 (N_15158,N_13802,N_12690);
nor U15159 (N_15159,N_14476,N_12538);
nor U15160 (N_15160,N_12893,N_14998);
or U15161 (N_15161,N_14724,N_13440);
and U15162 (N_15162,N_13195,N_13720);
xnor U15163 (N_15163,N_14794,N_13354);
and U15164 (N_15164,N_14781,N_12579);
xnor U15165 (N_15165,N_14808,N_14835);
xnor U15166 (N_15166,N_14066,N_13594);
and U15167 (N_15167,N_12933,N_14407);
and U15168 (N_15168,N_14246,N_14285);
and U15169 (N_15169,N_13470,N_14799);
nor U15170 (N_15170,N_13532,N_14941);
or U15171 (N_15171,N_13076,N_14504);
and U15172 (N_15172,N_14668,N_13098);
or U15173 (N_15173,N_14211,N_14217);
or U15174 (N_15174,N_13412,N_14455);
or U15175 (N_15175,N_13177,N_13453);
nor U15176 (N_15176,N_13492,N_14994);
nand U15177 (N_15177,N_13515,N_14124);
and U15178 (N_15178,N_12849,N_13114);
nand U15179 (N_15179,N_12609,N_13066);
and U15180 (N_15180,N_14563,N_13844);
nand U15181 (N_15181,N_14480,N_14078);
and U15182 (N_15182,N_14500,N_13707);
nor U15183 (N_15183,N_12951,N_12808);
xor U15184 (N_15184,N_14731,N_14271);
nand U15185 (N_15185,N_13757,N_14992);
or U15186 (N_15186,N_13108,N_13348);
nand U15187 (N_15187,N_14971,N_14696);
or U15188 (N_15188,N_14626,N_14943);
nand U15189 (N_15189,N_12524,N_14048);
and U15190 (N_15190,N_13046,N_12794);
or U15191 (N_15191,N_14917,N_14725);
or U15192 (N_15192,N_12873,N_13387);
or U15193 (N_15193,N_13682,N_13914);
and U15194 (N_15194,N_13989,N_14914);
nor U15195 (N_15195,N_13189,N_14818);
or U15196 (N_15196,N_14667,N_14312);
xnor U15197 (N_15197,N_14558,N_14876);
and U15198 (N_15198,N_14705,N_13243);
nand U15199 (N_15199,N_14467,N_14142);
nand U15200 (N_15200,N_13672,N_13717);
and U15201 (N_15201,N_13376,N_14635);
nor U15202 (N_15202,N_14269,N_13615);
xor U15203 (N_15203,N_14057,N_12792);
nor U15204 (N_15204,N_14950,N_14683);
nand U15205 (N_15205,N_12950,N_14362);
nor U15206 (N_15206,N_14420,N_13949);
nor U15207 (N_15207,N_14628,N_13705);
nand U15208 (N_15208,N_13641,N_13146);
nor U15209 (N_15209,N_13841,N_12631);
nand U15210 (N_15210,N_14497,N_13606);
xnor U15211 (N_15211,N_14281,N_13421);
or U15212 (N_15212,N_13033,N_13430);
xnor U15213 (N_15213,N_12779,N_14845);
or U15214 (N_15214,N_13383,N_12696);
and U15215 (N_15215,N_13083,N_12580);
nor U15216 (N_15216,N_13983,N_12818);
and U15217 (N_15217,N_13193,N_14423);
nand U15218 (N_15218,N_14734,N_14162);
nand U15219 (N_15219,N_12561,N_14175);
nor U15220 (N_15220,N_13498,N_13612);
or U15221 (N_15221,N_13171,N_14873);
or U15222 (N_15222,N_12954,N_13758);
nor U15223 (N_15223,N_14029,N_14410);
and U15224 (N_15224,N_13293,N_14548);
and U15225 (N_15225,N_12539,N_14068);
xor U15226 (N_15226,N_14713,N_12506);
nand U15227 (N_15227,N_12784,N_13356);
or U15228 (N_15228,N_13374,N_13648);
and U15229 (N_15229,N_13392,N_14918);
nor U15230 (N_15230,N_13433,N_14005);
nor U15231 (N_15231,N_13769,N_12526);
nand U15232 (N_15232,N_14800,N_14018);
xor U15233 (N_15233,N_12984,N_13886);
nand U15234 (N_15234,N_14870,N_12747);
xor U15235 (N_15235,N_14518,N_14191);
nor U15236 (N_15236,N_14976,N_14842);
or U15237 (N_15237,N_13536,N_14666);
and U15238 (N_15238,N_12947,N_13737);
xor U15239 (N_15239,N_13379,N_14278);
xor U15240 (N_15240,N_14702,N_14274);
xnor U15241 (N_15241,N_13918,N_12902);
nand U15242 (N_15242,N_12505,N_13264);
nor U15243 (N_15243,N_14010,N_13730);
xnor U15244 (N_15244,N_13958,N_12584);
or U15245 (N_15245,N_14637,N_12544);
and U15246 (N_15246,N_14926,N_13832);
or U15247 (N_15247,N_14111,N_13851);
or U15248 (N_15248,N_14710,N_12857);
nand U15249 (N_15249,N_14791,N_14765);
nand U15250 (N_15250,N_14906,N_14302);
and U15251 (N_15251,N_12718,N_13223);
xnor U15252 (N_15252,N_13785,N_12674);
and U15253 (N_15253,N_12766,N_14916);
nor U15254 (N_15254,N_14602,N_13449);
and U15255 (N_15255,N_13265,N_14601);
or U15256 (N_15256,N_13724,N_14159);
or U15257 (N_15257,N_14757,N_14711);
and U15258 (N_15258,N_14657,N_13710);
and U15259 (N_15259,N_13858,N_12536);
nand U15260 (N_15260,N_14661,N_12644);
xor U15261 (N_15261,N_14929,N_13216);
and U15262 (N_15262,N_13263,N_14035);
xnor U15263 (N_15263,N_14828,N_13691);
nand U15264 (N_15264,N_14314,N_14884);
and U15265 (N_15265,N_13038,N_13927);
or U15266 (N_15266,N_13614,N_13116);
nor U15267 (N_15267,N_13965,N_12734);
and U15268 (N_15268,N_13284,N_14295);
xnor U15269 (N_15269,N_13968,N_13917);
and U15270 (N_15270,N_14888,N_13300);
or U15271 (N_15271,N_13472,N_13398);
and U15272 (N_15272,N_14655,N_12512);
or U15273 (N_15273,N_14405,N_13198);
or U15274 (N_15274,N_12714,N_12645);
and U15275 (N_15275,N_14861,N_12744);
or U15276 (N_15276,N_14999,N_13400);
or U15277 (N_15277,N_12879,N_13607);
nor U15278 (N_15278,N_12594,N_13570);
and U15279 (N_15279,N_14433,N_13663);
and U15280 (N_15280,N_12559,N_12762);
nor U15281 (N_15281,N_12960,N_14774);
and U15282 (N_15282,N_14233,N_14446);
xnor U15283 (N_15283,N_12797,N_13683);
and U15284 (N_15284,N_12790,N_13362);
and U15285 (N_15285,N_13107,N_14100);
and U15286 (N_15286,N_13244,N_13595);
nor U15287 (N_15287,N_13181,N_13239);
xnor U15288 (N_15288,N_12817,N_12838);
nand U15289 (N_15289,N_14566,N_13397);
nand U15290 (N_15290,N_13701,N_14143);
xnor U15291 (N_15291,N_13719,N_14921);
xnor U15292 (N_15292,N_13913,N_12702);
or U15293 (N_15293,N_14040,N_12751);
or U15294 (N_15294,N_14228,N_13011);
nor U15295 (N_15295,N_12596,N_14586);
nor U15296 (N_15296,N_12895,N_13585);
nor U15297 (N_15297,N_14154,N_12912);
xnor U15298 (N_15298,N_13227,N_14198);
xor U15299 (N_15299,N_13008,N_14937);
nand U15300 (N_15300,N_14297,N_13553);
nand U15301 (N_15301,N_14125,N_14449);
nand U15302 (N_15302,N_14913,N_13299);
nand U15303 (N_15303,N_14825,N_13298);
nor U15304 (N_15304,N_13089,N_13058);
xor U15305 (N_15305,N_12962,N_14807);
or U15306 (N_15306,N_12920,N_14569);
nand U15307 (N_15307,N_14978,N_12578);
or U15308 (N_15308,N_13875,N_13665);
and U15309 (N_15309,N_14495,N_13870);
nor U15310 (N_15310,N_12666,N_12982);
xnor U15311 (N_15311,N_12974,N_14908);
nand U15312 (N_15312,N_13745,N_13026);
and U15313 (N_15313,N_14568,N_14551);
and U15314 (N_15314,N_13056,N_14844);
xor U15315 (N_15315,N_14946,N_13964);
xnor U15316 (N_15316,N_13932,N_13950);
and U15317 (N_15317,N_13995,N_14855);
xor U15318 (N_15318,N_13732,N_13600);
or U15319 (N_15319,N_13039,N_14786);
or U15320 (N_15320,N_14378,N_13273);
or U15321 (N_15321,N_13411,N_14418);
nand U15322 (N_15322,N_12994,N_13550);
or U15323 (N_15323,N_12919,N_14308);
and U15324 (N_15324,N_13805,N_14092);
xor U15325 (N_15325,N_12883,N_14676);
nor U15326 (N_15326,N_13403,N_13773);
or U15327 (N_15327,N_14440,N_12990);
nor U15328 (N_15328,N_13912,N_14621);
nor U15329 (N_15329,N_14310,N_13036);
xnor U15330 (N_15330,N_14582,N_14508);
nor U15331 (N_15331,N_13248,N_13369);
nor U15332 (N_15332,N_12608,N_13460);
nand U15333 (N_15333,N_12736,N_14401);
and U15334 (N_15334,N_14901,N_14140);
or U15335 (N_15335,N_14795,N_14121);
or U15336 (N_15336,N_14479,N_12843);
and U15337 (N_15337,N_14967,N_14391);
nor U15338 (N_15338,N_14947,N_13652);
nand U15339 (N_15339,N_13956,N_13676);
xnor U15340 (N_15340,N_14096,N_13945);
nand U15341 (N_15341,N_13895,N_14132);
xor U15342 (N_15342,N_14014,N_13303);
or U15343 (N_15343,N_14339,N_13767);
nor U15344 (N_15344,N_14287,N_13901);
or U15345 (N_15345,N_13558,N_14979);
xnor U15346 (N_15346,N_12708,N_14892);
nor U15347 (N_15347,N_14299,N_13431);
xor U15348 (N_15348,N_13503,N_14212);
xnor U15349 (N_15349,N_13101,N_13071);
xor U15350 (N_15350,N_13023,N_13697);
nand U15351 (N_15351,N_13155,N_13133);
nand U15352 (N_15352,N_14755,N_14270);
nand U15353 (N_15353,N_12560,N_12529);
nor U15354 (N_15354,N_12807,N_13365);
nor U15355 (N_15355,N_13139,N_13013);
or U15356 (N_15356,N_12839,N_12664);
nand U15357 (N_15357,N_14816,N_12656);
and U15358 (N_15358,N_14260,N_14254);
and U15359 (N_15359,N_13222,N_13541);
nor U15360 (N_15360,N_14638,N_14307);
or U15361 (N_15361,N_14325,N_13262);
nor U15362 (N_15362,N_13138,N_13179);
or U15363 (N_15363,N_14644,N_13507);
xnor U15364 (N_15364,N_13489,N_13476);
and U15365 (N_15365,N_13260,N_14642);
or U15366 (N_15366,N_13286,N_14365);
or U15367 (N_15367,N_13324,N_13554);
and U15368 (N_15368,N_14031,N_14462);
nand U15369 (N_15369,N_14894,N_14546);
and U15370 (N_15370,N_13725,N_14954);
xor U15371 (N_15371,N_13686,N_12595);
nor U15372 (N_15372,N_14323,N_14394);
or U15373 (N_15373,N_14496,N_13632);
nand U15374 (N_15374,N_14751,N_14039);
and U15375 (N_15375,N_14131,N_14396);
or U15376 (N_15376,N_14253,N_12746);
and U15377 (N_15377,N_14133,N_13660);
xor U15378 (N_15378,N_13249,N_12574);
xnor U15379 (N_15379,N_12997,N_13128);
or U15380 (N_15380,N_13734,N_12996);
nor U15381 (N_15381,N_13176,N_12819);
nand U15382 (N_15382,N_12850,N_13130);
xor U15383 (N_15383,N_13828,N_13372);
nand U15384 (N_15384,N_14531,N_14058);
or U15385 (N_15385,N_13367,N_13051);
xor U15386 (N_15386,N_14098,N_12868);
and U15387 (N_15387,N_14215,N_13291);
or U15388 (N_15388,N_14598,N_13831);
xnor U15389 (N_15389,N_14772,N_13140);
xor U15390 (N_15390,N_13342,N_14050);
xnor U15391 (N_15391,N_13281,N_13105);
and U15392 (N_15392,N_14895,N_12914);
nor U15393 (N_15393,N_14735,N_14354);
xnor U15394 (N_15394,N_13429,N_14338);
or U15395 (N_15395,N_14044,N_12756);
and U15396 (N_15396,N_12867,N_13978);
and U15397 (N_15397,N_13065,N_14248);
or U15398 (N_15398,N_12643,N_13350);
xnor U15399 (N_15399,N_13092,N_14754);
nand U15400 (N_15400,N_12581,N_14358);
and U15401 (N_15401,N_13338,N_13224);
nand U15402 (N_15402,N_13396,N_13233);
and U15403 (N_15403,N_14458,N_14452);
nor U15404 (N_15404,N_13382,N_14414);
xor U15405 (N_15405,N_14036,N_14684);
or U15406 (N_15406,N_13706,N_13333);
nand U15407 (N_15407,N_14206,N_13811);
nor U15408 (N_15408,N_14963,N_14813);
nand U15409 (N_15409,N_13557,N_13336);
xnor U15410 (N_15410,N_13054,N_12525);
nor U15411 (N_15411,N_13235,N_13282);
and U15412 (N_15412,N_12840,N_13115);
nand U15413 (N_15413,N_12802,N_14606);
and U15414 (N_15414,N_13752,N_13608);
or U15415 (N_15415,N_14619,N_12783);
or U15416 (N_15416,N_14273,N_14032);
nor U15417 (N_15417,N_14822,N_13974);
and U15418 (N_15418,N_14406,N_13199);
or U15419 (N_15419,N_12550,N_13535);
and U15420 (N_15420,N_14072,N_13168);
or U15421 (N_15421,N_13471,N_14760);
xor U15422 (N_15422,N_12815,N_14613);
or U15423 (N_15423,N_13994,N_13015);
or U15424 (N_15424,N_13238,N_12886);
nor U15425 (N_15425,N_13768,N_13037);
nand U15426 (N_15426,N_12942,N_14700);
nand U15427 (N_15427,N_14594,N_13474);
nor U15428 (N_15428,N_13869,N_14289);
nand U15429 (N_15429,N_13731,N_14445);
or U15430 (N_15430,N_13100,N_12823);
and U15431 (N_15431,N_13016,N_12552);
nor U15432 (N_15432,N_12824,N_12973);
nand U15433 (N_15433,N_13006,N_13821);
or U15434 (N_15434,N_12809,N_14703);
or U15435 (N_15435,N_12787,N_14377);
and U15436 (N_15436,N_13694,N_13040);
and U15437 (N_15437,N_14171,N_13590);
xor U15438 (N_15438,N_14009,N_14443);
and U15439 (N_15439,N_13909,N_13709);
nand U15440 (N_15440,N_12507,N_13824);
nand U15441 (N_15441,N_13505,N_14062);
or U15442 (N_15442,N_14369,N_14292);
xor U15443 (N_15443,N_13748,N_14471);
xor U15444 (N_15444,N_12862,N_12958);
nand U15445 (N_15445,N_13564,N_13360);
nand U15446 (N_15446,N_13559,N_13225);
nand U15447 (N_15447,N_12855,N_12978);
nor U15448 (N_15448,N_13201,N_13217);
or U15449 (N_15449,N_14958,N_13539);
and U15450 (N_15450,N_13935,N_12588);
nor U15451 (N_15451,N_12998,N_14197);
and U15452 (N_15452,N_12602,N_14662);
and U15453 (N_15453,N_13316,N_13771);
and U15454 (N_15454,N_14169,N_14775);
nor U15455 (N_15455,N_12813,N_13772);
nand U15456 (N_15456,N_13887,N_13584);
or U15457 (N_15457,N_14245,N_14167);
nand U15458 (N_15458,N_13055,N_14514);
xnor U15459 (N_15459,N_14128,N_12992);
or U15460 (N_15460,N_14022,N_14244);
xnor U15461 (N_15461,N_14483,N_12798);
nand U15462 (N_15462,N_13416,N_13921);
and U15463 (N_15463,N_12949,N_14395);
nor U15464 (N_15464,N_14434,N_14831);
xnor U15465 (N_15465,N_14328,N_13254);
xor U15466 (N_15466,N_13629,N_13414);
and U15467 (N_15467,N_14919,N_14416);
or U15468 (N_15468,N_12615,N_12713);
or U15469 (N_15469,N_12654,N_13838);
xnor U15470 (N_15470,N_14087,N_13088);
xnor U15471 (N_15471,N_14837,N_14475);
or U15472 (N_15472,N_14534,N_14798);
xor U15473 (N_15473,N_12875,N_14091);
xor U15474 (N_15474,N_14466,N_14489);
nor U15475 (N_15475,N_13587,N_14298);
nand U15476 (N_15476,N_14424,N_14344);
xor U15477 (N_15477,N_14451,N_13508);
or U15478 (N_15478,N_14412,N_13528);
nand U15479 (N_15479,N_14848,N_14612);
nor U15480 (N_15480,N_12930,N_13389);
xor U15481 (N_15481,N_14675,N_13762);
xnor U15482 (N_15482,N_14153,N_12677);
and U15483 (N_15483,N_13631,N_13799);
nor U15484 (N_15484,N_14712,N_12943);
or U15485 (N_15485,N_12934,N_14617);
or U15486 (N_15486,N_13031,N_13969);
or U15487 (N_15487,N_14176,N_13269);
nor U15488 (N_15488,N_14106,N_13788);
and U15489 (N_15489,N_14893,N_12810);
nor U15490 (N_15490,N_12676,N_12557);
and U15491 (N_15491,N_12546,N_14021);
or U15492 (N_15492,N_14674,N_14905);
nand U15493 (N_15493,N_14204,N_13650);
xnor U15494 (N_15494,N_12806,N_12881);
nand U15495 (N_15495,N_14592,N_13211);
or U15496 (N_15496,N_14043,N_14588);
nand U15497 (N_15497,N_13746,N_14052);
nand U15498 (N_15498,N_14706,N_13977);
nand U15499 (N_15499,N_14166,N_14232);
and U15500 (N_15500,N_12793,N_12649);
xnor U15501 (N_15501,N_13794,N_14507);
or U15502 (N_15502,N_13125,N_14311);
xor U15503 (N_15503,N_13075,N_14524);
nand U15504 (N_15504,N_13653,N_13586);
nor U15505 (N_15505,N_12607,N_13647);
nor U15506 (N_15506,N_14408,N_13712);
xnor U15507 (N_15507,N_13473,N_13319);
nand U15508 (N_15508,N_13544,N_13796);
xnor U15509 (N_15509,N_14687,N_13551);
nand U15510 (N_15510,N_12628,N_14847);
or U15511 (N_15511,N_12966,N_13070);
nor U15512 (N_15512,N_14871,N_14745);
nand U15513 (N_15513,N_12616,N_12926);
or U15514 (N_15514,N_14017,N_14360);
nand U15515 (N_15515,N_13902,N_13680);
nand U15516 (N_15516,N_12832,N_14766);
or U15517 (N_15517,N_12500,N_14793);
nand U15518 (N_15518,N_13504,N_13352);
nand U15519 (N_15519,N_12922,N_14962);
nand U15520 (N_15520,N_14960,N_13847);
or U15521 (N_15521,N_12972,N_13659);
or U15522 (N_15522,N_12911,N_14538);
or U15523 (N_15523,N_14819,N_13361);
nand U15524 (N_15524,N_14055,N_14746);
nand U15525 (N_15525,N_14860,N_14714);
and U15526 (N_15526,N_14404,N_14575);
xor U15527 (N_15527,N_13159,N_14136);
nand U15528 (N_15528,N_13776,N_14202);
nor U15529 (N_15529,N_13860,N_12624);
nor U15530 (N_15530,N_12692,N_12983);
or U15531 (N_15531,N_14510,N_14368);
nor U15532 (N_15532,N_13020,N_13723);
and U15533 (N_15533,N_13104,N_14977);
or U15534 (N_15534,N_14948,N_14079);
xnor U15535 (N_15535,N_14151,N_14134);
nor U15536 (N_15536,N_14526,N_13543);
and U15537 (N_15537,N_14207,N_14749);
or U15538 (N_15538,N_13990,N_12629);
and U15539 (N_15539,N_12551,N_13378);
and U15540 (N_15540,N_14540,N_12976);
nand U15541 (N_15541,N_12605,N_13915);
nand U15542 (N_15542,N_14255,N_14743);
nand U15543 (N_15543,N_13980,N_13761);
nor U15544 (N_15544,N_13708,N_12516);
xnor U15545 (N_15545,N_14350,N_14672);
xor U15546 (N_15546,N_13703,N_12742);
nand U15547 (N_15547,N_13923,N_14220);
nor U15548 (N_15548,N_13864,N_14883);
nor U15549 (N_15549,N_13736,N_13247);
nor U15550 (N_15550,N_13329,N_12623);
or U15551 (N_15551,N_14477,N_12598);
xor U15552 (N_15552,N_13405,N_13582);
nand U15553 (N_15553,N_14002,N_13654);
or U15554 (N_15554,N_14618,N_14478);
nand U15555 (N_15555,N_12547,N_13381);
xor U15556 (N_15556,N_14516,N_13250);
or U15557 (N_15557,N_14996,N_13261);
or U15558 (N_15558,N_12924,N_13085);
xor U15559 (N_15559,N_14317,N_12828);
xor U15560 (N_15560,N_13292,N_13390);
xnor U15561 (N_15561,N_14099,N_13861);
and U15562 (N_15562,N_14796,N_12891);
or U15563 (N_15563,N_14730,N_14552);
xnor U15564 (N_15564,N_14320,N_13213);
nor U15565 (N_15565,N_13347,N_12937);
xor U15566 (N_15566,N_13258,N_12622);
or U15567 (N_15567,N_13666,N_14388);
and U15568 (N_15568,N_12503,N_14422);
xnor U15569 (N_15569,N_14624,N_13642);
xor U15570 (N_15570,N_14047,N_13891);
nor U15571 (N_15571,N_14523,N_14294);
xnor U15572 (N_15572,N_12786,N_12765);
xnor U15573 (N_15573,N_12599,N_14923);
nor U15574 (N_15574,N_12804,N_12957);
or U15575 (N_15575,N_12768,N_13237);
and U15576 (N_15576,N_13141,N_14322);
and U15577 (N_15577,N_12864,N_13874);
xnor U15578 (N_15578,N_13328,N_14903);
xnor U15579 (N_15579,N_12858,N_12936);
nor U15580 (N_15580,N_12753,N_13161);
nand U15581 (N_15581,N_13704,N_14083);
nand U15582 (N_15582,N_14707,N_13452);
and U15583 (N_15583,N_13332,N_13552);
and U15584 (N_15584,N_14373,N_13003);
and U15585 (N_15585,N_13542,N_14093);
xnor U15586 (N_15586,N_13009,N_13072);
xor U15587 (N_15587,N_14069,N_13304);
nor U15588 (N_15588,N_13546,N_14145);
nor U15589 (N_15589,N_12636,N_13059);
or U15590 (N_15590,N_13651,N_13308);
xnor U15591 (N_15591,N_14758,N_14852);
nand U15592 (N_15592,N_12754,N_14004);
xnor U15593 (N_15593,N_14955,N_14669);
or U15594 (N_15594,N_14838,N_12898);
and U15595 (N_15595,N_12811,N_14417);
or U15596 (N_15596,N_13760,N_12688);
nand U15597 (N_15597,N_14331,N_14150);
nor U15598 (N_15598,N_13275,N_14236);
or U15599 (N_15599,N_13530,N_14024);
and U15600 (N_15600,N_13512,N_14103);
nor U15601 (N_15601,N_14193,N_12728);
nor U15602 (N_15602,N_14425,N_14506);
and U15603 (N_15603,N_14752,N_14665);
nor U15604 (N_15604,N_13279,N_14957);
nand U15605 (N_15605,N_13206,N_13893);
xor U15606 (N_15606,N_13418,N_13533);
or U15607 (N_15607,N_13135,N_14649);
nand U15608 (N_15608,N_14243,N_13363);
or U15609 (N_15609,N_12646,N_14525);
nor U15610 (N_15610,N_13700,N_13482);
nor U15611 (N_15611,N_14609,N_13880);
xor U15612 (N_15612,N_12748,N_14866);
and U15613 (N_15613,N_14104,N_14850);
and U15614 (N_15614,N_12711,N_13005);
and U15615 (N_15615,N_14597,N_13813);
xor U15616 (N_15616,N_13465,N_13925);
or U15617 (N_15617,N_13988,N_12884);
nand U15618 (N_15618,N_13754,N_13859);
xnor U15619 (N_15619,N_14580,N_14629);
and U15620 (N_15620,N_14363,N_13529);
or U15621 (N_15621,N_14263,N_14450);
nand U15622 (N_15622,N_12985,N_14487);
and U15623 (N_15623,N_14330,N_12575);
nor U15624 (N_15624,N_13823,N_14723);
or U15625 (N_15625,N_14900,N_14019);
nand U15626 (N_15626,N_13854,N_14726);
nor U15627 (N_15627,N_13455,N_14279);
and U15628 (N_15628,N_14280,N_13803);
nor U15629 (N_15629,N_12725,N_14013);
xor U15630 (N_15630,N_12511,N_12603);
nor U15631 (N_15631,N_12772,N_13355);
xor U15632 (N_15632,N_12504,N_13936);
nor U15633 (N_15633,N_14411,N_13593);
nand U15634 (N_15634,N_14301,N_12658);
nand U15635 (N_15635,N_14315,N_12952);
and U15636 (N_15636,N_14304,N_13226);
nand U15637 (N_15637,N_14988,N_13167);
and U15638 (N_15638,N_12841,N_13395);
nor U15639 (N_15639,N_13693,N_13126);
xnor U15640 (N_15640,N_14801,N_13749);
nor U15641 (N_15641,N_14985,N_13894);
nor U15642 (N_15642,N_13792,N_12721);
nor U15643 (N_15643,N_13044,N_14041);
nand U15644 (N_15644,N_14234,N_12777);
nor U15645 (N_15645,N_12993,N_14074);
nand U15646 (N_15646,N_13144,N_13698);
and U15647 (N_15647,N_13976,N_12763);
nor U15648 (N_15648,N_13537,N_12767);
nand U15649 (N_15649,N_14251,N_14158);
nor U15650 (N_15650,N_12929,N_14332);
and U15651 (N_15651,N_13954,N_13842);
nor U15652 (N_15652,N_12567,N_13345);
and U15653 (N_15653,N_13910,N_14738);
xor U15654 (N_15654,N_13408,N_13163);
or U15655 (N_15655,N_12866,N_13245);
nand U15656 (N_15656,N_14869,N_12639);
nor U15657 (N_15657,N_13798,N_14222);
or U15658 (N_15658,N_14195,N_13002);
nor U15659 (N_15659,N_13671,N_14006);
and U15660 (N_15660,N_14995,N_13322);
and U15661 (N_15661,N_14067,N_14762);
or U15662 (N_15662,N_13572,N_14095);
and U15663 (N_15663,N_12715,N_14610);
and U15664 (N_15664,N_14102,N_12641);
nor U15665 (N_15665,N_13853,N_14316);
nand U15666 (N_15666,N_12870,N_13905);
nand U15667 (N_15667,N_12627,N_14177);
and U15668 (N_15668,N_12689,N_14178);
or U15669 (N_15669,N_14741,N_13728);
nor U15670 (N_15670,N_13380,N_13399);
xor U15671 (N_15671,N_13320,N_14390);
xor U15672 (N_15672,N_14763,N_14239);
xnor U15673 (N_15673,N_13829,N_14398);
nor U15674 (N_15674,N_12745,N_13491);
and U15675 (N_15675,N_14737,N_14896);
or U15676 (N_15676,N_13280,N_13145);
nand U15677 (N_15677,N_13457,N_14345);
or U15678 (N_15678,N_13866,N_13747);
nand U15679 (N_15679,N_14951,N_14353);
and U15680 (N_15680,N_13053,N_13973);
xor U15681 (N_15681,N_12528,N_13450);
nand U15682 (N_15682,N_14226,N_14073);
and U15683 (N_15683,N_14447,N_14770);
or U15684 (N_15684,N_14583,N_13568);
xor U15685 (N_15685,N_13836,N_14023);
nor U15686 (N_15686,N_13049,N_13943);
or U15687 (N_15687,N_14472,N_14841);
or U15688 (N_15688,N_12761,N_12903);
or U15689 (N_15689,N_13797,N_13510);
or U15690 (N_15690,N_13742,N_13596);
nand U15691 (N_15691,N_13787,N_13021);
and U15692 (N_15692,N_13643,N_14928);
or U15693 (N_15693,N_13565,N_14932);
or U15694 (N_15694,N_14352,N_13394);
nand U15695 (N_15695,N_13649,N_14386);
or U15696 (N_15696,N_14864,N_14779);
xor U15697 (N_15697,N_14097,N_12845);
xnor U15698 (N_15698,N_13097,N_13930);
and U15699 (N_15699,N_13129,N_13446);
xor U15700 (N_15700,N_12859,N_14084);
xnor U15701 (N_15701,N_12521,N_14016);
or U15702 (N_15702,N_13566,N_13667);
nor U15703 (N_15703,N_14293,N_12821);
xnor U15704 (N_15704,N_13207,N_13743);
and U15705 (N_15705,N_13555,N_13611);
and U15706 (N_15706,N_14987,N_13311);
nand U15707 (N_15707,N_13353,N_12612);
nor U15708 (N_15708,N_13276,N_14081);
nor U15709 (N_15709,N_13845,N_13407);
nand U15710 (N_15710,N_14634,N_13940);
nor U15711 (N_15711,N_12851,N_13624);
or U15712 (N_15712,N_14826,N_14403);
and U15713 (N_15713,N_14812,N_14415);
nand U15714 (N_15714,N_13609,N_13034);
and U15715 (N_15715,N_14061,N_14584);
xor U15716 (N_15716,N_14636,N_12738);
and U15717 (N_15717,N_13493,N_13583);
or U15718 (N_15718,N_14521,N_14219);
and U15719 (N_15719,N_14997,N_13461);
nor U15720 (N_15720,N_14930,N_13357);
and U15721 (N_15721,N_12965,N_14944);
xnor U15722 (N_15722,N_14491,N_13625);
and U15723 (N_15723,N_13781,N_12963);
nor U15724 (N_15724,N_13318,N_12825);
and U15725 (N_15725,N_13789,N_14231);
or U15726 (N_15726,N_12871,N_12619);
nor U15727 (N_15727,N_14327,N_14241);
or U15728 (N_15728,N_13855,N_14604);
and U15729 (N_15729,N_14753,N_14615);
or U15730 (N_15730,N_14740,N_14677);
xnor U15731 (N_15731,N_13093,N_13563);
nand U15732 (N_15732,N_13884,N_14532);
nand U15733 (N_15733,N_12673,N_13830);
nand U15734 (N_15734,N_14938,N_14722);
xnor U15735 (N_15735,N_14460,N_13236);
xor U15736 (N_15736,N_14953,N_13645);
nor U15737 (N_15737,N_13696,N_12592);
nor U15738 (N_15738,N_14587,N_14482);
and U15739 (N_15739,N_14326,N_12837);
and U15740 (N_15740,N_13295,N_14283);
nor U15741 (N_15741,N_13981,N_13131);
xnor U15742 (N_15742,N_13444,N_14110);
and U15743 (N_15743,N_12953,N_13137);
nor U15744 (N_15744,N_13778,N_14459);
or U15745 (N_15745,N_12848,N_13739);
nor U15746 (N_15746,N_14129,N_13868);
xnor U15747 (N_15747,N_12759,N_13928);
or U15748 (N_15748,N_14519,N_13057);
nor U15749 (N_15749,N_12774,N_13992);
nand U15750 (N_15750,N_12659,N_13818);
xnor U15751 (N_15751,N_14645,N_13934);
and U15752 (N_15752,N_13755,N_13714);
and U15753 (N_15753,N_13516,N_13509);
nand U15754 (N_15754,N_12827,N_14940);
and U15755 (N_15755,N_14509,N_14520);
nor U15756 (N_15756,N_14640,N_13871);
nor U15757 (N_15757,N_12687,N_12569);
nor U15758 (N_15758,N_13306,N_14681);
nand U15759 (N_15759,N_13192,N_13636);
nor U15760 (N_15760,N_12716,N_13160);
nand U15761 (N_15761,N_14015,N_13795);
and U15762 (N_15762,N_13240,N_12508);
xor U15763 (N_15763,N_14042,N_14868);
nor U15764 (N_15764,N_14593,N_14690);
xor U15765 (N_15765,N_13873,N_14915);
nor U15766 (N_15766,N_13196,N_12853);
nor U15767 (N_15767,N_13074,N_14830);
nor U15768 (N_15768,N_13294,N_14622);
and U15769 (N_15769,N_14370,N_14364);
xor U15770 (N_15770,N_14879,N_13946);
or U15771 (N_15771,N_12709,N_13099);
nor U15772 (N_15772,N_14194,N_14114);
nand U15773 (N_15773,N_13339,N_14744);
nor U15774 (N_15774,N_14909,N_13257);
and U15775 (N_15775,N_13947,N_13061);
nand U15776 (N_15776,N_14623,N_12939);
and U15777 (N_15777,N_13916,N_13616);
and U15778 (N_15778,N_13152,N_14119);
xnor U15779 (N_15779,N_14468,N_14956);
nor U15780 (N_15780,N_12655,N_13343);
nand U15781 (N_15781,N_13191,N_14671);
nor U15782 (N_15782,N_13373,N_13944);
and U15783 (N_15783,N_12737,N_13970);
or U15784 (N_15784,N_14268,N_13948);
nor U15785 (N_15785,N_14933,N_14257);
xnor U15786 (N_15786,N_13991,N_14109);
xnor U15787 (N_15787,N_14969,N_12733);
and U15788 (N_15788,N_12969,N_14564);
nand U15789 (N_15789,N_12820,N_13113);
xnor U15790 (N_15790,N_13428,N_13766);
or U15791 (N_15791,N_14902,N_14356);
nor U15792 (N_15792,N_13527,N_13166);
nor U15793 (N_15793,N_12948,N_13426);
nor U15794 (N_15794,N_12980,N_13230);
and U15795 (N_15795,N_14699,N_14115);
nand U15796 (N_15796,N_13084,N_13232);
xnor U15797 (N_15797,N_14501,N_12816);
xor U15798 (N_15798,N_14343,N_14046);
or U15799 (N_15799,N_14562,N_14815);
or U15800 (N_15800,N_13722,N_13172);
nor U15801 (N_15801,N_14502,N_12695);
or U15802 (N_15802,N_14965,N_14814);
or U15803 (N_15803,N_14993,N_12722);
nor U15804 (N_15804,N_13127,N_14288);
and U15805 (N_15805,N_13892,N_12693);
nand U15806 (N_15806,N_14827,N_14682);
and U15807 (N_15807,N_13547,N_13435);
and U15808 (N_15808,N_14007,N_13906);
xnor U15809 (N_15809,N_13627,N_13079);
nand U15810 (N_15810,N_12701,N_12915);
nor U15811 (N_15811,N_13183,N_14484);
or U15812 (N_15812,N_14464,N_14608);
and U15813 (N_15813,N_13346,N_14727);
and U15814 (N_15814,N_14790,N_13143);
or U15815 (N_15815,N_14565,N_14397);
nor U15816 (N_15816,N_14887,N_13630);
and U15817 (N_15817,N_14340,N_12913);
or U15818 (N_15818,N_13639,N_14719);
or U15819 (N_15819,N_12591,N_14120);
xnor U15820 (N_15820,N_13780,N_12630);
xnor U15821 (N_15821,N_12842,N_13882);
xor U15822 (N_15822,N_14012,N_14064);
and U15823 (N_15823,N_12833,N_13103);
xor U15824 (N_15824,N_14867,N_12791);
nor U15825 (N_15825,N_14567,N_13520);
nor U15826 (N_15826,N_13173,N_13751);
nand U15827 (N_15827,N_14553,N_14804);
nand U15828 (N_15828,N_14473,N_13086);
and U15829 (N_15829,N_12932,N_14493);
and U15830 (N_15830,N_13580,N_12897);
nand U15831 (N_15831,N_12847,N_14179);
nor U15832 (N_15832,N_13784,N_12651);
or U15833 (N_15833,N_14784,N_14148);
xor U15834 (N_15834,N_13911,N_14716);
xnor U15835 (N_15835,N_14431,N_13715);
xor U15836 (N_15836,N_13960,N_14759);
xor U15837 (N_15837,N_14783,N_13815);
or U15838 (N_15838,N_14335,N_13951);
nand U15839 (N_15839,N_13241,N_13806);
and U15840 (N_15840,N_13617,N_13765);
and U15841 (N_15841,N_12938,N_14695);
nor U15842 (N_15842,N_13848,N_14750);
and U15843 (N_15843,N_12719,N_14708);
nor U15844 (N_15844,N_12712,N_12617);
or U15845 (N_15845,N_14152,N_13415);
nand U15846 (N_15846,N_13330,N_13782);
and U15847 (N_15847,N_13574,N_14276);
xnor U15848 (N_15848,N_13063,N_14296);
or U15849 (N_15849,N_14899,N_14261);
nor U15850 (N_15850,N_12589,N_14924);
nor U15851 (N_15851,N_14981,N_14454);
and U15852 (N_15852,N_12558,N_14607);
or U15853 (N_15853,N_13638,N_13404);
xor U15854 (N_15854,N_12675,N_13111);
nand U15855 (N_15855,N_14183,N_13229);
nor U15856 (N_15856,N_14313,N_13569);
or U15857 (N_15857,N_13197,N_13106);
nand U15858 (N_15858,N_14437,N_14547);
nand U15859 (N_15859,N_14165,N_14660);
nor U15860 (N_15860,N_13047,N_12941);
nand U15861 (N_15861,N_13359,N_14399);
and U15862 (N_15862,N_13231,N_13285);
nor U15863 (N_15863,N_13863,N_13817);
or U15864 (N_15864,N_12899,N_13190);
nand U15865 (N_15865,N_14190,N_12799);
and U15866 (N_15866,N_14968,N_14208);
nand U15867 (N_15867,N_13274,N_12835);
xor U15868 (N_15868,N_14959,N_14400);
nor U15869 (N_15869,N_13840,N_14223);
nor U15870 (N_15870,N_13786,N_12650);
nand U15871 (N_15871,N_13017,N_14964);
and U15872 (N_15872,N_13985,N_13048);
and U15873 (N_15873,N_12517,N_13497);
nand U15874 (N_15874,N_13808,N_13307);
nor U15875 (N_15875,N_13979,N_12770);
nand U15876 (N_15876,N_13290,N_12844);
or U15877 (N_15877,N_14351,N_13735);
nand U15878 (N_15878,N_12520,N_13121);
and U15879 (N_15879,N_12968,N_14589);
xnor U15880 (N_15880,N_14059,N_14515);
xor U15881 (N_15881,N_14785,N_12634);
and U15882 (N_15882,N_13200,N_12614);
nand U15883 (N_15883,N_14945,N_12758);
xnor U15884 (N_15884,N_13432,N_14367);
or U15885 (N_15885,N_12545,N_12682);
xor U15886 (N_15886,N_12890,N_14488);
or U15887 (N_15887,N_13165,N_12795);
and U15888 (N_15888,N_13317,N_13519);
nand U15889 (N_15889,N_14126,N_13538);
or U15890 (N_15890,N_13571,N_13525);
or U15891 (N_15891,N_14817,N_12812);
or U15892 (N_15892,N_14380,N_14026);
xnor U15893 (N_15893,N_14528,N_14761);
xnor U15894 (N_15894,N_14155,N_13327);
and U15895 (N_15895,N_14633,N_12600);
nor U15896 (N_15896,N_14931,N_14910);
nor U15897 (N_15897,N_13313,N_13521);
xnor U15898 (N_15898,N_13825,N_12780);
nand U15899 (N_15899,N_12921,N_13214);
xor U15900 (N_15900,N_13562,N_13656);
nor U15901 (N_15901,N_14366,N_12501);
or U15902 (N_15902,N_14164,N_12987);
or U15903 (N_15903,N_14897,N_14486);
xor U15904 (N_15904,N_14627,N_13331);
xor U15905 (N_15905,N_14843,N_13366);
nor U15906 (N_15906,N_14625,N_14453);
and U15907 (N_15907,N_13208,N_14144);
and U15908 (N_15908,N_13637,N_13069);
nor U15909 (N_15909,N_12836,N_13955);
nand U15910 (N_15910,N_14620,N_12679);
and U15911 (N_15911,N_12729,N_13657);
nand U15912 (N_15912,N_13422,N_13677);
or U15913 (N_15913,N_14122,N_13479);
nor U15914 (N_15914,N_13982,N_12775);
or U15915 (N_15915,N_14911,N_12710);
nand U15916 (N_15916,N_13903,N_12667);
nand U15917 (N_15917,N_12778,N_14393);
nor U15918 (N_15918,N_14780,N_13987);
and U15919 (N_15919,N_13644,N_13926);
nor U15920 (N_15920,N_13305,N_14441);
nor U15921 (N_15921,N_14376,N_12830);
nor U15922 (N_15922,N_13613,N_13164);
and U15923 (N_15923,N_12597,N_14782);
or U15924 (N_15924,N_12760,N_14135);
nand U15925 (N_15925,N_13534,N_13834);
and U15926 (N_15926,N_12986,N_12800);
or U15927 (N_15927,N_13277,N_13827);
or U15928 (N_15928,N_13581,N_12562);
xnor U15929 (N_15929,N_13862,N_14229);
nor U15930 (N_15930,N_13496,N_14108);
or U15931 (N_15931,N_12727,N_12882);
xnor U15932 (N_15932,N_14334,N_14991);
nand U15933 (N_15933,N_14141,N_12586);
and U15934 (N_15934,N_12704,N_13178);
or U15935 (N_15935,N_13154,N_13494);
nor U15936 (N_15936,N_14778,N_13800);
or U15937 (N_15937,N_14834,N_13975);
nor U15938 (N_15938,N_13633,N_12571);
and U15939 (N_15939,N_13019,N_13091);
nand U15940 (N_15940,N_14777,N_14550);
xor U15941 (N_15941,N_12522,N_13879);
or U15942 (N_15942,N_14641,N_12731);
and U15943 (N_15943,N_14318,N_12670);
or U15944 (N_15944,N_13325,N_13358);
or U15945 (N_15945,N_14284,N_13120);
nand U15946 (N_15946,N_12955,N_13256);
nand U15947 (N_15947,N_13441,N_13628);
or U15948 (N_15948,N_14823,N_14107);
or U15949 (N_15949,N_12752,N_14748);
nor U15950 (N_15950,N_13219,N_14336);
nor U15951 (N_15951,N_14986,N_13242);
and U15952 (N_15952,N_13486,N_13684);
nor U15953 (N_15953,N_12678,N_14184);
or U15954 (N_15954,N_12652,N_14186);
nand U15955 (N_15955,N_13312,N_14498);
or U15956 (N_15956,N_14925,N_13149);
nor U15957 (N_15957,N_13576,N_14578);
nand U15958 (N_15958,N_13966,N_13014);
and U15959 (N_15959,N_12570,N_13314);
nor U15960 (N_15960,N_13618,N_14118);
or U15961 (N_15961,N_12720,N_14413);
or U15962 (N_15962,N_13888,N_12863);
nor U15963 (N_15963,N_13518,N_13062);
xnor U15964 (N_15964,N_12872,N_13124);
and U15965 (N_15965,N_14574,N_13032);
or U15966 (N_15966,N_12665,N_12621);
nand U15967 (N_15967,N_12540,N_13678);
and U15968 (N_15968,N_12685,N_13658);
nand U15969 (N_15969,N_12964,N_14579);
nand U15970 (N_15970,N_14853,N_13876);
or U15971 (N_15971,N_14277,N_12730);
or U15972 (N_15972,N_12537,N_14659);
or U15973 (N_15973,N_13468,N_12632);
nand U15974 (N_15974,N_13375,N_12834);
nor U15975 (N_15975,N_14881,N_12604);
xor U15976 (N_15976,N_14034,N_14187);
xnor U15977 (N_15977,N_13738,N_14833);
xnor U15978 (N_15978,N_12553,N_14387);
nand U15979 (N_15979,N_14982,N_13302);
nand U15980 (N_15980,N_12657,N_13439);
xnor U15981 (N_15981,N_13150,N_14658);
nand U15982 (N_15982,N_14213,N_12946);
or U15983 (N_15983,N_14419,N_12887);
nand U15984 (N_15984,N_14077,N_14086);
and U15985 (N_15985,N_12523,N_13599);
nor U15986 (N_15986,N_14632,N_12707);
and U15987 (N_15987,N_14182,N_12945);
nand U15988 (N_15988,N_13673,N_14355);
xnor U15989 (N_15989,N_14889,N_13485);
nand U15990 (N_15990,N_14349,N_12977);
nand U15991 (N_15991,N_13702,N_14882);
nor U15992 (N_15992,N_14849,N_12970);
and U15993 (N_15993,N_12541,N_13931);
nand U15994 (N_15994,N_14630,N_12900);
nand U15995 (N_15995,N_12530,N_14576);
nor U15996 (N_15996,N_14573,N_14037);
nor U15997 (N_15997,N_13655,N_14732);
or U15998 (N_15998,N_14839,N_12894);
and U15999 (N_15999,N_13220,N_13883);
nand U16000 (N_16000,N_14359,N_13517);
xor U16001 (N_16001,N_13939,N_14912);
xor U16002 (N_16002,N_13341,N_14256);
or U16003 (N_16003,N_13462,N_13640);
and U16004 (N_16004,N_12717,N_13899);
or U16005 (N_16005,N_14262,N_13060);
nor U16006 (N_16006,N_14776,N_13344);
nand U16007 (N_16007,N_14461,N_14071);
and U16008 (N_16008,N_14698,N_14003);
and U16009 (N_16009,N_12502,N_12769);
nor U16010 (N_16010,N_13664,N_13007);
nor U16011 (N_16011,N_12995,N_13810);
nand U16012 (N_16012,N_13963,N_13783);
nor U16013 (N_16013,N_13597,N_13718);
and U16014 (N_16014,N_13484,N_14972);
or U16015 (N_16015,N_12889,N_14105);
or U16016 (N_16016,N_13775,N_13142);
xor U16017 (N_16017,N_14787,N_13933);
or U16018 (N_16018,N_14663,N_12822);
and U16019 (N_16019,N_14199,N_14238);
xor U16020 (N_16020,N_14577,N_13246);
nor U16021 (N_16021,N_13134,N_13259);
and U16022 (N_16022,N_12587,N_13839);
xor U16023 (N_16023,N_13619,N_14935);
or U16024 (N_16024,N_13406,N_13205);
and U16025 (N_16025,N_14898,N_13890);
nand U16026 (N_16026,N_13523,N_13522);
and U16027 (N_16027,N_13402,N_13623);
xnor U16028 (N_16028,N_14485,N_12896);
and U16029 (N_16029,N_14265,N_13289);
xor U16030 (N_16030,N_14904,N_14160);
xor U16031 (N_16031,N_14113,N_14266);
xor U16032 (N_16032,N_13456,N_13687);
nor U16033 (N_16033,N_14688,N_13843);
or U16034 (N_16034,N_13052,N_14149);
and U16035 (N_16035,N_13549,N_13592);
or U16036 (N_16036,N_14011,N_13865);
xor U16037 (N_16037,N_14678,N_13110);
and U16038 (N_16038,N_14768,N_14444);
xnor U16039 (N_16039,N_13050,N_12514);
and U16040 (N_16040,N_13370,N_14196);
or U16041 (N_16041,N_13924,N_14020);
xnor U16042 (N_16042,N_12576,N_12999);
xnor U16043 (N_16043,N_14130,N_13690);
and U16044 (N_16044,N_13271,N_14820);
nor U16045 (N_16045,N_12705,N_14200);
nor U16046 (N_16046,N_14347,N_13695);
xnor U16047 (N_16047,N_12513,N_14872);
nand U16048 (N_16048,N_14733,N_13621);
xnor U16049 (N_16049,N_13180,N_12861);
and U16050 (N_16050,N_12961,N_12805);
nand U16051 (N_16051,N_13610,N_14492);
nor U16052 (N_16052,N_13996,N_14856);
or U16053 (N_16053,N_13561,N_14747);
or U16054 (N_16054,N_12956,N_12885);
nand U16055 (N_16055,N_13929,N_13896);
nand U16056 (N_16056,N_14181,N_12573);
and U16057 (N_16057,N_13475,N_14025);
xnor U16058 (N_16058,N_13986,N_13025);
or U16059 (N_16059,N_12981,N_13080);
xnor U16060 (N_16060,N_14209,N_14156);
or U16061 (N_16061,N_14237,N_12698);
nor U16062 (N_16062,N_14382,N_13997);
xor U16063 (N_16063,N_14952,N_14596);
nand U16064 (N_16064,N_13156,N_12625);
nor U16065 (N_16065,N_14218,N_14721);
nor U16066 (N_16066,N_13920,N_13488);
nor U16067 (N_16067,N_13502,N_13941);
nand U16068 (N_16068,N_14247,N_14174);
nor U16069 (N_16069,N_14554,N_14697);
or U16070 (N_16070,N_14664,N_13123);
nor U16071 (N_16071,N_12874,N_13041);
and U16072 (N_16072,N_14309,N_13215);
nor U16073 (N_16073,N_14788,N_13907);
or U16074 (N_16074,N_13556,N_13162);
nor U16075 (N_16075,N_14792,N_12518);
or U16076 (N_16076,N_14290,N_12869);
nand U16077 (N_16077,N_13391,N_13500);
and U16078 (N_16078,N_13251,N_14805);
xor U16079 (N_16079,N_12735,N_13790);
nand U16080 (N_16080,N_13669,N_14427);
xnor U16081 (N_16081,N_13801,N_14877);
or U16082 (N_16082,N_14189,N_13867);
nand U16083 (N_16083,N_13000,N_14880);
and U16084 (N_16084,N_14258,N_13540);
and U16085 (N_16085,N_13726,N_12694);
and U16086 (N_16086,N_13727,N_13309);
nand U16087 (N_16087,N_12647,N_14090);
xnor U16088 (N_16088,N_13315,N_13740);
nor U16089 (N_16089,N_13268,N_12831);
nor U16090 (N_16090,N_13560,N_13067);
xor U16091 (N_16091,N_13506,N_12611);
and U16092 (N_16092,N_13481,N_13024);
nand U16093 (N_16093,N_14173,N_14639);
and U16094 (N_16094,N_13816,N_12927);
nand U16095 (N_16095,N_13288,N_13427);
nor U16096 (N_16096,N_12613,N_13210);
and U16097 (N_16097,N_12878,N_13812);
nor U16098 (N_16098,N_14300,N_14739);
and U16099 (N_16099,N_13511,N_13445);
nor U16100 (N_16100,N_14811,N_14384);
and U16101 (N_16101,N_14494,N_13267);
xnor U16102 (N_16102,N_14082,N_13384);
nand U16103 (N_16103,N_13228,N_13297);
xor U16104 (N_16104,N_14729,N_13635);
xnor U16105 (N_16105,N_14137,N_14878);
nor U16106 (N_16106,N_14920,N_13662);
nand U16107 (N_16107,N_12509,N_12739);
xor U16108 (N_16108,N_13756,N_14585);
nor U16109 (N_16109,N_13681,N_14205);
nand U16110 (N_16110,N_14539,N_14927);
and U16111 (N_16111,N_13323,N_14536);
nor U16112 (N_16112,N_13972,N_12931);
and U16113 (N_16113,N_13763,N_13287);
or U16114 (N_16114,N_14648,N_14541);
or U16115 (N_16115,N_13218,N_13467);
and U16116 (N_16116,N_13203,N_13278);
nor U16117 (N_16117,N_13436,N_12700);
nor U16118 (N_16118,N_13351,N_14840);
nand U16119 (N_16119,N_12542,N_14653);
xor U16120 (N_16120,N_12776,N_13959);
or U16121 (N_16121,N_12880,N_13849);
or U16122 (N_16122,N_12764,N_13035);
xnor U16123 (N_16123,N_13575,N_13598);
or U16124 (N_16124,N_13194,N_14974);
nor U16125 (N_16125,N_13187,N_14513);
nor U16126 (N_16126,N_14650,N_12703);
xor U16127 (N_16127,N_14806,N_12662);
or U16128 (N_16128,N_13759,N_13030);
nand U16129 (N_16129,N_13393,N_13004);
xor U16130 (N_16130,N_14027,N_13620);
or U16131 (N_16131,N_12801,N_13018);
or U16132 (N_16132,N_13283,N_14803);
nand U16133 (N_16133,N_14890,N_14249);
nand U16134 (N_16134,N_12543,N_13424);
nand U16135 (N_16135,N_14693,N_13967);
nor U16136 (N_16136,N_13028,N_14647);
nand U16137 (N_16137,N_14192,N_14127);
or U16138 (N_16138,N_12706,N_14874);
and U16139 (N_16139,N_14857,N_13270);
xor U16140 (N_16140,N_12755,N_14652);
or U16141 (N_16141,N_14381,N_13326);
or U16142 (N_16142,N_14984,N_13814);
nor U16143 (N_16143,N_12892,N_13478);
nor U16144 (N_16144,N_13501,N_14934);
xor U16145 (N_16145,N_14428,N_12989);
and U16146 (N_16146,N_13463,N_14505);
nand U16147 (N_16147,N_13688,N_12637);
or U16148 (N_16148,N_13764,N_14537);
nand U16149 (N_16149,N_14163,N_14767);
nor U16150 (N_16150,N_14556,N_13602);
and U16151 (N_16151,N_14692,N_12671);
and U16152 (N_16152,N_14357,N_13443);
or U16153 (N_16153,N_13094,N_12691);
and U16154 (N_16154,N_13119,N_14614);
xnor U16155 (N_16155,N_13898,N_12568);
and U16156 (N_16156,N_12620,N_13699);
or U16157 (N_16157,N_13668,N_13634);
nand U16158 (N_16158,N_12564,N_14170);
and U16159 (N_16159,N_14436,N_14764);
xnor U16160 (N_16160,N_13588,N_14147);
or U16161 (N_16161,N_13820,N_14689);
xnor U16162 (N_16162,N_14691,N_14530);
or U16163 (N_16163,N_13513,N_12988);
xor U16164 (N_16164,N_14701,N_13791);
nand U16165 (N_16165,N_13188,N_14970);
or U16166 (N_16166,N_13850,N_14527);
xor U16167 (N_16167,N_13661,N_12740);
nor U16168 (N_16168,N_13410,N_12519);
and U16169 (N_16169,N_12906,N_13495);
nor U16170 (N_16170,N_13090,N_14463);
xor U16171 (N_16171,N_13148,N_12668);
nor U16172 (N_16172,N_14535,N_13881);
xnor U16173 (N_16173,N_12971,N_14094);
or U16174 (N_16174,N_13908,N_12918);
and U16175 (N_16175,N_14000,N_12907);
nand U16176 (N_16176,N_12533,N_14088);
nor U16177 (N_16177,N_13578,N_14435);
xor U16178 (N_16178,N_14989,N_12663);
or U16179 (N_16179,N_13454,N_12699);
xnor U16180 (N_16180,N_13809,N_12633);
nand U16181 (N_16181,N_12726,N_13029);
and U16182 (N_16182,N_14465,N_13266);
xor U16183 (N_16183,N_13253,N_13984);
and U16184 (N_16184,N_13234,N_12923);
nand U16185 (N_16185,N_12781,N_13102);
xnor U16186 (N_16186,N_14490,N_14112);
and U16187 (N_16187,N_14291,N_13957);
and U16188 (N_16188,N_14581,N_14324);
or U16189 (N_16189,N_14939,N_14922);
and U16190 (N_16190,N_13364,N_13209);
nand U16191 (N_16191,N_12549,N_12741);
nand U16192 (N_16192,N_13852,N_14529);
nor U16193 (N_16193,N_12925,N_12917);
and U16194 (N_16194,N_14756,N_14329);
or U16195 (N_16195,N_12697,N_13027);
nand U16196 (N_16196,N_13459,N_14773);
and U16197 (N_16197,N_14679,N_14603);
xnor U16198 (N_16198,N_13448,N_14555);
nor U16199 (N_16199,N_13856,N_13158);
nor U16200 (N_16200,N_13716,N_14259);
nor U16201 (N_16201,N_14511,N_14891);
nand U16202 (N_16202,N_13073,N_14600);
nand U16203 (N_16203,N_14654,N_13729);
nor U16204 (N_16204,N_12554,N_13877);
xnor U16205 (N_16205,N_13169,N_14517);
and U16206 (N_16206,N_12901,N_14961);
nor U16207 (N_16207,N_14966,N_12660);
xor U16208 (N_16208,N_14306,N_13548);
nor U16209 (N_16209,N_13603,N_14242);
and U16210 (N_16210,N_14341,N_12723);
and U16211 (N_16211,N_13096,N_13750);
and U16212 (N_16212,N_13310,N_13804);
or U16213 (N_16213,N_12534,N_13833);
xor U16214 (N_16214,N_12959,N_12583);
xnor U16215 (N_16215,N_13147,N_14321);
or U16216 (N_16216,N_14836,N_14718);
xor U16217 (N_16217,N_14590,N_14216);
and U16218 (N_16218,N_13081,N_12749);
xnor U16219 (N_16219,N_14230,N_14474);
nor U16220 (N_16220,N_14264,N_12642);
or U16221 (N_16221,N_13490,N_12789);
or U16222 (N_16222,N_14203,N_14846);
nor U16223 (N_16223,N_13321,N_14862);
or U16224 (N_16224,N_13337,N_13837);
and U16225 (N_16225,N_14389,N_12556);
or U16226 (N_16226,N_13296,N_12852);
and U16227 (N_16227,N_14481,N_14670);
nand U16228 (N_16228,N_14117,N_14185);
nand U16229 (N_16229,N_13001,N_14161);
nor U16230 (N_16230,N_14797,N_13753);
and U16231 (N_16231,N_14379,N_12555);
or U16232 (N_16232,N_13524,N_12909);
and U16233 (N_16233,N_14560,N_12829);
or U16234 (N_16234,N_14975,N_13999);
and U16235 (N_16235,N_13713,N_12888);
nor U16236 (N_16236,N_12905,N_14051);
nor U16237 (N_16237,N_14146,N_14303);
nor U16238 (N_16238,N_14980,N_13589);
or U16239 (N_16239,N_14227,N_13409);
or U16240 (N_16240,N_13117,N_13136);
xor U16241 (N_16241,N_13423,N_12593);
nor U16242 (N_16242,N_12648,N_13835);
or U16243 (N_16243,N_14045,N_13692);
or U16244 (N_16244,N_14643,N_14053);
or U16245 (N_16245,N_14374,N_13082);
and U16246 (N_16246,N_14907,N_14139);
and U16247 (N_16247,N_12515,N_14235);
or U16248 (N_16248,N_12854,N_14685);
nor U16249 (N_16249,N_14720,N_12910);
or U16250 (N_16250,N_14701,N_13159);
and U16251 (N_16251,N_14260,N_13645);
and U16252 (N_16252,N_14188,N_14441);
and U16253 (N_16253,N_13528,N_14032);
xnor U16254 (N_16254,N_14481,N_12590);
nand U16255 (N_16255,N_14836,N_13885);
xor U16256 (N_16256,N_13342,N_12631);
nor U16257 (N_16257,N_14463,N_14060);
or U16258 (N_16258,N_13933,N_14778);
nand U16259 (N_16259,N_13981,N_14164);
or U16260 (N_16260,N_12513,N_12803);
or U16261 (N_16261,N_13268,N_12553);
and U16262 (N_16262,N_13957,N_14340);
nand U16263 (N_16263,N_12653,N_13434);
xnor U16264 (N_16264,N_14587,N_13579);
and U16265 (N_16265,N_13184,N_14561);
nor U16266 (N_16266,N_14805,N_13962);
and U16267 (N_16267,N_13922,N_12567);
xnor U16268 (N_16268,N_14057,N_13628);
nand U16269 (N_16269,N_13807,N_13437);
nor U16270 (N_16270,N_13428,N_14545);
or U16271 (N_16271,N_13626,N_13894);
and U16272 (N_16272,N_13493,N_13115);
or U16273 (N_16273,N_13300,N_12534);
nand U16274 (N_16274,N_13924,N_12854);
or U16275 (N_16275,N_12789,N_13590);
or U16276 (N_16276,N_13362,N_13621);
xnor U16277 (N_16277,N_13080,N_13345);
nor U16278 (N_16278,N_14459,N_14991);
xnor U16279 (N_16279,N_12669,N_13151);
and U16280 (N_16280,N_14136,N_13518);
nand U16281 (N_16281,N_14554,N_13716);
or U16282 (N_16282,N_14879,N_14946);
xnor U16283 (N_16283,N_14161,N_13808);
or U16284 (N_16284,N_14644,N_13185);
xor U16285 (N_16285,N_14023,N_13975);
nand U16286 (N_16286,N_14435,N_14885);
or U16287 (N_16287,N_12645,N_14417);
and U16288 (N_16288,N_14103,N_13671);
nand U16289 (N_16289,N_13694,N_13890);
or U16290 (N_16290,N_13367,N_14597);
nor U16291 (N_16291,N_13232,N_12729);
nand U16292 (N_16292,N_14773,N_13876);
and U16293 (N_16293,N_13800,N_13962);
nand U16294 (N_16294,N_13188,N_13379);
nor U16295 (N_16295,N_13592,N_13337);
nand U16296 (N_16296,N_14606,N_12843);
or U16297 (N_16297,N_12568,N_14384);
and U16298 (N_16298,N_14192,N_14357);
nand U16299 (N_16299,N_13552,N_13661);
or U16300 (N_16300,N_13960,N_12798);
nand U16301 (N_16301,N_12900,N_13411);
and U16302 (N_16302,N_12699,N_14460);
and U16303 (N_16303,N_12671,N_12814);
and U16304 (N_16304,N_14715,N_14499);
xor U16305 (N_16305,N_13732,N_14169);
nand U16306 (N_16306,N_14431,N_13263);
and U16307 (N_16307,N_13487,N_13283);
or U16308 (N_16308,N_14614,N_13434);
nor U16309 (N_16309,N_13470,N_12895);
nor U16310 (N_16310,N_14992,N_14041);
xnor U16311 (N_16311,N_13528,N_13924);
or U16312 (N_16312,N_13991,N_14742);
nor U16313 (N_16313,N_13432,N_12811);
nor U16314 (N_16314,N_14843,N_14851);
nor U16315 (N_16315,N_14203,N_14599);
nand U16316 (N_16316,N_13010,N_13057);
or U16317 (N_16317,N_14873,N_14348);
xnor U16318 (N_16318,N_12765,N_13297);
nand U16319 (N_16319,N_14759,N_12983);
xnor U16320 (N_16320,N_14174,N_13315);
nor U16321 (N_16321,N_13997,N_13976);
and U16322 (N_16322,N_14377,N_12513);
or U16323 (N_16323,N_13234,N_13959);
or U16324 (N_16324,N_14769,N_14982);
or U16325 (N_16325,N_14338,N_13171);
nor U16326 (N_16326,N_12588,N_13171);
nand U16327 (N_16327,N_13125,N_13059);
and U16328 (N_16328,N_13701,N_14941);
or U16329 (N_16329,N_14675,N_14972);
nand U16330 (N_16330,N_14927,N_14479);
nand U16331 (N_16331,N_14012,N_14123);
nor U16332 (N_16332,N_14573,N_13222);
nor U16333 (N_16333,N_13050,N_14794);
xor U16334 (N_16334,N_14777,N_14976);
and U16335 (N_16335,N_14857,N_13974);
or U16336 (N_16336,N_14198,N_13651);
xnor U16337 (N_16337,N_13880,N_14496);
nand U16338 (N_16338,N_14080,N_13331);
and U16339 (N_16339,N_12699,N_14747);
or U16340 (N_16340,N_14415,N_14600);
or U16341 (N_16341,N_13110,N_14846);
or U16342 (N_16342,N_12924,N_14473);
xnor U16343 (N_16343,N_14885,N_14991);
or U16344 (N_16344,N_13200,N_12898);
and U16345 (N_16345,N_13568,N_12516);
or U16346 (N_16346,N_12912,N_13375);
nor U16347 (N_16347,N_12733,N_12864);
or U16348 (N_16348,N_14768,N_13046);
and U16349 (N_16349,N_14219,N_12933);
nor U16350 (N_16350,N_12828,N_13258);
xnor U16351 (N_16351,N_12632,N_13891);
or U16352 (N_16352,N_14250,N_12917);
nand U16353 (N_16353,N_13220,N_14359);
and U16354 (N_16354,N_12977,N_14684);
and U16355 (N_16355,N_12996,N_14770);
nand U16356 (N_16356,N_14136,N_14973);
or U16357 (N_16357,N_14347,N_13108);
xnor U16358 (N_16358,N_14284,N_12602);
and U16359 (N_16359,N_14328,N_13738);
nor U16360 (N_16360,N_13783,N_14613);
and U16361 (N_16361,N_13267,N_13541);
xor U16362 (N_16362,N_13168,N_12521);
nor U16363 (N_16363,N_14469,N_14512);
or U16364 (N_16364,N_13227,N_13143);
or U16365 (N_16365,N_12619,N_14294);
and U16366 (N_16366,N_13527,N_13012);
or U16367 (N_16367,N_13733,N_14371);
nor U16368 (N_16368,N_12632,N_13546);
nor U16369 (N_16369,N_14941,N_13638);
xor U16370 (N_16370,N_14809,N_13505);
xnor U16371 (N_16371,N_14582,N_12809);
xnor U16372 (N_16372,N_14216,N_12953);
and U16373 (N_16373,N_14015,N_12813);
nand U16374 (N_16374,N_13256,N_13527);
xor U16375 (N_16375,N_13433,N_13594);
nor U16376 (N_16376,N_14121,N_13928);
or U16377 (N_16377,N_13046,N_12713);
or U16378 (N_16378,N_12518,N_13190);
xnor U16379 (N_16379,N_12837,N_12980);
nor U16380 (N_16380,N_13849,N_13367);
nand U16381 (N_16381,N_13063,N_12936);
nand U16382 (N_16382,N_13810,N_13382);
nand U16383 (N_16383,N_12976,N_12778);
nand U16384 (N_16384,N_12730,N_13806);
nand U16385 (N_16385,N_14385,N_12791);
nor U16386 (N_16386,N_14472,N_14186);
nor U16387 (N_16387,N_14091,N_14078);
nand U16388 (N_16388,N_14336,N_14051);
and U16389 (N_16389,N_13652,N_13825);
nand U16390 (N_16390,N_14588,N_13803);
xor U16391 (N_16391,N_13493,N_13453);
or U16392 (N_16392,N_14765,N_14980);
nor U16393 (N_16393,N_13582,N_14757);
and U16394 (N_16394,N_13422,N_12578);
nand U16395 (N_16395,N_14884,N_13846);
nor U16396 (N_16396,N_12946,N_13620);
xor U16397 (N_16397,N_14139,N_14049);
nand U16398 (N_16398,N_14481,N_14824);
and U16399 (N_16399,N_12539,N_13361);
xor U16400 (N_16400,N_14582,N_13637);
nand U16401 (N_16401,N_12726,N_13357);
or U16402 (N_16402,N_13641,N_14914);
xor U16403 (N_16403,N_12868,N_14241);
xor U16404 (N_16404,N_14611,N_13033);
xor U16405 (N_16405,N_12522,N_14053);
xnor U16406 (N_16406,N_13203,N_12621);
nor U16407 (N_16407,N_14750,N_14357);
and U16408 (N_16408,N_12620,N_13200);
xnor U16409 (N_16409,N_14825,N_13000);
nor U16410 (N_16410,N_13959,N_13016);
nor U16411 (N_16411,N_14181,N_13504);
and U16412 (N_16412,N_13150,N_13693);
or U16413 (N_16413,N_13947,N_14982);
or U16414 (N_16414,N_14643,N_13805);
and U16415 (N_16415,N_12548,N_12878);
nand U16416 (N_16416,N_13668,N_14609);
nand U16417 (N_16417,N_14012,N_13126);
nor U16418 (N_16418,N_13935,N_14615);
and U16419 (N_16419,N_13253,N_13890);
nor U16420 (N_16420,N_12546,N_13100);
nor U16421 (N_16421,N_13443,N_13177);
nand U16422 (N_16422,N_14479,N_12933);
or U16423 (N_16423,N_13967,N_12777);
or U16424 (N_16424,N_14294,N_14850);
nor U16425 (N_16425,N_13087,N_14249);
and U16426 (N_16426,N_12896,N_14802);
xor U16427 (N_16427,N_14362,N_13875);
nor U16428 (N_16428,N_14925,N_12647);
nand U16429 (N_16429,N_13088,N_13412);
and U16430 (N_16430,N_12637,N_13727);
nand U16431 (N_16431,N_14742,N_12758);
nand U16432 (N_16432,N_14903,N_14473);
nand U16433 (N_16433,N_14001,N_14245);
and U16434 (N_16434,N_14593,N_12536);
xnor U16435 (N_16435,N_14828,N_12906);
xnor U16436 (N_16436,N_14889,N_14769);
and U16437 (N_16437,N_14341,N_13824);
xor U16438 (N_16438,N_13098,N_14573);
or U16439 (N_16439,N_14047,N_13938);
or U16440 (N_16440,N_12717,N_14146);
nor U16441 (N_16441,N_14335,N_12888);
and U16442 (N_16442,N_14727,N_13655);
and U16443 (N_16443,N_12730,N_13542);
nor U16444 (N_16444,N_13464,N_14624);
nand U16445 (N_16445,N_12608,N_14280);
and U16446 (N_16446,N_12906,N_13415);
or U16447 (N_16447,N_14562,N_13990);
nand U16448 (N_16448,N_14690,N_14857);
nand U16449 (N_16449,N_13430,N_14630);
nor U16450 (N_16450,N_14497,N_14649);
nor U16451 (N_16451,N_14491,N_13147);
or U16452 (N_16452,N_13727,N_13421);
or U16453 (N_16453,N_12916,N_13687);
and U16454 (N_16454,N_14213,N_14927);
or U16455 (N_16455,N_12782,N_14743);
xnor U16456 (N_16456,N_14352,N_13652);
and U16457 (N_16457,N_14300,N_13555);
nor U16458 (N_16458,N_13313,N_13497);
nor U16459 (N_16459,N_13352,N_13330);
or U16460 (N_16460,N_12971,N_13701);
nor U16461 (N_16461,N_14531,N_13291);
nand U16462 (N_16462,N_13013,N_13339);
nor U16463 (N_16463,N_14479,N_14960);
and U16464 (N_16464,N_12682,N_14003);
or U16465 (N_16465,N_12555,N_14817);
nor U16466 (N_16466,N_13130,N_12970);
nor U16467 (N_16467,N_13728,N_14954);
xnor U16468 (N_16468,N_13001,N_14147);
xnor U16469 (N_16469,N_14438,N_12510);
nor U16470 (N_16470,N_13470,N_13562);
and U16471 (N_16471,N_13766,N_13346);
or U16472 (N_16472,N_14463,N_13961);
or U16473 (N_16473,N_13196,N_13929);
or U16474 (N_16474,N_14322,N_13189);
nand U16475 (N_16475,N_14295,N_14033);
xnor U16476 (N_16476,N_14155,N_13622);
nor U16477 (N_16477,N_13384,N_13414);
nor U16478 (N_16478,N_12724,N_13056);
or U16479 (N_16479,N_13989,N_13951);
nor U16480 (N_16480,N_14439,N_13481);
nor U16481 (N_16481,N_14313,N_14561);
and U16482 (N_16482,N_13420,N_13047);
nor U16483 (N_16483,N_13331,N_14581);
and U16484 (N_16484,N_13111,N_13508);
and U16485 (N_16485,N_14700,N_14937);
or U16486 (N_16486,N_14570,N_13378);
xnor U16487 (N_16487,N_14665,N_12597);
nor U16488 (N_16488,N_13945,N_12950);
xnor U16489 (N_16489,N_13370,N_14161);
nor U16490 (N_16490,N_14817,N_13758);
xor U16491 (N_16491,N_14288,N_12923);
nand U16492 (N_16492,N_13488,N_14040);
nor U16493 (N_16493,N_14829,N_13855);
xor U16494 (N_16494,N_12783,N_12533);
and U16495 (N_16495,N_13756,N_13878);
nor U16496 (N_16496,N_13962,N_13451);
nor U16497 (N_16497,N_13076,N_13557);
or U16498 (N_16498,N_13629,N_12830);
or U16499 (N_16499,N_14807,N_14571);
xor U16500 (N_16500,N_13257,N_14252);
and U16501 (N_16501,N_14420,N_14509);
nor U16502 (N_16502,N_12675,N_13543);
nand U16503 (N_16503,N_14325,N_14917);
or U16504 (N_16504,N_13826,N_12785);
nor U16505 (N_16505,N_13078,N_13721);
xnor U16506 (N_16506,N_14735,N_14213);
or U16507 (N_16507,N_13865,N_13182);
nor U16508 (N_16508,N_14710,N_12685);
nand U16509 (N_16509,N_14289,N_14703);
or U16510 (N_16510,N_12602,N_13623);
nand U16511 (N_16511,N_14134,N_13650);
or U16512 (N_16512,N_14401,N_13713);
nor U16513 (N_16513,N_14489,N_12966);
or U16514 (N_16514,N_13806,N_14541);
nor U16515 (N_16515,N_14381,N_14292);
nand U16516 (N_16516,N_14799,N_14540);
and U16517 (N_16517,N_14719,N_14005);
and U16518 (N_16518,N_14808,N_13801);
and U16519 (N_16519,N_14522,N_14417);
or U16520 (N_16520,N_12556,N_12889);
xnor U16521 (N_16521,N_13718,N_14340);
xor U16522 (N_16522,N_12758,N_12582);
nor U16523 (N_16523,N_12602,N_14020);
xor U16524 (N_16524,N_12984,N_14255);
nand U16525 (N_16525,N_12876,N_14087);
xor U16526 (N_16526,N_13819,N_13144);
nor U16527 (N_16527,N_12711,N_13355);
nand U16528 (N_16528,N_12826,N_14487);
or U16529 (N_16529,N_13530,N_12722);
or U16530 (N_16530,N_14683,N_14922);
or U16531 (N_16531,N_14598,N_13222);
xor U16532 (N_16532,N_13122,N_13740);
nand U16533 (N_16533,N_14684,N_14434);
or U16534 (N_16534,N_14935,N_13594);
nand U16535 (N_16535,N_13830,N_12823);
nand U16536 (N_16536,N_14303,N_14908);
xor U16537 (N_16537,N_14951,N_12603);
or U16538 (N_16538,N_14830,N_13130);
xnor U16539 (N_16539,N_13019,N_12546);
and U16540 (N_16540,N_12809,N_13214);
xnor U16541 (N_16541,N_13883,N_14604);
or U16542 (N_16542,N_13894,N_13663);
or U16543 (N_16543,N_14110,N_14653);
nand U16544 (N_16544,N_14402,N_14712);
and U16545 (N_16545,N_14213,N_14083);
nor U16546 (N_16546,N_14094,N_12941);
and U16547 (N_16547,N_13627,N_14958);
nor U16548 (N_16548,N_14312,N_13288);
nor U16549 (N_16549,N_13545,N_13453);
xor U16550 (N_16550,N_13619,N_12767);
nand U16551 (N_16551,N_13925,N_14808);
and U16552 (N_16552,N_14681,N_13176);
and U16553 (N_16553,N_13521,N_14686);
nor U16554 (N_16554,N_14717,N_12811);
xnor U16555 (N_16555,N_12784,N_13926);
nor U16556 (N_16556,N_13812,N_14461);
nand U16557 (N_16557,N_14369,N_13916);
nand U16558 (N_16558,N_13431,N_12713);
and U16559 (N_16559,N_14669,N_14498);
nand U16560 (N_16560,N_13583,N_13795);
or U16561 (N_16561,N_13811,N_14035);
xnor U16562 (N_16562,N_13043,N_14536);
nand U16563 (N_16563,N_14938,N_14805);
nor U16564 (N_16564,N_13608,N_12679);
nand U16565 (N_16565,N_14233,N_14861);
or U16566 (N_16566,N_14232,N_13881);
nor U16567 (N_16567,N_14306,N_14529);
nor U16568 (N_16568,N_13557,N_13487);
xnor U16569 (N_16569,N_12629,N_13000);
nand U16570 (N_16570,N_14086,N_13522);
nor U16571 (N_16571,N_13654,N_13966);
xor U16572 (N_16572,N_14613,N_12718);
and U16573 (N_16573,N_14979,N_14316);
and U16574 (N_16574,N_14287,N_12581);
nand U16575 (N_16575,N_14498,N_14558);
xnor U16576 (N_16576,N_13066,N_12527);
and U16577 (N_16577,N_13570,N_14123);
nand U16578 (N_16578,N_14101,N_13814);
and U16579 (N_16579,N_13703,N_14750);
nor U16580 (N_16580,N_14519,N_12568);
or U16581 (N_16581,N_12980,N_14317);
and U16582 (N_16582,N_14013,N_14121);
nand U16583 (N_16583,N_13036,N_14231);
or U16584 (N_16584,N_14494,N_13828);
nor U16585 (N_16585,N_13292,N_13831);
xnor U16586 (N_16586,N_13088,N_12556);
nand U16587 (N_16587,N_13651,N_13552);
nand U16588 (N_16588,N_14043,N_14640);
and U16589 (N_16589,N_12665,N_14008);
nor U16590 (N_16590,N_13885,N_14496);
xnor U16591 (N_16591,N_14286,N_12633);
xnor U16592 (N_16592,N_14933,N_14878);
nor U16593 (N_16593,N_14705,N_13914);
nand U16594 (N_16594,N_14205,N_12800);
nand U16595 (N_16595,N_14619,N_12838);
and U16596 (N_16596,N_13060,N_13632);
nand U16597 (N_16597,N_14413,N_14874);
and U16598 (N_16598,N_12527,N_13228);
nand U16599 (N_16599,N_14438,N_14427);
and U16600 (N_16600,N_13322,N_14342);
and U16601 (N_16601,N_12922,N_12695);
or U16602 (N_16602,N_14713,N_13179);
and U16603 (N_16603,N_14011,N_12938);
xor U16604 (N_16604,N_12832,N_14581);
nor U16605 (N_16605,N_14539,N_13550);
xnor U16606 (N_16606,N_14212,N_14345);
and U16607 (N_16607,N_14972,N_12750);
nand U16608 (N_16608,N_14605,N_14141);
and U16609 (N_16609,N_13726,N_14875);
or U16610 (N_16610,N_13674,N_12673);
nor U16611 (N_16611,N_12566,N_13437);
xnor U16612 (N_16612,N_13232,N_13271);
xnor U16613 (N_16613,N_14781,N_13891);
xor U16614 (N_16614,N_14855,N_14247);
nand U16615 (N_16615,N_13447,N_13418);
and U16616 (N_16616,N_12638,N_13722);
nand U16617 (N_16617,N_14892,N_14881);
and U16618 (N_16618,N_14052,N_14354);
nand U16619 (N_16619,N_14481,N_14215);
or U16620 (N_16620,N_13274,N_14637);
nor U16621 (N_16621,N_13159,N_12948);
nand U16622 (N_16622,N_13942,N_12724);
xor U16623 (N_16623,N_13642,N_14826);
xnor U16624 (N_16624,N_13935,N_12993);
xor U16625 (N_16625,N_14701,N_14304);
xnor U16626 (N_16626,N_12667,N_14153);
and U16627 (N_16627,N_14434,N_14537);
nand U16628 (N_16628,N_14949,N_14961);
or U16629 (N_16629,N_13904,N_14956);
and U16630 (N_16630,N_13114,N_13660);
and U16631 (N_16631,N_12958,N_12857);
and U16632 (N_16632,N_13803,N_13751);
nor U16633 (N_16633,N_14735,N_14210);
or U16634 (N_16634,N_13957,N_13094);
and U16635 (N_16635,N_13738,N_12742);
and U16636 (N_16636,N_12777,N_14467);
xnor U16637 (N_16637,N_14317,N_12745);
nand U16638 (N_16638,N_14645,N_12847);
nor U16639 (N_16639,N_13743,N_14405);
and U16640 (N_16640,N_14497,N_13531);
xor U16641 (N_16641,N_13940,N_14990);
nor U16642 (N_16642,N_13654,N_14230);
or U16643 (N_16643,N_12612,N_12787);
nand U16644 (N_16644,N_13854,N_13456);
nand U16645 (N_16645,N_14228,N_12791);
nand U16646 (N_16646,N_12712,N_13369);
xnor U16647 (N_16647,N_13288,N_13289);
nand U16648 (N_16648,N_13750,N_13220);
or U16649 (N_16649,N_14323,N_12927);
and U16650 (N_16650,N_14618,N_13998);
nand U16651 (N_16651,N_14933,N_13895);
nor U16652 (N_16652,N_13094,N_13588);
or U16653 (N_16653,N_14287,N_12684);
nand U16654 (N_16654,N_13309,N_14080);
and U16655 (N_16655,N_14192,N_12828);
xnor U16656 (N_16656,N_13137,N_12604);
nand U16657 (N_16657,N_14096,N_12582);
nand U16658 (N_16658,N_13549,N_13603);
xor U16659 (N_16659,N_13892,N_13318);
xor U16660 (N_16660,N_12823,N_13017);
xnor U16661 (N_16661,N_13371,N_14785);
nor U16662 (N_16662,N_14554,N_12828);
or U16663 (N_16663,N_13532,N_13297);
or U16664 (N_16664,N_12678,N_14618);
or U16665 (N_16665,N_14727,N_14185);
and U16666 (N_16666,N_13780,N_12901);
and U16667 (N_16667,N_12710,N_13441);
xnor U16668 (N_16668,N_14258,N_14751);
or U16669 (N_16669,N_14609,N_13895);
nand U16670 (N_16670,N_14568,N_14538);
xor U16671 (N_16671,N_13631,N_13141);
nor U16672 (N_16672,N_14363,N_13638);
and U16673 (N_16673,N_12547,N_13579);
nand U16674 (N_16674,N_13766,N_14292);
xor U16675 (N_16675,N_13210,N_13381);
and U16676 (N_16676,N_14869,N_13433);
nand U16677 (N_16677,N_13449,N_14365);
nor U16678 (N_16678,N_13556,N_13925);
nand U16679 (N_16679,N_13011,N_14415);
nor U16680 (N_16680,N_14515,N_12958);
xor U16681 (N_16681,N_13766,N_14188);
nand U16682 (N_16682,N_14659,N_13038);
nor U16683 (N_16683,N_12561,N_14656);
nor U16684 (N_16684,N_14500,N_13369);
nor U16685 (N_16685,N_14002,N_13023);
nor U16686 (N_16686,N_14660,N_13535);
and U16687 (N_16687,N_14620,N_13308);
or U16688 (N_16688,N_12517,N_13430);
and U16689 (N_16689,N_13557,N_14396);
or U16690 (N_16690,N_12526,N_14229);
nor U16691 (N_16691,N_14726,N_13830);
nand U16692 (N_16692,N_14018,N_13038);
nand U16693 (N_16693,N_13101,N_14904);
nand U16694 (N_16694,N_12761,N_12784);
nand U16695 (N_16695,N_14524,N_13625);
or U16696 (N_16696,N_14144,N_13849);
and U16697 (N_16697,N_14522,N_13428);
xnor U16698 (N_16698,N_14484,N_13149);
or U16699 (N_16699,N_12940,N_14672);
xnor U16700 (N_16700,N_13266,N_13429);
or U16701 (N_16701,N_14593,N_13459);
and U16702 (N_16702,N_13591,N_12711);
xnor U16703 (N_16703,N_13293,N_14022);
nor U16704 (N_16704,N_14898,N_14482);
or U16705 (N_16705,N_14820,N_14221);
and U16706 (N_16706,N_14004,N_13713);
and U16707 (N_16707,N_13648,N_13683);
xnor U16708 (N_16708,N_14248,N_14484);
nor U16709 (N_16709,N_13139,N_14060);
and U16710 (N_16710,N_13565,N_14770);
and U16711 (N_16711,N_12503,N_14856);
and U16712 (N_16712,N_14801,N_14592);
and U16713 (N_16713,N_13881,N_14565);
and U16714 (N_16714,N_13865,N_14866);
xor U16715 (N_16715,N_13334,N_13282);
and U16716 (N_16716,N_12700,N_14593);
xnor U16717 (N_16717,N_12719,N_14908);
and U16718 (N_16718,N_13366,N_14316);
nor U16719 (N_16719,N_13833,N_12657);
or U16720 (N_16720,N_14905,N_14812);
xor U16721 (N_16721,N_13772,N_13062);
nor U16722 (N_16722,N_13498,N_14774);
or U16723 (N_16723,N_12847,N_13307);
and U16724 (N_16724,N_14760,N_14081);
or U16725 (N_16725,N_13928,N_12921);
or U16726 (N_16726,N_12671,N_13958);
nand U16727 (N_16727,N_14348,N_13698);
xor U16728 (N_16728,N_13210,N_13833);
and U16729 (N_16729,N_12977,N_13148);
xor U16730 (N_16730,N_13875,N_14289);
or U16731 (N_16731,N_14740,N_13908);
or U16732 (N_16732,N_13223,N_13375);
nor U16733 (N_16733,N_14327,N_14774);
or U16734 (N_16734,N_13625,N_12658);
xor U16735 (N_16735,N_14492,N_12799);
nor U16736 (N_16736,N_13669,N_13158);
or U16737 (N_16737,N_14963,N_13416);
and U16738 (N_16738,N_14540,N_14042);
xor U16739 (N_16739,N_12801,N_12800);
and U16740 (N_16740,N_13715,N_12773);
and U16741 (N_16741,N_12870,N_13626);
nand U16742 (N_16742,N_13330,N_14535);
xnor U16743 (N_16743,N_13338,N_14675);
nand U16744 (N_16744,N_13525,N_14957);
and U16745 (N_16745,N_14508,N_13188);
nand U16746 (N_16746,N_14779,N_13093);
or U16747 (N_16747,N_14627,N_14200);
nor U16748 (N_16748,N_13502,N_14102);
and U16749 (N_16749,N_13605,N_13764);
or U16750 (N_16750,N_13282,N_14012);
nand U16751 (N_16751,N_12780,N_14801);
xor U16752 (N_16752,N_13615,N_14005);
and U16753 (N_16753,N_14919,N_12631);
and U16754 (N_16754,N_13107,N_14644);
or U16755 (N_16755,N_13265,N_14452);
nand U16756 (N_16756,N_13999,N_12665);
or U16757 (N_16757,N_13368,N_14488);
and U16758 (N_16758,N_13038,N_12609);
nand U16759 (N_16759,N_14493,N_14957);
and U16760 (N_16760,N_13706,N_13009);
or U16761 (N_16761,N_14782,N_14738);
xor U16762 (N_16762,N_14262,N_13664);
xnor U16763 (N_16763,N_14205,N_12824);
and U16764 (N_16764,N_13895,N_14210);
nand U16765 (N_16765,N_14887,N_13516);
or U16766 (N_16766,N_13180,N_14105);
xor U16767 (N_16767,N_14941,N_13242);
nor U16768 (N_16768,N_14232,N_12918);
xnor U16769 (N_16769,N_13493,N_12814);
nor U16770 (N_16770,N_14265,N_14848);
or U16771 (N_16771,N_12530,N_14651);
and U16772 (N_16772,N_13695,N_14891);
nand U16773 (N_16773,N_12693,N_13022);
nor U16774 (N_16774,N_12771,N_14378);
and U16775 (N_16775,N_14822,N_13675);
xnor U16776 (N_16776,N_13378,N_13561);
xor U16777 (N_16777,N_14713,N_13262);
nand U16778 (N_16778,N_14627,N_12537);
xnor U16779 (N_16779,N_14435,N_13627);
nand U16780 (N_16780,N_14815,N_13365);
nor U16781 (N_16781,N_14761,N_14261);
xnor U16782 (N_16782,N_14215,N_13496);
xor U16783 (N_16783,N_13757,N_14920);
or U16784 (N_16784,N_13350,N_14992);
nor U16785 (N_16785,N_14275,N_13205);
nand U16786 (N_16786,N_14021,N_13224);
nand U16787 (N_16787,N_13840,N_14251);
xor U16788 (N_16788,N_13201,N_12794);
xor U16789 (N_16789,N_14446,N_14695);
and U16790 (N_16790,N_12967,N_13743);
nand U16791 (N_16791,N_14669,N_13160);
and U16792 (N_16792,N_14950,N_13080);
and U16793 (N_16793,N_13848,N_13613);
nand U16794 (N_16794,N_14623,N_13598);
or U16795 (N_16795,N_13152,N_12580);
or U16796 (N_16796,N_12811,N_13003);
nor U16797 (N_16797,N_13305,N_13427);
nand U16798 (N_16798,N_13984,N_14259);
and U16799 (N_16799,N_14600,N_13323);
and U16800 (N_16800,N_12836,N_13087);
xor U16801 (N_16801,N_14715,N_12722);
nor U16802 (N_16802,N_13907,N_14365);
and U16803 (N_16803,N_14794,N_13211);
xnor U16804 (N_16804,N_12583,N_12946);
nor U16805 (N_16805,N_14770,N_12769);
nor U16806 (N_16806,N_12537,N_12684);
nand U16807 (N_16807,N_13551,N_13621);
nor U16808 (N_16808,N_14678,N_13367);
xor U16809 (N_16809,N_14263,N_13802);
and U16810 (N_16810,N_14049,N_12814);
nor U16811 (N_16811,N_13457,N_14000);
and U16812 (N_16812,N_12816,N_13845);
nand U16813 (N_16813,N_14645,N_13343);
or U16814 (N_16814,N_12609,N_13360);
nor U16815 (N_16815,N_13285,N_13829);
nor U16816 (N_16816,N_13040,N_12579);
or U16817 (N_16817,N_13307,N_12586);
or U16818 (N_16818,N_13904,N_13300);
nand U16819 (N_16819,N_13646,N_14304);
nand U16820 (N_16820,N_13503,N_14218);
and U16821 (N_16821,N_13198,N_13147);
xnor U16822 (N_16822,N_14316,N_14984);
nand U16823 (N_16823,N_12896,N_14062);
nor U16824 (N_16824,N_12855,N_14251);
and U16825 (N_16825,N_14192,N_13788);
and U16826 (N_16826,N_12733,N_14133);
nor U16827 (N_16827,N_12854,N_12676);
xor U16828 (N_16828,N_13245,N_14220);
xnor U16829 (N_16829,N_13194,N_13115);
nor U16830 (N_16830,N_13039,N_12618);
and U16831 (N_16831,N_14523,N_14733);
or U16832 (N_16832,N_14496,N_13586);
nand U16833 (N_16833,N_14342,N_12722);
xnor U16834 (N_16834,N_13152,N_12930);
or U16835 (N_16835,N_14555,N_13071);
nor U16836 (N_16836,N_14763,N_14264);
nand U16837 (N_16837,N_14362,N_14703);
nand U16838 (N_16838,N_14093,N_13517);
nor U16839 (N_16839,N_14787,N_12745);
nor U16840 (N_16840,N_14026,N_13731);
nand U16841 (N_16841,N_14965,N_13469);
and U16842 (N_16842,N_14327,N_14049);
xor U16843 (N_16843,N_14116,N_13289);
and U16844 (N_16844,N_13229,N_14226);
and U16845 (N_16845,N_13912,N_12994);
nand U16846 (N_16846,N_13706,N_13439);
or U16847 (N_16847,N_14406,N_13956);
or U16848 (N_16848,N_13824,N_14592);
nand U16849 (N_16849,N_12924,N_13945);
xnor U16850 (N_16850,N_12506,N_14284);
nor U16851 (N_16851,N_14562,N_14914);
nand U16852 (N_16852,N_13842,N_14493);
nor U16853 (N_16853,N_14465,N_14034);
and U16854 (N_16854,N_14686,N_12637);
and U16855 (N_16855,N_12856,N_14992);
nand U16856 (N_16856,N_13120,N_13100);
and U16857 (N_16857,N_13670,N_14234);
xnor U16858 (N_16858,N_13867,N_14226);
xor U16859 (N_16859,N_13517,N_14999);
xor U16860 (N_16860,N_13643,N_14871);
nor U16861 (N_16861,N_14081,N_13212);
nand U16862 (N_16862,N_13904,N_14382);
nand U16863 (N_16863,N_12680,N_13059);
and U16864 (N_16864,N_14452,N_13879);
xnor U16865 (N_16865,N_14376,N_12636);
or U16866 (N_16866,N_14934,N_13675);
nand U16867 (N_16867,N_14554,N_13537);
nor U16868 (N_16868,N_14002,N_14605);
nor U16869 (N_16869,N_13554,N_13275);
xor U16870 (N_16870,N_12543,N_12975);
and U16871 (N_16871,N_13585,N_14112);
and U16872 (N_16872,N_12607,N_12955);
xnor U16873 (N_16873,N_13025,N_13680);
nor U16874 (N_16874,N_12902,N_14981);
xor U16875 (N_16875,N_14797,N_14036);
nor U16876 (N_16876,N_14562,N_12839);
and U16877 (N_16877,N_14946,N_13761);
xor U16878 (N_16878,N_13244,N_14126);
nand U16879 (N_16879,N_13935,N_13788);
or U16880 (N_16880,N_14257,N_13603);
or U16881 (N_16881,N_14142,N_13320);
xnor U16882 (N_16882,N_14459,N_14410);
and U16883 (N_16883,N_14902,N_12521);
or U16884 (N_16884,N_13025,N_13348);
nor U16885 (N_16885,N_14203,N_12550);
xor U16886 (N_16886,N_14120,N_13295);
or U16887 (N_16887,N_13979,N_13776);
xnor U16888 (N_16888,N_13438,N_13732);
nand U16889 (N_16889,N_12647,N_12908);
and U16890 (N_16890,N_13606,N_13234);
nand U16891 (N_16891,N_13465,N_13193);
and U16892 (N_16892,N_13024,N_13464);
or U16893 (N_16893,N_13038,N_14501);
xor U16894 (N_16894,N_13804,N_13726);
nand U16895 (N_16895,N_13633,N_12622);
or U16896 (N_16896,N_13361,N_13379);
xor U16897 (N_16897,N_13175,N_13521);
and U16898 (N_16898,N_14885,N_14465);
xnor U16899 (N_16899,N_13764,N_13772);
nand U16900 (N_16900,N_14896,N_13050);
nand U16901 (N_16901,N_13688,N_14893);
and U16902 (N_16902,N_12655,N_14479);
and U16903 (N_16903,N_12565,N_13303);
xnor U16904 (N_16904,N_13013,N_12557);
or U16905 (N_16905,N_12793,N_14529);
or U16906 (N_16906,N_13511,N_13774);
nand U16907 (N_16907,N_13854,N_14984);
nor U16908 (N_16908,N_13186,N_13710);
nor U16909 (N_16909,N_14316,N_14768);
xnor U16910 (N_16910,N_14124,N_14290);
nand U16911 (N_16911,N_14331,N_12724);
or U16912 (N_16912,N_13070,N_13908);
xor U16913 (N_16913,N_12786,N_13326);
xor U16914 (N_16914,N_12983,N_13678);
xnor U16915 (N_16915,N_14014,N_13121);
nand U16916 (N_16916,N_12644,N_14338);
nor U16917 (N_16917,N_12731,N_12630);
xor U16918 (N_16918,N_14788,N_13632);
xnor U16919 (N_16919,N_13065,N_13775);
and U16920 (N_16920,N_13594,N_13291);
nand U16921 (N_16921,N_14656,N_13467);
nor U16922 (N_16922,N_13048,N_12523);
and U16923 (N_16923,N_12792,N_13944);
nand U16924 (N_16924,N_14023,N_14254);
or U16925 (N_16925,N_12927,N_12621);
nand U16926 (N_16926,N_12815,N_14014);
nor U16927 (N_16927,N_14961,N_13477);
xnor U16928 (N_16928,N_13876,N_14774);
xnor U16929 (N_16929,N_12843,N_13417);
or U16930 (N_16930,N_13694,N_14121);
or U16931 (N_16931,N_12998,N_13436);
xor U16932 (N_16932,N_13970,N_12948);
nor U16933 (N_16933,N_13194,N_14197);
or U16934 (N_16934,N_13807,N_14850);
and U16935 (N_16935,N_13840,N_14390);
nor U16936 (N_16936,N_13511,N_14289);
nand U16937 (N_16937,N_13323,N_13515);
nor U16938 (N_16938,N_12688,N_14851);
nand U16939 (N_16939,N_12694,N_14715);
nand U16940 (N_16940,N_12640,N_13748);
or U16941 (N_16941,N_13259,N_13332);
xnor U16942 (N_16942,N_13498,N_12819);
xor U16943 (N_16943,N_14531,N_13906);
nor U16944 (N_16944,N_13510,N_13260);
nor U16945 (N_16945,N_14565,N_14461);
nand U16946 (N_16946,N_13046,N_12642);
nand U16947 (N_16947,N_12833,N_13019);
xor U16948 (N_16948,N_13534,N_14076);
or U16949 (N_16949,N_14100,N_12982);
xnor U16950 (N_16950,N_14090,N_13594);
xor U16951 (N_16951,N_14546,N_12842);
or U16952 (N_16952,N_14620,N_12738);
xnor U16953 (N_16953,N_14557,N_12959);
xnor U16954 (N_16954,N_13421,N_14170);
nor U16955 (N_16955,N_14645,N_13705);
xor U16956 (N_16956,N_14822,N_12543);
nand U16957 (N_16957,N_14048,N_13440);
xnor U16958 (N_16958,N_13841,N_13787);
nand U16959 (N_16959,N_13255,N_12533);
and U16960 (N_16960,N_14336,N_12539);
nor U16961 (N_16961,N_12839,N_13412);
nor U16962 (N_16962,N_13670,N_14641);
and U16963 (N_16963,N_13335,N_14924);
xor U16964 (N_16964,N_12672,N_13771);
or U16965 (N_16965,N_13820,N_12619);
or U16966 (N_16966,N_13531,N_14054);
xnor U16967 (N_16967,N_13832,N_14511);
or U16968 (N_16968,N_13614,N_13727);
xor U16969 (N_16969,N_12808,N_13548);
xor U16970 (N_16970,N_12801,N_14715);
or U16971 (N_16971,N_13575,N_14631);
nor U16972 (N_16972,N_13058,N_14990);
or U16973 (N_16973,N_13702,N_14382);
nand U16974 (N_16974,N_14503,N_13857);
or U16975 (N_16975,N_13639,N_12938);
nor U16976 (N_16976,N_12503,N_13308);
nor U16977 (N_16977,N_12741,N_14139);
nand U16978 (N_16978,N_13645,N_14031);
nand U16979 (N_16979,N_14694,N_14493);
and U16980 (N_16980,N_12993,N_12645);
xor U16981 (N_16981,N_12868,N_13733);
xnor U16982 (N_16982,N_12639,N_12599);
nor U16983 (N_16983,N_14673,N_13455);
nand U16984 (N_16984,N_13319,N_13990);
or U16985 (N_16985,N_13528,N_13300);
and U16986 (N_16986,N_12873,N_14566);
xor U16987 (N_16987,N_12591,N_13411);
nand U16988 (N_16988,N_13069,N_13530);
or U16989 (N_16989,N_14516,N_13996);
nor U16990 (N_16990,N_13604,N_14809);
xor U16991 (N_16991,N_14120,N_13175);
xnor U16992 (N_16992,N_13355,N_13460);
xnor U16993 (N_16993,N_14020,N_12782);
or U16994 (N_16994,N_12802,N_12998);
and U16995 (N_16995,N_13373,N_12698);
and U16996 (N_16996,N_14558,N_14878);
xnor U16997 (N_16997,N_14463,N_14841);
nand U16998 (N_16998,N_13702,N_12753);
nand U16999 (N_16999,N_14761,N_14983);
or U17000 (N_17000,N_13646,N_12850);
and U17001 (N_17001,N_13669,N_14955);
nor U17002 (N_17002,N_14188,N_14766);
and U17003 (N_17003,N_12833,N_14857);
or U17004 (N_17004,N_14773,N_14076);
and U17005 (N_17005,N_12772,N_12650);
and U17006 (N_17006,N_13918,N_14805);
or U17007 (N_17007,N_12959,N_14835);
nand U17008 (N_17008,N_12783,N_14365);
and U17009 (N_17009,N_13149,N_13824);
and U17010 (N_17010,N_14182,N_13273);
nand U17011 (N_17011,N_14636,N_13429);
xnor U17012 (N_17012,N_14944,N_13855);
or U17013 (N_17013,N_14947,N_12871);
and U17014 (N_17014,N_13301,N_14973);
and U17015 (N_17015,N_14764,N_13375);
nand U17016 (N_17016,N_12661,N_13391);
and U17017 (N_17017,N_13946,N_14010);
xnor U17018 (N_17018,N_13280,N_13126);
or U17019 (N_17019,N_13449,N_12663);
nand U17020 (N_17020,N_13905,N_13275);
and U17021 (N_17021,N_14316,N_12520);
nor U17022 (N_17022,N_13142,N_13258);
nand U17023 (N_17023,N_14194,N_14608);
nand U17024 (N_17024,N_13443,N_14214);
and U17025 (N_17025,N_12922,N_13107);
nor U17026 (N_17026,N_14673,N_14114);
and U17027 (N_17027,N_13524,N_12716);
and U17028 (N_17028,N_14543,N_13420);
xnor U17029 (N_17029,N_13711,N_12850);
or U17030 (N_17030,N_14076,N_13101);
or U17031 (N_17031,N_12742,N_14916);
or U17032 (N_17032,N_13919,N_13880);
nor U17033 (N_17033,N_14397,N_12689);
xor U17034 (N_17034,N_14246,N_14805);
nand U17035 (N_17035,N_14129,N_12510);
xnor U17036 (N_17036,N_12610,N_13421);
and U17037 (N_17037,N_14010,N_14355);
and U17038 (N_17038,N_14843,N_14520);
nor U17039 (N_17039,N_12843,N_13276);
xnor U17040 (N_17040,N_12818,N_14571);
nor U17041 (N_17041,N_12592,N_14398);
or U17042 (N_17042,N_12617,N_13286);
nor U17043 (N_17043,N_14953,N_14197);
nand U17044 (N_17044,N_13445,N_14292);
and U17045 (N_17045,N_13179,N_13150);
or U17046 (N_17046,N_13263,N_14530);
or U17047 (N_17047,N_13780,N_14936);
and U17048 (N_17048,N_14830,N_13398);
or U17049 (N_17049,N_14479,N_13869);
nor U17050 (N_17050,N_13431,N_12930);
and U17051 (N_17051,N_14565,N_13024);
nand U17052 (N_17052,N_13877,N_14109);
or U17053 (N_17053,N_14150,N_12781);
or U17054 (N_17054,N_13644,N_13137);
xnor U17055 (N_17055,N_14434,N_12545);
nand U17056 (N_17056,N_13113,N_12597);
or U17057 (N_17057,N_12861,N_13672);
nor U17058 (N_17058,N_13758,N_13281);
nand U17059 (N_17059,N_13122,N_13617);
and U17060 (N_17060,N_13877,N_14668);
nor U17061 (N_17061,N_12851,N_13618);
and U17062 (N_17062,N_13746,N_12638);
xor U17063 (N_17063,N_12917,N_14324);
nand U17064 (N_17064,N_12793,N_12841);
and U17065 (N_17065,N_13413,N_13922);
nand U17066 (N_17066,N_13769,N_13613);
or U17067 (N_17067,N_14387,N_13059);
xor U17068 (N_17068,N_14925,N_13093);
and U17069 (N_17069,N_13291,N_12510);
xnor U17070 (N_17070,N_14774,N_14872);
or U17071 (N_17071,N_14565,N_13027);
nor U17072 (N_17072,N_13760,N_14753);
nand U17073 (N_17073,N_14709,N_14928);
nor U17074 (N_17074,N_13877,N_14776);
nand U17075 (N_17075,N_14006,N_14218);
nor U17076 (N_17076,N_13363,N_13555);
xor U17077 (N_17077,N_13507,N_14421);
xnor U17078 (N_17078,N_14968,N_13766);
xor U17079 (N_17079,N_14394,N_12900);
and U17080 (N_17080,N_14315,N_13501);
or U17081 (N_17081,N_14297,N_14247);
nor U17082 (N_17082,N_13745,N_14926);
or U17083 (N_17083,N_13394,N_13617);
nor U17084 (N_17084,N_13068,N_13185);
xnor U17085 (N_17085,N_14147,N_13534);
nand U17086 (N_17086,N_14406,N_14904);
xnor U17087 (N_17087,N_14703,N_12954);
or U17088 (N_17088,N_12789,N_13518);
nor U17089 (N_17089,N_13912,N_12843);
nor U17090 (N_17090,N_14509,N_13193);
nor U17091 (N_17091,N_12639,N_14252);
nor U17092 (N_17092,N_14184,N_14327);
nor U17093 (N_17093,N_12788,N_14689);
nand U17094 (N_17094,N_13705,N_12555);
and U17095 (N_17095,N_12865,N_14128);
nor U17096 (N_17096,N_13885,N_12880);
or U17097 (N_17097,N_12781,N_14390);
xnor U17098 (N_17098,N_14564,N_13025);
xnor U17099 (N_17099,N_12705,N_14042);
and U17100 (N_17100,N_14853,N_12634);
or U17101 (N_17101,N_12744,N_12929);
or U17102 (N_17102,N_12955,N_14820);
nand U17103 (N_17103,N_14682,N_14405);
xor U17104 (N_17104,N_13526,N_14077);
or U17105 (N_17105,N_13738,N_14910);
xnor U17106 (N_17106,N_13297,N_14567);
or U17107 (N_17107,N_14690,N_14119);
nor U17108 (N_17108,N_12625,N_14406);
nand U17109 (N_17109,N_12506,N_13531);
and U17110 (N_17110,N_12954,N_13218);
xnor U17111 (N_17111,N_13503,N_14737);
and U17112 (N_17112,N_14926,N_13598);
and U17113 (N_17113,N_13572,N_14675);
xor U17114 (N_17114,N_14546,N_13513);
nand U17115 (N_17115,N_12865,N_13272);
and U17116 (N_17116,N_13521,N_14782);
nand U17117 (N_17117,N_14381,N_14603);
nor U17118 (N_17118,N_13886,N_13820);
or U17119 (N_17119,N_13470,N_12883);
nor U17120 (N_17120,N_14582,N_13591);
nor U17121 (N_17121,N_13044,N_13522);
or U17122 (N_17122,N_13954,N_13844);
or U17123 (N_17123,N_12929,N_13885);
xor U17124 (N_17124,N_12680,N_14963);
nor U17125 (N_17125,N_14680,N_13773);
or U17126 (N_17126,N_13452,N_12906);
nand U17127 (N_17127,N_14071,N_14958);
and U17128 (N_17128,N_12561,N_13454);
and U17129 (N_17129,N_12768,N_13332);
xnor U17130 (N_17130,N_14525,N_14380);
xnor U17131 (N_17131,N_14062,N_12980);
and U17132 (N_17132,N_13995,N_12515);
nor U17133 (N_17133,N_13473,N_14879);
xnor U17134 (N_17134,N_12604,N_12904);
xor U17135 (N_17135,N_14473,N_14132);
xor U17136 (N_17136,N_14967,N_14455);
nor U17137 (N_17137,N_12958,N_14358);
or U17138 (N_17138,N_12848,N_12578);
or U17139 (N_17139,N_12782,N_13046);
nand U17140 (N_17140,N_13158,N_14375);
and U17141 (N_17141,N_14832,N_12828);
nor U17142 (N_17142,N_13829,N_14705);
and U17143 (N_17143,N_14962,N_13443);
and U17144 (N_17144,N_13094,N_14106);
or U17145 (N_17145,N_13803,N_13206);
and U17146 (N_17146,N_12692,N_14061);
xor U17147 (N_17147,N_13797,N_13708);
xnor U17148 (N_17148,N_14472,N_14558);
nor U17149 (N_17149,N_13572,N_14310);
nor U17150 (N_17150,N_14549,N_14201);
nand U17151 (N_17151,N_14168,N_12936);
nor U17152 (N_17152,N_14948,N_13495);
xor U17153 (N_17153,N_14101,N_13388);
and U17154 (N_17154,N_13325,N_14167);
xor U17155 (N_17155,N_13508,N_14257);
and U17156 (N_17156,N_14281,N_12664);
and U17157 (N_17157,N_12966,N_12870);
or U17158 (N_17158,N_14401,N_13782);
nand U17159 (N_17159,N_13808,N_12693);
and U17160 (N_17160,N_14970,N_14258);
or U17161 (N_17161,N_12771,N_13445);
xnor U17162 (N_17162,N_14256,N_13817);
nor U17163 (N_17163,N_14709,N_13005);
nor U17164 (N_17164,N_14928,N_14829);
nor U17165 (N_17165,N_14280,N_14044);
xnor U17166 (N_17166,N_14141,N_13895);
and U17167 (N_17167,N_13326,N_12829);
and U17168 (N_17168,N_13560,N_13041);
xor U17169 (N_17169,N_14974,N_12666);
nand U17170 (N_17170,N_14893,N_14082);
or U17171 (N_17171,N_14599,N_13563);
nor U17172 (N_17172,N_14415,N_14418);
nand U17173 (N_17173,N_14267,N_13549);
xor U17174 (N_17174,N_12765,N_14016);
and U17175 (N_17175,N_12787,N_13960);
xnor U17176 (N_17176,N_12729,N_13341);
or U17177 (N_17177,N_13914,N_14431);
nor U17178 (N_17178,N_13460,N_13774);
xor U17179 (N_17179,N_14445,N_14992);
nand U17180 (N_17180,N_14379,N_13457);
nand U17181 (N_17181,N_12931,N_13431);
nand U17182 (N_17182,N_12572,N_14927);
and U17183 (N_17183,N_14505,N_12506);
xnor U17184 (N_17184,N_12671,N_14892);
or U17185 (N_17185,N_12916,N_14339);
or U17186 (N_17186,N_14149,N_14852);
nand U17187 (N_17187,N_13729,N_14997);
or U17188 (N_17188,N_14054,N_14602);
nor U17189 (N_17189,N_13809,N_14168);
nor U17190 (N_17190,N_14236,N_14750);
or U17191 (N_17191,N_12596,N_14049);
or U17192 (N_17192,N_14820,N_12808);
nand U17193 (N_17193,N_13184,N_12731);
or U17194 (N_17194,N_13675,N_14067);
and U17195 (N_17195,N_13159,N_13130);
or U17196 (N_17196,N_14518,N_14536);
nor U17197 (N_17197,N_12906,N_14831);
nor U17198 (N_17198,N_13662,N_14229);
xor U17199 (N_17199,N_14887,N_14810);
nor U17200 (N_17200,N_14906,N_14750);
nor U17201 (N_17201,N_13733,N_13366);
nor U17202 (N_17202,N_12642,N_14169);
and U17203 (N_17203,N_12563,N_13051);
nor U17204 (N_17204,N_12611,N_14877);
nand U17205 (N_17205,N_13447,N_13446);
nor U17206 (N_17206,N_14288,N_13777);
and U17207 (N_17207,N_14782,N_13538);
nor U17208 (N_17208,N_13569,N_14909);
and U17209 (N_17209,N_14708,N_13734);
and U17210 (N_17210,N_13437,N_14899);
nand U17211 (N_17211,N_14782,N_13838);
nor U17212 (N_17212,N_12525,N_14802);
nand U17213 (N_17213,N_14529,N_13257);
xor U17214 (N_17214,N_14151,N_14314);
or U17215 (N_17215,N_13676,N_13329);
or U17216 (N_17216,N_13669,N_13988);
xor U17217 (N_17217,N_13604,N_13690);
xor U17218 (N_17218,N_12886,N_13038);
and U17219 (N_17219,N_13821,N_12638);
nor U17220 (N_17220,N_14960,N_14618);
and U17221 (N_17221,N_13076,N_14147);
nand U17222 (N_17222,N_14074,N_13129);
nand U17223 (N_17223,N_14840,N_14647);
nand U17224 (N_17224,N_14062,N_14216);
nand U17225 (N_17225,N_13850,N_14529);
nand U17226 (N_17226,N_13023,N_13075);
nor U17227 (N_17227,N_14855,N_14579);
nand U17228 (N_17228,N_12701,N_14524);
and U17229 (N_17229,N_13988,N_13665);
and U17230 (N_17230,N_13913,N_12821);
and U17231 (N_17231,N_14230,N_13166);
xnor U17232 (N_17232,N_13561,N_12536);
and U17233 (N_17233,N_14804,N_13296);
or U17234 (N_17234,N_12795,N_14999);
and U17235 (N_17235,N_14131,N_12738);
nand U17236 (N_17236,N_14570,N_13685);
or U17237 (N_17237,N_14099,N_14185);
nand U17238 (N_17238,N_12555,N_13139);
nor U17239 (N_17239,N_13497,N_13548);
or U17240 (N_17240,N_14457,N_13007);
or U17241 (N_17241,N_12995,N_14729);
nor U17242 (N_17242,N_14975,N_14175);
or U17243 (N_17243,N_14217,N_14459);
nor U17244 (N_17244,N_12506,N_14523);
or U17245 (N_17245,N_13604,N_13951);
or U17246 (N_17246,N_12831,N_13876);
nand U17247 (N_17247,N_14227,N_14810);
or U17248 (N_17248,N_12764,N_13149);
or U17249 (N_17249,N_13152,N_13112);
and U17250 (N_17250,N_12809,N_14423);
nand U17251 (N_17251,N_13364,N_13081);
and U17252 (N_17252,N_13129,N_14183);
nor U17253 (N_17253,N_12693,N_13781);
nor U17254 (N_17254,N_14708,N_12766);
nand U17255 (N_17255,N_13935,N_14937);
or U17256 (N_17256,N_14377,N_13094);
nand U17257 (N_17257,N_14514,N_13321);
nor U17258 (N_17258,N_12828,N_12758);
nand U17259 (N_17259,N_14887,N_13585);
nand U17260 (N_17260,N_13478,N_14885);
and U17261 (N_17261,N_13183,N_14840);
and U17262 (N_17262,N_14725,N_13657);
and U17263 (N_17263,N_14453,N_13370);
xor U17264 (N_17264,N_13981,N_14743);
nor U17265 (N_17265,N_14485,N_12885);
or U17266 (N_17266,N_13621,N_14265);
nand U17267 (N_17267,N_12611,N_14372);
and U17268 (N_17268,N_13458,N_13474);
or U17269 (N_17269,N_13582,N_12581);
and U17270 (N_17270,N_12581,N_13846);
xnor U17271 (N_17271,N_13006,N_12759);
nor U17272 (N_17272,N_12718,N_13880);
xnor U17273 (N_17273,N_13354,N_13062);
nor U17274 (N_17274,N_14283,N_13503);
or U17275 (N_17275,N_13752,N_13424);
nor U17276 (N_17276,N_13420,N_12669);
or U17277 (N_17277,N_13067,N_13005);
nand U17278 (N_17278,N_13800,N_14774);
or U17279 (N_17279,N_12666,N_12636);
nor U17280 (N_17280,N_14938,N_14223);
xor U17281 (N_17281,N_14538,N_12881);
nand U17282 (N_17282,N_14101,N_14483);
or U17283 (N_17283,N_13902,N_13352);
and U17284 (N_17284,N_14359,N_13540);
nand U17285 (N_17285,N_13303,N_14705);
nand U17286 (N_17286,N_13475,N_13029);
and U17287 (N_17287,N_14223,N_13621);
or U17288 (N_17288,N_14192,N_13621);
or U17289 (N_17289,N_14535,N_13519);
and U17290 (N_17290,N_13698,N_14681);
and U17291 (N_17291,N_14483,N_14012);
or U17292 (N_17292,N_12907,N_14469);
nor U17293 (N_17293,N_14836,N_12991);
nand U17294 (N_17294,N_14485,N_12585);
nor U17295 (N_17295,N_13258,N_14432);
or U17296 (N_17296,N_12952,N_14426);
nor U17297 (N_17297,N_13986,N_12760);
nand U17298 (N_17298,N_14039,N_13066);
nor U17299 (N_17299,N_13800,N_13636);
nor U17300 (N_17300,N_13013,N_12572);
nor U17301 (N_17301,N_13091,N_12725);
or U17302 (N_17302,N_14282,N_12739);
and U17303 (N_17303,N_13887,N_12906);
xor U17304 (N_17304,N_14827,N_12713);
nor U17305 (N_17305,N_12896,N_13703);
nand U17306 (N_17306,N_14035,N_12823);
nor U17307 (N_17307,N_12581,N_14516);
or U17308 (N_17308,N_14753,N_13272);
xnor U17309 (N_17309,N_14776,N_14000);
xnor U17310 (N_17310,N_12606,N_14003);
or U17311 (N_17311,N_14267,N_14377);
and U17312 (N_17312,N_13579,N_13499);
xor U17313 (N_17313,N_14627,N_12508);
nor U17314 (N_17314,N_14844,N_14620);
or U17315 (N_17315,N_14450,N_14743);
and U17316 (N_17316,N_12682,N_14423);
nand U17317 (N_17317,N_12661,N_14469);
xnor U17318 (N_17318,N_13911,N_13244);
nor U17319 (N_17319,N_14671,N_13467);
or U17320 (N_17320,N_13464,N_13765);
xor U17321 (N_17321,N_13940,N_12584);
nand U17322 (N_17322,N_14177,N_12710);
and U17323 (N_17323,N_14680,N_14182);
or U17324 (N_17324,N_13635,N_14237);
xor U17325 (N_17325,N_13091,N_13935);
xnor U17326 (N_17326,N_13123,N_13679);
nor U17327 (N_17327,N_12812,N_14871);
nand U17328 (N_17328,N_14007,N_14157);
nand U17329 (N_17329,N_14230,N_13050);
xor U17330 (N_17330,N_13717,N_14820);
and U17331 (N_17331,N_14152,N_13160);
nand U17332 (N_17332,N_13965,N_13778);
and U17333 (N_17333,N_13964,N_13540);
or U17334 (N_17334,N_13486,N_13491);
nor U17335 (N_17335,N_12708,N_12653);
nand U17336 (N_17336,N_12880,N_14085);
nand U17337 (N_17337,N_13257,N_14598);
nand U17338 (N_17338,N_13792,N_12636);
xnor U17339 (N_17339,N_13087,N_14266);
nand U17340 (N_17340,N_13294,N_13384);
xnor U17341 (N_17341,N_12536,N_13190);
nor U17342 (N_17342,N_12982,N_13177);
or U17343 (N_17343,N_13338,N_14195);
xnor U17344 (N_17344,N_12556,N_14037);
and U17345 (N_17345,N_13815,N_14200);
and U17346 (N_17346,N_13992,N_14704);
nor U17347 (N_17347,N_12613,N_13112);
xor U17348 (N_17348,N_12722,N_12637);
or U17349 (N_17349,N_14877,N_14241);
or U17350 (N_17350,N_14983,N_14643);
xor U17351 (N_17351,N_12995,N_13243);
nand U17352 (N_17352,N_14490,N_14722);
and U17353 (N_17353,N_13895,N_14535);
nor U17354 (N_17354,N_12796,N_13067);
xnor U17355 (N_17355,N_13403,N_14460);
xnor U17356 (N_17356,N_13683,N_13279);
and U17357 (N_17357,N_14702,N_13728);
nor U17358 (N_17358,N_14868,N_13068);
nand U17359 (N_17359,N_14612,N_13568);
and U17360 (N_17360,N_13792,N_14644);
xnor U17361 (N_17361,N_14245,N_12865);
nor U17362 (N_17362,N_12757,N_14989);
xnor U17363 (N_17363,N_13545,N_13469);
nand U17364 (N_17364,N_13577,N_14221);
or U17365 (N_17365,N_14540,N_13398);
or U17366 (N_17366,N_13462,N_12897);
xnor U17367 (N_17367,N_14956,N_14503);
nor U17368 (N_17368,N_12945,N_13838);
nor U17369 (N_17369,N_12785,N_13243);
xnor U17370 (N_17370,N_14545,N_12876);
xnor U17371 (N_17371,N_12548,N_14355);
nand U17372 (N_17372,N_14654,N_14802);
nand U17373 (N_17373,N_13395,N_14444);
nor U17374 (N_17374,N_14536,N_13575);
and U17375 (N_17375,N_14645,N_12801);
or U17376 (N_17376,N_13988,N_13743);
or U17377 (N_17377,N_13302,N_13159);
nand U17378 (N_17378,N_13486,N_13364);
xnor U17379 (N_17379,N_14504,N_12871);
nor U17380 (N_17380,N_14911,N_13609);
xnor U17381 (N_17381,N_13894,N_12938);
or U17382 (N_17382,N_12511,N_14099);
nor U17383 (N_17383,N_14104,N_14652);
xnor U17384 (N_17384,N_14163,N_14762);
and U17385 (N_17385,N_12891,N_14865);
nor U17386 (N_17386,N_13322,N_12921);
and U17387 (N_17387,N_12821,N_12775);
nand U17388 (N_17388,N_13296,N_13915);
nand U17389 (N_17389,N_13299,N_13551);
xor U17390 (N_17390,N_12580,N_14520);
or U17391 (N_17391,N_13333,N_14893);
nand U17392 (N_17392,N_14801,N_14618);
nand U17393 (N_17393,N_12569,N_12760);
nand U17394 (N_17394,N_14373,N_12782);
or U17395 (N_17395,N_13870,N_12857);
and U17396 (N_17396,N_13946,N_13992);
xor U17397 (N_17397,N_13034,N_13103);
or U17398 (N_17398,N_13059,N_13038);
nand U17399 (N_17399,N_13332,N_13083);
or U17400 (N_17400,N_13654,N_14851);
nor U17401 (N_17401,N_14082,N_14537);
xor U17402 (N_17402,N_14842,N_14278);
or U17403 (N_17403,N_13767,N_14885);
nor U17404 (N_17404,N_13334,N_12886);
nor U17405 (N_17405,N_13918,N_13189);
or U17406 (N_17406,N_14970,N_13297);
and U17407 (N_17407,N_12926,N_12861);
and U17408 (N_17408,N_14672,N_14446);
nand U17409 (N_17409,N_14900,N_12602);
and U17410 (N_17410,N_14490,N_14315);
xnor U17411 (N_17411,N_13158,N_14007);
nor U17412 (N_17412,N_13064,N_14515);
nor U17413 (N_17413,N_13406,N_12545);
nand U17414 (N_17414,N_13892,N_12821);
nor U17415 (N_17415,N_13724,N_13981);
nor U17416 (N_17416,N_13708,N_12827);
nor U17417 (N_17417,N_14354,N_12974);
or U17418 (N_17418,N_13625,N_13940);
xnor U17419 (N_17419,N_12762,N_12565);
or U17420 (N_17420,N_13424,N_14630);
or U17421 (N_17421,N_14934,N_14278);
and U17422 (N_17422,N_14277,N_13277);
nand U17423 (N_17423,N_13985,N_14411);
xnor U17424 (N_17424,N_13818,N_14986);
and U17425 (N_17425,N_14250,N_14016);
or U17426 (N_17426,N_13466,N_14107);
and U17427 (N_17427,N_14960,N_13596);
nand U17428 (N_17428,N_13625,N_13929);
and U17429 (N_17429,N_13530,N_12501);
nor U17430 (N_17430,N_13253,N_12805);
nor U17431 (N_17431,N_14879,N_14983);
nor U17432 (N_17432,N_14465,N_12861);
nand U17433 (N_17433,N_13008,N_13427);
nor U17434 (N_17434,N_13685,N_13357);
nand U17435 (N_17435,N_13268,N_14058);
xnor U17436 (N_17436,N_14486,N_14850);
nand U17437 (N_17437,N_13080,N_14931);
or U17438 (N_17438,N_13636,N_13208);
nand U17439 (N_17439,N_13629,N_12619);
xnor U17440 (N_17440,N_14942,N_14055);
and U17441 (N_17441,N_12570,N_14843);
nand U17442 (N_17442,N_14030,N_13006);
nand U17443 (N_17443,N_14922,N_14411);
xor U17444 (N_17444,N_12740,N_14140);
xor U17445 (N_17445,N_13403,N_12883);
nand U17446 (N_17446,N_14560,N_12795);
or U17447 (N_17447,N_14261,N_14131);
or U17448 (N_17448,N_13543,N_14763);
and U17449 (N_17449,N_14964,N_13083);
xnor U17450 (N_17450,N_14759,N_12862);
nand U17451 (N_17451,N_14264,N_14625);
or U17452 (N_17452,N_14151,N_12794);
or U17453 (N_17453,N_13445,N_14427);
xnor U17454 (N_17454,N_14242,N_13811);
nand U17455 (N_17455,N_14568,N_14010);
nand U17456 (N_17456,N_13567,N_14321);
nand U17457 (N_17457,N_13564,N_13205);
xnor U17458 (N_17458,N_13057,N_14802);
or U17459 (N_17459,N_14647,N_13039);
and U17460 (N_17460,N_12607,N_14691);
or U17461 (N_17461,N_14657,N_13585);
nand U17462 (N_17462,N_13906,N_12561);
and U17463 (N_17463,N_13587,N_14393);
and U17464 (N_17464,N_14158,N_14198);
or U17465 (N_17465,N_14728,N_12901);
and U17466 (N_17466,N_14963,N_12887);
or U17467 (N_17467,N_12564,N_14931);
nand U17468 (N_17468,N_14826,N_12751);
xnor U17469 (N_17469,N_13691,N_14033);
nor U17470 (N_17470,N_14454,N_13796);
xor U17471 (N_17471,N_14646,N_13146);
nand U17472 (N_17472,N_14556,N_13050);
and U17473 (N_17473,N_12946,N_14296);
nand U17474 (N_17474,N_13813,N_12543);
xnor U17475 (N_17475,N_14085,N_12519);
nand U17476 (N_17476,N_12500,N_14299);
nand U17477 (N_17477,N_12922,N_12958);
nor U17478 (N_17478,N_13141,N_13924);
and U17479 (N_17479,N_13477,N_13275);
nand U17480 (N_17480,N_14189,N_13525);
xnor U17481 (N_17481,N_13061,N_13869);
nor U17482 (N_17482,N_13680,N_14247);
nor U17483 (N_17483,N_14070,N_14841);
nand U17484 (N_17484,N_13887,N_13956);
or U17485 (N_17485,N_14951,N_12650);
or U17486 (N_17486,N_14955,N_13577);
xor U17487 (N_17487,N_13145,N_14498);
and U17488 (N_17488,N_14788,N_14913);
or U17489 (N_17489,N_13654,N_12978);
nand U17490 (N_17490,N_14789,N_12886);
xor U17491 (N_17491,N_14618,N_12997);
and U17492 (N_17492,N_14135,N_13087);
xnor U17493 (N_17493,N_13411,N_14976);
or U17494 (N_17494,N_12525,N_12586);
xnor U17495 (N_17495,N_14183,N_12810);
nand U17496 (N_17496,N_12923,N_12929);
xor U17497 (N_17497,N_13809,N_13462);
nor U17498 (N_17498,N_13809,N_12594);
xnor U17499 (N_17499,N_12615,N_13426);
nor U17500 (N_17500,N_15607,N_16747);
nor U17501 (N_17501,N_15989,N_15099);
nor U17502 (N_17502,N_16234,N_15817);
or U17503 (N_17503,N_16423,N_15695);
nor U17504 (N_17504,N_16185,N_17311);
nand U17505 (N_17505,N_16861,N_15257);
nand U17506 (N_17506,N_17203,N_15545);
and U17507 (N_17507,N_15045,N_17373);
nor U17508 (N_17508,N_16481,N_15402);
nand U17509 (N_17509,N_17446,N_17222);
nand U17510 (N_17510,N_17286,N_15575);
xor U17511 (N_17511,N_15993,N_16233);
or U17512 (N_17512,N_15332,N_17452);
nor U17513 (N_17513,N_16199,N_15300);
xnor U17514 (N_17514,N_15723,N_16084);
or U17515 (N_17515,N_16552,N_16476);
or U17516 (N_17516,N_16532,N_17433);
nand U17517 (N_17517,N_15017,N_15763);
and U17518 (N_17518,N_17183,N_17475);
nand U17519 (N_17519,N_16804,N_15442);
nand U17520 (N_17520,N_15736,N_17482);
nor U17521 (N_17521,N_15034,N_16181);
and U17522 (N_17522,N_15433,N_15251);
xnor U17523 (N_17523,N_15363,N_17226);
nor U17524 (N_17524,N_16628,N_15127);
xor U17525 (N_17525,N_17239,N_16895);
nand U17526 (N_17526,N_16375,N_15120);
nor U17527 (N_17527,N_16820,N_15177);
and U17528 (N_17528,N_16781,N_16283);
xor U17529 (N_17529,N_15183,N_15794);
and U17530 (N_17530,N_15956,N_16454);
or U17531 (N_17531,N_15893,N_16878);
and U17532 (N_17532,N_16665,N_15046);
xnor U17533 (N_17533,N_15854,N_16852);
nand U17534 (N_17534,N_16396,N_15002);
nand U17535 (N_17535,N_16395,N_16633);
and U17536 (N_17536,N_16831,N_16240);
xnor U17537 (N_17537,N_15862,N_16042);
and U17538 (N_17538,N_17251,N_16179);
nand U17539 (N_17539,N_16510,N_17093);
nor U17540 (N_17540,N_15281,N_16448);
nor U17541 (N_17541,N_17212,N_17437);
or U17542 (N_17542,N_15542,N_16700);
and U17543 (N_17543,N_16856,N_17380);
nand U17544 (N_17544,N_17220,N_17229);
xor U17545 (N_17545,N_15303,N_15248);
xnor U17546 (N_17546,N_16288,N_16349);
and U17547 (N_17547,N_15319,N_16818);
or U17548 (N_17548,N_15296,N_17237);
or U17549 (N_17549,N_15440,N_17135);
nand U17550 (N_17550,N_16620,N_15239);
and U17551 (N_17551,N_16544,N_15153);
nor U17552 (N_17552,N_17090,N_15829);
and U17553 (N_17553,N_17391,N_15224);
nand U17554 (N_17554,N_15881,N_16365);
xnor U17555 (N_17555,N_16276,N_16488);
or U17556 (N_17556,N_17315,N_15681);
xnor U17557 (N_17557,N_15385,N_17271);
or U17558 (N_17558,N_15636,N_15826);
nand U17559 (N_17559,N_17454,N_17416);
nand U17560 (N_17560,N_16703,N_16829);
nor U17561 (N_17561,N_15538,N_15503);
xor U17562 (N_17562,N_16340,N_16063);
nand U17563 (N_17563,N_15596,N_16688);
or U17564 (N_17564,N_15412,N_16145);
nand U17565 (N_17565,N_16428,N_15949);
and U17566 (N_17566,N_15320,N_15137);
nor U17567 (N_17567,N_15079,N_15330);
and U17568 (N_17568,N_16743,N_15197);
nand U17569 (N_17569,N_17221,N_16260);
xor U17570 (N_17570,N_15124,N_16641);
or U17571 (N_17571,N_15109,N_16668);
nor U17572 (N_17572,N_17146,N_16192);
and U17573 (N_17573,N_17334,N_15738);
nand U17574 (N_17574,N_17164,N_16606);
nor U17575 (N_17575,N_17044,N_15876);
nor U17576 (N_17576,N_15858,N_15229);
nor U17577 (N_17577,N_15592,N_15312);
or U17578 (N_17578,N_16092,N_17361);
xnor U17579 (N_17579,N_16971,N_16989);
nor U17580 (N_17580,N_16549,N_17127);
and U17581 (N_17581,N_15253,N_17255);
nand U17582 (N_17582,N_17425,N_16733);
xor U17583 (N_17583,N_16027,N_15050);
nor U17584 (N_17584,N_15992,N_17245);
and U17585 (N_17585,N_15907,N_15613);
nand U17586 (N_17586,N_15806,N_16422);
xnor U17587 (N_17587,N_16585,N_15689);
nand U17588 (N_17588,N_17216,N_17342);
xor U17589 (N_17589,N_16958,N_15174);
nor U17590 (N_17590,N_16296,N_16386);
nor U17591 (N_17591,N_16931,N_16754);
and U17592 (N_17592,N_16123,N_17075);
nor U17593 (N_17593,N_17247,N_17148);
nand U17594 (N_17594,N_16963,N_15697);
nand U17595 (N_17595,N_17491,N_16498);
nor U17596 (N_17596,N_16011,N_15435);
nor U17597 (N_17597,N_15105,N_17029);
nand U17598 (N_17598,N_16095,N_16682);
and U17599 (N_17599,N_16307,N_17483);
or U17600 (N_17600,N_16281,N_15717);
xnor U17601 (N_17601,N_16290,N_16492);
or U17602 (N_17602,N_15390,N_16387);
nor U17603 (N_17603,N_15485,N_15850);
or U17604 (N_17604,N_15111,N_15539);
and U17605 (N_17605,N_17367,N_15737);
and U17606 (N_17606,N_17206,N_15928);
or U17607 (N_17607,N_16675,N_15874);
or U17608 (N_17608,N_15983,N_16566);
and U17609 (N_17609,N_15943,N_17412);
nor U17610 (N_17610,N_16035,N_16659);
xnor U17611 (N_17611,N_15525,N_17041);
nand U17612 (N_17612,N_15375,N_17473);
nand U17613 (N_17613,N_17072,N_15166);
xnor U17614 (N_17614,N_15511,N_15128);
nand U17615 (N_17615,N_17031,N_16917);
xnor U17616 (N_17616,N_15527,N_17046);
or U17617 (N_17617,N_15643,N_15811);
nor U17618 (N_17618,N_16681,N_16266);
xor U17619 (N_17619,N_15703,N_15916);
xnor U17620 (N_17620,N_17336,N_17394);
or U17621 (N_17621,N_17295,N_17376);
nand U17622 (N_17622,N_15043,N_17118);
xnor U17623 (N_17623,N_16708,N_16982);
nor U17624 (N_17624,N_15199,N_16564);
and U17625 (N_17625,N_16643,N_17460);
xnor U17626 (N_17626,N_16467,N_15944);
and U17627 (N_17627,N_16978,N_16739);
or U17628 (N_17628,N_15634,N_17094);
or U17629 (N_17629,N_15600,N_15213);
and U17630 (N_17630,N_16038,N_16022);
nand U17631 (N_17631,N_16079,N_16049);
nand U17632 (N_17632,N_17038,N_17018);
xor U17633 (N_17633,N_15187,N_17450);
nor U17634 (N_17634,N_15740,N_15221);
and U17635 (N_17635,N_17474,N_16600);
nor U17636 (N_17636,N_15752,N_16134);
xnor U17637 (N_17637,N_15730,N_15981);
nand U17638 (N_17638,N_17154,N_15479);
and U17639 (N_17639,N_15360,N_16830);
xor U17640 (N_17640,N_15204,N_17250);
nand U17641 (N_17641,N_15914,N_16112);
or U17642 (N_17642,N_15472,N_16166);
and U17643 (N_17643,N_17443,N_16259);
nor U17644 (N_17644,N_15147,N_17277);
nor U17645 (N_17645,N_16937,N_15578);
and U17646 (N_17646,N_16823,N_17264);
nor U17647 (N_17647,N_15693,N_16440);
and U17648 (N_17648,N_17400,N_17134);
or U17649 (N_17649,N_15387,N_15875);
or U17650 (N_17650,N_17370,N_16973);
xnor U17651 (N_17651,N_15522,N_17301);
nor U17652 (N_17652,N_16378,N_16923);
nand U17653 (N_17653,N_15136,N_16886);
or U17654 (N_17654,N_17177,N_15181);
and U17655 (N_17655,N_15800,N_15805);
nor U17656 (N_17656,N_16920,N_15910);
or U17657 (N_17657,N_15945,N_17346);
or U17658 (N_17658,N_15408,N_15236);
nor U17659 (N_17659,N_16197,N_17492);
nor U17660 (N_17660,N_17257,N_16508);
nor U17661 (N_17661,N_15097,N_17432);
xnor U17662 (N_17662,N_15658,N_15698);
nor U17663 (N_17663,N_16985,N_17019);
xnor U17664 (N_17664,N_15477,N_16983);
xnor U17665 (N_17665,N_15597,N_16790);
or U17666 (N_17666,N_15628,N_16556);
or U17667 (N_17667,N_15941,N_16252);
nand U17668 (N_17668,N_16175,N_15947);
or U17669 (N_17669,N_16597,N_16928);
nand U17670 (N_17670,N_15116,N_15107);
nand U17671 (N_17671,N_15190,N_15306);
xor U17672 (N_17672,N_16466,N_15062);
xor U17673 (N_17673,N_16486,N_16418);
or U17674 (N_17674,N_16086,N_17055);
xnor U17675 (N_17675,N_16315,N_16726);
and U17676 (N_17676,N_15683,N_15798);
xnor U17677 (N_17677,N_15238,N_15401);
nand U17678 (N_17678,N_16356,N_16059);
nor U17679 (N_17679,N_16594,N_15568);
nor U17680 (N_17680,N_15760,N_16222);
xnor U17681 (N_17681,N_16940,N_16780);
nand U17682 (N_17682,N_16526,N_15548);
or U17683 (N_17683,N_16507,N_17372);
and U17684 (N_17684,N_16026,N_15140);
or U17685 (N_17685,N_17084,N_16696);
nor U17686 (N_17686,N_16225,N_16490);
or U17687 (N_17687,N_16727,N_15513);
or U17688 (N_17688,N_16713,N_16006);
xor U17689 (N_17689,N_16002,N_17179);
nor U17690 (N_17690,N_16817,N_15493);
xor U17691 (N_17691,N_17027,N_15583);
xor U17692 (N_17692,N_16915,N_16875);
nand U17693 (N_17693,N_17100,N_16005);
or U17694 (N_17694,N_16216,N_17086);
nand U17695 (N_17695,N_15845,N_17371);
nor U17696 (N_17696,N_15599,N_15973);
nor U17697 (N_17697,N_16630,N_16207);
nand U17698 (N_17698,N_15155,N_15103);
xor U17699 (N_17699,N_16200,N_16567);
nor U17700 (N_17700,N_15749,N_16913);
or U17701 (N_17701,N_16907,N_17061);
nor U17702 (N_17702,N_16114,N_15096);
nor U17703 (N_17703,N_16081,N_16598);
or U17704 (N_17704,N_15788,N_16047);
xnor U17705 (N_17705,N_15486,N_15610);
and U17706 (N_17706,N_17350,N_17248);
nand U17707 (N_17707,N_17362,N_16029);
and U17708 (N_17708,N_16221,N_16496);
xor U17709 (N_17709,N_16096,N_17211);
and U17710 (N_17710,N_15781,N_17276);
and U17711 (N_17711,N_16772,N_16477);
or U17712 (N_17712,N_16401,N_15235);
nand U17713 (N_17713,N_15972,N_15500);
nand U17714 (N_17714,N_15092,N_17014);
nor U17715 (N_17715,N_17244,N_16310);
or U17716 (N_17716,N_15008,N_17156);
nand U17717 (N_17717,N_15333,N_16309);
xor U17718 (N_17718,N_16004,N_17291);
and U17719 (N_17719,N_16302,N_17403);
and U17720 (N_17720,N_17411,N_16765);
and U17721 (N_17721,N_15203,N_16586);
and U17722 (N_17722,N_16250,N_15437);
and U17723 (N_17723,N_16948,N_16720);
and U17724 (N_17724,N_16226,N_16794);
xor U17725 (N_17725,N_16832,N_16445);
nor U17726 (N_17726,N_17321,N_15428);
xor U17727 (N_17727,N_17360,N_15612);
nand U17728 (N_17728,N_16909,N_16455);
and U17729 (N_17729,N_16009,N_16548);
nor U17730 (N_17730,N_17102,N_17444);
xor U17731 (N_17731,N_16591,N_17363);
nor U17732 (N_17732,N_15378,N_16786);
nor U17733 (N_17733,N_16358,N_15819);
and U17734 (N_17734,N_17340,N_16361);
xor U17735 (N_17735,N_16242,N_16291);
or U17736 (N_17736,N_17149,N_16570);
and U17737 (N_17737,N_15812,N_15409);
xor U17738 (N_17738,N_15744,N_15556);
or U17739 (N_17739,N_16057,N_15519);
nand U17740 (N_17740,N_17457,N_16524);
and U17741 (N_17741,N_17185,N_16795);
and U17742 (N_17742,N_17083,N_15460);
nand U17743 (N_17743,N_17407,N_15368);
nand U17744 (N_17744,N_15001,N_16874);
nor U17745 (N_17745,N_16205,N_15345);
nand U17746 (N_17746,N_15842,N_15344);
or U17747 (N_17747,N_16579,N_15158);
or U17748 (N_17748,N_15160,N_15976);
nand U17749 (N_17749,N_15671,N_17181);
nand U17750 (N_17750,N_16131,N_16328);
or U17751 (N_17751,N_15362,N_17263);
nor U17752 (N_17752,N_15739,N_15093);
and U17753 (N_17753,N_17007,N_15807);
xor U17754 (N_17754,N_16887,N_16629);
xnor U17755 (N_17755,N_17304,N_15899);
nand U17756 (N_17756,N_15751,N_17485);
and U17757 (N_17757,N_16483,N_16609);
or U17758 (N_17758,N_16984,N_17498);
nand U17759 (N_17759,N_15870,N_16213);
xnor U17760 (N_17760,N_15076,N_16655);
or U17761 (N_17761,N_17218,N_17104);
or U17762 (N_17762,N_16834,N_16130);
xnor U17763 (N_17763,N_17115,N_16974);
nor U17764 (N_17764,N_16761,N_15066);
nand U17765 (N_17765,N_17385,N_16154);
nor U17766 (N_17766,N_15650,N_15929);
xnor U17767 (N_17767,N_17223,N_16444);
or U17768 (N_17768,N_17052,N_15787);
or U17769 (N_17769,N_16561,N_15821);
nor U17770 (N_17770,N_17441,N_16229);
or U17771 (N_17771,N_17172,N_15492);
xnor U17772 (N_17772,N_16404,N_16788);
nand U17773 (N_17773,N_16777,N_17284);
and U17774 (N_17774,N_15586,N_16402);
xor U17775 (N_17775,N_16683,N_17314);
and U17776 (N_17776,N_16731,N_15713);
nor U17777 (N_17777,N_16415,N_15524);
xnor U17778 (N_17778,N_15595,N_17410);
nand U17779 (N_17779,N_15172,N_15232);
nor U17780 (N_17780,N_15655,N_16419);
nand U17781 (N_17781,N_16413,N_16089);
nand U17782 (N_17782,N_16452,N_15497);
and U17783 (N_17783,N_16209,N_15543);
nor U17784 (N_17784,N_15252,N_16749);
nor U17785 (N_17785,N_16143,N_15380);
nor U17786 (N_17786,N_16577,N_17236);
xor U17787 (N_17787,N_15642,N_16157);
xor U17788 (N_17788,N_17010,N_17274);
nor U17789 (N_17789,N_16345,N_15678);
xor U17790 (N_17790,N_17493,N_16075);
nor U17791 (N_17791,N_16730,N_16919);
xor U17792 (N_17792,N_17106,N_16922);
and U17793 (N_17793,N_17117,N_16491);
nand U17794 (N_17794,N_15413,N_15579);
and U17795 (N_17795,N_17005,N_16450);
and U17796 (N_17796,N_16278,N_16468);
nand U17797 (N_17797,N_15459,N_16254);
and U17798 (N_17798,N_16124,N_17289);
and U17799 (N_17799,N_16836,N_16531);
xor U17800 (N_17800,N_17316,N_15509);
nand U17801 (N_17801,N_15178,N_16107);
and U17802 (N_17802,N_16397,N_15660);
and U17803 (N_17803,N_15036,N_15661);
nand U17804 (N_17804,N_17079,N_16693);
and U17805 (N_17805,N_15602,N_15733);
nand U17806 (N_17806,N_17024,N_17144);
or U17807 (N_17807,N_17310,N_15209);
or U17808 (N_17808,N_15028,N_15264);
nor U17809 (N_17809,N_17298,N_16332);
nand U17810 (N_17810,N_17497,N_16458);
xnor U17811 (N_17811,N_15039,N_16146);
nor U17812 (N_17812,N_15631,N_17208);
nor U17813 (N_17813,N_15756,N_17200);
or U17814 (N_17814,N_16333,N_15984);
or U17815 (N_17815,N_15016,N_15145);
xor U17816 (N_17816,N_15887,N_15063);
nand U17817 (N_17817,N_16778,N_16479);
and U17818 (N_17818,N_16545,N_17260);
nand U17819 (N_17819,N_17068,N_16807);
nor U17820 (N_17820,N_17365,N_15827);
or U17821 (N_17821,N_17309,N_15102);
or U17822 (N_17822,N_17125,N_16992);
nand U17823 (N_17823,N_16416,N_15786);
nand U17824 (N_17824,N_17012,N_16742);
and U17825 (N_17825,N_15889,N_15902);
xor U17826 (N_17826,N_15393,N_17170);
nor U17827 (N_17827,N_15975,N_15216);
nand U17828 (N_17828,N_16306,N_15569);
or U17829 (N_17829,N_15732,N_15215);
nor U17830 (N_17830,N_17300,N_17327);
xor U17831 (N_17831,N_16624,N_16286);
xnor U17832 (N_17832,N_17477,N_15270);
nand U17833 (N_17833,N_17252,N_15741);
nor U17834 (N_17834,N_15852,N_16910);
nor U17835 (N_17835,N_16582,N_16756);
xnor U17836 (N_17836,N_17230,N_15377);
and U17837 (N_17837,N_17002,N_15423);
nor U17838 (N_17838,N_16824,N_16964);
nor U17839 (N_17839,N_15449,N_17338);
xnor U17840 (N_17840,N_16251,N_17076);
and U17841 (N_17841,N_16892,N_17234);
nor U17842 (N_17842,N_15226,N_15243);
nor U17843 (N_17843,N_15272,N_15411);
and U17844 (N_17844,N_17466,N_16784);
or U17845 (N_17845,N_15011,N_17349);
xor U17846 (N_17846,N_16344,N_17312);
xnor U17847 (N_17847,N_16826,N_17313);
or U17848 (N_17848,N_15255,N_16870);
nand U17849 (N_17849,N_17438,N_17069);
xnor U17850 (N_17850,N_15588,N_15835);
and U17851 (N_17851,N_16596,N_16246);
and U17852 (N_17852,N_15946,N_16966);
or U17853 (N_17853,N_15635,N_16300);
nor U17854 (N_17854,N_16894,N_16190);
nor U17855 (N_17855,N_15774,N_15657);
xor U17856 (N_17856,N_16899,N_16627);
and U17857 (N_17857,N_15026,N_16076);
and U17858 (N_17858,N_17000,N_16243);
nor U17859 (N_17859,N_15978,N_15968);
nor U17860 (N_17860,N_16196,N_15911);
nor U17861 (N_17861,N_16269,N_17063);
and U17862 (N_17862,N_16798,N_15388);
or U17863 (N_17863,N_16712,N_15591);
xor U17864 (N_17864,N_16433,N_17131);
nor U17865 (N_17865,N_17130,N_16939);
or U17866 (N_17866,N_15176,N_15715);
xor U17867 (N_17867,N_16563,N_15258);
xnor U17868 (N_17868,N_16789,N_15626);
and U17869 (N_17869,N_16019,N_16580);
or U17870 (N_17870,N_17455,N_16148);
xnor U17871 (N_17871,N_16253,N_15397);
nand U17872 (N_17872,N_15623,N_16980);
and U17873 (N_17873,N_16745,N_17337);
nand U17874 (N_17874,N_15982,N_15095);
nand U17875 (N_17875,N_16204,N_15572);
nand U17876 (N_17876,N_17070,N_16847);
or U17877 (N_17877,N_16128,N_16295);
or U17878 (N_17878,N_15188,N_17384);
and U17879 (N_17879,N_15815,N_16871);
xnor U17880 (N_17880,N_16334,N_15672);
or U17881 (N_17881,N_15173,N_16429);
and U17882 (N_17882,N_16136,N_15259);
xnor U17883 (N_17883,N_16152,N_15206);
or U17884 (N_17884,N_17352,N_17249);
xor U17885 (N_17885,N_16317,N_15339);
and U17886 (N_17886,N_16523,N_16631);
nor U17887 (N_17887,N_15718,N_17341);
xor U17888 (N_17888,N_16129,N_16318);
and U17889 (N_17889,N_15919,N_16319);
nor U17890 (N_17890,N_17199,N_17173);
xor U17891 (N_17891,N_17267,N_16719);
nand U17892 (N_17892,N_15376,N_16881);
or U17893 (N_17893,N_15802,N_16037);
nor U17894 (N_17894,N_16137,N_15381);
and U17895 (N_17895,N_16374,N_15784);
nor U17896 (N_17896,N_15777,N_17382);
xor U17897 (N_17897,N_15405,N_15117);
and U17898 (N_17898,N_17458,N_17030);
or U17899 (N_17899,N_17499,N_16670);
xor U17900 (N_17900,N_15824,N_17241);
or U17901 (N_17901,N_15957,N_16069);
nand U17902 (N_17902,N_16686,N_15419);
and U17903 (N_17903,N_17461,N_17140);
nand U17904 (N_17904,N_15645,N_16028);
nor U17905 (N_17905,N_15220,N_15669);
xnor U17906 (N_17906,N_16372,N_17355);
and U17907 (N_17907,N_16411,N_16993);
or U17908 (N_17908,N_15065,N_15906);
nand U17909 (N_17909,N_16487,N_16064);
nor U17910 (N_17910,N_17123,N_15663);
nand U17911 (N_17911,N_15013,N_15310);
and U17912 (N_17912,N_16149,N_15284);
xnor U17913 (N_17913,N_15892,N_15585);
or U17914 (N_17914,N_15084,N_16692);
and U17915 (N_17915,N_16275,N_16336);
nor U17916 (N_17916,N_16439,N_15304);
nand U17917 (N_17917,N_16048,N_16799);
and U17918 (N_17918,N_16421,N_16967);
xnor U17919 (N_17919,N_16043,N_16465);
nor U17920 (N_17920,N_15776,N_16088);
nand U17921 (N_17921,N_15044,N_15951);
and U17922 (N_17922,N_15133,N_15307);
or U17923 (N_17923,N_15652,N_17465);
xnor U17924 (N_17924,N_15894,N_15508);
nand U17925 (N_17925,N_16759,N_16768);
xor U17926 (N_17926,N_16592,N_15233);
nand U17927 (N_17927,N_16844,N_17353);
nand U17928 (N_17928,N_16188,N_15465);
nor U17929 (N_17929,N_17449,N_15048);
nand U17930 (N_17930,N_17469,N_15901);
or U17931 (N_17931,N_16257,N_16431);
xnor U17932 (N_17932,N_15438,N_15980);
and U17933 (N_17933,N_15474,N_15654);
and U17934 (N_17934,N_17377,N_15020);
and U17935 (N_17935,N_15676,N_15125);
nand U17936 (N_17936,N_15990,N_15955);
and U17937 (N_17937,N_16678,N_15922);
nand U17938 (N_17938,N_16626,N_16699);
xnor U17939 (N_17939,N_16791,N_15799);
and U17940 (N_17940,N_15603,N_16947);
nor U17941 (N_17941,N_16868,N_15491);
xor U17942 (N_17942,N_15856,N_16156);
xor U17943 (N_17943,N_15974,N_17167);
nand U17944 (N_17944,N_17393,N_16827);
or U17945 (N_17945,N_16877,N_15115);
xnor U17946 (N_17946,N_15078,N_16173);
and U17947 (N_17947,N_16371,N_16031);
and U17948 (N_17948,N_15534,N_17472);
xor U17949 (N_17949,N_15407,N_16648);
nand U17950 (N_17950,N_17097,N_15970);
or U17951 (N_17951,N_17378,N_17111);
or U17952 (N_17952,N_15242,N_16554);
nor U17953 (N_17953,N_16614,N_17490);
or U17954 (N_17954,N_16998,N_16674);
xnor U17955 (N_17955,N_16521,N_16108);
nand U17956 (N_17956,N_15447,N_15085);
nand U17957 (N_17957,N_15694,N_15606);
nand U17958 (N_17958,N_17120,N_16697);
xnor U17959 (N_17959,N_16835,N_16932);
or U17960 (N_17960,N_16459,N_15262);
nor U17961 (N_17961,N_16390,N_15753);
or U17962 (N_17962,N_16441,N_16559);
and U17963 (N_17963,N_17109,N_16325);
nor U17964 (N_17964,N_16119,N_16921);
or U17965 (N_17965,N_16294,N_16640);
and U17966 (N_17966,N_16093,N_17161);
nor U17967 (N_17967,N_17088,N_16695);
and U17968 (N_17968,N_15818,N_15561);
or U17969 (N_17969,N_16438,N_15415);
nand U17970 (N_17970,N_16228,N_15836);
and U17971 (N_17971,N_15189,N_16535);
xor U17972 (N_17972,N_17166,N_15100);
nor U17973 (N_17973,N_17045,N_15987);
nor U17974 (N_17974,N_15536,N_17113);
xnor U17975 (N_17975,N_16258,N_15716);
nand U17976 (N_17976,N_16007,N_15927);
nand U17977 (N_17977,N_15832,N_16127);
nand U17978 (N_17978,N_17348,N_16273);
nor U17979 (N_17979,N_17253,N_16198);
nand U17980 (N_17980,N_15179,N_17470);
and U17981 (N_17981,N_16808,N_15466);
nor U17982 (N_17982,N_15131,N_17488);
and U17983 (N_17983,N_15988,N_15454);
nor U17984 (N_17984,N_16469,N_16694);
xor U17985 (N_17985,N_17194,N_16351);
nand U17986 (N_17986,N_17142,N_16320);
nand U17987 (N_17987,N_15195,N_16572);
xnor U17988 (N_17988,N_15544,N_17379);
and U17989 (N_17989,N_17098,N_16854);
and U17990 (N_17990,N_16812,N_17035);
nand U17991 (N_17991,N_15727,N_17178);
nand U17992 (N_17992,N_15614,N_16965);
nor U17993 (N_17993,N_16426,N_15418);
and U17994 (N_17994,N_15487,N_16977);
and U17995 (N_17995,N_15468,N_15664);
xor U17996 (N_17996,N_16999,N_15374);
nor U17997 (N_17997,N_15331,N_15383);
or U17998 (N_17998,N_15847,N_15604);
nor U17999 (N_17999,N_17463,N_16389);
or U18000 (N_18000,N_16480,N_15015);
nor U18001 (N_18001,N_16359,N_16509);
nor U18002 (N_18002,N_16212,N_16217);
nand U18003 (N_18003,N_15322,N_17165);
nand U18004 (N_18004,N_16357,N_17112);
nor U18005 (N_18005,N_16806,N_16470);
nor U18006 (N_18006,N_16083,N_16908);
nor U18007 (N_18007,N_16153,N_17282);
and U18008 (N_18008,N_15040,N_15343);
nor U18009 (N_18009,N_17395,N_17037);
nor U18010 (N_18010,N_15139,N_16132);
xor U18011 (N_18011,N_16734,N_16863);
or U18012 (N_18012,N_15848,N_17272);
nor U18013 (N_18013,N_16355,N_16970);
nand U18014 (N_18014,N_16018,N_15638);
nor U18015 (N_18015,N_15594,N_16403);
xnor U18016 (N_18016,N_16430,N_15969);
and U18017 (N_18017,N_15593,N_17413);
or U18018 (N_18018,N_16723,N_15882);
nor U18019 (N_18019,N_15478,N_15677);
nor U18020 (N_18020,N_15762,N_16612);
nor U18021 (N_18021,N_15152,N_15735);
or U18022 (N_18022,N_16698,N_16056);
nand U18023 (N_18023,N_16534,N_15900);
or U18024 (N_18024,N_15210,N_15324);
and U18025 (N_18025,N_17332,N_16193);
xnor U18026 (N_18026,N_17296,N_15425);
and U18027 (N_18027,N_17042,N_15617);
or U18028 (N_18028,N_16822,N_15912);
xnor U18029 (N_18029,N_15072,N_16638);
xnor U18030 (N_18030,N_17190,N_17462);
nor U18031 (N_18031,N_16391,N_16417);
or U18032 (N_18032,N_15682,N_16451);
nor U18033 (N_18033,N_16044,N_16800);
and U18034 (N_18034,N_17459,N_16410);
or U18035 (N_18035,N_15861,N_15532);
or U18036 (N_18036,N_16223,N_16161);
and U18037 (N_18037,N_15649,N_17006);
nor U18038 (N_18038,N_15445,N_15632);
and U18039 (N_18039,N_15446,N_17331);
xor U18040 (N_18040,N_15049,N_17453);
xnor U18041 (N_18041,N_15554,N_15742);
xor U18042 (N_18042,N_17189,N_15456);
xor U18043 (N_18043,N_17417,N_16456);
nor U18044 (N_18044,N_15728,N_15481);
and U18045 (N_18045,N_16017,N_15184);
nor U18046 (N_18046,N_15247,N_17081);
xor U18047 (N_18047,N_16851,N_15926);
or U18048 (N_18048,N_15104,N_15334);
or U18049 (N_18049,N_16715,N_16343);
nand U18050 (N_18050,N_17424,N_17442);
and U18051 (N_18051,N_16741,N_16218);
and U18052 (N_18052,N_17383,N_17387);
and U18053 (N_18053,N_15641,N_16687);
nor U18054 (N_18054,N_16764,N_17124);
or U18055 (N_18055,N_16008,N_16380);
nand U18056 (N_18056,N_15119,N_16537);
and U18057 (N_18057,N_15504,N_16383);
or U18058 (N_18058,N_16194,N_16377);
and U18059 (N_18059,N_15526,N_15081);
or U18060 (N_18060,N_15879,N_17427);
xnor U18061 (N_18061,N_15337,N_15782);
nand U18062 (N_18062,N_15406,N_15867);
nand U18063 (N_18063,N_16840,N_17242);
nor U18064 (N_18064,N_15458,N_16603);
or U18065 (N_18065,N_15212,N_17155);
nor U18066 (N_18066,N_16805,N_16976);
and U18067 (N_18067,N_16282,N_16652);
nor U18068 (N_18068,N_15773,N_15358);
nand U18069 (N_18069,N_17126,N_16639);
and U18070 (N_18070,N_16144,N_15436);
nand U18071 (N_18071,N_16872,N_17481);
and U18072 (N_18072,N_15961,N_15483);
nand U18073 (N_18073,N_15341,N_16335);
xnor U18074 (N_18074,N_15414,N_16503);
or U18075 (N_18075,N_15535,N_15692);
and U18076 (N_18076,N_16657,N_15808);
xnor U18077 (N_18077,N_15625,N_17033);
or U18078 (N_18078,N_16065,N_16901);
or U18079 (N_18079,N_15953,N_15938);
nand U18080 (N_18080,N_17333,N_16885);
or U18081 (N_18081,N_15529,N_16530);
nand U18082 (N_18082,N_16816,N_17133);
nand U18083 (N_18083,N_16943,N_16360);
nor U18084 (N_18084,N_17404,N_15790);
and U18085 (N_18085,N_15971,N_16925);
or U18086 (N_18086,N_16617,N_15132);
and U18087 (N_18087,N_16055,N_17065);
or U18088 (N_18088,N_16529,N_16547);
and U18089 (N_18089,N_16850,N_16116);
nand U18090 (N_18090,N_17448,N_16608);
or U18091 (N_18091,N_15090,N_15336);
and U18092 (N_18092,N_15688,N_15091);
nor U18093 (N_18093,N_16171,N_16717);
nand U18094 (N_18094,N_16539,N_16672);
and U18095 (N_18095,N_16289,N_16244);
or U18096 (N_18096,N_17145,N_16284);
and U18097 (N_18097,N_15315,N_15142);
and U18098 (N_18098,N_17408,N_17246);
nand U18099 (N_18099,N_16685,N_16513);
xnor U18100 (N_18100,N_16471,N_16954);
and U18101 (N_18101,N_15164,N_15114);
or U18102 (N_18102,N_15211,N_16904);
nand U18103 (N_18103,N_15791,N_16691);
and U18104 (N_18104,N_17426,N_16701);
xnor U18105 (N_18105,N_15553,N_16679);
nor U18106 (N_18106,N_16736,N_15005);
or U18107 (N_18107,N_16542,N_16271);
xor U18108 (N_18108,N_15340,N_16995);
xnor U18109 (N_18109,N_15217,N_16301);
or U18110 (N_18110,N_16636,N_17008);
nor U18111 (N_18111,N_15202,N_15382);
and U18112 (N_18112,N_16990,N_16893);
or U18113 (N_18113,N_15675,N_16658);
nor U18114 (N_18114,N_15059,N_15659);
xor U18115 (N_18115,N_15779,N_16436);
and U18116 (N_18116,N_15857,N_16750);
or U18117 (N_18117,N_15038,N_16074);
nand U18118 (N_18118,N_16400,N_16766);
or U18119 (N_18119,N_15290,N_15869);
nand U18120 (N_18120,N_17233,N_16039);
nand U18121 (N_18121,N_15293,N_16499);
nor U18122 (N_18122,N_17231,N_16814);
and U18123 (N_18123,N_16460,N_15335);
nor U18124 (N_18124,N_16177,N_16769);
and U18125 (N_18125,N_15156,N_17205);
nand U18126 (N_18126,N_17209,N_15823);
xor U18127 (N_18127,N_16595,N_15621);
and U18128 (N_18128,N_15704,N_17089);
nor U18129 (N_18129,N_17103,N_16138);
or U18130 (N_18130,N_17238,N_15750);
xnor U18131 (N_18131,N_16115,N_16500);
nand U18132 (N_18132,N_15191,N_16574);
nand U18133 (N_18133,N_17269,N_15007);
xor U18134 (N_18134,N_16060,N_17293);
and U18135 (N_18135,N_16803,N_15584);
or U18136 (N_18136,N_16381,N_15410);
or U18137 (N_18137,N_16034,N_17091);
and U18138 (N_18138,N_15403,N_16362);
nand U18139 (N_18139,N_17132,N_15069);
nor U18140 (N_18140,N_15547,N_15758);
nand U18141 (N_18141,N_16514,N_15495);
and U18142 (N_18142,N_16167,N_17150);
xnor U18143 (N_18143,N_17036,N_16905);
xor U18144 (N_18144,N_15168,N_16045);
and U18145 (N_18145,N_17047,N_16366);
nand U18146 (N_18146,N_15551,N_16853);
xor U18147 (N_18147,N_16024,N_16959);
nand U18148 (N_18148,N_16565,N_17476);
xnor U18149 (N_18149,N_15761,N_15205);
nor U18150 (N_18150,N_16555,N_16656);
xnor U18151 (N_18151,N_16819,N_15917);
and U18152 (N_18152,N_17215,N_16330);
and U18153 (N_18153,N_16159,N_15711);
nor U18154 (N_18154,N_15814,N_15866);
and U18155 (N_18155,N_16247,N_16821);
or U18156 (N_18156,N_15283,N_16649);
nor U18157 (N_18157,N_16100,N_15985);
or U18158 (N_18158,N_17324,N_15457);
nor U18159 (N_18159,N_16916,N_16867);
nor U18160 (N_18160,N_16779,N_15121);
nand U18161 (N_18161,N_16182,N_16770);
nor U18162 (N_18162,N_15269,N_15288);
or U18163 (N_18163,N_15357,N_16013);
or U18164 (N_18164,N_15348,N_15499);
and U18165 (N_18165,N_15473,N_15510);
xnor U18166 (N_18166,N_16292,N_16996);
xnor U18167 (N_18167,N_15708,N_16053);
xnor U18168 (N_18168,N_16813,N_15420);
and U18169 (N_18169,N_16139,N_16710);
nor U18170 (N_18170,N_17354,N_16453);
nor U18171 (N_18171,N_15921,N_15937);
nand U18172 (N_18172,N_15450,N_15371);
or U18173 (N_18173,N_16170,N_15843);
xnor U18174 (N_18174,N_16504,N_17389);
nand U18175 (N_18175,N_16279,N_17270);
nor U18176 (N_18176,N_15769,N_15171);
xor U18177 (N_18177,N_15516,N_16164);
nand U18178 (N_18178,N_17356,N_15877);
nor U18179 (N_18179,N_16261,N_17414);
and U18180 (N_18180,N_17435,N_16903);
nor U18181 (N_18181,N_15110,N_17478);
xnor U18182 (N_18182,N_15469,N_15666);
or U18183 (N_18183,N_16398,N_15143);
nor U18184 (N_18184,N_17159,N_16716);
and U18185 (N_18185,N_16012,N_15317);
and U18186 (N_18186,N_15389,N_17428);
xor U18187 (N_18187,N_16515,N_16771);
and U18188 (N_18188,N_17095,N_16957);
or U18189 (N_18189,N_16729,N_15369);
nor U18190 (N_18190,N_16825,N_17279);
nand U18191 (N_18191,N_17307,N_15590);
or U18192 (N_18192,N_15995,N_15289);
xor U18193 (N_18193,N_15721,N_16030);
and U18194 (N_18194,N_15895,N_15608);
nor U18195 (N_18195,N_15537,N_15193);
xor U18196 (N_18196,N_16297,N_17480);
and U18197 (N_18197,N_17213,N_15844);
xnor U18198 (N_18198,N_15860,N_15463);
xnor U18199 (N_18199,N_15214,N_17160);
nand U18200 (N_18200,N_16382,N_15301);
nand U18201 (N_18201,N_15261,N_16126);
xor U18202 (N_18202,N_15986,N_16960);
nor U18203 (N_18203,N_16793,N_17217);
nand U18204 (N_18204,N_17487,N_15506);
nand U18205 (N_18205,N_15563,N_17082);
or U18206 (N_18206,N_16558,N_16517);
xnor U18207 (N_18207,N_15453,N_15129);
nand U18208 (N_18208,N_15977,N_15230);
and U18209 (N_18209,N_15032,N_15146);
xnor U18210 (N_18210,N_16324,N_15923);
or U18211 (N_18211,N_16224,N_17051);
xnor U18212 (N_18212,N_16274,N_16815);
or U18213 (N_18213,N_15913,N_15674);
nor U18214 (N_18214,N_15699,N_16299);
or U18215 (N_18215,N_15577,N_16125);
xor U18216 (N_18216,N_17191,N_16802);
nor U18217 (N_18217,N_15925,N_15010);
and U18218 (N_18218,N_16950,N_15268);
xor U18219 (N_18219,N_15801,N_16446);
and U18220 (N_18220,N_16176,N_16763);
and U18221 (N_18221,N_17471,N_15170);
nand U18222 (N_18222,N_16680,N_17243);
or U18223 (N_18223,N_15154,N_17306);
nor U18224 (N_18224,N_15006,N_15089);
nand U18225 (N_18225,N_15196,N_15839);
nand U18226 (N_18226,N_16991,N_16186);
nor U18227 (N_18227,N_15354,N_16399);
and U18228 (N_18228,N_17302,N_15630);
nand U18229 (N_18229,N_17325,N_15662);
or U18230 (N_18230,N_15873,N_16187);
and U18231 (N_18231,N_16121,N_16707);
or U18232 (N_18232,N_17434,N_16557);
or U18233 (N_18233,N_17025,N_15803);
xnor U18234 (N_18234,N_16512,N_16120);
or U18235 (N_18235,N_15615,N_15325);
nand U18236 (N_18236,N_15047,N_17479);
xnor U18237 (N_18237,N_16379,N_17105);
and U18238 (N_18238,N_17305,N_16010);
nand U18239 (N_18239,N_16787,N_16873);
and U18240 (N_18240,N_17174,N_15668);
and U18241 (N_18241,N_16669,N_15646);
and U18242 (N_18242,N_17176,N_15783);
and U18243 (N_18243,N_16702,N_15275);
and U18244 (N_18244,N_15314,N_16714);
nor U18245 (N_18245,N_15083,N_16986);
or U18246 (N_18246,N_15633,N_17138);
nor U18247 (N_18247,N_16677,N_15872);
nor U18248 (N_18248,N_17322,N_16902);
nor U18249 (N_18249,N_15080,N_15396);
and U18250 (N_18250,N_15151,N_17020);
or U18251 (N_18251,N_16613,N_15328);
nor U18252 (N_18252,N_15605,N_15759);
nand U18253 (N_18253,N_16792,N_16067);
nand U18254 (N_18254,N_15890,N_17297);
and U18255 (N_18255,N_16172,N_16810);
nor U18256 (N_18256,N_16201,N_15426);
and U18257 (N_18257,N_16409,N_17345);
nor U18258 (N_18258,N_16796,N_15897);
nand U18259 (N_18259,N_15056,N_16666);
or U18260 (N_18260,N_16828,N_17224);
nand U18261 (N_18261,N_15748,N_17328);
or U18262 (N_18262,N_16023,N_16599);
nand U18263 (N_18263,N_15766,N_16111);
nor U18264 (N_18264,N_15019,N_15498);
nor U18265 (N_18265,N_16876,N_17285);
or U18266 (N_18266,N_16265,N_16541);
or U18267 (N_18267,N_15765,N_16896);
nor U18268 (N_18268,N_15430,N_15880);
and U18269 (N_18269,N_16236,N_17141);
nor U18270 (N_18270,N_16082,N_15709);
and U18271 (N_18271,N_16929,N_17096);
nor U18272 (N_18272,N_15952,N_17261);
and U18273 (N_18273,N_16058,N_16890);
and U18274 (N_18274,N_16938,N_16298);
nor U18275 (N_18275,N_17015,N_16020);
nor U18276 (N_18276,N_15555,N_16979);
or U18277 (N_18277,N_16846,N_15667);
or U18278 (N_18278,N_15541,N_17323);
or U18279 (N_18279,N_16762,N_16906);
xor U18280 (N_18280,N_16040,N_15082);
nor U18281 (N_18281,N_15734,N_16953);
or U18282 (N_18282,N_15014,N_15558);
xnor U18283 (N_18283,N_17184,N_15186);
nor U18284 (N_18284,N_15141,N_16046);
nand U18285 (N_18285,N_15309,N_15505);
nor U18286 (N_18286,N_16263,N_15768);
and U18287 (N_18287,N_15077,N_17366);
or U18288 (N_18288,N_16041,N_16774);
xnor U18289 (N_18289,N_16968,N_16384);
nand U18290 (N_18290,N_16150,N_15939);
xnor U18291 (N_18291,N_17107,N_15000);
or U18292 (N_18292,N_15051,N_16489);
nor U18293 (N_18293,N_15451,N_16464);
nor U18294 (N_18294,N_15313,N_17464);
and U18295 (N_18295,N_16773,N_15853);
xor U18296 (N_18296,N_16927,N_15582);
and U18297 (N_18297,N_16245,N_15169);
and U18298 (N_18298,N_15640,N_16883);
and U18299 (N_18299,N_16036,N_16783);
nand U18300 (N_18300,N_16434,N_15180);
and U18301 (N_18301,N_16272,N_15346);
nor U18302 (N_18302,N_16647,N_15298);
nand U18303 (N_18303,N_15998,N_17329);
xnor U18304 (N_18304,N_16248,N_15710);
or U18305 (N_18305,N_16482,N_15514);
or U18306 (N_18306,N_15567,N_15429);
xnor U18307 (N_18307,N_15851,N_15775);
and U18308 (N_18308,N_17347,N_17290);
and U18309 (N_18309,N_17430,N_17057);
nor U18310 (N_18310,N_16147,N_16744);
nand U18311 (N_18311,N_17158,N_16728);
and U18312 (N_18312,N_15329,N_15455);
or U18313 (N_18313,N_16516,N_16106);
nor U18314 (N_18314,N_17058,N_16619);
nand U18315 (N_18315,N_16033,N_16935);
or U18316 (N_18316,N_16208,N_16849);
and U18317 (N_18317,N_15448,N_16215);
nor U18318 (N_18318,N_16109,N_15338);
nor U18319 (N_18319,N_15462,N_16443);
nand U18320 (N_18320,N_17129,N_16449);
nand U18321 (N_18321,N_16220,N_16267);
and U18322 (N_18322,N_16662,N_15885);
nand U18323 (N_18323,N_17273,N_16506);
xor U18324 (N_18324,N_15057,N_15277);
nand U18325 (N_18325,N_15227,N_15546);
or U18326 (N_18326,N_16238,N_15157);
and U18327 (N_18327,N_15316,N_15291);
or U18328 (N_18328,N_15932,N_15182);
xnor U18329 (N_18329,N_17067,N_17339);
xnor U18330 (N_18330,N_17420,N_15295);
and U18331 (N_18331,N_15962,N_17137);
and U18332 (N_18332,N_15991,N_15959);
and U18333 (N_18333,N_16623,N_16231);
and U18334 (N_18334,N_16311,N_16933);
nand U18335 (N_18335,N_15427,N_15035);
and U18336 (N_18336,N_15265,N_15651);
nor U18337 (N_18337,N_16961,N_16191);
xnor U18338 (N_18338,N_16232,N_15282);
nor U18339 (N_18339,N_15706,N_16651);
or U18340 (N_18340,N_16424,N_16866);
nand U18341 (N_18341,N_16178,N_17040);
xnor U18342 (N_18342,N_15098,N_16615);
and U18343 (N_18343,N_16900,N_15849);
and U18344 (N_18344,N_15326,N_15223);
xor U18345 (N_18345,N_15502,N_15702);
xnor U18346 (N_18346,N_15162,N_15122);
nand U18347 (N_18347,N_17288,N_16348);
nand U18348 (N_18348,N_16551,N_15496);
nor U18349 (N_18349,N_17225,N_17026);
xor U18350 (N_18350,N_17401,N_16195);
nand U18351 (N_18351,N_17021,N_16105);
or U18352 (N_18352,N_16412,N_15237);
nor U18353 (N_18353,N_16000,N_16016);
or U18354 (N_18354,N_16752,N_16661);
nand U18355 (N_18355,N_16497,N_17318);
nand U18356 (N_18356,N_15618,N_15398);
and U18357 (N_18357,N_15644,N_15373);
or U18358 (N_18358,N_16981,N_15022);
nor U18359 (N_18359,N_17364,N_16475);
nand U18360 (N_18360,N_15395,N_15816);
nand U18361 (N_18361,N_16767,N_15163);
or U18362 (N_18362,N_15722,N_15581);
xnor U18363 (N_18363,N_17467,N_15909);
nor U18364 (N_18364,N_15770,N_15624);
or U18365 (N_18365,N_16425,N_15267);
nand U18366 (N_18366,N_16664,N_16637);
and U18367 (N_18367,N_17278,N_16884);
nor U18368 (N_18368,N_15627,N_17062);
nand U18369 (N_18369,N_16955,N_16462);
xor U18370 (N_18370,N_16353,N_15094);
xor U18371 (N_18371,N_15725,N_17399);
and U18372 (N_18372,N_15837,N_15809);
nand U18373 (N_18373,N_16393,N_16533);
nor U18374 (N_18374,N_16072,N_16635);
or U18375 (N_18375,N_16994,N_16369);
xor U18376 (N_18376,N_17445,N_15855);
nor U18377 (N_18377,N_15686,N_15241);
nor U18378 (N_18378,N_16485,N_15075);
or U18379 (N_18379,N_16087,N_15767);
xnor U18380 (N_18380,N_15745,N_15088);
nor U18381 (N_18381,N_17101,N_16924);
or U18382 (N_18382,N_16110,N_16782);
nand U18383 (N_18383,N_16180,N_16407);
nand U18384 (N_18384,N_15521,N_16888);
and U18385 (N_18385,N_16280,N_15772);
nand U18386 (N_18386,N_16025,N_15647);
or U18387 (N_18387,N_15144,N_15053);
nand U18388 (N_18388,N_16312,N_15562);
nand U18389 (N_18389,N_16394,N_15351);
nor U18390 (N_18390,N_16859,N_15432);
nand U18391 (N_18391,N_16339,N_17195);
nor U18392 (N_18392,N_16376,N_16571);
xor U18393 (N_18393,N_15531,N_15687);
or U18394 (N_18394,N_16879,N_15935);
xnor U18395 (N_18395,N_15883,N_17182);
nor U18396 (N_18396,N_16474,N_16942);
nor U18397 (N_18397,N_15323,N_15372);
xnor U18398 (N_18398,N_15731,N_16842);
or U18399 (N_18399,N_15271,N_15994);
nor U18400 (N_18400,N_17227,N_15108);
nor U18401 (N_18401,N_15135,N_16562);
nor U18402 (N_18402,N_16189,N_15384);
xnor U18403 (N_18403,N_15517,N_16080);
nor U18404 (N_18404,N_16077,N_16689);
xor U18405 (N_18405,N_15476,N_15754);
xor U18406 (N_18406,N_15086,N_15691);
xor U18407 (N_18407,N_16653,N_15560);
and U18408 (N_18408,N_16202,N_16569);
or U18409 (N_18409,N_15112,N_17119);
xnor U18410 (N_18410,N_15391,N_17415);
nor U18411 (N_18411,N_16519,N_15365);
xnor U18412 (N_18412,N_16420,N_16001);
or U18413 (N_18413,N_16841,N_16094);
nor U18414 (N_18414,N_15518,N_17152);
nor U18415 (N_18415,N_15931,N_16862);
and U18416 (N_18416,N_16625,N_15347);
or U18417 (N_18417,N_15490,N_15940);
or U18418 (N_18418,N_16809,N_15863);
or U18419 (N_18419,N_17180,N_15670);
or U18420 (N_18420,N_15185,N_16350);
nor U18421 (N_18421,N_16032,N_17219);
and U18422 (N_18422,N_16408,N_15942);
nand U18423 (N_18423,N_17175,N_15101);
nor U18424 (N_18424,N_15755,N_15838);
and U18425 (N_18425,N_15996,N_15274);
nand U18426 (N_18426,N_15370,N_17032);
nand U18427 (N_18427,N_17303,N_17085);
and U18428 (N_18428,N_17259,N_15489);
xnor U18429 (N_18429,N_16936,N_15218);
or U18430 (N_18430,N_17421,N_17121);
nand U18431 (N_18431,N_15746,N_15865);
or U18432 (N_18432,N_16538,N_15399);
nor U18433 (N_18433,N_17335,N_16014);
and U18434 (N_18434,N_16654,N_15720);
or U18435 (N_18435,N_15488,N_15589);
or U18436 (N_18436,N_16560,N_15979);
nand U18437 (N_18437,N_16494,N_15222);
xnor U18438 (N_18438,N_17204,N_16256);
and U18439 (N_18439,N_15830,N_15366);
and U18440 (N_18440,N_15825,N_15149);
xor U18441 (N_18441,N_17495,N_15778);
xnor U18442 (N_18442,N_16587,N_16650);
nand U18443 (N_18443,N_16785,N_17494);
nand U18444 (N_18444,N_16323,N_17011);
nand U18445 (N_18445,N_17214,N_15648);
and U18446 (N_18446,N_15240,N_17357);
and U18447 (N_18447,N_17028,N_15208);
nand U18448 (N_18448,N_15064,N_15574);
nor U18449 (N_18449,N_16801,N_16435);
and U18450 (N_18450,N_17143,N_15201);
or U18451 (N_18451,N_17110,N_16528);
nor U18452 (N_18452,N_15920,N_16952);
or U18453 (N_18453,N_15785,N_15286);
xor U18454 (N_18454,N_15452,N_17080);
nor U18455 (N_18455,N_16740,N_16341);
or U18456 (N_18456,N_15822,N_16287);
xnor U18457 (N_18457,N_17381,N_15297);
or U18458 (N_18458,N_16975,N_16671);
and U18459 (N_18459,N_16709,N_16406);
nor U18460 (N_18460,N_17358,N_15719);
nand U18461 (N_18461,N_15292,N_15846);
xor U18462 (N_18462,N_16314,N_16214);
nand U18463 (N_18463,N_15009,N_15106);
nand U18464 (N_18464,N_16003,N_15087);
and U18465 (N_18465,N_16364,N_16811);
nor U18466 (N_18466,N_17368,N_17489);
xor U18467 (N_18467,N_15494,N_15564);
nor U18468 (N_18468,N_16354,N_15552);
nor U18469 (N_18469,N_17193,N_15165);
or U18470 (N_18470,N_16432,N_17071);
xnor U18471 (N_18471,N_16663,N_16071);
or U18472 (N_18472,N_16437,N_17060);
or U18473 (N_18473,N_15394,N_15705);
xor U18474 (N_18474,N_17054,N_15359);
nor U18475 (N_18475,N_16797,N_15933);
xor U18476 (N_18476,N_15609,N_16321);
nor U18477 (N_18477,N_16463,N_17197);
nor U18478 (N_18478,N_17043,N_16505);
or U18479 (N_18479,N_16206,N_15461);
and U18480 (N_18480,N_15318,N_16484);
nor U18481 (N_18481,N_15576,N_16501);
nand U18482 (N_18482,N_17258,N_16104);
or U18483 (N_18483,N_16237,N_15367);
nor U18484 (N_18484,N_17281,N_16262);
and U18485 (N_18485,N_16174,N_15639);
and U18486 (N_18486,N_15550,N_15967);
nor U18487 (N_18487,N_16385,N_17108);
and U18488 (N_18488,N_16388,N_15470);
nand U18489 (N_18489,N_16473,N_16331);
xor U18490 (N_18490,N_15150,N_15515);
nand U18491 (N_18491,N_16718,N_15965);
xor U18492 (N_18492,N_15278,N_17308);
and U18493 (N_18493,N_16078,N_16601);
or U18494 (N_18494,N_15244,N_17039);
and U18495 (N_18495,N_15792,N_15031);
or U18496 (N_18496,N_16607,N_15665);
nor U18497 (N_18497,N_16140,N_16304);
or U18498 (N_18498,N_16898,N_16645);
nor U18499 (N_18499,N_16308,N_16543);
nor U18500 (N_18500,N_15598,N_15954);
nand U18501 (N_18501,N_16051,N_15680);
and U18502 (N_18502,N_17268,N_17275);
or U18503 (N_18503,N_15918,N_17073);
and U18504 (N_18504,N_15060,N_16097);
nand U18505 (N_18505,N_15789,N_17451);
nand U18506 (N_18506,N_17022,N_15225);
xor U18507 (N_18507,N_15023,N_15930);
nor U18508 (N_18508,N_16553,N_17440);
or U18509 (N_18509,N_15254,N_15245);
xor U18510 (N_18510,N_15250,N_17016);
or U18511 (N_18511,N_15167,N_15828);
nor U18512 (N_18512,N_15061,N_15138);
nand U18513 (N_18513,N_15025,N_16277);
nand U18514 (N_18514,N_16117,N_16520);
or U18515 (N_18515,N_17398,N_16634);
and U18516 (N_18516,N_16405,N_16346);
xor U18517 (N_18517,N_17283,N_15471);
and U18518 (N_18518,N_15404,N_15342);
and U18519 (N_18519,N_16725,N_16293);
xor U18520 (N_18520,N_16370,N_17319);
nor U18521 (N_18521,N_17187,N_16865);
or U18522 (N_18522,N_16021,N_15629);
xor U18523 (N_18523,N_15966,N_17003);
and U18524 (N_18524,N_16751,N_15673);
nand U18525 (N_18525,N_16880,N_16211);
or U18526 (N_18526,N_15528,N_17397);
nand U18527 (N_18527,N_15520,N_16930);
xor U18528 (N_18528,N_15908,N_16118);
nor U18529 (N_18529,N_15422,N_15898);
xor U18530 (N_18530,N_17386,N_17013);
nand U18531 (N_18531,N_16493,N_17210);
nand U18532 (N_18532,N_17265,N_15018);
xnor U18533 (N_18533,N_17326,N_17330);
and U18534 (N_18534,N_17344,N_16568);
xor U18535 (N_18535,N_15997,N_16518);
and U18536 (N_18536,N_16427,N_16838);
nand U18537 (N_18537,N_15434,N_16101);
or U18538 (N_18538,N_17114,N_16169);
nor U18539 (N_18539,N_17254,N_16073);
and U18540 (N_18540,N_16525,N_16511);
or U18541 (N_18541,N_15780,N_16611);
nand U18542 (N_18542,N_16593,N_17202);
and U18543 (N_18543,N_17153,N_17287);
nor U18544 (N_18544,N_16618,N_15037);
nand U18545 (N_18545,N_16536,N_16578);
and U18546 (N_18546,N_17405,N_16684);
nor U18547 (N_18547,N_15729,N_15684);
xnor U18548 (N_18548,N_15707,N_16162);
xor U18549 (N_18549,N_15033,N_16941);
xor U18550 (N_18550,N_16676,N_16054);
nor U18551 (N_18551,N_15400,N_17023);
or U18552 (N_18552,N_16502,N_15549);
nand U18553 (N_18553,N_16442,N_15764);
nor U18554 (N_18554,N_15557,N_16066);
nand U18555 (N_18555,N_16326,N_15198);
nand U18556 (N_18556,N_15042,N_16495);
or U18557 (N_18557,N_17009,N_16721);
and U18558 (N_18558,N_16098,N_16882);
xor U18559 (N_18559,N_17390,N_16848);
or U18560 (N_18560,N_15234,N_16581);
xnor U18561 (N_18561,N_15068,N_17439);
and U18562 (N_18562,N_16891,N_16113);
nand U18563 (N_18563,N_16239,N_17320);
and U18564 (N_18564,N_17048,N_16230);
and U18565 (N_18565,N_15565,N_16183);
nor U18566 (N_18566,N_15041,N_15507);
xor U18567 (N_18567,N_15859,N_15891);
nand U18568 (N_18568,N_15958,N_15352);
or U18569 (N_18569,N_15566,N_17496);
nand U18570 (N_18570,N_15964,N_16588);
or U18571 (N_18571,N_15305,N_16522);
nand U18572 (N_18572,N_17232,N_17359);
and U18573 (N_18573,N_15948,N_16347);
nor U18574 (N_18574,N_17256,N_16062);
or U18575 (N_18575,N_15726,N_17077);
or U18576 (N_18576,N_16338,N_16264);
nand U18577 (N_18577,N_15868,N_17128);
and U18578 (N_18578,N_17423,N_17409);
nor U18579 (N_18579,N_16737,N_15444);
xor U18580 (N_18580,N_15884,N_16091);
nor U18581 (N_18581,N_15058,N_16163);
xnor U18582 (N_18582,N_15071,N_15439);
nand U18583 (N_18583,N_15417,N_15637);
or U18584 (N_18584,N_15027,N_15249);
xor U18585 (N_18585,N_15353,N_15793);
and U18586 (N_18586,N_16926,N_15055);
nor U18587 (N_18587,N_16457,N_15653);
nand U18588 (N_18588,N_16911,N_17078);
or U18589 (N_18589,N_16642,N_17049);
nor U18590 (N_18590,N_17196,N_16843);
xnor U18591 (N_18591,N_15159,N_15207);
and U18592 (N_18592,N_16583,N_15219);
and U18593 (N_18593,N_15364,N_15724);
nand U18594 (N_18594,N_17001,N_17396);
or U18595 (N_18595,N_16621,N_17188);
nor U18596 (N_18596,N_17447,N_16255);
and U18597 (N_18597,N_16249,N_17262);
nand U18598 (N_18598,N_15148,N_15379);
or U18599 (N_18599,N_15587,N_17402);
nand U18600 (N_18600,N_16755,N_16151);
nand U18601 (N_18601,N_17064,N_16753);
xnor U18602 (N_18602,N_15690,N_15361);
nor U18603 (N_18603,N_16590,N_16776);
xnor U18604 (N_18604,N_15915,N_15841);
xor U18605 (N_18605,N_16951,N_15421);
xnor U18606 (N_18606,N_15441,N_15021);
xnor U18607 (N_18607,N_16285,N_16392);
xnor U18608 (N_18608,N_15611,N_16478);
and U18609 (N_18609,N_15355,N_16732);
nor U18610 (N_18610,N_16575,N_16644);
nor U18611 (N_18611,N_16550,N_17280);
nor U18612 (N_18612,N_15392,N_16690);
xor U18613 (N_18613,N_15302,N_16738);
xor U18614 (N_18614,N_15712,N_16858);
or U18615 (N_18615,N_15743,N_16632);
nand U18616 (N_18616,N_16610,N_16184);
or U18617 (N_18617,N_15246,N_15386);
nand U18618 (N_18618,N_15573,N_16337);
nand U18619 (N_18619,N_15263,N_16168);
or U18620 (N_18620,N_16305,N_15656);
xor U18621 (N_18621,N_17171,N_16748);
xor U18622 (N_18622,N_16546,N_16912);
or U18623 (N_18623,N_15747,N_16705);
or U18624 (N_18624,N_16322,N_16141);
or U18625 (N_18625,N_15934,N_15194);
nor U18626 (N_18626,N_16722,N_15024);
or U18627 (N_18627,N_17192,N_17004);
nand U18628 (N_18628,N_16155,N_17162);
and U18629 (N_18629,N_17186,N_17343);
xor U18630 (N_18630,N_16158,N_15533);
nand U18631 (N_18631,N_15523,N_17235);
xnor U18632 (N_18632,N_15134,N_17429);
or U18633 (N_18633,N_16329,N_16133);
and U18634 (N_18634,N_15831,N_17087);
xor U18635 (N_18635,N_16268,N_16373);
and U18636 (N_18636,N_17201,N_16472);
and U18637 (N_18637,N_16673,N_15161);
and U18638 (N_18638,N_15356,N_16972);
and U18639 (N_18639,N_15714,N_16527);
or U18640 (N_18640,N_15840,N_15113);
xnor U18641 (N_18641,N_16757,N_15029);
and U18642 (N_18642,N_15701,N_17074);
nor U18643 (N_18643,N_16061,N_16363);
nand U18644 (N_18644,N_15622,N_15464);
and U18645 (N_18645,N_15810,N_17486);
xnor U18646 (N_18646,N_16122,N_16758);
nand U18647 (N_18647,N_15886,N_16997);
and U18648 (N_18648,N_17484,N_16622);
xnor U18649 (N_18649,N_15294,N_16342);
xnor U18650 (N_18650,N_16165,N_16946);
nor U18651 (N_18651,N_17431,N_17198);
nand U18652 (N_18652,N_16352,N_16327);
or U18653 (N_18653,N_16845,N_15936);
nor U18654 (N_18654,N_16227,N_15896);
and U18655 (N_18655,N_15311,N_15287);
nand U18656 (N_18656,N_15999,N_15276);
or U18657 (N_18657,N_15475,N_15067);
and U18658 (N_18658,N_15797,N_16860);
and U18659 (N_18659,N_16210,N_15530);
or U18660 (N_18660,N_17169,N_16746);
nor U18661 (N_18661,N_15228,N_15700);
and U18662 (N_18662,N_16735,N_17116);
and U18663 (N_18663,N_17122,N_15685);
nand U18664 (N_18664,N_16969,N_15004);
xor U18665 (N_18665,N_16368,N_17375);
xnor U18666 (N_18666,N_16897,N_15963);
nor U18667 (N_18667,N_17456,N_15540);
xor U18668 (N_18668,N_16303,N_16135);
and U18669 (N_18669,N_16099,N_15443);
or U18670 (N_18670,N_15260,N_17228);
xor U18671 (N_18671,N_16711,N_17436);
and U18672 (N_18672,N_16052,N_17240);
xnor U18673 (N_18673,N_17050,N_16988);
nor U18674 (N_18674,N_17147,N_15327);
or U18675 (N_18675,N_16589,N_16949);
and U18676 (N_18676,N_15570,N_15118);
nand U18677 (N_18677,N_16918,N_15501);
or U18678 (N_18678,N_16914,N_15192);
or U18679 (N_18679,N_16102,N_17056);
nor U18680 (N_18680,N_16576,N_15888);
xnor U18681 (N_18681,N_16869,N_17034);
xnor U18682 (N_18682,N_15416,N_17163);
nand U18683 (N_18683,N_15620,N_17207);
nand U18684 (N_18684,N_17351,N_16142);
and U18685 (N_18685,N_16160,N_16934);
or U18686 (N_18686,N_16944,N_15619);
nand U18687 (N_18687,N_15903,N_16839);
xor U18688 (N_18688,N_17468,N_15273);
nor U18689 (N_18689,N_15321,N_16367);
xnor U18690 (N_18690,N_16857,N_15960);
and U18691 (N_18691,N_16235,N_17059);
xnor U18692 (N_18692,N_17294,N_16945);
nor U18693 (N_18693,N_17369,N_16090);
and U18694 (N_18694,N_16667,N_16313);
or U18695 (N_18695,N_16602,N_16447);
xor U18696 (N_18696,N_16962,N_16414);
xor U18697 (N_18697,N_15559,N_15571);
nor U18698 (N_18698,N_16616,N_16203);
xor U18699 (N_18699,N_16050,N_16070);
nand U18700 (N_18700,N_16573,N_17053);
nor U18701 (N_18701,N_15299,N_17151);
or U18702 (N_18702,N_15073,N_15012);
nor U18703 (N_18703,N_15580,N_17374);
nand U18704 (N_18704,N_16241,N_15074);
nor U18705 (N_18705,N_16015,N_15123);
or U18706 (N_18706,N_16219,N_17092);
and U18707 (N_18707,N_16855,N_16704);
and U18708 (N_18708,N_16085,N_17392);
and U18709 (N_18709,N_16775,N_15200);
xnor U18710 (N_18710,N_15480,N_15796);
and U18711 (N_18711,N_15126,N_15285);
and U18712 (N_18712,N_15484,N_15757);
or U18713 (N_18713,N_16103,N_17168);
and U18714 (N_18714,N_15070,N_15864);
or U18715 (N_18715,N_16604,N_16837);
xnor U18716 (N_18716,N_17292,N_17299);
nor U18717 (N_18717,N_16540,N_15279);
nand U18718 (N_18718,N_15231,N_15482);
xor U18719 (N_18719,N_16660,N_17406);
and U18720 (N_18720,N_16461,N_15924);
xor U18721 (N_18721,N_15266,N_15813);
nand U18722 (N_18722,N_15424,N_17422);
and U18723 (N_18723,N_17099,N_15054);
nor U18724 (N_18724,N_16584,N_17266);
and U18725 (N_18725,N_15030,N_16889);
nor U18726 (N_18726,N_16864,N_15616);
xnor U18727 (N_18727,N_16270,N_15349);
xor U18728 (N_18728,N_16956,N_16706);
xnor U18729 (N_18729,N_15795,N_15512);
or U18730 (N_18730,N_16316,N_15256);
and U18731 (N_18731,N_15003,N_16760);
and U18732 (N_18732,N_15350,N_17419);
or U18733 (N_18733,N_15771,N_15878);
nor U18734 (N_18734,N_15280,N_16646);
nand U18735 (N_18735,N_15130,N_17139);
and U18736 (N_18736,N_15834,N_17017);
and U18737 (N_18737,N_17388,N_16605);
xor U18738 (N_18738,N_15833,N_16724);
xnor U18739 (N_18739,N_17136,N_15904);
xnor U18740 (N_18740,N_15679,N_15696);
nand U18741 (N_18741,N_15804,N_15467);
xnor U18742 (N_18742,N_15905,N_15820);
xor U18743 (N_18743,N_15175,N_15601);
or U18744 (N_18744,N_15308,N_16833);
nor U18745 (N_18745,N_17066,N_16987);
or U18746 (N_18746,N_17317,N_17157);
or U18747 (N_18747,N_17418,N_15950);
nand U18748 (N_18748,N_15431,N_15052);
or U18749 (N_18749,N_15871,N_16068);
or U18750 (N_18750,N_15059,N_16856);
nor U18751 (N_18751,N_17458,N_15661);
nor U18752 (N_18752,N_15966,N_16654);
and U18753 (N_18753,N_15126,N_16042);
nor U18754 (N_18754,N_17242,N_16754);
xor U18755 (N_18755,N_15068,N_17371);
xor U18756 (N_18756,N_16450,N_15461);
or U18757 (N_18757,N_15163,N_17084);
nor U18758 (N_18758,N_15766,N_15997);
or U18759 (N_18759,N_15717,N_16176);
or U18760 (N_18760,N_17144,N_15998);
nor U18761 (N_18761,N_17320,N_16491);
nor U18762 (N_18762,N_15118,N_16552);
or U18763 (N_18763,N_15595,N_15647);
or U18764 (N_18764,N_16987,N_16731);
nand U18765 (N_18765,N_16016,N_16611);
nor U18766 (N_18766,N_15371,N_15143);
and U18767 (N_18767,N_16293,N_16630);
and U18768 (N_18768,N_15046,N_16605);
xor U18769 (N_18769,N_15344,N_16616);
xnor U18770 (N_18770,N_16116,N_16639);
xnor U18771 (N_18771,N_16942,N_15511);
or U18772 (N_18772,N_15652,N_16568);
nand U18773 (N_18773,N_15422,N_15168);
and U18774 (N_18774,N_15895,N_17380);
nand U18775 (N_18775,N_16929,N_16678);
nor U18776 (N_18776,N_16876,N_16027);
nor U18777 (N_18777,N_15387,N_16973);
nor U18778 (N_18778,N_15920,N_16721);
and U18779 (N_18779,N_15439,N_15273);
xor U18780 (N_18780,N_15006,N_16457);
or U18781 (N_18781,N_16529,N_16783);
or U18782 (N_18782,N_15254,N_16680);
nor U18783 (N_18783,N_16253,N_15126);
or U18784 (N_18784,N_15777,N_16337);
nor U18785 (N_18785,N_15563,N_15119);
nand U18786 (N_18786,N_16066,N_16853);
xor U18787 (N_18787,N_16245,N_16721);
and U18788 (N_18788,N_17079,N_16396);
nor U18789 (N_18789,N_16825,N_15704);
xor U18790 (N_18790,N_16185,N_15342);
and U18791 (N_18791,N_15048,N_15777);
xor U18792 (N_18792,N_15882,N_17358);
xnor U18793 (N_18793,N_15368,N_15643);
xnor U18794 (N_18794,N_16510,N_16875);
and U18795 (N_18795,N_16175,N_16553);
nor U18796 (N_18796,N_17420,N_15782);
nand U18797 (N_18797,N_16733,N_16680);
and U18798 (N_18798,N_16355,N_16795);
or U18799 (N_18799,N_15554,N_16723);
nor U18800 (N_18800,N_17051,N_16325);
and U18801 (N_18801,N_15374,N_17064);
or U18802 (N_18802,N_17275,N_15055);
nand U18803 (N_18803,N_17290,N_15015);
nor U18804 (N_18804,N_17074,N_15270);
and U18805 (N_18805,N_15420,N_15708);
nor U18806 (N_18806,N_16490,N_16526);
nor U18807 (N_18807,N_15890,N_16123);
nor U18808 (N_18808,N_15619,N_15636);
and U18809 (N_18809,N_15127,N_15538);
or U18810 (N_18810,N_15234,N_16372);
nand U18811 (N_18811,N_16675,N_15356);
nor U18812 (N_18812,N_17175,N_17087);
nor U18813 (N_18813,N_17224,N_15186);
and U18814 (N_18814,N_16831,N_16227);
or U18815 (N_18815,N_15681,N_15635);
nor U18816 (N_18816,N_17275,N_17129);
nor U18817 (N_18817,N_17305,N_16455);
xnor U18818 (N_18818,N_15508,N_17157);
xor U18819 (N_18819,N_15418,N_15992);
nor U18820 (N_18820,N_15622,N_17440);
nor U18821 (N_18821,N_16446,N_15227);
nor U18822 (N_18822,N_15501,N_15913);
xnor U18823 (N_18823,N_15593,N_17114);
or U18824 (N_18824,N_15454,N_15372);
nand U18825 (N_18825,N_15957,N_16174);
and U18826 (N_18826,N_15366,N_16886);
nand U18827 (N_18827,N_15606,N_17052);
nor U18828 (N_18828,N_17289,N_16469);
nand U18829 (N_18829,N_15678,N_15304);
and U18830 (N_18830,N_16977,N_15600);
nor U18831 (N_18831,N_16345,N_15758);
xor U18832 (N_18832,N_17314,N_15088);
nor U18833 (N_18833,N_16739,N_16335);
and U18834 (N_18834,N_16204,N_16723);
nand U18835 (N_18835,N_15501,N_15405);
nor U18836 (N_18836,N_16917,N_15706);
or U18837 (N_18837,N_16654,N_16979);
xor U18838 (N_18838,N_17209,N_15562);
nor U18839 (N_18839,N_17248,N_16193);
nand U18840 (N_18840,N_16848,N_15751);
or U18841 (N_18841,N_16714,N_17387);
xor U18842 (N_18842,N_16922,N_15121);
or U18843 (N_18843,N_16571,N_17224);
and U18844 (N_18844,N_16227,N_16572);
xor U18845 (N_18845,N_15694,N_15897);
and U18846 (N_18846,N_15735,N_17000);
and U18847 (N_18847,N_15811,N_17462);
nand U18848 (N_18848,N_15286,N_16383);
xnor U18849 (N_18849,N_17091,N_17002);
nand U18850 (N_18850,N_16026,N_15782);
and U18851 (N_18851,N_17382,N_16887);
xnor U18852 (N_18852,N_16472,N_17233);
nor U18853 (N_18853,N_15143,N_15685);
and U18854 (N_18854,N_16954,N_15349);
nand U18855 (N_18855,N_15934,N_16975);
or U18856 (N_18856,N_16537,N_16575);
and U18857 (N_18857,N_16644,N_16175);
and U18858 (N_18858,N_15898,N_15779);
nor U18859 (N_18859,N_15630,N_15620);
or U18860 (N_18860,N_16814,N_15258);
and U18861 (N_18861,N_16233,N_15888);
and U18862 (N_18862,N_15278,N_15948);
xor U18863 (N_18863,N_15158,N_16251);
nor U18864 (N_18864,N_17276,N_15192);
nor U18865 (N_18865,N_15698,N_15325);
and U18866 (N_18866,N_16312,N_15066);
and U18867 (N_18867,N_17083,N_15535);
nand U18868 (N_18868,N_15681,N_16027);
xor U18869 (N_18869,N_17374,N_15178);
nand U18870 (N_18870,N_15361,N_16124);
nor U18871 (N_18871,N_16271,N_16282);
nor U18872 (N_18872,N_15957,N_16490);
nor U18873 (N_18873,N_16920,N_16205);
xor U18874 (N_18874,N_16928,N_16045);
xor U18875 (N_18875,N_16367,N_15903);
nor U18876 (N_18876,N_15018,N_16565);
nor U18877 (N_18877,N_15500,N_15372);
nor U18878 (N_18878,N_16322,N_17327);
nor U18879 (N_18879,N_16958,N_16969);
or U18880 (N_18880,N_16489,N_15753);
and U18881 (N_18881,N_15972,N_16177);
nor U18882 (N_18882,N_15277,N_16620);
and U18883 (N_18883,N_15333,N_15179);
or U18884 (N_18884,N_15566,N_15541);
nor U18885 (N_18885,N_17299,N_17034);
xor U18886 (N_18886,N_15977,N_16996);
nand U18887 (N_18887,N_15827,N_17222);
nor U18888 (N_18888,N_16166,N_15781);
xnor U18889 (N_18889,N_16803,N_15609);
and U18890 (N_18890,N_15506,N_17363);
or U18891 (N_18891,N_15068,N_17262);
nor U18892 (N_18892,N_16538,N_16107);
xnor U18893 (N_18893,N_15797,N_16061);
nor U18894 (N_18894,N_15031,N_16075);
or U18895 (N_18895,N_17104,N_15363);
or U18896 (N_18896,N_15596,N_16476);
and U18897 (N_18897,N_15085,N_15434);
and U18898 (N_18898,N_16383,N_15321);
and U18899 (N_18899,N_15346,N_16534);
xnor U18900 (N_18900,N_15332,N_15059);
xnor U18901 (N_18901,N_16791,N_16066);
nand U18902 (N_18902,N_17392,N_17116);
or U18903 (N_18903,N_15276,N_15720);
nand U18904 (N_18904,N_15120,N_15255);
nor U18905 (N_18905,N_16944,N_16952);
and U18906 (N_18906,N_17045,N_16846);
nor U18907 (N_18907,N_15289,N_16268);
or U18908 (N_18908,N_16943,N_16308);
nor U18909 (N_18909,N_17190,N_16355);
and U18910 (N_18910,N_17220,N_17222);
nand U18911 (N_18911,N_16239,N_16947);
xnor U18912 (N_18912,N_16941,N_17412);
nor U18913 (N_18913,N_15206,N_16639);
xor U18914 (N_18914,N_15413,N_16556);
nand U18915 (N_18915,N_16876,N_17118);
nand U18916 (N_18916,N_15234,N_15946);
nand U18917 (N_18917,N_17222,N_15980);
or U18918 (N_18918,N_15590,N_15160);
or U18919 (N_18919,N_16592,N_16372);
nand U18920 (N_18920,N_16806,N_17276);
nand U18921 (N_18921,N_15060,N_15321);
nand U18922 (N_18922,N_17200,N_16324);
xnor U18923 (N_18923,N_15859,N_17331);
or U18924 (N_18924,N_15262,N_17150);
and U18925 (N_18925,N_15365,N_15723);
nor U18926 (N_18926,N_15156,N_17496);
or U18927 (N_18927,N_15872,N_17115);
nand U18928 (N_18928,N_15634,N_16826);
xnor U18929 (N_18929,N_16086,N_16480);
xor U18930 (N_18930,N_15520,N_16426);
nand U18931 (N_18931,N_16516,N_15428);
nor U18932 (N_18932,N_15046,N_15240);
nor U18933 (N_18933,N_15063,N_16608);
and U18934 (N_18934,N_16180,N_16925);
nand U18935 (N_18935,N_15946,N_16728);
nand U18936 (N_18936,N_17325,N_16390);
or U18937 (N_18937,N_15803,N_16673);
xnor U18938 (N_18938,N_16698,N_16546);
nand U18939 (N_18939,N_17161,N_15835);
nor U18940 (N_18940,N_16977,N_16194);
and U18941 (N_18941,N_15579,N_16205);
nand U18942 (N_18942,N_15134,N_16372);
nand U18943 (N_18943,N_17414,N_16089);
nand U18944 (N_18944,N_16867,N_16141);
or U18945 (N_18945,N_15538,N_15056);
and U18946 (N_18946,N_15126,N_16911);
and U18947 (N_18947,N_16967,N_16058);
and U18948 (N_18948,N_16316,N_17046);
xor U18949 (N_18949,N_16179,N_16591);
and U18950 (N_18950,N_17005,N_16514);
nor U18951 (N_18951,N_15974,N_15595);
nor U18952 (N_18952,N_15433,N_17290);
xnor U18953 (N_18953,N_15845,N_17389);
nand U18954 (N_18954,N_15702,N_15736);
nand U18955 (N_18955,N_15842,N_15171);
xnor U18956 (N_18956,N_16815,N_17000);
nor U18957 (N_18957,N_15507,N_16658);
xnor U18958 (N_18958,N_15039,N_15572);
xnor U18959 (N_18959,N_15255,N_16565);
xnor U18960 (N_18960,N_15354,N_16609);
or U18961 (N_18961,N_16563,N_15298);
nand U18962 (N_18962,N_17384,N_17086);
nand U18963 (N_18963,N_16884,N_17211);
or U18964 (N_18964,N_15462,N_16739);
and U18965 (N_18965,N_15216,N_16191);
and U18966 (N_18966,N_15530,N_16143);
nor U18967 (N_18967,N_15666,N_16153);
or U18968 (N_18968,N_16208,N_16618);
and U18969 (N_18969,N_16799,N_16738);
and U18970 (N_18970,N_15823,N_16796);
xor U18971 (N_18971,N_17456,N_16513);
or U18972 (N_18972,N_16423,N_16841);
nand U18973 (N_18973,N_15653,N_16147);
xor U18974 (N_18974,N_15536,N_15866);
xor U18975 (N_18975,N_17346,N_16535);
xnor U18976 (N_18976,N_17210,N_16354);
xnor U18977 (N_18977,N_15496,N_15364);
and U18978 (N_18978,N_15942,N_16409);
xor U18979 (N_18979,N_15580,N_16631);
or U18980 (N_18980,N_15428,N_15261);
or U18981 (N_18981,N_16520,N_16940);
nor U18982 (N_18982,N_16539,N_17094);
and U18983 (N_18983,N_15589,N_15769);
or U18984 (N_18984,N_15220,N_17093);
xor U18985 (N_18985,N_15471,N_15179);
nor U18986 (N_18986,N_15837,N_16540);
xnor U18987 (N_18987,N_16935,N_16115);
xnor U18988 (N_18988,N_15822,N_15674);
nand U18989 (N_18989,N_15929,N_16828);
xor U18990 (N_18990,N_16634,N_15828);
or U18991 (N_18991,N_16287,N_16615);
xor U18992 (N_18992,N_15633,N_15190);
nor U18993 (N_18993,N_16190,N_16288);
or U18994 (N_18994,N_15454,N_15878);
xnor U18995 (N_18995,N_16256,N_15854);
nand U18996 (N_18996,N_15717,N_16384);
or U18997 (N_18997,N_15784,N_17370);
nand U18998 (N_18998,N_16177,N_16478);
xnor U18999 (N_18999,N_16192,N_17036);
nand U19000 (N_19000,N_17051,N_15175);
or U19001 (N_19001,N_15141,N_16172);
nand U19002 (N_19002,N_17360,N_16963);
and U19003 (N_19003,N_16652,N_16214);
nand U19004 (N_19004,N_16113,N_17404);
xor U19005 (N_19005,N_15513,N_16006);
nand U19006 (N_19006,N_17235,N_16713);
nor U19007 (N_19007,N_16079,N_16174);
or U19008 (N_19008,N_15207,N_16180);
or U19009 (N_19009,N_16530,N_17094);
xor U19010 (N_19010,N_16577,N_15227);
nor U19011 (N_19011,N_15243,N_16793);
nor U19012 (N_19012,N_17362,N_16439);
nand U19013 (N_19013,N_15890,N_15249);
nor U19014 (N_19014,N_15418,N_15479);
or U19015 (N_19015,N_16835,N_16416);
nor U19016 (N_19016,N_15485,N_15524);
nor U19017 (N_19017,N_16687,N_16464);
and U19018 (N_19018,N_16636,N_15282);
nand U19019 (N_19019,N_15609,N_16466);
nand U19020 (N_19020,N_16994,N_15669);
nand U19021 (N_19021,N_16237,N_17131);
nand U19022 (N_19022,N_15255,N_16833);
nand U19023 (N_19023,N_15643,N_16369);
nand U19024 (N_19024,N_15663,N_17423);
or U19025 (N_19025,N_16123,N_15122);
and U19026 (N_19026,N_15477,N_15967);
xor U19027 (N_19027,N_16320,N_16706);
xnor U19028 (N_19028,N_17447,N_15122);
and U19029 (N_19029,N_16113,N_15888);
and U19030 (N_19030,N_16190,N_15387);
or U19031 (N_19031,N_17105,N_17332);
nand U19032 (N_19032,N_16487,N_15583);
nor U19033 (N_19033,N_16358,N_17375);
and U19034 (N_19034,N_17476,N_15028);
or U19035 (N_19035,N_16073,N_15624);
or U19036 (N_19036,N_16930,N_17110);
and U19037 (N_19037,N_16491,N_15807);
nor U19038 (N_19038,N_16754,N_16131);
nor U19039 (N_19039,N_15876,N_16825);
and U19040 (N_19040,N_16307,N_17186);
or U19041 (N_19041,N_17095,N_15471);
nand U19042 (N_19042,N_17430,N_16979);
xnor U19043 (N_19043,N_16182,N_16400);
or U19044 (N_19044,N_17266,N_15876);
or U19045 (N_19045,N_15597,N_15764);
or U19046 (N_19046,N_16116,N_15241);
and U19047 (N_19047,N_16820,N_16074);
nor U19048 (N_19048,N_16372,N_16525);
and U19049 (N_19049,N_15035,N_17099);
and U19050 (N_19050,N_16697,N_17337);
and U19051 (N_19051,N_16955,N_15241);
and U19052 (N_19052,N_16865,N_16959);
nand U19053 (N_19053,N_17363,N_17410);
nand U19054 (N_19054,N_16193,N_15773);
xor U19055 (N_19055,N_16415,N_15112);
nor U19056 (N_19056,N_15431,N_16903);
and U19057 (N_19057,N_15137,N_16340);
nor U19058 (N_19058,N_16239,N_15005);
and U19059 (N_19059,N_17076,N_16540);
or U19060 (N_19060,N_16807,N_15967);
xor U19061 (N_19061,N_16649,N_15940);
or U19062 (N_19062,N_15386,N_16078);
xnor U19063 (N_19063,N_16951,N_16436);
and U19064 (N_19064,N_15812,N_17102);
nand U19065 (N_19065,N_15870,N_17371);
nor U19066 (N_19066,N_15436,N_16663);
or U19067 (N_19067,N_16808,N_15936);
nand U19068 (N_19068,N_17162,N_16083);
and U19069 (N_19069,N_15645,N_15886);
nand U19070 (N_19070,N_16529,N_16273);
nor U19071 (N_19071,N_17121,N_16653);
and U19072 (N_19072,N_16574,N_16519);
nor U19073 (N_19073,N_16651,N_17177);
nand U19074 (N_19074,N_16986,N_16533);
or U19075 (N_19075,N_15462,N_17199);
nand U19076 (N_19076,N_15667,N_17074);
and U19077 (N_19077,N_15744,N_16558);
xnor U19078 (N_19078,N_17276,N_17111);
nor U19079 (N_19079,N_16944,N_16696);
xnor U19080 (N_19080,N_17305,N_16957);
and U19081 (N_19081,N_17425,N_15780);
or U19082 (N_19082,N_15338,N_16865);
or U19083 (N_19083,N_15062,N_17453);
or U19084 (N_19084,N_15974,N_16181);
nor U19085 (N_19085,N_15005,N_16225);
xnor U19086 (N_19086,N_15734,N_17341);
and U19087 (N_19087,N_17274,N_15331);
nor U19088 (N_19088,N_16431,N_17297);
and U19089 (N_19089,N_15695,N_15656);
nand U19090 (N_19090,N_15605,N_15481);
nor U19091 (N_19091,N_16140,N_15420);
nand U19092 (N_19092,N_15978,N_16306);
xnor U19093 (N_19093,N_16633,N_16101);
xor U19094 (N_19094,N_16663,N_16668);
nand U19095 (N_19095,N_15046,N_15027);
nor U19096 (N_19096,N_15983,N_16947);
and U19097 (N_19097,N_15747,N_15305);
and U19098 (N_19098,N_16750,N_15694);
nand U19099 (N_19099,N_16169,N_16111);
nor U19100 (N_19100,N_17470,N_16928);
or U19101 (N_19101,N_16439,N_16474);
xnor U19102 (N_19102,N_15857,N_16606);
nand U19103 (N_19103,N_16435,N_16322);
xnor U19104 (N_19104,N_15053,N_16469);
or U19105 (N_19105,N_16960,N_15455);
nor U19106 (N_19106,N_16809,N_15907);
xnor U19107 (N_19107,N_15430,N_17172);
or U19108 (N_19108,N_16482,N_16848);
xnor U19109 (N_19109,N_15570,N_17367);
nor U19110 (N_19110,N_16092,N_16950);
xnor U19111 (N_19111,N_15759,N_16917);
and U19112 (N_19112,N_15842,N_15860);
nor U19113 (N_19113,N_15921,N_17330);
and U19114 (N_19114,N_16170,N_15733);
nand U19115 (N_19115,N_17472,N_16221);
xnor U19116 (N_19116,N_15492,N_16845);
or U19117 (N_19117,N_16659,N_16221);
xnor U19118 (N_19118,N_15939,N_15532);
and U19119 (N_19119,N_17486,N_15314);
and U19120 (N_19120,N_15327,N_16119);
or U19121 (N_19121,N_16779,N_16648);
and U19122 (N_19122,N_16249,N_17204);
nand U19123 (N_19123,N_17384,N_15113);
xor U19124 (N_19124,N_17202,N_15070);
nand U19125 (N_19125,N_15859,N_17222);
nor U19126 (N_19126,N_15710,N_16124);
nand U19127 (N_19127,N_15256,N_16709);
xnor U19128 (N_19128,N_17261,N_17203);
or U19129 (N_19129,N_17023,N_17151);
or U19130 (N_19130,N_17259,N_15865);
xnor U19131 (N_19131,N_17443,N_16597);
and U19132 (N_19132,N_16097,N_16254);
nor U19133 (N_19133,N_16778,N_15786);
nand U19134 (N_19134,N_15815,N_16422);
xor U19135 (N_19135,N_15231,N_15265);
or U19136 (N_19136,N_15315,N_15273);
nor U19137 (N_19137,N_17390,N_16527);
xor U19138 (N_19138,N_16818,N_15862);
and U19139 (N_19139,N_16414,N_16376);
nand U19140 (N_19140,N_15477,N_17102);
and U19141 (N_19141,N_15403,N_16260);
or U19142 (N_19142,N_15465,N_17312);
xor U19143 (N_19143,N_16150,N_15873);
and U19144 (N_19144,N_15554,N_15820);
xnor U19145 (N_19145,N_15994,N_16149);
or U19146 (N_19146,N_16826,N_16627);
and U19147 (N_19147,N_16604,N_16814);
xnor U19148 (N_19148,N_17125,N_16637);
xor U19149 (N_19149,N_16996,N_16019);
or U19150 (N_19150,N_16619,N_16336);
xnor U19151 (N_19151,N_16147,N_16022);
or U19152 (N_19152,N_15545,N_15348);
nand U19153 (N_19153,N_17047,N_16720);
and U19154 (N_19154,N_16527,N_15101);
xnor U19155 (N_19155,N_15864,N_15955);
and U19156 (N_19156,N_16578,N_16375);
xnor U19157 (N_19157,N_15721,N_15606);
nor U19158 (N_19158,N_16691,N_15149);
xnor U19159 (N_19159,N_17196,N_17289);
nand U19160 (N_19160,N_17326,N_15753);
or U19161 (N_19161,N_17419,N_16004);
or U19162 (N_19162,N_16116,N_17312);
xnor U19163 (N_19163,N_15092,N_15093);
or U19164 (N_19164,N_15417,N_16955);
xor U19165 (N_19165,N_15932,N_17147);
or U19166 (N_19166,N_15478,N_16507);
nor U19167 (N_19167,N_15430,N_15138);
and U19168 (N_19168,N_16752,N_15993);
nand U19169 (N_19169,N_15671,N_16648);
nor U19170 (N_19170,N_17411,N_16953);
xor U19171 (N_19171,N_16703,N_15234);
nor U19172 (N_19172,N_15189,N_15266);
nor U19173 (N_19173,N_15475,N_16193);
xor U19174 (N_19174,N_15292,N_16732);
nor U19175 (N_19175,N_15742,N_15751);
nor U19176 (N_19176,N_16211,N_16318);
nand U19177 (N_19177,N_16718,N_15778);
nor U19178 (N_19178,N_16438,N_16572);
xnor U19179 (N_19179,N_16492,N_17031);
and U19180 (N_19180,N_16865,N_15465);
xor U19181 (N_19181,N_16642,N_15036);
and U19182 (N_19182,N_15394,N_15204);
or U19183 (N_19183,N_15926,N_15160);
xnor U19184 (N_19184,N_15504,N_15695);
or U19185 (N_19185,N_15656,N_16713);
and U19186 (N_19186,N_15252,N_15261);
xnor U19187 (N_19187,N_16903,N_15950);
nand U19188 (N_19188,N_15129,N_16240);
nand U19189 (N_19189,N_16560,N_16568);
or U19190 (N_19190,N_16801,N_15207);
nor U19191 (N_19191,N_15079,N_17229);
and U19192 (N_19192,N_16038,N_15435);
nor U19193 (N_19193,N_16785,N_15727);
nand U19194 (N_19194,N_16570,N_17423);
and U19195 (N_19195,N_17449,N_15204);
or U19196 (N_19196,N_17493,N_17199);
xnor U19197 (N_19197,N_17254,N_17302);
nor U19198 (N_19198,N_16817,N_17348);
nor U19199 (N_19199,N_17298,N_15026);
xor U19200 (N_19200,N_16843,N_15070);
xnor U19201 (N_19201,N_15875,N_17273);
and U19202 (N_19202,N_15316,N_15487);
and U19203 (N_19203,N_17318,N_15975);
or U19204 (N_19204,N_15462,N_16890);
xor U19205 (N_19205,N_16616,N_16632);
or U19206 (N_19206,N_15117,N_16203);
nor U19207 (N_19207,N_16571,N_15040);
nand U19208 (N_19208,N_15121,N_17093);
or U19209 (N_19209,N_17304,N_16825);
nor U19210 (N_19210,N_15896,N_16059);
xor U19211 (N_19211,N_17180,N_15334);
nand U19212 (N_19212,N_17246,N_15472);
xnor U19213 (N_19213,N_15333,N_15586);
xnor U19214 (N_19214,N_15526,N_15774);
or U19215 (N_19215,N_16385,N_17378);
xnor U19216 (N_19216,N_16886,N_15120);
nand U19217 (N_19217,N_16408,N_16044);
nor U19218 (N_19218,N_15050,N_16849);
nand U19219 (N_19219,N_15554,N_16183);
nand U19220 (N_19220,N_15647,N_17101);
xnor U19221 (N_19221,N_17264,N_17126);
or U19222 (N_19222,N_15946,N_16575);
nand U19223 (N_19223,N_16248,N_15456);
and U19224 (N_19224,N_15312,N_15165);
or U19225 (N_19225,N_15100,N_16068);
and U19226 (N_19226,N_16207,N_17430);
xnor U19227 (N_19227,N_15546,N_16100);
xor U19228 (N_19228,N_16513,N_17397);
nand U19229 (N_19229,N_16091,N_16228);
nand U19230 (N_19230,N_16238,N_15000);
and U19231 (N_19231,N_16252,N_16473);
nand U19232 (N_19232,N_16189,N_15816);
nand U19233 (N_19233,N_15569,N_17384);
nand U19234 (N_19234,N_16630,N_15236);
or U19235 (N_19235,N_15191,N_17227);
or U19236 (N_19236,N_16470,N_15696);
or U19237 (N_19237,N_16700,N_17091);
nand U19238 (N_19238,N_15795,N_15716);
nand U19239 (N_19239,N_16259,N_16882);
xor U19240 (N_19240,N_15961,N_15094);
or U19241 (N_19241,N_16573,N_16519);
xnor U19242 (N_19242,N_16034,N_15209);
xnor U19243 (N_19243,N_15022,N_16293);
nor U19244 (N_19244,N_17462,N_15157);
and U19245 (N_19245,N_16555,N_16585);
or U19246 (N_19246,N_15703,N_17364);
and U19247 (N_19247,N_16378,N_16028);
xnor U19248 (N_19248,N_16062,N_15668);
or U19249 (N_19249,N_17251,N_16273);
nor U19250 (N_19250,N_15865,N_17096);
xnor U19251 (N_19251,N_16300,N_16412);
or U19252 (N_19252,N_16155,N_15494);
xor U19253 (N_19253,N_15939,N_17014);
xnor U19254 (N_19254,N_17384,N_15984);
nor U19255 (N_19255,N_17316,N_15453);
and U19256 (N_19256,N_15746,N_15337);
and U19257 (N_19257,N_17466,N_16338);
or U19258 (N_19258,N_15453,N_16577);
xor U19259 (N_19259,N_17183,N_15412);
nand U19260 (N_19260,N_17309,N_16629);
xor U19261 (N_19261,N_16960,N_15978);
xor U19262 (N_19262,N_15218,N_15262);
xnor U19263 (N_19263,N_17277,N_16101);
or U19264 (N_19264,N_17480,N_16000);
nor U19265 (N_19265,N_15695,N_16346);
nor U19266 (N_19266,N_15066,N_17394);
and U19267 (N_19267,N_17270,N_17298);
nor U19268 (N_19268,N_16786,N_16166);
or U19269 (N_19269,N_15412,N_17149);
nand U19270 (N_19270,N_16169,N_15733);
or U19271 (N_19271,N_17283,N_16076);
xor U19272 (N_19272,N_16158,N_16978);
and U19273 (N_19273,N_16817,N_16471);
or U19274 (N_19274,N_17452,N_16947);
or U19275 (N_19275,N_17336,N_15296);
nor U19276 (N_19276,N_15026,N_16403);
nand U19277 (N_19277,N_15764,N_16272);
xnor U19278 (N_19278,N_16199,N_16278);
and U19279 (N_19279,N_17280,N_15716);
nor U19280 (N_19280,N_16320,N_16611);
nor U19281 (N_19281,N_15569,N_17073);
nor U19282 (N_19282,N_15134,N_15391);
nand U19283 (N_19283,N_15590,N_15098);
or U19284 (N_19284,N_17034,N_16354);
xor U19285 (N_19285,N_17197,N_15991);
and U19286 (N_19286,N_15767,N_15031);
nor U19287 (N_19287,N_15418,N_16918);
and U19288 (N_19288,N_16849,N_16075);
nor U19289 (N_19289,N_15202,N_16567);
or U19290 (N_19290,N_16703,N_15328);
nand U19291 (N_19291,N_15361,N_17080);
and U19292 (N_19292,N_15372,N_16441);
and U19293 (N_19293,N_15716,N_16820);
nor U19294 (N_19294,N_15870,N_15642);
and U19295 (N_19295,N_16402,N_15864);
nor U19296 (N_19296,N_15655,N_16741);
nor U19297 (N_19297,N_15621,N_15049);
nor U19298 (N_19298,N_16829,N_16405);
nand U19299 (N_19299,N_15141,N_15014);
and U19300 (N_19300,N_15011,N_16117);
xor U19301 (N_19301,N_15473,N_15998);
or U19302 (N_19302,N_16616,N_15146);
nor U19303 (N_19303,N_16445,N_16719);
nand U19304 (N_19304,N_16478,N_15679);
nand U19305 (N_19305,N_17012,N_16641);
or U19306 (N_19306,N_15947,N_15744);
or U19307 (N_19307,N_17236,N_15748);
nor U19308 (N_19308,N_15737,N_17449);
nor U19309 (N_19309,N_17310,N_17009);
nand U19310 (N_19310,N_16140,N_16398);
and U19311 (N_19311,N_17027,N_17075);
nor U19312 (N_19312,N_16462,N_15427);
nor U19313 (N_19313,N_16956,N_15215);
nand U19314 (N_19314,N_15339,N_17085);
nor U19315 (N_19315,N_15031,N_15088);
and U19316 (N_19316,N_16752,N_16566);
nand U19317 (N_19317,N_17160,N_15753);
and U19318 (N_19318,N_16927,N_16367);
and U19319 (N_19319,N_15803,N_15380);
and U19320 (N_19320,N_17300,N_16200);
and U19321 (N_19321,N_16308,N_16358);
and U19322 (N_19322,N_15304,N_15129);
or U19323 (N_19323,N_15289,N_15182);
nor U19324 (N_19324,N_17206,N_16764);
nand U19325 (N_19325,N_17280,N_17348);
nor U19326 (N_19326,N_17487,N_16216);
xnor U19327 (N_19327,N_15991,N_15781);
or U19328 (N_19328,N_16311,N_17433);
xnor U19329 (N_19329,N_16309,N_15261);
nor U19330 (N_19330,N_16558,N_17128);
nand U19331 (N_19331,N_15087,N_17470);
nand U19332 (N_19332,N_15664,N_15452);
or U19333 (N_19333,N_15291,N_15404);
nand U19334 (N_19334,N_16945,N_15868);
xor U19335 (N_19335,N_15888,N_15255);
nor U19336 (N_19336,N_15069,N_17054);
and U19337 (N_19337,N_15306,N_16666);
or U19338 (N_19338,N_15294,N_15934);
nand U19339 (N_19339,N_16766,N_16683);
or U19340 (N_19340,N_15609,N_15499);
xnor U19341 (N_19341,N_16478,N_16237);
nor U19342 (N_19342,N_17346,N_16385);
nand U19343 (N_19343,N_16449,N_15909);
nor U19344 (N_19344,N_16045,N_16117);
and U19345 (N_19345,N_16120,N_15746);
xor U19346 (N_19346,N_16672,N_16063);
nand U19347 (N_19347,N_15537,N_16280);
xnor U19348 (N_19348,N_17247,N_15989);
or U19349 (N_19349,N_16998,N_15861);
or U19350 (N_19350,N_15982,N_17403);
nor U19351 (N_19351,N_15740,N_17244);
nor U19352 (N_19352,N_15503,N_17100);
nor U19353 (N_19353,N_16576,N_15830);
nor U19354 (N_19354,N_16330,N_16191);
xor U19355 (N_19355,N_16248,N_15673);
or U19356 (N_19356,N_15605,N_16709);
and U19357 (N_19357,N_17365,N_16787);
xnor U19358 (N_19358,N_16536,N_16890);
nor U19359 (N_19359,N_16161,N_17000);
nor U19360 (N_19360,N_15338,N_16363);
nor U19361 (N_19361,N_16993,N_17002);
nand U19362 (N_19362,N_16376,N_15188);
and U19363 (N_19363,N_17003,N_16933);
and U19364 (N_19364,N_17002,N_16698);
nor U19365 (N_19365,N_15334,N_16287);
or U19366 (N_19366,N_16639,N_15297);
and U19367 (N_19367,N_15249,N_15872);
nand U19368 (N_19368,N_16951,N_16241);
and U19369 (N_19369,N_17241,N_17156);
xor U19370 (N_19370,N_17335,N_15391);
xnor U19371 (N_19371,N_15126,N_15296);
and U19372 (N_19372,N_17425,N_17251);
nand U19373 (N_19373,N_16823,N_15071);
xor U19374 (N_19374,N_15910,N_15703);
xor U19375 (N_19375,N_16835,N_15390);
nor U19376 (N_19376,N_15181,N_16331);
or U19377 (N_19377,N_16842,N_16715);
and U19378 (N_19378,N_15385,N_16023);
nand U19379 (N_19379,N_16471,N_17107);
or U19380 (N_19380,N_17078,N_15191);
and U19381 (N_19381,N_16840,N_15687);
xnor U19382 (N_19382,N_17383,N_16559);
nand U19383 (N_19383,N_16567,N_16139);
xnor U19384 (N_19384,N_15919,N_15714);
nor U19385 (N_19385,N_16898,N_15412);
and U19386 (N_19386,N_15807,N_17065);
nor U19387 (N_19387,N_15442,N_16001);
nor U19388 (N_19388,N_15492,N_15853);
xnor U19389 (N_19389,N_15467,N_17013);
nand U19390 (N_19390,N_16376,N_17238);
xor U19391 (N_19391,N_16449,N_15542);
nor U19392 (N_19392,N_15692,N_15178);
nor U19393 (N_19393,N_16872,N_15422);
nor U19394 (N_19394,N_15198,N_17479);
xor U19395 (N_19395,N_17027,N_15274);
xor U19396 (N_19396,N_16630,N_16973);
nor U19397 (N_19397,N_15712,N_16160);
xor U19398 (N_19398,N_17004,N_17088);
nor U19399 (N_19399,N_15210,N_15118);
or U19400 (N_19400,N_16205,N_16561);
xor U19401 (N_19401,N_17349,N_16148);
xnor U19402 (N_19402,N_16904,N_15651);
xor U19403 (N_19403,N_16306,N_17064);
or U19404 (N_19404,N_17321,N_16611);
and U19405 (N_19405,N_16180,N_16186);
xor U19406 (N_19406,N_16190,N_15288);
or U19407 (N_19407,N_15319,N_17162);
nor U19408 (N_19408,N_15373,N_16793);
nand U19409 (N_19409,N_16970,N_17160);
nand U19410 (N_19410,N_15922,N_17231);
and U19411 (N_19411,N_17490,N_16697);
nor U19412 (N_19412,N_15298,N_16012);
nor U19413 (N_19413,N_15684,N_16835);
nor U19414 (N_19414,N_16113,N_16947);
nor U19415 (N_19415,N_15676,N_15047);
and U19416 (N_19416,N_15766,N_16337);
nor U19417 (N_19417,N_16219,N_17411);
nor U19418 (N_19418,N_16722,N_15960);
or U19419 (N_19419,N_15521,N_16844);
xnor U19420 (N_19420,N_16917,N_16801);
and U19421 (N_19421,N_16530,N_15454);
or U19422 (N_19422,N_16586,N_17348);
xor U19423 (N_19423,N_15310,N_16148);
xor U19424 (N_19424,N_17225,N_15810);
nor U19425 (N_19425,N_15540,N_16801);
nor U19426 (N_19426,N_17261,N_17016);
xnor U19427 (N_19427,N_15590,N_15633);
or U19428 (N_19428,N_15932,N_15346);
or U19429 (N_19429,N_16680,N_15386);
nand U19430 (N_19430,N_15951,N_16547);
and U19431 (N_19431,N_15298,N_15353);
xor U19432 (N_19432,N_17369,N_17228);
xnor U19433 (N_19433,N_16489,N_15301);
nand U19434 (N_19434,N_16851,N_16079);
nand U19435 (N_19435,N_16052,N_17091);
and U19436 (N_19436,N_15758,N_16514);
nand U19437 (N_19437,N_17098,N_16275);
nor U19438 (N_19438,N_16332,N_15252);
and U19439 (N_19439,N_16783,N_17417);
or U19440 (N_19440,N_15332,N_16259);
xor U19441 (N_19441,N_15897,N_15754);
xnor U19442 (N_19442,N_17249,N_16530);
or U19443 (N_19443,N_15527,N_15009);
nand U19444 (N_19444,N_16488,N_15826);
and U19445 (N_19445,N_17162,N_16429);
nor U19446 (N_19446,N_16277,N_17226);
nand U19447 (N_19447,N_16999,N_16520);
and U19448 (N_19448,N_17327,N_16115);
or U19449 (N_19449,N_16359,N_16192);
nand U19450 (N_19450,N_15860,N_15586);
nor U19451 (N_19451,N_17061,N_15188);
nand U19452 (N_19452,N_15751,N_16423);
or U19453 (N_19453,N_15171,N_16149);
nand U19454 (N_19454,N_15197,N_17499);
nor U19455 (N_19455,N_15045,N_15196);
and U19456 (N_19456,N_15818,N_17277);
nand U19457 (N_19457,N_15661,N_15011);
nor U19458 (N_19458,N_16752,N_16754);
or U19459 (N_19459,N_15728,N_15581);
xnor U19460 (N_19460,N_16062,N_15448);
nor U19461 (N_19461,N_16068,N_16177);
xor U19462 (N_19462,N_16787,N_15468);
xnor U19463 (N_19463,N_15542,N_16948);
and U19464 (N_19464,N_17045,N_16673);
or U19465 (N_19465,N_16255,N_15808);
nor U19466 (N_19466,N_15776,N_15925);
xor U19467 (N_19467,N_16661,N_16261);
nor U19468 (N_19468,N_15890,N_17249);
and U19469 (N_19469,N_15441,N_16327);
or U19470 (N_19470,N_16339,N_15745);
and U19471 (N_19471,N_16713,N_16455);
nor U19472 (N_19472,N_15037,N_17487);
or U19473 (N_19473,N_16441,N_16432);
nand U19474 (N_19474,N_15822,N_17279);
nor U19475 (N_19475,N_17111,N_16707);
xnor U19476 (N_19476,N_16931,N_15460);
or U19477 (N_19477,N_15112,N_16240);
nor U19478 (N_19478,N_16139,N_16094);
nor U19479 (N_19479,N_15931,N_16811);
or U19480 (N_19480,N_15005,N_15134);
xor U19481 (N_19481,N_16821,N_15513);
or U19482 (N_19482,N_15363,N_16307);
and U19483 (N_19483,N_17264,N_16948);
nand U19484 (N_19484,N_15021,N_16954);
nand U19485 (N_19485,N_15670,N_15052);
nor U19486 (N_19486,N_16579,N_16940);
or U19487 (N_19487,N_15246,N_16200);
xor U19488 (N_19488,N_17100,N_17009);
and U19489 (N_19489,N_16389,N_15079);
nor U19490 (N_19490,N_17275,N_15597);
and U19491 (N_19491,N_15346,N_16171);
nand U19492 (N_19492,N_16326,N_15397);
nand U19493 (N_19493,N_17482,N_16218);
nor U19494 (N_19494,N_15361,N_16594);
nand U19495 (N_19495,N_16383,N_16978);
and U19496 (N_19496,N_15396,N_16272);
and U19497 (N_19497,N_15107,N_15715);
and U19498 (N_19498,N_16413,N_16382);
nand U19499 (N_19499,N_16625,N_17350);
nand U19500 (N_19500,N_17309,N_17205);
and U19501 (N_19501,N_16118,N_17301);
and U19502 (N_19502,N_15557,N_15873);
xnor U19503 (N_19503,N_15858,N_17142);
or U19504 (N_19504,N_16077,N_16313);
xor U19505 (N_19505,N_17354,N_15864);
nand U19506 (N_19506,N_17193,N_16462);
or U19507 (N_19507,N_16943,N_16140);
nor U19508 (N_19508,N_16066,N_16718);
nor U19509 (N_19509,N_15986,N_15209);
or U19510 (N_19510,N_16031,N_15385);
nor U19511 (N_19511,N_17390,N_16667);
nor U19512 (N_19512,N_15851,N_16373);
xnor U19513 (N_19513,N_15805,N_17352);
or U19514 (N_19514,N_16295,N_15766);
or U19515 (N_19515,N_15599,N_16862);
nand U19516 (N_19516,N_15685,N_17082);
xor U19517 (N_19517,N_15937,N_15613);
and U19518 (N_19518,N_16319,N_15119);
xnor U19519 (N_19519,N_15409,N_16848);
xnor U19520 (N_19520,N_15027,N_16974);
xor U19521 (N_19521,N_15403,N_15559);
nand U19522 (N_19522,N_15813,N_15539);
and U19523 (N_19523,N_15325,N_17106);
nor U19524 (N_19524,N_16055,N_17177);
nand U19525 (N_19525,N_15179,N_15638);
or U19526 (N_19526,N_16837,N_16104);
or U19527 (N_19527,N_15997,N_17078);
nor U19528 (N_19528,N_15891,N_17351);
xnor U19529 (N_19529,N_15959,N_15527);
or U19530 (N_19530,N_16674,N_16834);
and U19531 (N_19531,N_16609,N_16924);
and U19532 (N_19532,N_17462,N_17368);
xor U19533 (N_19533,N_16690,N_16958);
xnor U19534 (N_19534,N_16677,N_15432);
nor U19535 (N_19535,N_15449,N_16134);
xor U19536 (N_19536,N_16765,N_16570);
or U19537 (N_19537,N_16606,N_15353);
nor U19538 (N_19538,N_17223,N_16741);
or U19539 (N_19539,N_17458,N_16922);
or U19540 (N_19540,N_16718,N_16478);
xor U19541 (N_19541,N_17483,N_16971);
and U19542 (N_19542,N_15979,N_15971);
nand U19543 (N_19543,N_15411,N_15738);
and U19544 (N_19544,N_15165,N_15529);
xor U19545 (N_19545,N_15989,N_17072);
nand U19546 (N_19546,N_15088,N_16323);
or U19547 (N_19547,N_17178,N_15166);
or U19548 (N_19548,N_15411,N_15479);
nor U19549 (N_19549,N_15985,N_16727);
nor U19550 (N_19550,N_16670,N_15497);
nor U19551 (N_19551,N_17147,N_15529);
and U19552 (N_19552,N_15071,N_16267);
xor U19553 (N_19553,N_16204,N_15566);
or U19554 (N_19554,N_15054,N_17135);
nand U19555 (N_19555,N_16660,N_15761);
nor U19556 (N_19556,N_16704,N_16358);
or U19557 (N_19557,N_17330,N_17238);
or U19558 (N_19558,N_15484,N_16956);
nor U19559 (N_19559,N_16985,N_17129);
xor U19560 (N_19560,N_16764,N_16102);
nand U19561 (N_19561,N_16770,N_16353);
and U19562 (N_19562,N_15742,N_15295);
and U19563 (N_19563,N_15697,N_15332);
nand U19564 (N_19564,N_15341,N_17440);
and U19565 (N_19565,N_17443,N_15145);
or U19566 (N_19566,N_16279,N_16111);
nor U19567 (N_19567,N_15287,N_17362);
nor U19568 (N_19568,N_15806,N_17147);
nand U19569 (N_19569,N_17190,N_16168);
nor U19570 (N_19570,N_15970,N_15517);
nor U19571 (N_19571,N_17433,N_16765);
or U19572 (N_19572,N_15424,N_15255);
and U19573 (N_19573,N_15202,N_17249);
xor U19574 (N_19574,N_16579,N_15848);
nor U19575 (N_19575,N_15113,N_15640);
nand U19576 (N_19576,N_15863,N_15923);
nor U19577 (N_19577,N_16632,N_16026);
and U19578 (N_19578,N_17265,N_15305);
nor U19579 (N_19579,N_15289,N_16210);
nor U19580 (N_19580,N_16326,N_15358);
or U19581 (N_19581,N_16864,N_16575);
nor U19582 (N_19582,N_17179,N_15871);
nor U19583 (N_19583,N_17241,N_16268);
and U19584 (N_19584,N_16196,N_17209);
and U19585 (N_19585,N_16541,N_15419);
xor U19586 (N_19586,N_16468,N_15299);
nand U19587 (N_19587,N_15430,N_17415);
or U19588 (N_19588,N_15919,N_16465);
and U19589 (N_19589,N_15260,N_15008);
nand U19590 (N_19590,N_15877,N_16732);
nand U19591 (N_19591,N_15458,N_17205);
nand U19592 (N_19592,N_17157,N_16772);
nor U19593 (N_19593,N_15437,N_15482);
nand U19594 (N_19594,N_17222,N_15113);
nor U19595 (N_19595,N_16165,N_16851);
xnor U19596 (N_19596,N_17177,N_16193);
nor U19597 (N_19597,N_16080,N_15311);
nand U19598 (N_19598,N_16579,N_15692);
xnor U19599 (N_19599,N_16584,N_16024);
xor U19600 (N_19600,N_15182,N_15526);
nand U19601 (N_19601,N_15522,N_16482);
or U19602 (N_19602,N_15735,N_15568);
nor U19603 (N_19603,N_17475,N_15241);
nor U19604 (N_19604,N_16466,N_16854);
xnor U19605 (N_19605,N_16241,N_15746);
and U19606 (N_19606,N_15166,N_15427);
nor U19607 (N_19607,N_16727,N_15328);
xnor U19608 (N_19608,N_17265,N_17069);
nand U19609 (N_19609,N_15015,N_15870);
or U19610 (N_19610,N_15900,N_15895);
nand U19611 (N_19611,N_16307,N_16653);
or U19612 (N_19612,N_15996,N_15356);
and U19613 (N_19613,N_16520,N_15057);
xnor U19614 (N_19614,N_16292,N_16840);
xor U19615 (N_19615,N_16365,N_15830);
or U19616 (N_19616,N_16938,N_15133);
or U19617 (N_19617,N_15928,N_17334);
nor U19618 (N_19618,N_15957,N_16698);
nand U19619 (N_19619,N_15181,N_15870);
nor U19620 (N_19620,N_17298,N_15137);
nor U19621 (N_19621,N_16231,N_15227);
nand U19622 (N_19622,N_17185,N_16415);
nand U19623 (N_19623,N_17102,N_17131);
or U19624 (N_19624,N_16850,N_15085);
nor U19625 (N_19625,N_15264,N_16693);
and U19626 (N_19626,N_15437,N_16423);
nand U19627 (N_19627,N_15236,N_15638);
and U19628 (N_19628,N_15737,N_17310);
nor U19629 (N_19629,N_16290,N_16929);
nand U19630 (N_19630,N_16590,N_16088);
and U19631 (N_19631,N_16052,N_16421);
nand U19632 (N_19632,N_17423,N_16551);
nand U19633 (N_19633,N_16888,N_15094);
xnor U19634 (N_19634,N_17496,N_17308);
nor U19635 (N_19635,N_15322,N_15819);
or U19636 (N_19636,N_15864,N_15873);
nand U19637 (N_19637,N_15271,N_16756);
xnor U19638 (N_19638,N_16977,N_15476);
xor U19639 (N_19639,N_17159,N_15180);
xnor U19640 (N_19640,N_15613,N_16114);
xnor U19641 (N_19641,N_15521,N_15927);
xor U19642 (N_19642,N_15484,N_15666);
or U19643 (N_19643,N_15359,N_16724);
nand U19644 (N_19644,N_17194,N_16579);
or U19645 (N_19645,N_16274,N_15033);
or U19646 (N_19646,N_15480,N_17432);
nand U19647 (N_19647,N_15395,N_15327);
and U19648 (N_19648,N_15909,N_15796);
or U19649 (N_19649,N_15825,N_15333);
and U19650 (N_19650,N_16484,N_17212);
or U19651 (N_19651,N_17395,N_15939);
xor U19652 (N_19652,N_17147,N_16990);
xor U19653 (N_19653,N_16337,N_16016);
or U19654 (N_19654,N_15797,N_15923);
xor U19655 (N_19655,N_16698,N_16033);
nor U19656 (N_19656,N_15812,N_15756);
and U19657 (N_19657,N_17025,N_16765);
nand U19658 (N_19658,N_15362,N_16704);
nand U19659 (N_19659,N_15534,N_16985);
xor U19660 (N_19660,N_16884,N_17445);
xnor U19661 (N_19661,N_16266,N_15171);
xnor U19662 (N_19662,N_15923,N_15493);
or U19663 (N_19663,N_15764,N_17007);
or U19664 (N_19664,N_16049,N_16793);
nand U19665 (N_19665,N_17388,N_17135);
xor U19666 (N_19666,N_16964,N_15955);
nor U19667 (N_19667,N_16042,N_16602);
and U19668 (N_19668,N_17424,N_16904);
and U19669 (N_19669,N_15327,N_15921);
or U19670 (N_19670,N_15012,N_15443);
nor U19671 (N_19671,N_15355,N_15794);
and U19672 (N_19672,N_16641,N_15659);
nor U19673 (N_19673,N_15413,N_17359);
xnor U19674 (N_19674,N_15192,N_15781);
or U19675 (N_19675,N_15041,N_15353);
nor U19676 (N_19676,N_16520,N_17027);
nor U19677 (N_19677,N_17002,N_15572);
and U19678 (N_19678,N_17165,N_15817);
xnor U19679 (N_19679,N_17122,N_15274);
nand U19680 (N_19680,N_16031,N_17211);
or U19681 (N_19681,N_17357,N_16463);
and U19682 (N_19682,N_16324,N_16411);
xnor U19683 (N_19683,N_16994,N_15767);
nand U19684 (N_19684,N_17252,N_16939);
nand U19685 (N_19685,N_16425,N_17387);
nor U19686 (N_19686,N_15493,N_15692);
xnor U19687 (N_19687,N_16977,N_15619);
xor U19688 (N_19688,N_16584,N_15751);
or U19689 (N_19689,N_17383,N_15827);
xnor U19690 (N_19690,N_15550,N_16450);
xnor U19691 (N_19691,N_15843,N_16958);
or U19692 (N_19692,N_17403,N_16377);
or U19693 (N_19693,N_16354,N_15786);
and U19694 (N_19694,N_16598,N_15276);
and U19695 (N_19695,N_15023,N_16166);
and U19696 (N_19696,N_17104,N_15266);
nor U19697 (N_19697,N_15010,N_16841);
or U19698 (N_19698,N_17235,N_15749);
and U19699 (N_19699,N_15695,N_16445);
xnor U19700 (N_19700,N_15965,N_15674);
and U19701 (N_19701,N_16519,N_16187);
or U19702 (N_19702,N_17134,N_15132);
and U19703 (N_19703,N_15646,N_17365);
nor U19704 (N_19704,N_16545,N_16296);
or U19705 (N_19705,N_17361,N_16572);
and U19706 (N_19706,N_15148,N_16010);
xnor U19707 (N_19707,N_16526,N_17056);
nor U19708 (N_19708,N_15554,N_15942);
nor U19709 (N_19709,N_17152,N_17277);
nand U19710 (N_19710,N_15683,N_16318);
or U19711 (N_19711,N_16239,N_15428);
or U19712 (N_19712,N_16259,N_16491);
nand U19713 (N_19713,N_16806,N_17012);
nor U19714 (N_19714,N_16025,N_17349);
and U19715 (N_19715,N_15537,N_15791);
and U19716 (N_19716,N_16872,N_17297);
nor U19717 (N_19717,N_16872,N_16100);
and U19718 (N_19718,N_15466,N_15651);
nand U19719 (N_19719,N_16263,N_15153);
or U19720 (N_19720,N_15265,N_16553);
or U19721 (N_19721,N_16791,N_15123);
xnor U19722 (N_19722,N_15407,N_17415);
xor U19723 (N_19723,N_16178,N_15811);
and U19724 (N_19724,N_15755,N_17314);
and U19725 (N_19725,N_16549,N_15355);
or U19726 (N_19726,N_15403,N_15040);
nand U19727 (N_19727,N_15963,N_17394);
xnor U19728 (N_19728,N_16040,N_16128);
or U19729 (N_19729,N_16847,N_17160);
nor U19730 (N_19730,N_16525,N_17310);
or U19731 (N_19731,N_16721,N_17318);
xor U19732 (N_19732,N_16259,N_17269);
xor U19733 (N_19733,N_16544,N_16639);
or U19734 (N_19734,N_17205,N_15670);
or U19735 (N_19735,N_15080,N_16735);
or U19736 (N_19736,N_15973,N_16782);
or U19737 (N_19737,N_15804,N_16757);
xnor U19738 (N_19738,N_15874,N_16105);
nand U19739 (N_19739,N_16566,N_15022);
xnor U19740 (N_19740,N_15839,N_16042);
and U19741 (N_19741,N_15577,N_16827);
nor U19742 (N_19742,N_16679,N_16550);
xor U19743 (N_19743,N_17176,N_17062);
nand U19744 (N_19744,N_17081,N_16279);
xor U19745 (N_19745,N_15752,N_15733);
xnor U19746 (N_19746,N_17403,N_16565);
and U19747 (N_19747,N_16106,N_16154);
xnor U19748 (N_19748,N_17317,N_16711);
xor U19749 (N_19749,N_16957,N_15000);
and U19750 (N_19750,N_15863,N_15990);
xor U19751 (N_19751,N_15790,N_15026);
xor U19752 (N_19752,N_16428,N_16110);
or U19753 (N_19753,N_16360,N_16206);
or U19754 (N_19754,N_15693,N_15117);
nand U19755 (N_19755,N_17288,N_16367);
or U19756 (N_19756,N_17082,N_16403);
nor U19757 (N_19757,N_15204,N_16336);
or U19758 (N_19758,N_15975,N_15610);
and U19759 (N_19759,N_16456,N_15422);
nor U19760 (N_19760,N_16699,N_17386);
xnor U19761 (N_19761,N_15122,N_15570);
and U19762 (N_19762,N_16822,N_17000);
or U19763 (N_19763,N_15017,N_17112);
nand U19764 (N_19764,N_15968,N_16324);
nand U19765 (N_19765,N_15834,N_16314);
or U19766 (N_19766,N_16764,N_15363);
nor U19767 (N_19767,N_17436,N_15200);
nor U19768 (N_19768,N_16767,N_15009);
nor U19769 (N_19769,N_17290,N_15880);
nor U19770 (N_19770,N_16825,N_15961);
and U19771 (N_19771,N_15715,N_15370);
nor U19772 (N_19772,N_15011,N_15072);
and U19773 (N_19773,N_15124,N_16055);
and U19774 (N_19774,N_15859,N_16336);
nand U19775 (N_19775,N_16344,N_16929);
and U19776 (N_19776,N_17029,N_17119);
xor U19777 (N_19777,N_15276,N_15653);
xnor U19778 (N_19778,N_17420,N_15098);
or U19779 (N_19779,N_17150,N_16682);
and U19780 (N_19780,N_17258,N_16083);
or U19781 (N_19781,N_16603,N_16468);
and U19782 (N_19782,N_15492,N_17367);
nand U19783 (N_19783,N_16072,N_15884);
or U19784 (N_19784,N_17029,N_15072);
nand U19785 (N_19785,N_15832,N_15924);
nand U19786 (N_19786,N_17197,N_16010);
nand U19787 (N_19787,N_16282,N_16032);
and U19788 (N_19788,N_16095,N_15472);
nand U19789 (N_19789,N_16038,N_15208);
nand U19790 (N_19790,N_16492,N_15116);
xor U19791 (N_19791,N_15237,N_16171);
or U19792 (N_19792,N_15809,N_16409);
and U19793 (N_19793,N_15379,N_16094);
or U19794 (N_19794,N_15553,N_16502);
or U19795 (N_19795,N_16096,N_16316);
or U19796 (N_19796,N_16219,N_16732);
and U19797 (N_19797,N_15387,N_17085);
nor U19798 (N_19798,N_16347,N_15200);
nand U19799 (N_19799,N_16058,N_16740);
nand U19800 (N_19800,N_15051,N_16808);
xnor U19801 (N_19801,N_16298,N_15655);
nor U19802 (N_19802,N_16916,N_15964);
nand U19803 (N_19803,N_15367,N_15206);
or U19804 (N_19804,N_15239,N_16073);
xnor U19805 (N_19805,N_15222,N_15431);
nor U19806 (N_19806,N_16709,N_16163);
and U19807 (N_19807,N_16362,N_15166);
xor U19808 (N_19808,N_16126,N_15813);
xnor U19809 (N_19809,N_15988,N_16634);
and U19810 (N_19810,N_15794,N_16955);
xor U19811 (N_19811,N_16554,N_15164);
or U19812 (N_19812,N_16820,N_16728);
nand U19813 (N_19813,N_16196,N_17036);
nand U19814 (N_19814,N_16830,N_17403);
nand U19815 (N_19815,N_15886,N_15126);
or U19816 (N_19816,N_15908,N_16159);
nand U19817 (N_19817,N_16779,N_16502);
or U19818 (N_19818,N_15264,N_15837);
and U19819 (N_19819,N_17025,N_17215);
xnor U19820 (N_19820,N_16157,N_17113);
nor U19821 (N_19821,N_17426,N_15788);
or U19822 (N_19822,N_15178,N_15739);
nand U19823 (N_19823,N_16319,N_15121);
nand U19824 (N_19824,N_15148,N_15319);
nor U19825 (N_19825,N_15340,N_16099);
or U19826 (N_19826,N_17458,N_15432);
xor U19827 (N_19827,N_15674,N_17123);
nor U19828 (N_19828,N_15391,N_16011);
or U19829 (N_19829,N_16582,N_16523);
or U19830 (N_19830,N_16412,N_17134);
and U19831 (N_19831,N_15435,N_15952);
xor U19832 (N_19832,N_15867,N_15634);
or U19833 (N_19833,N_15440,N_15143);
or U19834 (N_19834,N_16616,N_15795);
and U19835 (N_19835,N_15708,N_16757);
and U19836 (N_19836,N_17148,N_16913);
nand U19837 (N_19837,N_16818,N_16514);
nand U19838 (N_19838,N_15334,N_15146);
and U19839 (N_19839,N_15886,N_15118);
and U19840 (N_19840,N_15389,N_17314);
and U19841 (N_19841,N_15282,N_17304);
xor U19842 (N_19842,N_15367,N_17307);
nand U19843 (N_19843,N_15380,N_16729);
xor U19844 (N_19844,N_17413,N_16867);
and U19845 (N_19845,N_15205,N_15199);
nor U19846 (N_19846,N_15732,N_17425);
xnor U19847 (N_19847,N_17085,N_15869);
nor U19848 (N_19848,N_15547,N_16754);
nor U19849 (N_19849,N_16923,N_15524);
or U19850 (N_19850,N_15021,N_15288);
xnor U19851 (N_19851,N_16290,N_17262);
nor U19852 (N_19852,N_15107,N_17130);
or U19853 (N_19853,N_17193,N_15330);
nand U19854 (N_19854,N_16456,N_17480);
and U19855 (N_19855,N_15291,N_15267);
nand U19856 (N_19856,N_15978,N_16152);
and U19857 (N_19857,N_15438,N_15834);
xnor U19858 (N_19858,N_15973,N_16783);
or U19859 (N_19859,N_15456,N_15307);
or U19860 (N_19860,N_15332,N_16597);
nand U19861 (N_19861,N_17434,N_16737);
xor U19862 (N_19862,N_15452,N_15022);
xor U19863 (N_19863,N_16319,N_16605);
xnor U19864 (N_19864,N_17248,N_16348);
and U19865 (N_19865,N_15295,N_15675);
and U19866 (N_19866,N_16549,N_16805);
and U19867 (N_19867,N_17157,N_16649);
nand U19868 (N_19868,N_15564,N_16866);
and U19869 (N_19869,N_15578,N_15925);
or U19870 (N_19870,N_15832,N_15592);
xor U19871 (N_19871,N_16684,N_16774);
nand U19872 (N_19872,N_15483,N_15615);
and U19873 (N_19873,N_16749,N_16138);
nand U19874 (N_19874,N_15067,N_16005);
or U19875 (N_19875,N_15065,N_17337);
xor U19876 (N_19876,N_16027,N_16019);
xnor U19877 (N_19877,N_15430,N_15100);
nor U19878 (N_19878,N_16414,N_15818);
or U19879 (N_19879,N_17446,N_16688);
xnor U19880 (N_19880,N_17108,N_16162);
nor U19881 (N_19881,N_16404,N_15649);
xnor U19882 (N_19882,N_15310,N_15343);
nor U19883 (N_19883,N_17179,N_17389);
nand U19884 (N_19884,N_15920,N_17161);
and U19885 (N_19885,N_16604,N_15594);
or U19886 (N_19886,N_15057,N_17011);
nor U19887 (N_19887,N_16993,N_16008);
or U19888 (N_19888,N_15824,N_16537);
nand U19889 (N_19889,N_15434,N_16250);
or U19890 (N_19890,N_17012,N_16669);
nand U19891 (N_19891,N_15047,N_17232);
nor U19892 (N_19892,N_17045,N_16953);
and U19893 (N_19893,N_16738,N_15098);
xor U19894 (N_19894,N_16740,N_16187);
nand U19895 (N_19895,N_16736,N_15098);
xor U19896 (N_19896,N_16290,N_15341);
nand U19897 (N_19897,N_15109,N_16720);
xnor U19898 (N_19898,N_15837,N_17054);
nand U19899 (N_19899,N_16346,N_15419);
nor U19900 (N_19900,N_15329,N_16545);
and U19901 (N_19901,N_16546,N_15291);
xor U19902 (N_19902,N_15014,N_15247);
nand U19903 (N_19903,N_17156,N_15474);
or U19904 (N_19904,N_16252,N_15082);
and U19905 (N_19905,N_16636,N_17278);
and U19906 (N_19906,N_16354,N_16692);
and U19907 (N_19907,N_17283,N_16414);
and U19908 (N_19908,N_15198,N_16823);
nand U19909 (N_19909,N_16797,N_15865);
or U19910 (N_19910,N_16815,N_15714);
xor U19911 (N_19911,N_17471,N_15435);
xor U19912 (N_19912,N_17032,N_15196);
nand U19913 (N_19913,N_15933,N_17132);
and U19914 (N_19914,N_15256,N_15447);
and U19915 (N_19915,N_16535,N_16739);
xnor U19916 (N_19916,N_15831,N_16955);
and U19917 (N_19917,N_16200,N_17148);
or U19918 (N_19918,N_15483,N_15278);
and U19919 (N_19919,N_15668,N_15038);
nor U19920 (N_19920,N_15256,N_17448);
and U19921 (N_19921,N_16545,N_17232);
nand U19922 (N_19922,N_17143,N_15558);
or U19923 (N_19923,N_16686,N_16920);
xor U19924 (N_19924,N_16960,N_17367);
nor U19925 (N_19925,N_15209,N_16995);
xor U19926 (N_19926,N_15718,N_15198);
xor U19927 (N_19927,N_17446,N_15676);
nand U19928 (N_19928,N_16054,N_15978);
nor U19929 (N_19929,N_17140,N_15791);
xnor U19930 (N_19930,N_16871,N_17158);
nor U19931 (N_19931,N_17073,N_15632);
and U19932 (N_19932,N_16080,N_16444);
nor U19933 (N_19933,N_15795,N_16926);
xnor U19934 (N_19934,N_15545,N_16867);
nor U19935 (N_19935,N_15437,N_16348);
nand U19936 (N_19936,N_17395,N_16614);
nand U19937 (N_19937,N_16893,N_16405);
and U19938 (N_19938,N_16205,N_15063);
or U19939 (N_19939,N_15971,N_16589);
or U19940 (N_19940,N_16846,N_17042);
nand U19941 (N_19941,N_16895,N_16132);
nand U19942 (N_19942,N_16166,N_16278);
xnor U19943 (N_19943,N_17185,N_17081);
nor U19944 (N_19944,N_15357,N_16641);
nand U19945 (N_19945,N_16907,N_15507);
or U19946 (N_19946,N_16487,N_15964);
or U19947 (N_19947,N_16155,N_16487);
or U19948 (N_19948,N_15311,N_16000);
and U19949 (N_19949,N_16566,N_15265);
xnor U19950 (N_19950,N_16630,N_15229);
or U19951 (N_19951,N_15348,N_15746);
xor U19952 (N_19952,N_16774,N_15228);
nor U19953 (N_19953,N_17407,N_17329);
or U19954 (N_19954,N_16611,N_16987);
xnor U19955 (N_19955,N_15444,N_17122);
xnor U19956 (N_19956,N_16060,N_16004);
and U19957 (N_19957,N_15013,N_16653);
and U19958 (N_19958,N_15000,N_16837);
nand U19959 (N_19959,N_16791,N_17282);
xor U19960 (N_19960,N_15228,N_15371);
nor U19961 (N_19961,N_15634,N_16992);
nand U19962 (N_19962,N_15891,N_15990);
nand U19963 (N_19963,N_15763,N_16096);
or U19964 (N_19964,N_17239,N_16405);
or U19965 (N_19965,N_15982,N_16622);
nand U19966 (N_19966,N_16825,N_17198);
and U19967 (N_19967,N_16585,N_15020);
nor U19968 (N_19968,N_15680,N_16504);
xor U19969 (N_19969,N_15455,N_15478);
nor U19970 (N_19970,N_15842,N_17448);
or U19971 (N_19971,N_15889,N_15624);
and U19972 (N_19972,N_15901,N_15403);
xor U19973 (N_19973,N_16380,N_15340);
and U19974 (N_19974,N_17028,N_16048);
nand U19975 (N_19975,N_16061,N_17007);
nand U19976 (N_19976,N_16996,N_15160);
or U19977 (N_19977,N_17037,N_16452);
nand U19978 (N_19978,N_17317,N_15704);
nor U19979 (N_19979,N_15257,N_17174);
xor U19980 (N_19980,N_15764,N_16811);
and U19981 (N_19981,N_16380,N_16531);
and U19982 (N_19982,N_16532,N_17090);
nand U19983 (N_19983,N_15856,N_17260);
and U19984 (N_19984,N_17254,N_15101);
xor U19985 (N_19985,N_15620,N_16688);
nand U19986 (N_19986,N_17376,N_15238);
and U19987 (N_19987,N_16192,N_16504);
xor U19988 (N_19988,N_16690,N_15447);
nand U19989 (N_19989,N_16405,N_15605);
or U19990 (N_19990,N_15719,N_16386);
and U19991 (N_19991,N_15629,N_17131);
xor U19992 (N_19992,N_15933,N_16920);
nand U19993 (N_19993,N_15328,N_16475);
nand U19994 (N_19994,N_15751,N_16977);
and U19995 (N_19995,N_16571,N_17478);
xnor U19996 (N_19996,N_16008,N_15593);
nor U19997 (N_19997,N_17176,N_15601);
xnor U19998 (N_19998,N_17023,N_17187);
and U19999 (N_19999,N_16151,N_16596);
nor U20000 (N_20000,N_19132,N_17914);
xnor U20001 (N_20001,N_17609,N_19761);
or U20002 (N_20002,N_19297,N_19335);
nand U20003 (N_20003,N_18218,N_18166);
xnor U20004 (N_20004,N_17989,N_19515);
nand U20005 (N_20005,N_19381,N_19180);
or U20006 (N_20006,N_19193,N_18376);
and U20007 (N_20007,N_18138,N_18472);
xor U20008 (N_20008,N_19800,N_18751);
or U20009 (N_20009,N_18824,N_17710);
nand U20010 (N_20010,N_18651,N_17675);
or U20011 (N_20011,N_18168,N_18474);
nor U20012 (N_20012,N_19284,N_18086);
nand U20013 (N_20013,N_19007,N_18446);
or U20014 (N_20014,N_17698,N_18089);
or U20015 (N_20015,N_19799,N_17712);
nor U20016 (N_20016,N_19118,N_19313);
nand U20017 (N_20017,N_18359,N_17629);
or U20018 (N_20018,N_19862,N_18702);
nand U20019 (N_20019,N_18003,N_18793);
and U20020 (N_20020,N_18906,N_19221);
nand U20021 (N_20021,N_19172,N_19576);
xor U20022 (N_20022,N_19927,N_17970);
nand U20023 (N_20023,N_18554,N_18189);
nand U20024 (N_20024,N_19601,N_19101);
xor U20025 (N_20025,N_19818,N_17669);
xor U20026 (N_20026,N_19616,N_19873);
or U20027 (N_20027,N_19588,N_18722);
xnor U20028 (N_20028,N_18642,N_19569);
nand U20029 (N_20029,N_19706,N_19508);
nor U20030 (N_20030,N_19342,N_18210);
nand U20031 (N_20031,N_17800,N_19655);
and U20032 (N_20032,N_17895,N_17876);
and U20033 (N_20033,N_17967,N_18071);
nand U20034 (N_20034,N_18338,N_17590);
and U20035 (N_20035,N_19806,N_17718);
nor U20036 (N_20036,N_18820,N_18082);
nor U20037 (N_20037,N_19143,N_19306);
and U20038 (N_20038,N_17846,N_19715);
nand U20039 (N_20039,N_19861,N_18303);
nand U20040 (N_20040,N_18779,N_17690);
nor U20041 (N_20041,N_19982,N_18070);
or U20042 (N_20042,N_19201,N_18840);
xor U20043 (N_20043,N_17924,N_18146);
and U20044 (N_20044,N_19496,N_19675);
nor U20045 (N_20045,N_18783,N_18899);
and U20046 (N_20046,N_19840,N_19446);
nor U20047 (N_20047,N_19415,N_19980);
nand U20048 (N_20048,N_17742,N_17950);
xnor U20049 (N_20049,N_19159,N_19499);
xnor U20050 (N_20050,N_19764,N_19234);
xnor U20051 (N_20051,N_18269,N_18099);
xor U20052 (N_20052,N_19832,N_17975);
xor U20053 (N_20053,N_19164,N_17603);
nor U20054 (N_20054,N_18100,N_18666);
nand U20055 (N_20055,N_18664,N_17550);
nand U20056 (N_20056,N_17642,N_17785);
nor U20057 (N_20057,N_18630,N_19393);
or U20058 (N_20058,N_19334,N_19626);
xor U20059 (N_20059,N_18998,N_19236);
xnor U20060 (N_20060,N_18067,N_17582);
and U20061 (N_20061,N_17891,N_18533);
and U20062 (N_20062,N_18774,N_18952);
and U20063 (N_20063,N_18813,N_19040);
or U20064 (N_20064,N_19605,N_19489);
or U20065 (N_20065,N_19188,N_18075);
or U20066 (N_20066,N_18718,N_18128);
nand U20067 (N_20067,N_19788,N_19509);
or U20068 (N_20068,N_19753,N_17608);
nand U20069 (N_20069,N_18234,N_19198);
xor U20070 (N_20070,N_18827,N_19526);
xor U20071 (N_20071,N_18291,N_19329);
nor U20072 (N_20072,N_18018,N_19822);
nand U20073 (N_20073,N_18668,N_19653);
and U20074 (N_20074,N_19875,N_19893);
xnor U20075 (N_20075,N_19562,N_19519);
nand U20076 (N_20076,N_19116,N_18069);
or U20077 (N_20077,N_18419,N_19249);
nand U20078 (N_20078,N_18029,N_19561);
nor U20079 (N_20079,N_19106,N_18851);
xnor U20080 (N_20080,N_17646,N_17734);
or U20081 (N_20081,N_18962,N_19196);
xor U20082 (N_20082,N_19014,N_19583);
or U20083 (N_20083,N_19537,N_18406);
nor U20084 (N_20084,N_18611,N_18917);
nand U20085 (N_20085,N_17663,N_19389);
nand U20086 (N_20086,N_19787,N_19487);
nand U20087 (N_20087,N_18053,N_19896);
nor U20088 (N_20088,N_18312,N_17702);
nor U20089 (N_20089,N_18966,N_19093);
nand U20090 (N_20090,N_17579,N_19360);
nor U20091 (N_20091,N_19936,N_18402);
nor U20092 (N_20092,N_17701,N_18842);
nand U20093 (N_20093,N_18014,N_19940);
and U20094 (N_20094,N_17858,N_17833);
and U20095 (N_20095,N_18500,N_19190);
nand U20096 (N_20096,N_18949,N_17904);
or U20097 (N_20097,N_19433,N_18978);
nand U20098 (N_20098,N_19044,N_19812);
nor U20099 (N_20099,N_19957,N_19482);
and U20100 (N_20100,N_18788,N_18366);
or U20101 (N_20101,N_17761,N_19318);
nand U20102 (N_20102,N_19866,N_19039);
or U20103 (N_20103,N_19974,N_18864);
and U20104 (N_20104,N_17847,N_19837);
xnor U20105 (N_20105,N_18434,N_17659);
nand U20106 (N_20106,N_17720,N_17747);
or U20107 (N_20107,N_18423,N_19557);
nand U20108 (N_20108,N_18823,N_19632);
nand U20109 (N_20109,N_19046,N_18881);
nand U20110 (N_20110,N_18551,N_18797);
and U20111 (N_20111,N_18244,N_18095);
or U20112 (N_20112,N_18729,N_18608);
nor U20113 (N_20113,N_18943,N_17738);
and U20114 (N_20114,N_18490,N_19993);
nor U20115 (N_20115,N_17694,N_18343);
xnor U20116 (N_20116,N_18714,N_18931);
nand U20117 (N_20117,N_18114,N_19076);
nand U20118 (N_20118,N_17937,N_17886);
nand U20119 (N_20119,N_18846,N_17953);
xnor U20120 (N_20120,N_18353,N_18161);
xnor U20121 (N_20121,N_19219,N_17619);
nor U20122 (N_20122,N_19490,N_17898);
nor U20123 (N_20123,N_18932,N_17863);
and U20124 (N_20124,N_18557,N_18396);
xnor U20125 (N_20125,N_18122,N_19466);
nor U20126 (N_20126,N_19506,N_18290);
and U20127 (N_20127,N_17983,N_17523);
nand U20128 (N_20128,N_19793,N_18280);
or U20129 (N_20129,N_18461,N_18091);
nor U20130 (N_20130,N_17987,N_17888);
xnor U20131 (N_20131,N_18001,N_17957);
nor U20132 (N_20132,N_19006,N_19151);
nor U20133 (N_20133,N_18944,N_19992);
or U20134 (N_20134,N_19390,N_19384);
and U20135 (N_20135,N_17598,N_18103);
and U20136 (N_20136,N_19518,N_17796);
and U20137 (N_20137,N_19947,N_17614);
nand U20138 (N_20138,N_19803,N_17580);
and U20139 (N_20139,N_19447,N_18157);
nor U20140 (N_20140,N_19140,N_18717);
xnor U20141 (N_20141,N_18677,N_17963);
or U20142 (N_20142,N_19652,N_18653);
nand U20143 (N_20143,N_18242,N_17790);
nand U20144 (N_20144,N_19426,N_18828);
and U20145 (N_20145,N_18794,N_18921);
and U20146 (N_20146,N_17654,N_19063);
or U20147 (N_20147,N_19839,N_19386);
or U20148 (N_20148,N_18347,N_18395);
or U20149 (N_20149,N_17972,N_19780);
xnor U20150 (N_20150,N_17851,N_17620);
xor U20151 (N_20151,N_19609,N_19391);
and U20152 (N_20152,N_17695,N_18088);
nand U20153 (N_20153,N_18634,N_19035);
nand U20154 (N_20154,N_18129,N_19081);
nand U20155 (N_20155,N_19358,N_18473);
and U20156 (N_20156,N_17643,N_17996);
nand U20157 (N_20157,N_18044,N_19091);
xnor U20158 (N_20158,N_18649,N_18000);
or U20159 (N_20159,N_19842,N_19458);
and U20160 (N_20160,N_19952,N_18929);
nor U20161 (N_20161,N_19208,N_19829);
nand U20162 (N_20162,N_17520,N_18524);
nand U20163 (N_20163,N_18925,N_18509);
and U20164 (N_20164,N_19810,N_17705);
nand U20165 (N_20165,N_17573,N_17692);
nand U20166 (N_20166,N_17778,N_19410);
xnor U20167 (N_20167,N_19146,N_19846);
and U20168 (N_20168,N_18330,N_18937);
nor U20169 (N_20169,N_18809,N_17994);
and U20170 (N_20170,N_19621,N_17973);
nand U20171 (N_20171,N_19213,N_17799);
nor U20172 (N_20172,N_18172,N_18875);
or U20173 (N_20173,N_18764,N_19628);
xor U20174 (N_20174,N_19295,N_17716);
and U20175 (N_20175,N_17834,N_18391);
and U20176 (N_20176,N_19288,N_18156);
and U20177 (N_20177,N_19400,N_17507);
or U20178 (N_20178,N_19836,N_17991);
xnor U20179 (N_20179,N_19406,N_18999);
and U20180 (N_20180,N_19702,N_18352);
xor U20181 (N_20181,N_18380,N_19250);
xnor U20182 (N_20182,N_19773,N_18766);
or U20183 (N_20183,N_17636,N_17762);
xor U20184 (N_20184,N_18271,N_19905);
nand U20185 (N_20185,N_17805,N_18207);
nand U20186 (N_20186,N_19887,N_19918);
xor U20187 (N_20187,N_17911,N_18715);
and U20188 (N_20188,N_19034,N_18096);
xnor U20189 (N_20189,N_19928,N_19671);
xor U20190 (N_20190,N_19088,N_18215);
and U20191 (N_20191,N_17713,N_18455);
nor U20192 (N_20192,N_19082,N_17632);
nor U20193 (N_20193,N_19211,N_18744);
nand U20194 (N_20194,N_18682,N_19177);
nand U20195 (N_20195,N_17531,N_18553);
or U20196 (N_20196,N_19388,N_19405);
nor U20197 (N_20197,N_18394,N_17871);
and U20198 (N_20198,N_19454,N_19272);
xor U20199 (N_20199,N_18619,N_18017);
nor U20200 (N_20200,N_19871,N_18894);
xnor U20201 (N_20201,N_17770,N_19009);
nand U20202 (N_20202,N_19586,N_18205);
nor U20203 (N_20203,N_17666,N_19094);
nand U20204 (N_20204,N_18317,N_18769);
or U20205 (N_20205,N_18730,N_19951);
or U20206 (N_20206,N_19030,N_18361);
or U20207 (N_20207,N_18284,N_18226);
or U20208 (N_20208,N_18024,N_18540);
xnor U20209 (N_20209,N_19682,N_17848);
and U20210 (N_20210,N_18308,N_19054);
xor U20211 (N_20211,N_18115,N_18740);
nor U20212 (N_20212,N_18230,N_19817);
nor U20213 (N_20213,N_17645,N_19757);
nor U20214 (N_20214,N_18120,N_18439);
nor U20215 (N_20215,N_18165,N_17753);
nor U20216 (N_20216,N_18350,N_17901);
nand U20217 (N_20217,N_19192,N_18508);
and U20218 (N_20218,N_19680,N_19011);
xor U20219 (N_20219,N_18057,N_18325);
and U20220 (N_20220,N_19001,N_19550);
or U20221 (N_20221,N_17574,N_17586);
nand U20222 (N_20222,N_17611,N_18222);
nand U20223 (N_20223,N_18631,N_19921);
nor U20224 (N_20224,N_18424,N_19546);
and U20225 (N_20225,N_18883,N_19577);
xor U20226 (N_20226,N_19022,N_19794);
nor U20227 (N_20227,N_17992,N_18021);
xnor U20228 (N_20228,N_19536,N_17906);
xor U20229 (N_20229,N_19726,N_18311);
xor U20230 (N_20230,N_18538,N_18587);
and U20231 (N_20231,N_18983,N_17714);
or U20232 (N_20232,N_18351,N_19238);
nand U20233 (N_20233,N_18732,N_19748);
xnor U20234 (N_20234,N_18408,N_19950);
nand U20235 (N_20235,N_18371,N_17981);
and U20236 (N_20236,N_18652,N_19665);
or U20237 (N_20237,N_19606,N_19914);
and U20238 (N_20238,N_18151,N_18762);
nand U20239 (N_20239,N_18005,N_19455);
nand U20240 (N_20240,N_18042,N_18358);
xor U20241 (N_20241,N_19555,N_17926);
xor U20242 (N_20242,N_19777,N_17797);
xnor U20243 (N_20243,N_17978,N_18586);
nand U20244 (N_20244,N_19571,N_19813);
xor U20245 (N_20245,N_19811,N_18227);
nor U20246 (N_20246,N_17938,N_19684);
nand U20247 (N_20247,N_18695,N_19937);
and U20248 (N_20248,N_19805,N_19075);
or U20249 (N_20249,N_17791,N_19444);
and U20250 (N_20250,N_17649,N_18106);
nand U20251 (N_20251,N_19419,N_18759);
or U20252 (N_20252,N_18957,N_19638);
or U20253 (N_20253,N_19383,N_19268);
xor U20254 (N_20254,N_18958,N_19189);
nand U20255 (N_20255,N_17581,N_19195);
xor U20256 (N_20256,N_19868,N_18855);
and U20257 (N_20257,N_18585,N_17758);
or U20258 (N_20258,N_18671,N_19347);
xor U20259 (N_20259,N_19807,N_18985);
nor U20260 (N_20260,N_19567,N_19969);
nand U20261 (N_20261,N_18834,N_18987);
nor U20262 (N_20262,N_19549,N_17739);
nor U20263 (N_20263,N_18184,N_18140);
nor U20264 (N_20264,N_19949,N_18259);
or U20265 (N_20265,N_18485,N_18287);
and U20266 (N_20266,N_18041,N_19055);
nand U20267 (N_20267,N_19316,N_19654);
nand U20268 (N_20268,N_19804,N_18623);
and U20269 (N_20269,N_19084,N_19591);
and U20270 (N_20270,N_18690,N_18735);
or U20271 (N_20271,N_17741,N_18143);
and U20272 (N_20272,N_17831,N_18154);
or U20273 (N_20273,N_18697,N_19668);
xor U20274 (N_20274,N_19544,N_19791);
xor U20275 (N_20275,N_17672,N_17736);
and U20276 (N_20276,N_19120,N_19545);
or U20277 (N_20277,N_19850,N_17872);
nand U20278 (N_20278,N_19450,N_17638);
xor U20279 (N_20279,N_19319,N_19589);
xor U20280 (N_20280,N_18887,N_18970);
xnor U20281 (N_20281,N_19532,N_18570);
and U20282 (N_20282,N_18369,N_19279);
nand U20283 (N_20283,N_19476,N_18904);
or U20284 (N_20284,N_19721,N_18327);
nand U20285 (N_20285,N_18927,N_17612);
nor U20286 (N_20286,N_18491,N_18600);
nand U20287 (N_20287,N_19412,N_19963);
xor U20288 (N_20288,N_19864,N_18681);
or U20289 (N_20289,N_19237,N_17874);
nor U20290 (N_20290,N_19679,N_19163);
nand U20291 (N_20291,N_18795,N_18449);
nor U20292 (N_20292,N_18547,N_19428);
nor U20293 (N_20293,N_19340,N_18592);
and U20294 (N_20294,N_19833,N_17995);
nor U20295 (N_20295,N_19531,N_18436);
or U20296 (N_20296,N_18936,N_17766);
xnor U20297 (N_20297,N_19374,N_17516);
nand U20298 (N_20298,N_19994,N_17793);
nand U20299 (N_20299,N_19369,N_19475);
nor U20300 (N_20300,N_18986,N_17896);
or U20301 (N_20301,N_17711,N_18268);
xnor U20302 (N_20302,N_19965,N_19785);
nor U20303 (N_20303,N_17930,N_18701);
or U20304 (N_20304,N_17630,N_19286);
nor U20305 (N_20305,N_19263,N_17915);
xor U20306 (N_20306,N_18412,N_18833);
and U20307 (N_20307,N_17729,N_19112);
xnor U20308 (N_20308,N_18506,N_17674);
or U20309 (N_20309,N_17732,N_19573);
nand U20310 (N_20310,N_19227,N_18825);
nor U20311 (N_20311,N_19820,N_18784);
nor U20312 (N_20312,N_19988,N_19366);
nand U20313 (N_20313,N_18989,N_18415);
and U20314 (N_20314,N_18606,N_18847);
or U20315 (N_20315,N_18092,N_17999);
nor U20316 (N_20316,N_18401,N_18843);
nor U20317 (N_20317,N_18188,N_17775);
xnor U20318 (N_20318,N_19269,N_18922);
nor U20319 (N_20319,N_19888,N_18531);
or U20320 (N_20320,N_18563,N_17818);
nand U20321 (N_20321,N_19543,N_19534);
xor U20322 (N_20322,N_19498,N_18130);
and U20323 (N_20323,N_19321,N_19972);
xor U20324 (N_20324,N_18776,N_19397);
nand U20325 (N_20325,N_18738,N_18453);
xor U20326 (N_20326,N_17746,N_17866);
and U20327 (N_20327,N_18930,N_18572);
nor U20328 (N_20328,N_19470,N_19552);
and U20329 (N_20329,N_18422,N_19467);
nand U20330 (N_20330,N_18645,N_18495);
nor U20331 (N_20331,N_19870,N_19741);
nor U20332 (N_20332,N_19737,N_17777);
nand U20333 (N_20333,N_18583,N_18737);
nand U20334 (N_20334,N_19008,N_18216);
xor U20335 (N_20335,N_19853,N_19917);
or U20336 (N_20336,N_18054,N_19243);
and U20337 (N_20337,N_19540,N_19932);
nand U20338 (N_20338,N_19649,N_19713);
or U20339 (N_20339,N_19669,N_18329);
and U20340 (N_20340,N_19442,N_17942);
or U20341 (N_20341,N_17784,N_18074);
xnor U20342 (N_20342,N_17783,N_17668);
and U20343 (N_20343,N_18964,N_19041);
nor U20344 (N_20344,N_17884,N_19148);
nor U20345 (N_20345,N_18477,N_18426);
nor U20346 (N_20346,N_18909,N_18373);
nor U20347 (N_20347,N_19664,N_18065);
nand U20348 (N_20348,N_18535,N_19107);
or U20349 (N_20349,N_19194,N_18239);
xnor U20350 (N_20350,N_19233,N_19934);
or U20351 (N_20351,N_19368,N_18756);
nor U20352 (N_20352,N_18389,N_19987);
nor U20353 (N_20353,N_17838,N_17536);
nor U20354 (N_20354,N_19641,N_19058);
and U20355 (N_20355,N_18841,N_17706);
nor U20356 (N_20356,N_18322,N_18019);
nor U20357 (N_20357,N_18251,N_17526);
xor U20358 (N_20358,N_18267,N_19754);
and U20359 (N_20359,N_19309,N_18340);
xnor U20360 (N_20360,N_17887,N_18192);
xor U20361 (N_20361,N_17988,N_19123);
xnor U20362 (N_20362,N_18158,N_17869);
or U20363 (N_20363,N_18614,N_17843);
nand U20364 (N_20364,N_17860,N_19765);
or U20365 (N_20365,N_17745,N_18425);
and U20366 (N_20366,N_18736,N_19823);
or U20367 (N_20367,N_19050,N_18683);
nand U20368 (N_20368,N_18799,N_18755);
and U20369 (N_20369,N_17873,N_18597);
xor U20370 (N_20370,N_18852,N_18220);
and U20371 (N_20371,N_18107,N_19354);
xnor U20372 (N_20372,N_17859,N_17900);
nand U20373 (N_20373,N_18261,N_18386);
or U20374 (N_20374,N_19614,N_17689);
or U20375 (N_20375,N_17513,N_19109);
and U20376 (N_20376,N_18272,N_18298);
xor U20377 (N_20377,N_19398,N_19874);
nand U20378 (N_20378,N_18333,N_18118);
xor U20379 (N_20379,N_19202,N_19507);
xnor U20380 (N_20380,N_19261,N_19985);
nand U20381 (N_20381,N_18803,N_18475);
xnor U20382 (N_20382,N_19264,N_19124);
xnor U20383 (N_20383,N_19970,N_19967);
xor U20384 (N_20384,N_19005,N_18676);
nor U20385 (N_20385,N_17589,N_17837);
nor U20386 (N_20386,N_19372,N_19379);
nor U20387 (N_20387,N_18328,N_17677);
or U20388 (N_20388,N_19538,N_18432);
xnor U20389 (N_20389,N_18816,N_19625);
nor U20390 (N_20390,N_19954,N_17504);
xnor U20391 (N_20391,N_17708,N_17984);
and U20392 (N_20392,N_19572,N_19339);
and U20393 (N_20393,N_19239,N_18979);
nor U20394 (N_20394,N_19105,N_19979);
or U20395 (N_20395,N_19214,N_18526);
or U20396 (N_20396,N_18051,N_18617);
and U20397 (N_20397,N_18241,N_18076);
and U20398 (N_20398,N_19960,N_18097);
and U20399 (N_20399,N_18163,N_18160);
and U20400 (N_20400,N_19024,N_18741);
xnor U20401 (N_20401,N_19434,N_18973);
nand U20402 (N_20402,N_19341,N_17844);
or U20403 (N_20403,N_18915,N_17538);
and U20404 (N_20404,N_17765,N_19463);
nand U20405 (N_20405,N_19457,N_19998);
or U20406 (N_20406,N_19574,N_19436);
nand U20407 (N_20407,N_18926,N_17686);
and U20408 (N_20408,N_19302,N_18066);
and U20409 (N_20409,N_17618,N_19056);
and U20410 (N_20410,N_19471,N_18296);
or U20411 (N_20411,N_19530,N_18240);
nor U20412 (N_20412,N_17855,N_17658);
and U20413 (N_20413,N_18006,N_19171);
or U20414 (N_20414,N_17828,N_19184);
nand U20415 (N_20415,N_18421,N_19029);
nor U20416 (N_20416,N_19363,N_19139);
nor U20417 (N_20417,N_19078,N_18344);
or U20418 (N_20418,N_19150,N_19364);
xnor U20419 (N_20419,N_19373,N_17845);
nand U20420 (N_20420,N_18845,N_17652);
or U20421 (N_20421,N_19961,N_18031);
nand U20422 (N_20422,N_19714,N_18888);
or U20423 (N_20423,N_19396,N_19630);
or U20424 (N_20424,N_19413,N_19547);
nor U20425 (N_20425,N_19066,N_18615);
and U20426 (N_20426,N_17815,N_18302);
xnor U20427 (N_20427,N_17862,N_19964);
and U20428 (N_20428,N_19742,N_19941);
and U20429 (N_20429,N_19769,N_17902);
and U20430 (N_20430,N_18150,N_19634);
or U20431 (N_20431,N_19554,N_19663);
and U20432 (N_20432,N_18236,N_18913);
xor U20433 (N_20433,N_18233,N_17835);
nor U20434 (N_20434,N_18294,N_18213);
nor U20435 (N_20435,N_17546,N_17703);
xor U20436 (N_20436,N_19183,N_18780);
nand U20437 (N_20437,N_19445,N_19210);
xnor U20438 (N_20438,N_18636,N_18323);
and U20439 (N_20439,N_17759,N_19484);
or U20440 (N_20440,N_19835,N_17931);
and U20441 (N_20441,N_17685,N_18480);
xnor U20442 (N_20442,N_18669,N_18468);
and U20443 (N_20443,N_19289,N_19735);
or U20444 (N_20444,N_17565,N_18007);
nor U20445 (N_20445,N_17551,N_18518);
or U20446 (N_20446,N_18248,N_18775);
nand U20447 (N_20447,N_19182,N_17595);
or U20448 (N_20448,N_18658,N_19883);
nor U20449 (N_20449,N_19746,N_18628);
xnor U20450 (N_20450,N_18134,N_18428);
xor U20451 (N_20451,N_18257,N_18953);
or U20452 (N_20452,N_17757,N_18624);
nand U20453 (N_20453,N_19745,N_19459);
and U20454 (N_20454,N_19673,N_19204);
nand U20455 (N_20455,N_19414,N_19991);
and U20456 (N_20456,N_18043,N_19525);
nor U20457 (N_20457,N_19394,N_18754);
nand U20458 (N_20458,N_19904,N_18285);
nand U20459 (N_20459,N_19848,N_17564);
xnor U20460 (N_20460,N_18452,N_19324);
or U20461 (N_20461,N_18517,N_19271);
nor U20462 (N_20462,N_18602,N_19096);
and U20463 (N_20463,N_19395,N_19027);
or U20464 (N_20464,N_18719,N_18897);
xnor U20465 (N_20465,N_18886,N_19019);
nand U20466 (N_20466,N_17723,N_19215);
xor U20467 (N_20467,N_18721,N_19558);
or U20468 (N_20468,N_19077,N_19725);
nor U20469 (N_20469,N_18202,N_19175);
and U20470 (N_20470,N_19734,N_19580);
or U20471 (N_20471,N_19224,N_17570);
nor U20472 (N_20472,N_19352,N_17661);
nand U20473 (N_20473,N_18796,N_18772);
xor U20474 (N_20474,N_18955,N_17820);
xor U20475 (N_20475,N_18590,N_19062);
nand U20476 (N_20476,N_19326,N_19730);
xor U20477 (N_20477,N_18377,N_19185);
nand U20478 (N_20478,N_18574,N_18260);
nor U20479 (N_20479,N_19900,N_18594);
nor U20480 (N_20480,N_17958,N_17605);
nand U20481 (N_20481,N_18911,N_18871);
nor U20482 (N_20482,N_18621,N_18805);
or U20483 (N_20483,N_19042,N_18752);
nor U20484 (N_20484,N_19280,N_19104);
and U20485 (N_20485,N_19698,N_19167);
nand U20486 (N_20486,N_18061,N_18731);
or U20487 (N_20487,N_18250,N_19478);
nand U20488 (N_20488,N_17610,N_19281);
and U20489 (N_20489,N_18375,N_18219);
and U20490 (N_20490,N_18991,N_17946);
nand U20491 (N_20491,N_18374,N_19913);
or U20492 (N_20492,N_17607,N_19660);
nor U20493 (N_20493,N_18869,N_18607);
or U20494 (N_20494,N_18807,N_19662);
xor U20495 (N_20495,N_19432,N_19849);
or U20496 (N_20496,N_19517,N_19376);
or U20497 (N_20497,N_17679,N_18451);
and U20498 (N_20498,N_18555,N_19187);
nor U20499 (N_20499,N_19495,N_19242);
nor U20500 (N_20500,N_18893,N_17671);
xnor U20501 (N_20501,N_19130,N_19750);
or U20502 (N_20502,N_19253,N_19889);
nand U20503 (N_20503,N_19501,N_19494);
and U20504 (N_20504,N_18640,N_19119);
and U20505 (N_20505,N_18112,N_18703);
nor U20506 (N_20506,N_19997,N_18039);
nand U20507 (N_20507,N_18912,N_17774);
nor U20508 (N_20508,N_18960,N_19013);
nand U20509 (N_20509,N_19620,N_18638);
or U20510 (N_20510,N_18511,N_17728);
nand U20511 (N_20511,N_18387,N_19772);
nor U20512 (N_20512,N_19251,N_18898);
or U20513 (N_20513,N_19252,N_19497);
nand U20514 (N_20514,N_19778,N_17949);
nor U20515 (N_20515,N_18734,N_19824);
and U20516 (N_20516,N_18727,N_18811);
xnor U20517 (N_20517,N_18494,N_17576);
nor U20518 (N_20518,N_19385,N_19615);
xor U20519 (N_20519,N_19468,N_18810);
or U20520 (N_20520,N_17615,N_18968);
xnor U20521 (N_20521,N_17563,N_19877);
xnor U20522 (N_20522,N_18459,N_17506);
nand U20523 (N_20523,N_19303,N_19064);
and U20524 (N_20524,N_18032,N_17522);
and U20525 (N_20525,N_17724,N_19661);
and U20526 (N_20526,N_17616,N_18190);
xnor U20527 (N_20527,N_18224,N_19402);
and U20528 (N_20528,N_19080,N_19378);
nand U20529 (N_20529,N_19629,N_17764);
or U20530 (N_20530,N_17795,N_19144);
or U20531 (N_20531,N_19179,N_18782);
nor U20532 (N_20532,N_19923,N_19516);
nor U20533 (N_20533,N_19108,N_17748);
xnor U20534 (N_20534,N_19276,N_18080);
and U20535 (N_20535,N_18728,N_19431);
nor U20536 (N_20536,N_18193,N_18410);
or U20537 (N_20537,N_19821,N_18806);
nor U20538 (N_20538,N_19755,N_19959);
and U20539 (N_20539,N_18457,N_19311);
and U20540 (N_20540,N_17771,N_17647);
or U20541 (N_20541,N_18277,N_18237);
or U20542 (N_20542,N_18385,N_19097);
nor U20543 (N_20543,N_17656,N_19916);
and U20544 (N_20544,N_19018,N_18739);
nand U20545 (N_20545,N_17932,N_18433);
nand U20546 (N_20546,N_17596,N_17854);
nor U20547 (N_20547,N_19999,N_19375);
and U20548 (N_20548,N_19551,N_19350);
nand U20549 (N_20549,N_18050,N_18037);
nor U20550 (N_20550,N_19635,N_18132);
nand U20551 (N_20551,N_18513,N_18997);
xnor U20552 (N_20552,N_19984,N_18826);
nand U20553 (N_20553,N_17877,N_19502);
or U20554 (N_20554,N_19938,N_18141);
and U20555 (N_20555,N_18712,N_19881);
nor U20556 (N_20556,N_18147,N_18836);
nand U20557 (N_20557,N_19560,N_19217);
xor U20558 (N_20558,N_18882,N_18411);
xor U20559 (N_20559,N_19520,N_18503);
and U20560 (N_20560,N_18750,N_17559);
and U20561 (N_20561,N_18838,N_18418);
nor U20562 (N_20562,N_17832,N_19860);
nor U20563 (N_20563,N_18789,N_18467);
or U20564 (N_20564,N_18356,N_19440);
nor U20565 (N_20565,N_17907,N_18367);
or U20566 (N_20566,N_19377,N_19260);
xnor U20567 (N_20567,N_19724,N_18360);
or U20568 (N_20568,N_19453,N_19535);
xnor U20569 (N_20569,N_17809,N_19528);
nor U20570 (N_20570,N_19910,N_18315);
xnor U20571 (N_20571,N_18447,N_18209);
nand U20572 (N_20572,N_18108,N_17648);
or U20573 (N_20573,N_17707,N_19246);
xnor U20574 (N_20574,N_17641,N_18441);
nor U20575 (N_20575,N_18345,N_19869);
nand U20576 (N_20576,N_17628,N_18641);
xor U20577 (N_20577,N_19792,N_19325);
nor U20578 (N_20578,N_18497,N_18131);
or U20579 (N_20579,N_18346,N_18996);
nor U20580 (N_20580,N_18529,N_19656);
nor U20581 (N_20581,N_18116,N_19245);
or U20582 (N_20582,N_18048,N_17841);
xnor U20583 (N_20583,N_19863,N_18288);
and U20584 (N_20584,N_17974,N_19912);
nor U20585 (N_20585,N_19599,N_19529);
or U20586 (N_20586,N_18149,N_18357);
or U20587 (N_20587,N_19971,N_17788);
nand U20588 (N_20588,N_19565,N_17731);
xor U20589 (N_20589,N_18487,N_17966);
nand U20590 (N_20590,N_17639,N_18212);
xor U20591 (N_20591,N_18458,N_18264);
or U20592 (N_20592,N_19367,N_19085);
nor U20593 (N_20593,N_19989,N_18170);
or U20594 (N_20594,N_19323,N_18263);
or U20595 (N_20595,N_18648,N_18378);
and U20596 (N_20596,N_17673,N_19141);
or U20597 (N_20597,N_18765,N_18598);
nand U20598 (N_20598,N_18577,N_17700);
nand U20599 (N_20599,N_18026,N_18763);
or U20600 (N_20600,N_18903,N_18191);
nor U20601 (N_20601,N_18126,N_18382);
nand U20602 (N_20602,N_18365,N_18876);
xor U20603 (N_20603,N_19312,N_19801);
xnor U20604 (N_20604,N_17881,N_17567);
nor U20605 (N_20605,N_17971,N_17794);
xor U20606 (N_20606,N_17678,N_19624);
nand U20607 (N_20607,N_18873,N_19990);
or U20608 (N_20608,N_18228,N_19858);
or U20609 (N_20609,N_17763,N_19541);
and U20610 (N_20610,N_19462,N_19747);
and U20611 (N_20611,N_19958,N_19392);
nor U20612 (N_20612,N_19688,N_18924);
nor U20613 (N_20613,N_19071,N_19068);
or U20614 (N_20614,N_19645,N_17782);
and U20615 (N_20615,N_18084,N_19996);
nor U20616 (N_20616,N_18859,N_19283);
xor U20617 (N_20617,N_19717,N_18933);
nand U20618 (N_20618,N_18435,N_17917);
and U20619 (N_20619,N_17827,N_19165);
and U20620 (N_20620,N_18098,N_19784);
xor U20621 (N_20621,N_19169,N_18012);
or U20622 (N_20622,N_18354,N_19584);
or U20623 (N_20623,N_19481,N_18448);
nor U20624 (N_20624,N_18274,N_19493);
nand U20625 (N_20625,N_17534,N_17868);
nor U20626 (N_20626,N_19749,N_17976);
nand U20627 (N_20627,N_17542,N_17510);
or U20628 (N_20628,N_18232,N_18341);
nand U20629 (N_20629,N_17786,N_18767);
nor U20630 (N_20630,N_18148,N_17554);
and U20631 (N_20631,N_18297,N_18370);
and U20632 (N_20632,N_19524,N_17726);
and U20633 (N_20633,N_18445,N_17798);
nand U20634 (N_20634,N_19802,N_17735);
nand U20635 (N_20635,N_19568,N_19051);
xor U20636 (N_20636,N_19512,N_19149);
nand U20637 (N_20637,N_18085,N_18429);
and U20638 (N_20638,N_17553,N_19719);
and U20639 (N_20639,N_18866,N_19294);
nand U20640 (N_20640,N_18963,N_19258);
nand U20641 (N_20641,N_19948,N_18753);
or U20642 (N_20642,N_18543,N_18637);
xnor U20643 (N_20643,N_18593,N_18273);
nand U20644 (N_20644,N_17730,N_18409);
nor U20645 (N_20645,N_17676,N_18946);
nand U20646 (N_20646,N_19696,N_18591);
xnor U20647 (N_20647,N_18321,N_18660);
or U20648 (N_20648,N_19129,N_18542);
and U20649 (N_20649,N_19346,N_17861);
nor U20650 (N_20650,N_19943,N_17948);
nor U20651 (N_20651,N_18183,N_18708);
nor U20652 (N_20652,N_19158,N_17852);
nand U20653 (N_20653,N_18493,N_17592);
or U20654 (N_20654,N_19491,N_19639);
xnor U20655 (N_20655,N_18253,N_18090);
xor U20656 (N_20656,N_18525,N_18159);
nor U20657 (N_20657,N_18064,N_19089);
nor U20658 (N_20658,N_17889,N_18974);
and U20659 (N_20659,N_18046,N_19273);
nor U20660 (N_20660,N_19808,N_19667);
and U20661 (N_20661,N_19919,N_18123);
and U20662 (N_20662,N_19222,N_19727);
and U20663 (N_20663,N_18665,N_18510);
nand U20664 (N_20664,N_18180,N_19036);
or U20665 (N_20665,N_17830,N_18245);
nor U20666 (N_20666,N_17939,N_18397);
nand U20667 (N_20667,N_19338,N_17737);
and U20668 (N_20668,N_19845,N_18726);
and U20669 (N_20669,N_18186,N_19797);
nor U20670 (N_20670,N_17699,N_19371);
and U20671 (N_20671,N_19736,N_18889);
and U20672 (N_20672,N_19254,N_17959);
and U20673 (N_20673,N_17633,N_18830);
xor U20674 (N_20674,N_19240,N_19315);
or U20675 (N_20675,N_19733,N_18177);
xor U20676 (N_20676,N_17760,N_19774);
or U20677 (N_20677,N_18299,N_18733);
nor U20678 (N_20678,N_18860,N_19247);
and U20679 (N_20679,N_17560,N_18589);
nand U20680 (N_20680,N_19995,N_19045);
xnor U20681 (N_20681,N_18961,N_19191);
or U20682 (N_20682,N_19111,N_19403);
nor U20683 (N_20683,N_18289,N_19739);
or U20684 (N_20684,N_17529,N_18573);
nor U20685 (N_20685,N_19090,N_18646);
nor U20686 (N_20686,N_17836,N_17875);
nand U20687 (N_20687,N_18821,N_18546);
and U20688 (N_20688,N_19676,N_18596);
or U20689 (N_20689,N_18479,N_17594);
xnor U20690 (N_20690,N_19931,N_18450);
nor U20691 (N_20691,N_19244,N_19015);
nand U20692 (N_20692,N_17920,N_19703);
nor U20693 (N_20693,N_19816,N_19017);
and U20694 (N_20694,N_19890,N_19762);
nand U20695 (N_20695,N_17583,N_19083);
xor U20696 (N_20696,N_18301,N_18388);
or U20697 (N_20697,N_17865,N_19216);
or U20698 (N_20698,N_19197,N_18501);
or U20699 (N_20699,N_17768,N_18891);
and U20700 (N_20700,N_18742,N_19776);
xor U20701 (N_20701,N_18896,N_18778);
and U20702 (N_20702,N_19782,N_19631);
xor U20703 (N_20703,N_19740,N_17709);
or U20704 (N_20704,N_19648,N_17823);
or U20705 (N_20705,N_19830,N_19199);
nor U20706 (N_20706,N_18196,N_19170);
or U20707 (N_20707,N_19844,N_17593);
or U20708 (N_20708,N_18072,N_18880);
xnor U20709 (N_20709,N_18530,N_19908);
xnor U20710 (N_20710,N_18700,N_18094);
and U20711 (N_20711,N_17990,N_19865);
nand U20712 (N_20712,N_19065,N_18105);
nand U20713 (N_20713,N_17885,N_19899);
nand U20714 (N_20714,N_19032,N_18313);
nand U20715 (N_20715,N_19700,N_19708);
xor U20716 (N_20716,N_19570,N_17621);
xnor U20717 (N_20717,N_17547,N_17945);
nor U20718 (N_20718,N_18920,N_18400);
nand U20719 (N_20719,N_19637,N_17813);
and U20720 (N_20720,N_17955,N_19460);
and U20721 (N_20721,N_19929,N_18863);
and U20722 (N_20722,N_18379,N_19387);
xnor U20723 (N_20723,N_18610,N_17599);
or U20724 (N_20724,N_19646,N_18595);
or U20725 (N_20725,N_19153,N_18632);
nand U20726 (N_20726,N_19349,N_19137);
or U20727 (N_20727,N_19681,N_19795);
nor U20728 (N_20728,N_17817,N_18947);
nand U20729 (N_20729,N_19422,N_19920);
nor U20730 (N_20730,N_19465,N_18992);
xnor U20731 (N_20731,N_19308,N_18802);
or U20732 (N_20732,N_18015,N_17627);
and U20733 (N_20733,N_18870,N_19783);
and U20734 (N_20734,N_19622,N_19317);
or U20735 (N_20735,N_17776,N_19049);
nor U20736 (N_20736,N_17670,N_19026);
nor U20737 (N_20737,N_18460,N_19786);
nand U20738 (N_20738,N_17825,N_18609);
xor U20739 (N_20739,N_17928,N_19441);
nand U20740 (N_20740,N_18206,N_17752);
nand U20741 (N_20741,N_19355,N_18465);
nor U20742 (N_20742,N_19521,N_17982);
and U20743 (N_20743,N_17986,N_17631);
nor U20744 (N_20744,N_18197,N_17743);
xor U20745 (N_20745,N_19705,N_19203);
or U20746 (N_20746,N_17964,N_19469);
and U20747 (N_20747,N_19775,N_19435);
or U20748 (N_20748,N_18850,N_17625);
xor U20749 (N_20749,N_19651,N_19052);
nor U20750 (N_20750,N_18857,N_19607);
or U20751 (N_20751,N_17908,N_18901);
nor U20752 (N_20752,N_18635,N_17756);
or U20753 (N_20753,N_18713,N_18420);
xor U20754 (N_20754,N_18372,N_17502);
and U20755 (N_20755,N_18720,N_18124);
and U20756 (N_20756,N_18399,N_18940);
and U20757 (N_20757,N_18582,N_18694);
xnor U20758 (N_20758,N_19348,N_18173);
xor U20759 (N_20759,N_19956,N_17626);
and U20760 (N_20760,N_18010,N_17918);
or U20761 (N_20761,N_17772,N_19248);
nand U20762 (N_20762,N_18463,N_18438);
nand U20763 (N_20763,N_19595,N_18514);
xor U20764 (N_20764,N_17521,N_18104);
xnor U20765 (N_20765,N_19697,N_17511);
nor U20766 (N_20766,N_18620,N_17525);
or U20767 (N_20767,N_18879,N_18709);
and U20768 (N_20768,N_18521,N_18293);
and U20769 (N_20769,N_19070,N_19409);
xor U20770 (N_20770,N_19408,N_17503);
nor U20771 (N_20771,N_17587,N_18199);
nor U20772 (N_20772,N_19892,N_17960);
nand U20773 (N_20773,N_18622,N_18663);
nor U20774 (N_20774,N_18835,N_18578);
xor U20775 (N_20775,N_18654,N_17961);
and U20776 (N_20776,N_18238,N_17919);
and U20777 (N_20777,N_18994,N_17856);
and U20778 (N_20778,N_19331,N_18941);
and U20779 (N_20779,N_19826,N_19359);
or U20780 (N_20780,N_17696,N_18443);
nand U20781 (N_20781,N_18127,N_18198);
nor U20782 (N_20782,N_17512,N_19946);
nand U20783 (N_20783,N_17803,N_17808);
nor U20784 (N_20784,N_18431,N_18348);
nor U20785 (N_20785,N_19619,N_19053);
and U20786 (N_20786,N_19038,N_19126);
and U20787 (N_20787,N_19353,N_18532);
nor U20788 (N_20788,N_19300,N_17829);
and U20789 (N_20789,N_19712,N_17691);
or U20790 (N_20790,N_19973,N_18758);
or U20791 (N_20791,N_19880,N_19103);
and U20792 (N_20792,N_19365,N_18707);
and U20793 (N_20793,N_19650,N_18178);
nand U20794 (N_20794,N_19608,N_19113);
xor U20795 (N_20795,N_19933,N_18502);
or U20796 (N_20796,N_18316,N_17934);
nand U20797 (N_20797,N_18427,N_19344);
nand U20798 (N_20798,N_19265,N_18152);
nand U20799 (N_20799,N_17727,N_19581);
xor U20800 (N_20800,N_18928,N_18839);
xor U20801 (N_20801,N_18414,N_17840);
nor U20802 (N_20802,N_19449,N_18217);
or U20803 (N_20803,N_19598,N_17601);
nor U20804 (N_20804,N_18639,N_18035);
xor U20805 (N_20805,N_18033,N_18706);
or U20806 (N_20806,N_19290,N_19337);
or U20807 (N_20807,N_18004,N_18246);
xnor U20808 (N_20808,N_17826,N_17688);
and U20809 (N_20809,N_17537,N_17557);
and U20810 (N_20810,N_17842,N_18603);
and U20811 (N_20811,N_18162,N_19174);
xnor U20812 (N_20812,N_18907,N_19451);
nor U20813 (N_20813,N_19262,N_17922);
xnor U20814 (N_20814,N_18657,N_18680);
and U20815 (N_20815,N_19505,N_19796);
or U20816 (N_20816,N_19768,N_18483);
and U20817 (N_20817,N_18705,N_19897);
nor U20818 (N_20818,N_18384,N_17804);
nand U20819 (N_20819,N_17962,N_19689);
or U20820 (N_20820,N_18942,N_18938);
and U20821 (N_20821,N_19328,N_17811);
and U20822 (N_20822,N_19694,N_18307);
or U20823 (N_20823,N_17545,N_18175);
nand U20824 (N_20824,N_19548,N_19944);
nand U20825 (N_20825,N_17640,N_17544);
and U20826 (N_20826,N_18710,N_19437);
and U20827 (N_20827,N_17792,N_19670);
nand U20828 (N_20828,N_19575,N_18201);
and U20829 (N_20829,N_19692,N_18993);
and U20830 (N_20830,N_19966,N_19578);
xnor U20831 (N_20831,N_18073,N_18349);
xor U20832 (N_20832,N_18314,N_17956);
nor U20833 (N_20833,N_18413,N_19037);
or U20834 (N_20834,N_18588,N_18030);
xor U20835 (N_20835,N_19110,N_19566);
nor U20836 (N_20836,N_17527,N_19691);
nor U20837 (N_20837,N_18723,N_18895);
nand U20838 (N_20838,N_19456,N_18662);
or U20839 (N_20839,N_18456,N_19274);
xor U20840 (N_20840,N_18496,N_19304);
and U20841 (N_20841,N_18988,N_19582);
xor U20842 (N_20842,N_17501,N_18393);
and U20843 (N_20843,N_19488,N_18211);
nor U20844 (N_20844,N_18476,N_19709);
nand U20845 (N_20845,N_17634,N_18575);
xnor U20846 (N_20846,N_17635,N_18956);
nor U20847 (N_20847,N_18862,N_18892);
and U20848 (N_20848,N_17997,N_18692);
and U20849 (N_20849,N_18437,N_19332);
nand U20850 (N_20850,N_18691,N_18867);
or U20851 (N_20851,N_17993,N_18848);
nand U20852 (N_20852,N_19002,N_18698);
nor U20853 (N_20853,N_17890,N_19012);
xor U20854 (N_20854,N_19771,N_18109);
nand U20855 (N_20855,N_19228,N_18167);
xnor U20856 (N_20856,N_18036,N_18486);
nand U20857 (N_20857,N_19886,N_19542);
xor U20858 (N_20858,N_19307,N_18777);
and U20859 (N_20859,N_19500,N_18976);
and U20860 (N_20860,N_17806,N_17754);
nand U20861 (N_20861,N_19977,N_19299);
or U20862 (N_20862,N_19852,N_18101);
nand U20863 (N_20863,N_18258,N_18368);
xor U20864 (N_20864,N_18339,N_17936);
xor U20865 (N_20865,N_19640,N_17882);
or U20866 (N_20866,N_18068,N_18137);
nand U20867 (N_20867,N_17916,N_19115);
and U20868 (N_20868,N_18675,N_19060);
and U20869 (N_20869,N_19642,N_19121);
xnor U20870 (N_20870,N_18235,N_18275);
and U20871 (N_20871,N_18972,N_18398);
xor U20872 (N_20872,N_19145,N_17588);
nand U20873 (N_20873,N_18390,N_18616);
xnor U20874 (N_20874,N_17880,N_19851);
nor U20875 (N_20875,N_17721,N_19647);
xor U20876 (N_20876,N_18905,N_17505);
nand U20877 (N_20877,N_17617,N_19983);
nand U20878 (N_20878,N_18169,N_19162);
nand U20879 (N_20879,N_18625,N_17540);
or U20880 (N_20880,N_19010,N_19924);
nand U20881 (N_20881,N_19962,N_18056);
or U20882 (N_20882,N_18060,N_19539);
or U20883 (N_20883,N_17704,N_19942);
and U20884 (N_20884,N_17897,N_18541);
and U20885 (N_20885,N_19425,N_19935);
nand U20886 (N_20886,N_19592,N_18310);
and U20887 (N_20887,N_18854,N_19623);
xor U20888 (N_20888,N_19872,N_18552);
and U20889 (N_20889,N_18182,N_18471);
nand U20890 (N_20890,N_19152,N_18049);
nor U20891 (N_20891,N_19067,N_19760);
nor U20892 (N_20892,N_17552,N_18877);
xnor U20893 (N_20893,N_19100,N_19480);
xnor U20894 (N_20894,N_17548,N_17750);
nor U20895 (N_20895,N_18674,N_18761);
nand U20896 (N_20896,N_18009,N_19292);
xor U20897 (N_20897,N_17812,N_19483);
nor U20898 (N_20898,N_18945,N_18335);
nand U20899 (N_20899,N_19128,N_19168);
and U20900 (N_20900,N_18672,N_18504);
xor U20901 (N_20901,N_18643,N_18305);
nand U20902 (N_20902,N_18488,N_19915);
xor U20903 (N_20903,N_18364,N_18243);
nand U20904 (N_20904,N_18948,N_19361);
and U20905 (N_20905,N_19585,N_19023);
nand U20906 (N_20906,N_18135,N_18817);
or U20907 (N_20907,N_18599,N_17651);
nor U20908 (N_20908,N_19690,N_18950);
nor U20909 (N_20909,N_17539,N_19731);
or U20910 (N_20910,N_18849,N_18045);
nand U20911 (N_20911,N_19255,N_18667);
nand U20912 (N_20912,N_18278,N_18548);
or U20913 (N_20913,N_18083,N_19048);
or U20914 (N_20914,N_19362,N_19464);
nand U20915 (N_20915,N_18087,N_18536);
nand U20916 (N_20916,N_17751,N_18954);
or U20917 (N_20917,N_19207,N_18355);
xor U20918 (N_20918,N_17941,N_19738);
or U20919 (N_20919,N_19752,N_19429);
nand U20920 (N_20920,N_18560,N_18790);
and U20921 (N_20921,N_17532,N_18781);
xnor U20922 (N_20922,N_18362,N_19723);
nand U20923 (N_20923,N_18856,N_18516);
or U20924 (N_20924,N_18286,N_18874);
or U20925 (N_20925,N_18528,N_18815);
and U20926 (N_20926,N_17857,N_18808);
xnor U20927 (N_20927,N_18185,N_19593);
or U20928 (N_20928,N_18020,N_18885);
nor U20929 (N_20929,N_19072,N_19559);
nor U20930 (N_20930,N_19257,N_18965);
nor U20931 (N_20931,N_19282,N_18819);
nand U20932 (N_20932,N_17923,N_19701);
xnor U20933 (N_20933,N_18022,N_17883);
nor U20934 (N_20934,N_17667,N_19059);
and U20935 (N_20935,N_18295,N_18078);
and U20936 (N_20936,N_18760,N_19825);
xnor U20937 (N_20937,N_18469,N_18265);
and U20938 (N_20938,N_19685,N_18579);
and U20939 (N_20939,N_19025,N_19117);
and U20940 (N_20940,N_19838,N_17683);
and U20941 (N_20941,N_18661,N_17944);
nand U20942 (N_20942,N_18633,N_19232);
or U20943 (N_20943,N_19427,N_19086);
nand U20944 (N_20944,N_18673,N_17899);
nor U20945 (N_20945,N_17951,N_19278);
nor U20946 (N_20946,N_17910,N_19226);
and U20947 (N_20947,N_18951,N_19855);
nor U20948 (N_20948,N_19098,N_18725);
nand U20949 (N_20949,N_18139,N_18801);
xnor U20950 (N_20950,N_18102,N_18918);
nand U20951 (N_20951,N_18969,N_19907);
xor U20952 (N_20952,N_18093,N_19122);
and U20953 (N_20953,N_18462,N_18279);
or U20954 (N_20954,N_19430,N_19223);
xnor U20955 (N_20955,N_17681,N_18580);
nand U20956 (N_20956,N_17717,N_17849);
nand U20957 (N_20957,N_19922,N_19156);
and U20958 (N_20958,N_19043,N_19930);
nand U20959 (N_20959,N_17568,N_17566);
or U20960 (N_20960,N_18980,N_18336);
xnor U20961 (N_20961,N_19600,N_18685);
and U20962 (N_20962,N_17773,N_17541);
and U20963 (N_20963,N_19138,N_19330);
or U20964 (N_20964,N_19658,N_18934);
xnor U20965 (N_20965,N_17687,N_17965);
and U20966 (N_20966,N_18935,N_18266);
nand U20967 (N_20967,N_19411,N_19610);
nor U20968 (N_20968,N_19659,N_18522);
xnor U20969 (N_20969,N_18982,N_18868);
or U20970 (N_20970,N_19000,N_19926);
nor U20971 (N_20971,N_19275,N_18125);
nand U20972 (N_20972,N_18187,N_18440);
xor U20973 (N_20973,N_19485,N_18247);
nand U20974 (N_20974,N_19301,N_19418);
xor U20975 (N_20975,N_19953,N_19986);
and U20976 (N_20976,N_18417,N_19556);
xnor U20977 (N_20977,N_18786,N_19461);
nor U20978 (N_20978,N_19859,N_18484);
nand U20979 (N_20979,N_19176,N_18113);
and U20980 (N_20980,N_18647,N_18679);
nor U20981 (N_20981,N_19894,N_18686);
and U20982 (N_20982,N_19320,N_19770);
nor U20983 (N_20983,N_17528,N_19209);
nand U20984 (N_20984,N_18746,N_17952);
nand U20985 (N_20985,N_18792,N_19847);
or U20986 (N_20986,N_19683,N_17644);
nand U20987 (N_20987,N_18229,N_18804);
and U20988 (N_20988,N_18223,N_19277);
xor U20989 (N_20989,N_19472,N_19486);
xnor U20990 (N_20990,N_18858,N_18337);
nor U20991 (N_20991,N_19135,N_18770);
and U20992 (N_20992,N_19587,N_18047);
xnor U20993 (N_20993,N_18923,N_18136);
and U20994 (N_20994,N_18748,N_19004);
and U20995 (N_20995,N_17543,N_19477);
xor U20996 (N_20996,N_19155,N_19790);
nand U20997 (N_20997,N_18119,N_19230);
xor U20998 (N_20998,N_18990,N_19514);
and U20999 (N_20999,N_19073,N_17864);
nor U21000 (N_21000,N_19843,N_17602);
and U21001 (N_21001,N_18523,N_19718);
and U21002 (N_21002,N_19744,N_18208);
xnor U21003 (N_21003,N_18571,N_19270);
xor U21004 (N_21004,N_18696,N_19020);
nand U21005 (N_21005,N_19031,N_17802);
nand U21006 (N_21006,N_17584,N_17954);
nor U21007 (N_21007,N_19380,N_19220);
nand U21008 (N_21008,N_19021,N_19613);
nand U21009 (N_21009,N_17947,N_19597);
nor U21010 (N_21010,N_18392,N_17787);
nand U21011 (N_21011,N_18013,N_19310);
nand U21012 (N_21012,N_19438,N_17530);
nand U21013 (N_21013,N_18612,N_19759);
or U21014 (N_21014,N_18195,N_19612);
nor U21015 (N_21015,N_18077,N_18008);
nor U21016 (N_21016,N_19443,N_17892);
nor U21017 (N_21017,N_18300,N_17591);
nand U21018 (N_21018,N_18326,N_18281);
nor U21019 (N_21019,N_19322,N_18276);
and U21020 (N_21020,N_18383,N_19218);
or U21021 (N_21021,N_19028,N_17624);
xnor U21022 (N_21022,N_19114,N_18416);
and U21023 (N_21023,N_19200,N_19644);
and U21024 (N_21024,N_19743,N_19779);
and U21025 (N_21025,N_17816,N_19420);
xnor U21026 (N_21026,N_18342,N_19716);
xnor U21027 (N_21027,N_17569,N_19131);
nor U21028 (N_21028,N_18773,N_19161);
and U21029 (N_21029,N_17517,N_17500);
nand U21030 (N_21030,N_19452,N_17879);
xor U21031 (N_21031,N_17515,N_18482);
and U21032 (N_21032,N_19857,N_18204);
and U21033 (N_21033,N_18890,N_18430);
xnor U21034 (N_21034,N_18914,N_18505);
and U21035 (N_21035,N_17549,N_17903);
and U21036 (N_21036,N_19225,N_19636);
nor U21037 (N_21037,N_19879,N_19981);
nand U21038 (N_21038,N_17933,N_19259);
and U21039 (N_21039,N_18566,N_17749);
xnor U21040 (N_21040,N_19305,N_18304);
nand U21041 (N_21041,N_19212,N_18121);
nor U21042 (N_21042,N_18519,N_17912);
xnor U21043 (N_21043,N_18255,N_18498);
and U21044 (N_21044,N_17940,N_18559);
xnor U21045 (N_21045,N_18318,N_19678);
nor U21046 (N_21046,N_18878,N_17597);
and U21047 (N_21047,N_19617,N_18270);
nand U21048 (N_21048,N_18644,N_18768);
or U21049 (N_21049,N_17789,N_17744);
xor U21050 (N_21050,N_18153,N_19356);
nand U21051 (N_21051,N_19722,N_18214);
or U21052 (N_21052,N_18334,N_19160);
xnor U21053 (N_21053,N_18724,N_17913);
or U21054 (N_21054,N_19416,N_18900);
nor U21055 (N_21055,N_19417,N_18174);
nor U21056 (N_21056,N_19827,N_18743);
or U21057 (N_21057,N_19033,N_17571);
nand U21058 (N_21058,N_17807,N_18711);
or U21059 (N_21059,N_19166,N_19611);
and U21060 (N_21060,N_19333,N_18537);
nor U21061 (N_21061,N_18613,N_19594);
nand U21062 (N_21062,N_19401,N_18063);
nand U21063 (N_21063,N_19975,N_18919);
or U21064 (N_21064,N_19909,N_19814);
nand U21065 (N_21065,N_19911,N_18693);
nor U21066 (N_21066,N_19016,N_19142);
or U21067 (N_21067,N_17781,N_18038);
nand U21068 (N_21068,N_19533,N_18489);
nand U21069 (N_21069,N_19205,N_17810);
xor U21070 (N_21070,N_17556,N_19891);
and U21071 (N_21071,N_18829,N_19978);
nand U21072 (N_21072,N_19241,N_18749);
or U21073 (N_21073,N_19327,N_19127);
and U21074 (N_21074,N_19285,N_19069);
xor U21075 (N_21075,N_18282,N_17680);
nand U21076 (N_21076,N_19479,N_17769);
nor U21077 (N_21077,N_18454,N_18403);
and U21078 (N_21078,N_18837,N_19492);
and U21079 (N_21079,N_19178,N_19945);
nand U21080 (N_21080,N_18040,N_19674);
or U21081 (N_21081,N_18678,N_17665);
nor U21082 (N_21082,N_19229,N_18670);
nand U21083 (N_21083,N_19699,N_18684);
nand U21084 (N_21084,N_18254,N_18687);
xnor U21085 (N_21085,N_17968,N_18231);
nor U21086 (N_21086,N_18884,N_18466);
or U21087 (N_21087,N_17660,N_19789);
and U21088 (N_21088,N_17535,N_18200);
nor U21089 (N_21089,N_18822,N_19627);
or U21090 (N_21090,N_19099,N_19154);
and U21091 (N_21091,N_18626,N_18716);
or U21092 (N_21092,N_19968,N_19643);
or U21093 (N_21093,N_19903,N_19867);
or U21094 (N_21094,N_18902,N_17905);
nand U21095 (N_21095,N_18309,N_18110);
and U21096 (N_21096,N_17969,N_18481);
or U21097 (N_21097,N_19834,N_18967);
nand U21098 (N_21098,N_19856,N_17555);
nor U21099 (N_21099,N_19523,N_19345);
xor U21100 (N_21100,N_17819,N_18225);
nor U21101 (N_21101,N_17572,N_19092);
and U21102 (N_21102,N_17719,N_18256);
nand U21103 (N_21103,N_18520,N_19687);
xnor U21104 (N_21104,N_18027,N_18916);
xnor U21105 (N_21105,N_18133,N_19732);
nand U21106 (N_21106,N_17575,N_19399);
nor U21107 (N_21107,N_19291,N_19564);
nor U21108 (N_21108,N_17935,N_19157);
nand U21109 (N_21109,N_19604,N_18757);
and U21110 (N_21110,N_18194,N_18601);
xnor U21111 (N_21111,N_18405,N_19898);
xnor U21112 (N_21112,N_18568,N_17697);
or U21113 (N_21113,N_18629,N_18689);
nand U21114 (N_21114,N_17839,N_18176);
and U21115 (N_21115,N_19672,N_18556);
or U21116 (N_21116,N_18561,N_19287);
nand U21117 (N_21117,N_18512,N_17657);
and U21118 (N_21118,N_19815,N_17733);
nor U21119 (N_21119,N_17850,N_17779);
nand U21120 (N_21120,N_17509,N_18203);
nand U21121 (N_21121,N_17653,N_17577);
or U21122 (N_21122,N_17927,N_17514);
nand U21123 (N_21123,N_19473,N_18025);
or U21124 (N_21124,N_19057,N_18981);
nand U21125 (N_21125,N_18659,N_19125);
xnor U21126 (N_21126,N_17508,N_19423);
or U21127 (N_21127,N_17664,N_17780);
nor U21128 (N_21128,N_18688,N_18569);
xnor U21129 (N_21129,N_19231,N_18564);
xnor U21130 (N_21130,N_17725,N_18404);
or U21131 (N_21131,N_18016,N_18052);
xnor U21132 (N_21132,N_18959,N_18023);
or U21133 (N_21133,N_19876,N_19404);
or U21134 (N_21134,N_18444,N_18492);
xor U21135 (N_21135,N_17637,N_18331);
or U21136 (N_21136,N_19147,N_18650);
nand U21137 (N_21137,N_19235,N_18249);
nor U21138 (N_21138,N_18515,N_18910);
or U21139 (N_21139,N_19885,N_17878);
nor U21140 (N_21140,N_18062,N_19767);
or U21141 (N_21141,N_19720,N_19781);
xnor U21142 (N_21142,N_18798,N_18464);
or U21143 (N_21143,N_18283,N_17740);
nor U21144 (N_21144,N_17824,N_18787);
nor U21145 (N_21145,N_18081,N_19511);
xnor U21146 (N_21146,N_18699,N_19095);
nand U21147 (N_21147,N_19186,N_18576);
or U21148 (N_21148,N_17870,N_19424);
xnor U21149 (N_21149,N_17821,N_18984);
and U21150 (N_21150,N_17606,N_19448);
xnor U21151 (N_21151,N_18034,N_19854);
and U21152 (N_21152,N_19895,N_18144);
or U21153 (N_21153,N_18832,N_18971);
nand U21154 (N_21154,N_17822,N_19298);
nand U21155 (N_21155,N_18478,N_18995);
xnor U21156 (N_21156,N_19906,N_17893);
nand U21157 (N_21157,N_19267,N_17524);
xor U21158 (N_21158,N_17684,N_18584);
and U21159 (N_21159,N_19527,N_18604);
or U21160 (N_21160,N_19003,N_18164);
and U21161 (N_21161,N_18549,N_18262);
or U21162 (N_21162,N_19087,N_18605);
nand U21163 (N_21163,N_17767,N_19266);
and U21164 (N_21164,N_18853,N_17655);
nand U21165 (N_21165,N_18581,N_17558);
and U21166 (N_21166,N_18791,N_19711);
nand U21167 (N_21167,N_19173,N_19590);
and U21168 (N_21168,N_19133,N_19079);
and U21169 (N_21169,N_19407,N_19633);
xnor U21170 (N_21170,N_19370,N_19047);
xnor U21171 (N_21171,N_18320,N_18544);
or U21172 (N_21172,N_19293,N_19751);
xnor U21173 (N_21173,N_18002,N_18028);
nor U21174 (N_21174,N_17853,N_17801);
and U21175 (N_21175,N_18332,N_19504);
and U21176 (N_21176,N_19831,N_17519);
nor U21177 (N_21177,N_19579,N_17979);
nand U21178 (N_21178,N_18747,N_19707);
nor U21179 (N_21179,N_18507,N_19925);
nor U21180 (N_21180,N_18155,N_18618);
and U21181 (N_21181,N_18381,N_19728);
nor U21182 (N_21182,N_18252,N_18565);
nand U21183 (N_21183,N_18812,N_19351);
nand U21184 (N_21184,N_19256,N_18292);
and U21185 (N_21185,N_18844,N_17662);
nand U21186 (N_21186,N_18865,N_19503);
xor U21187 (N_21187,N_17693,N_19955);
and U21188 (N_21188,N_19657,N_19382);
nor U21189 (N_21189,N_18831,N_18534);
or U21190 (N_21190,N_18319,N_17977);
or U21191 (N_21191,N_17622,N_18407);
nand U21192 (N_21192,N_19819,N_19603);
or U21193 (N_21193,N_19074,N_18800);
nor U21194 (N_21194,N_19618,N_19693);
xnor U21195 (N_21195,N_18771,N_19421);
nand U21196 (N_21196,N_18655,N_19884);
nand U21197 (N_21197,N_18079,N_18324);
or U21198 (N_21198,N_18545,N_17604);
or U21199 (N_21199,N_19206,N_19882);
or U21200 (N_21200,N_19798,N_17650);
and U21201 (N_21201,N_17909,N_19695);
xor U21202 (N_21202,N_18704,N_18059);
and U21203 (N_21203,N_18011,N_17600);
or U21204 (N_21204,N_19976,N_18562);
or U21205 (N_21205,N_19563,N_17998);
nor U21206 (N_21206,N_18179,N_17578);
or U21207 (N_21207,N_17722,N_18539);
nor U21208 (N_21208,N_18470,N_19522);
xor U21209 (N_21209,N_19809,N_19902);
nor U21210 (N_21210,N_18058,N_18977);
nand U21211 (N_21211,N_19758,N_19901);
and U21212 (N_21212,N_19474,N_18142);
or U21213 (N_21213,N_19939,N_18527);
xor U21214 (N_21214,N_19756,N_18627);
nor U21215 (N_21215,N_18306,N_19677);
nand U21216 (N_21216,N_17561,N_18499);
or U21217 (N_21217,N_18442,N_17980);
nor U21218 (N_21218,N_17929,N_18861);
and U21219 (N_21219,N_19061,N_17613);
xor U21220 (N_21220,N_19314,N_19136);
nand U21221 (N_21221,N_18558,N_17533);
and U21222 (N_21222,N_17518,N_17985);
xnor U21223 (N_21223,N_17623,N_18656);
nand U21224 (N_21224,N_17715,N_19510);
or U21225 (N_21225,N_18814,N_18117);
nor U21226 (N_21226,N_18785,N_18567);
and U21227 (N_21227,N_18145,N_18975);
xor U21228 (N_21228,N_19553,N_18363);
nor U21229 (N_21229,N_19763,N_18221);
xor U21230 (N_21230,N_18550,N_19439);
and U21231 (N_21231,N_19878,N_19729);
xor U21232 (N_21232,N_17894,N_17585);
and U21233 (N_21233,N_18872,N_18055);
xnor U21234 (N_21234,N_18111,N_19686);
xor U21235 (N_21235,N_19602,N_18818);
xnor U21236 (N_21236,N_19828,N_19336);
and U21237 (N_21237,N_18939,N_19343);
nand U21238 (N_21238,N_17755,N_18908);
or U21239 (N_21239,N_18171,N_19766);
nand U21240 (N_21240,N_18181,N_17943);
and U21241 (N_21241,N_19181,N_19704);
nor U21242 (N_21242,N_19357,N_19710);
nor U21243 (N_21243,N_19596,N_18745);
nor U21244 (N_21244,N_17867,N_19841);
nor U21245 (N_21245,N_17682,N_17814);
xnor U21246 (N_21246,N_19134,N_19513);
xnor U21247 (N_21247,N_17562,N_19296);
nor U21248 (N_21248,N_19102,N_19666);
xor U21249 (N_21249,N_17925,N_17921);
and U21250 (N_21250,N_19918,N_19689);
and U21251 (N_21251,N_19060,N_19616);
or U21252 (N_21252,N_19484,N_19135);
nor U21253 (N_21253,N_17906,N_19352);
nor U21254 (N_21254,N_19197,N_18319);
nor U21255 (N_21255,N_18933,N_17749);
nor U21256 (N_21256,N_18806,N_19226);
or U21257 (N_21257,N_19771,N_17896);
nand U21258 (N_21258,N_19191,N_19949);
and U21259 (N_21259,N_19429,N_18020);
nand U21260 (N_21260,N_19978,N_19429);
xor U21261 (N_21261,N_17647,N_17911);
or U21262 (N_21262,N_19819,N_18619);
or U21263 (N_21263,N_18603,N_18453);
or U21264 (N_21264,N_18258,N_17516);
nand U21265 (N_21265,N_19555,N_18146);
nor U21266 (N_21266,N_19724,N_17524);
nand U21267 (N_21267,N_19705,N_17685);
xor U21268 (N_21268,N_19650,N_17531);
nand U21269 (N_21269,N_19620,N_17815);
nor U21270 (N_21270,N_18126,N_19230);
nor U21271 (N_21271,N_18063,N_17717);
nor U21272 (N_21272,N_19773,N_19319);
and U21273 (N_21273,N_17817,N_19132);
nand U21274 (N_21274,N_18677,N_19355);
or U21275 (N_21275,N_17738,N_19487);
nor U21276 (N_21276,N_17792,N_18807);
xor U21277 (N_21277,N_17908,N_18589);
or U21278 (N_21278,N_17689,N_19816);
nor U21279 (N_21279,N_19545,N_19390);
nor U21280 (N_21280,N_19999,N_19027);
nor U21281 (N_21281,N_19072,N_19768);
and U21282 (N_21282,N_19475,N_18924);
or U21283 (N_21283,N_18718,N_19333);
nand U21284 (N_21284,N_18218,N_18869);
nand U21285 (N_21285,N_17506,N_17537);
or U21286 (N_21286,N_19928,N_18386);
and U21287 (N_21287,N_18402,N_17998);
and U21288 (N_21288,N_18025,N_19100);
nand U21289 (N_21289,N_18190,N_19251);
xnor U21290 (N_21290,N_18072,N_18811);
nand U21291 (N_21291,N_17539,N_17727);
nor U21292 (N_21292,N_18807,N_18967);
xor U21293 (N_21293,N_19518,N_19419);
xnor U21294 (N_21294,N_18719,N_18584);
xor U21295 (N_21295,N_17638,N_18123);
nand U21296 (N_21296,N_18834,N_18612);
and U21297 (N_21297,N_19498,N_18278);
nor U21298 (N_21298,N_17607,N_18048);
nand U21299 (N_21299,N_18214,N_18766);
nand U21300 (N_21300,N_18531,N_19549);
or U21301 (N_21301,N_19270,N_19983);
or U21302 (N_21302,N_17745,N_18053);
xor U21303 (N_21303,N_18757,N_19244);
nor U21304 (N_21304,N_18572,N_17542);
nor U21305 (N_21305,N_19136,N_19502);
and U21306 (N_21306,N_18437,N_18830);
or U21307 (N_21307,N_19950,N_19342);
xnor U21308 (N_21308,N_17565,N_18076);
nor U21309 (N_21309,N_19539,N_17563);
xnor U21310 (N_21310,N_18089,N_18261);
xor U21311 (N_21311,N_19144,N_19355);
xor U21312 (N_21312,N_19168,N_19372);
xor U21313 (N_21313,N_19935,N_18349);
or U21314 (N_21314,N_18910,N_18464);
and U21315 (N_21315,N_18610,N_18570);
and U21316 (N_21316,N_17963,N_17785);
nand U21317 (N_21317,N_19439,N_17928);
and U21318 (N_21318,N_19868,N_19524);
xor U21319 (N_21319,N_19468,N_19323);
xnor U21320 (N_21320,N_18857,N_18029);
and U21321 (N_21321,N_19246,N_18565);
and U21322 (N_21322,N_18261,N_17738);
or U21323 (N_21323,N_17780,N_19578);
and U21324 (N_21324,N_18754,N_17798);
and U21325 (N_21325,N_19403,N_19514);
nand U21326 (N_21326,N_19752,N_17838);
xnor U21327 (N_21327,N_19364,N_18520);
and U21328 (N_21328,N_17717,N_19353);
or U21329 (N_21329,N_19813,N_19824);
nand U21330 (N_21330,N_18558,N_17909);
and U21331 (N_21331,N_18143,N_19991);
and U21332 (N_21332,N_17743,N_17535);
or U21333 (N_21333,N_19597,N_18710);
nor U21334 (N_21334,N_19132,N_18693);
nand U21335 (N_21335,N_17942,N_18422);
or U21336 (N_21336,N_19221,N_17644);
xnor U21337 (N_21337,N_17960,N_19033);
xor U21338 (N_21338,N_19290,N_18296);
nand U21339 (N_21339,N_18275,N_18732);
xnor U21340 (N_21340,N_17795,N_19067);
nor U21341 (N_21341,N_19424,N_18342);
nand U21342 (N_21342,N_17611,N_18405);
nand U21343 (N_21343,N_17821,N_19399);
nand U21344 (N_21344,N_19048,N_18979);
xnor U21345 (N_21345,N_19820,N_19036);
nor U21346 (N_21346,N_19463,N_17508);
or U21347 (N_21347,N_17705,N_19823);
or U21348 (N_21348,N_19639,N_19113);
xnor U21349 (N_21349,N_19331,N_18864);
nand U21350 (N_21350,N_18191,N_19171);
xor U21351 (N_21351,N_18899,N_19851);
nand U21352 (N_21352,N_17538,N_19933);
nand U21353 (N_21353,N_19712,N_17810);
or U21354 (N_21354,N_19163,N_17785);
or U21355 (N_21355,N_18130,N_17579);
xor U21356 (N_21356,N_18897,N_18846);
nor U21357 (N_21357,N_19116,N_18264);
xnor U21358 (N_21358,N_19369,N_19687);
xnor U21359 (N_21359,N_19163,N_19335);
nand U21360 (N_21360,N_18670,N_18460);
nor U21361 (N_21361,N_17864,N_18963);
nor U21362 (N_21362,N_19899,N_19694);
nor U21363 (N_21363,N_18669,N_18620);
nor U21364 (N_21364,N_18418,N_19975);
or U21365 (N_21365,N_17588,N_18508);
or U21366 (N_21366,N_18514,N_18440);
and U21367 (N_21367,N_18148,N_19318);
xnor U21368 (N_21368,N_19723,N_18431);
and U21369 (N_21369,N_19012,N_19234);
nor U21370 (N_21370,N_18972,N_19161);
nor U21371 (N_21371,N_19491,N_18835);
xnor U21372 (N_21372,N_19125,N_18857);
xor U21373 (N_21373,N_18275,N_18215);
xnor U21374 (N_21374,N_19118,N_19742);
nor U21375 (N_21375,N_18527,N_19306);
xnor U21376 (N_21376,N_18756,N_19834);
nor U21377 (N_21377,N_18538,N_19425);
nand U21378 (N_21378,N_17829,N_19316);
and U21379 (N_21379,N_19343,N_19083);
or U21380 (N_21380,N_19360,N_19082);
xnor U21381 (N_21381,N_18161,N_19186);
and U21382 (N_21382,N_17931,N_19942);
nor U21383 (N_21383,N_19635,N_18185);
xnor U21384 (N_21384,N_19323,N_17705);
and U21385 (N_21385,N_18191,N_18080);
or U21386 (N_21386,N_17940,N_17988);
or U21387 (N_21387,N_19410,N_17619);
xnor U21388 (N_21388,N_18096,N_17853);
xor U21389 (N_21389,N_17637,N_19058);
nand U21390 (N_21390,N_19018,N_18615);
or U21391 (N_21391,N_18686,N_18252);
nor U21392 (N_21392,N_19639,N_19923);
or U21393 (N_21393,N_17721,N_18801);
and U21394 (N_21394,N_18165,N_19507);
nand U21395 (N_21395,N_17781,N_17729);
nand U21396 (N_21396,N_19341,N_18273);
or U21397 (N_21397,N_19000,N_19813);
nand U21398 (N_21398,N_19129,N_19180);
xor U21399 (N_21399,N_19304,N_19622);
xor U21400 (N_21400,N_18325,N_19072);
nor U21401 (N_21401,N_18007,N_19928);
and U21402 (N_21402,N_18025,N_18252);
nand U21403 (N_21403,N_17754,N_19358);
nor U21404 (N_21404,N_19952,N_19333);
nor U21405 (N_21405,N_19500,N_19189);
or U21406 (N_21406,N_18677,N_19491);
xor U21407 (N_21407,N_17614,N_19687);
xnor U21408 (N_21408,N_19953,N_19857);
nor U21409 (N_21409,N_19453,N_18906);
xor U21410 (N_21410,N_19157,N_19769);
and U21411 (N_21411,N_17821,N_19172);
nand U21412 (N_21412,N_18690,N_18152);
or U21413 (N_21413,N_18204,N_17943);
nor U21414 (N_21414,N_17795,N_17571);
nor U21415 (N_21415,N_18371,N_18849);
nand U21416 (N_21416,N_18869,N_17586);
xnor U21417 (N_21417,N_19369,N_18237);
nor U21418 (N_21418,N_18128,N_17819);
nor U21419 (N_21419,N_17989,N_17962);
nand U21420 (N_21420,N_18694,N_17778);
xor U21421 (N_21421,N_18990,N_18947);
and U21422 (N_21422,N_19012,N_18779);
nand U21423 (N_21423,N_17963,N_18402);
and U21424 (N_21424,N_17590,N_18985);
nand U21425 (N_21425,N_19277,N_18702);
or U21426 (N_21426,N_19329,N_18206);
nand U21427 (N_21427,N_17922,N_19490);
nor U21428 (N_21428,N_18107,N_19289);
nor U21429 (N_21429,N_19443,N_19052);
xor U21430 (N_21430,N_17948,N_19791);
and U21431 (N_21431,N_19870,N_18266);
and U21432 (N_21432,N_18575,N_18595);
or U21433 (N_21433,N_17768,N_17692);
or U21434 (N_21434,N_19882,N_18719);
or U21435 (N_21435,N_19858,N_18020);
or U21436 (N_21436,N_19781,N_17910);
nand U21437 (N_21437,N_18765,N_18518);
nand U21438 (N_21438,N_18017,N_18319);
nand U21439 (N_21439,N_18928,N_17926);
or U21440 (N_21440,N_19130,N_17997);
or U21441 (N_21441,N_19137,N_19694);
or U21442 (N_21442,N_19978,N_19504);
xnor U21443 (N_21443,N_19343,N_18296);
nor U21444 (N_21444,N_17826,N_19929);
nor U21445 (N_21445,N_19241,N_18540);
xor U21446 (N_21446,N_19535,N_18581);
nand U21447 (N_21447,N_19764,N_18694);
nor U21448 (N_21448,N_18734,N_17803);
nand U21449 (N_21449,N_19892,N_19118);
xor U21450 (N_21450,N_19920,N_19503);
xor U21451 (N_21451,N_18871,N_19876);
nor U21452 (N_21452,N_19380,N_18841);
nor U21453 (N_21453,N_18022,N_19872);
xor U21454 (N_21454,N_19300,N_17941);
xnor U21455 (N_21455,N_19499,N_18074);
and U21456 (N_21456,N_19304,N_18844);
or U21457 (N_21457,N_18073,N_19831);
and U21458 (N_21458,N_18987,N_19255);
and U21459 (N_21459,N_18571,N_19753);
nand U21460 (N_21460,N_19149,N_18122);
nor U21461 (N_21461,N_19541,N_19613);
or U21462 (N_21462,N_18546,N_17807);
xor U21463 (N_21463,N_19593,N_17540);
nor U21464 (N_21464,N_18426,N_18637);
nor U21465 (N_21465,N_18137,N_19399);
and U21466 (N_21466,N_19459,N_19510);
xnor U21467 (N_21467,N_19079,N_18257);
nand U21468 (N_21468,N_18058,N_19708);
and U21469 (N_21469,N_19765,N_18687);
xor U21470 (N_21470,N_19134,N_18649);
xor U21471 (N_21471,N_18359,N_17714);
and U21472 (N_21472,N_18918,N_18089);
xnor U21473 (N_21473,N_19959,N_19188);
nand U21474 (N_21474,N_19082,N_17586);
and U21475 (N_21475,N_19377,N_19849);
nor U21476 (N_21476,N_19796,N_17689);
or U21477 (N_21477,N_17696,N_17655);
nor U21478 (N_21478,N_18659,N_19041);
xor U21479 (N_21479,N_19353,N_17861);
nand U21480 (N_21480,N_19883,N_19889);
or U21481 (N_21481,N_19560,N_18268);
and U21482 (N_21482,N_18293,N_18726);
xor U21483 (N_21483,N_19807,N_18764);
nor U21484 (N_21484,N_19242,N_18511);
and U21485 (N_21485,N_19704,N_18214);
or U21486 (N_21486,N_18999,N_18215);
xnor U21487 (N_21487,N_19542,N_19856);
and U21488 (N_21488,N_17656,N_18008);
or U21489 (N_21489,N_17621,N_19774);
nor U21490 (N_21490,N_19930,N_18619);
xnor U21491 (N_21491,N_19344,N_18941);
and U21492 (N_21492,N_18128,N_19222);
and U21493 (N_21493,N_19841,N_17721);
and U21494 (N_21494,N_19085,N_19190);
xor U21495 (N_21495,N_19183,N_18328);
or U21496 (N_21496,N_18659,N_17794);
nand U21497 (N_21497,N_18124,N_17646);
xor U21498 (N_21498,N_17670,N_18330);
xor U21499 (N_21499,N_18351,N_19299);
nand U21500 (N_21500,N_19443,N_17748);
xnor U21501 (N_21501,N_19908,N_19077);
nand U21502 (N_21502,N_19995,N_18966);
xnor U21503 (N_21503,N_19687,N_18960);
xnor U21504 (N_21504,N_19646,N_18876);
and U21505 (N_21505,N_18194,N_19245);
and U21506 (N_21506,N_19235,N_18349);
xnor U21507 (N_21507,N_18842,N_19070);
nor U21508 (N_21508,N_18593,N_17938);
nor U21509 (N_21509,N_18882,N_19086);
or U21510 (N_21510,N_18316,N_18994);
nand U21511 (N_21511,N_19969,N_18969);
or U21512 (N_21512,N_18221,N_18683);
nor U21513 (N_21513,N_17952,N_18216);
xnor U21514 (N_21514,N_17860,N_19535);
xnor U21515 (N_21515,N_19570,N_19802);
nor U21516 (N_21516,N_17681,N_19894);
nand U21517 (N_21517,N_18853,N_19688);
or U21518 (N_21518,N_17603,N_18203);
nor U21519 (N_21519,N_18326,N_19940);
xor U21520 (N_21520,N_18043,N_18542);
or U21521 (N_21521,N_19202,N_19336);
xor U21522 (N_21522,N_18287,N_18011);
or U21523 (N_21523,N_18926,N_19245);
or U21524 (N_21524,N_19238,N_19854);
and U21525 (N_21525,N_19461,N_17767);
nand U21526 (N_21526,N_19518,N_19550);
xor U21527 (N_21527,N_19139,N_18231);
and U21528 (N_21528,N_18981,N_19140);
and U21529 (N_21529,N_17581,N_18389);
nor U21530 (N_21530,N_18519,N_18050);
or U21531 (N_21531,N_19832,N_19009);
xor U21532 (N_21532,N_18318,N_18804);
nand U21533 (N_21533,N_19061,N_19188);
and U21534 (N_21534,N_17862,N_17538);
xnor U21535 (N_21535,N_19120,N_17995);
xor U21536 (N_21536,N_17885,N_19285);
nor U21537 (N_21537,N_19953,N_18482);
nand U21538 (N_21538,N_19193,N_19189);
xor U21539 (N_21539,N_19239,N_19757);
and U21540 (N_21540,N_17626,N_19279);
or U21541 (N_21541,N_18601,N_18637);
and U21542 (N_21542,N_18245,N_19716);
nand U21543 (N_21543,N_19838,N_19568);
xnor U21544 (N_21544,N_18008,N_19222);
nor U21545 (N_21545,N_18596,N_17514);
or U21546 (N_21546,N_18733,N_18768);
nor U21547 (N_21547,N_19330,N_19288);
xor U21548 (N_21548,N_18379,N_19064);
or U21549 (N_21549,N_18616,N_19043);
or U21550 (N_21550,N_19026,N_18129);
or U21551 (N_21551,N_19580,N_17704);
nor U21552 (N_21552,N_19415,N_18445);
nand U21553 (N_21553,N_18207,N_19315);
xnor U21554 (N_21554,N_18834,N_19599);
or U21555 (N_21555,N_17565,N_18942);
nor U21556 (N_21556,N_18258,N_18755);
xnor U21557 (N_21557,N_18509,N_19337);
nor U21558 (N_21558,N_17555,N_18391);
or U21559 (N_21559,N_17558,N_18735);
or U21560 (N_21560,N_19853,N_17594);
or U21561 (N_21561,N_18327,N_18893);
nor U21562 (N_21562,N_18157,N_18537);
nand U21563 (N_21563,N_19745,N_18079);
and U21564 (N_21564,N_18441,N_19362);
xor U21565 (N_21565,N_18281,N_17965);
and U21566 (N_21566,N_19090,N_18486);
xor U21567 (N_21567,N_19947,N_18862);
and U21568 (N_21568,N_18040,N_19097);
xor U21569 (N_21569,N_17867,N_19246);
or U21570 (N_21570,N_18532,N_18645);
nor U21571 (N_21571,N_18820,N_17645);
nor U21572 (N_21572,N_18803,N_18626);
or U21573 (N_21573,N_18425,N_18350);
and U21574 (N_21574,N_19693,N_17730);
nand U21575 (N_21575,N_19560,N_19876);
or U21576 (N_21576,N_18440,N_19341);
xor U21577 (N_21577,N_19068,N_19505);
nand U21578 (N_21578,N_19253,N_19082);
xnor U21579 (N_21579,N_17509,N_17642);
or U21580 (N_21580,N_18540,N_17842);
and U21581 (N_21581,N_18163,N_18112);
nor U21582 (N_21582,N_17780,N_19655);
xor U21583 (N_21583,N_19299,N_18043);
nand U21584 (N_21584,N_18667,N_18473);
nor U21585 (N_21585,N_17620,N_19558);
or U21586 (N_21586,N_19126,N_17688);
nand U21587 (N_21587,N_18473,N_19775);
nand U21588 (N_21588,N_18897,N_18981);
nand U21589 (N_21589,N_18739,N_18239);
xor U21590 (N_21590,N_19413,N_18515);
xor U21591 (N_21591,N_18158,N_17602);
and U21592 (N_21592,N_19098,N_18802);
and U21593 (N_21593,N_18269,N_19534);
nand U21594 (N_21594,N_19658,N_18176);
nor U21595 (N_21595,N_19596,N_19185);
or U21596 (N_21596,N_17898,N_18879);
nor U21597 (N_21597,N_19324,N_19577);
nor U21598 (N_21598,N_18806,N_19358);
nand U21599 (N_21599,N_18389,N_18783);
xor U21600 (N_21600,N_19582,N_18858);
xor U21601 (N_21601,N_19583,N_19212);
and U21602 (N_21602,N_18679,N_19862);
or U21603 (N_21603,N_18011,N_19187);
nor U21604 (N_21604,N_19286,N_18802);
nand U21605 (N_21605,N_18946,N_18471);
nand U21606 (N_21606,N_18751,N_18603);
nand U21607 (N_21607,N_19445,N_18280);
or U21608 (N_21608,N_18841,N_18075);
and U21609 (N_21609,N_19296,N_19889);
or U21610 (N_21610,N_19341,N_19636);
nor U21611 (N_21611,N_17766,N_19823);
nor U21612 (N_21612,N_17879,N_18148);
xor U21613 (N_21613,N_19959,N_19333);
xor U21614 (N_21614,N_19020,N_18099);
and U21615 (N_21615,N_18224,N_18127);
nor U21616 (N_21616,N_18927,N_17705);
or U21617 (N_21617,N_19855,N_18630);
nand U21618 (N_21618,N_19781,N_18246);
or U21619 (N_21619,N_18599,N_18156);
nand U21620 (N_21620,N_17679,N_19279);
nor U21621 (N_21621,N_19610,N_19342);
xor U21622 (N_21622,N_17883,N_17940);
nand U21623 (N_21623,N_18660,N_18548);
and U21624 (N_21624,N_19723,N_18242);
or U21625 (N_21625,N_19668,N_19744);
or U21626 (N_21626,N_18222,N_18258);
nand U21627 (N_21627,N_19658,N_18403);
nand U21628 (N_21628,N_19657,N_19629);
and U21629 (N_21629,N_18051,N_17739);
xor U21630 (N_21630,N_19778,N_18118);
xnor U21631 (N_21631,N_18840,N_18115);
xnor U21632 (N_21632,N_19755,N_19454);
nand U21633 (N_21633,N_18523,N_19478);
nand U21634 (N_21634,N_17742,N_18630);
nor U21635 (N_21635,N_18326,N_18199);
nand U21636 (N_21636,N_19655,N_18414);
nand U21637 (N_21637,N_19238,N_19195);
or U21638 (N_21638,N_18887,N_17509);
xor U21639 (N_21639,N_18228,N_18811);
or U21640 (N_21640,N_17563,N_17965);
nor U21641 (N_21641,N_17539,N_18881);
nor U21642 (N_21642,N_18100,N_19033);
xnor U21643 (N_21643,N_19937,N_19514);
nand U21644 (N_21644,N_19660,N_18169);
nand U21645 (N_21645,N_18245,N_19076);
and U21646 (N_21646,N_17608,N_17635);
xor U21647 (N_21647,N_18404,N_19773);
and U21648 (N_21648,N_19018,N_17970);
xor U21649 (N_21649,N_18967,N_17714);
nor U21650 (N_21650,N_19579,N_18928);
xnor U21651 (N_21651,N_18407,N_17940);
and U21652 (N_21652,N_18333,N_18105);
or U21653 (N_21653,N_18443,N_19931);
xor U21654 (N_21654,N_18348,N_17727);
xor U21655 (N_21655,N_18086,N_18190);
nor U21656 (N_21656,N_18742,N_19508);
nor U21657 (N_21657,N_19253,N_18575);
and U21658 (N_21658,N_18640,N_19460);
nand U21659 (N_21659,N_18475,N_19237);
xnor U21660 (N_21660,N_17596,N_18529);
or U21661 (N_21661,N_19594,N_17731);
or U21662 (N_21662,N_17759,N_17665);
nor U21663 (N_21663,N_17960,N_18485);
xor U21664 (N_21664,N_19284,N_18852);
nor U21665 (N_21665,N_18575,N_19897);
and U21666 (N_21666,N_17702,N_17557);
or U21667 (N_21667,N_19670,N_17533);
nand U21668 (N_21668,N_18104,N_19705);
or U21669 (N_21669,N_18821,N_19072);
nor U21670 (N_21670,N_17891,N_18419);
xor U21671 (N_21671,N_19576,N_17648);
and U21672 (N_21672,N_19345,N_18158);
and U21673 (N_21673,N_18186,N_17930);
xor U21674 (N_21674,N_19078,N_19720);
nand U21675 (N_21675,N_18527,N_19795);
nor U21676 (N_21676,N_19631,N_17772);
or U21677 (N_21677,N_18720,N_18727);
nand U21678 (N_21678,N_18227,N_19492);
nor U21679 (N_21679,N_17966,N_18915);
nand U21680 (N_21680,N_18762,N_18417);
or U21681 (N_21681,N_18397,N_19090);
or U21682 (N_21682,N_19772,N_19227);
nor U21683 (N_21683,N_19701,N_18399);
xnor U21684 (N_21684,N_18986,N_19259);
xnor U21685 (N_21685,N_17899,N_17916);
xor U21686 (N_21686,N_19798,N_18737);
nand U21687 (N_21687,N_19264,N_19153);
and U21688 (N_21688,N_18539,N_19398);
or U21689 (N_21689,N_19349,N_18682);
or U21690 (N_21690,N_19234,N_19090);
and U21691 (N_21691,N_19195,N_19827);
xnor U21692 (N_21692,N_18261,N_19983);
nor U21693 (N_21693,N_17877,N_17973);
or U21694 (N_21694,N_17942,N_19628);
nor U21695 (N_21695,N_19649,N_19895);
nor U21696 (N_21696,N_18725,N_18676);
nand U21697 (N_21697,N_19265,N_19640);
xnor U21698 (N_21698,N_17738,N_18183);
or U21699 (N_21699,N_18068,N_18415);
nand U21700 (N_21700,N_18870,N_17925);
nor U21701 (N_21701,N_19618,N_17507);
xor U21702 (N_21702,N_19149,N_18156);
or U21703 (N_21703,N_19715,N_19791);
nand U21704 (N_21704,N_19221,N_19078);
xnor U21705 (N_21705,N_18520,N_17599);
and U21706 (N_21706,N_17638,N_17994);
and U21707 (N_21707,N_19836,N_19853);
and U21708 (N_21708,N_19011,N_19714);
nand U21709 (N_21709,N_18346,N_19373);
xor U21710 (N_21710,N_17601,N_18202);
nor U21711 (N_21711,N_19558,N_17658);
nand U21712 (N_21712,N_18620,N_19664);
and U21713 (N_21713,N_17669,N_18099);
xnor U21714 (N_21714,N_18234,N_19709);
and U21715 (N_21715,N_18734,N_18969);
or U21716 (N_21716,N_17555,N_18913);
nor U21717 (N_21717,N_17902,N_17619);
and U21718 (N_21718,N_18746,N_17736);
nand U21719 (N_21719,N_19809,N_18545);
and U21720 (N_21720,N_19456,N_18215);
or U21721 (N_21721,N_17813,N_18213);
and U21722 (N_21722,N_19749,N_18008);
or U21723 (N_21723,N_17741,N_19339);
xnor U21724 (N_21724,N_19598,N_18989);
and U21725 (N_21725,N_17912,N_18349);
nor U21726 (N_21726,N_18757,N_19648);
xor U21727 (N_21727,N_19388,N_19566);
nor U21728 (N_21728,N_17627,N_19116);
and U21729 (N_21729,N_19626,N_18956);
xor U21730 (N_21730,N_18679,N_19818);
nor U21731 (N_21731,N_18639,N_18598);
xor U21732 (N_21732,N_18799,N_18971);
nand U21733 (N_21733,N_18950,N_18186);
xnor U21734 (N_21734,N_18212,N_17899);
nand U21735 (N_21735,N_18818,N_19633);
xor U21736 (N_21736,N_18677,N_19255);
nand U21737 (N_21737,N_19741,N_19847);
nand U21738 (N_21738,N_18327,N_18848);
or U21739 (N_21739,N_19457,N_18535);
or U21740 (N_21740,N_19296,N_17814);
and U21741 (N_21741,N_19390,N_17924);
xor U21742 (N_21742,N_18352,N_18670);
xnor U21743 (N_21743,N_18908,N_18886);
nand U21744 (N_21744,N_18769,N_19159);
nand U21745 (N_21745,N_19506,N_17880);
nand U21746 (N_21746,N_18033,N_19000);
or U21747 (N_21747,N_18930,N_18601);
nand U21748 (N_21748,N_18120,N_17636);
nor U21749 (N_21749,N_19364,N_18455);
nand U21750 (N_21750,N_19774,N_18901);
and U21751 (N_21751,N_19660,N_19736);
nor U21752 (N_21752,N_18126,N_18585);
nand U21753 (N_21753,N_19023,N_18952);
nor U21754 (N_21754,N_17845,N_18980);
nand U21755 (N_21755,N_18906,N_19490);
xnor U21756 (N_21756,N_19815,N_17925);
or U21757 (N_21757,N_18298,N_17894);
or U21758 (N_21758,N_17805,N_17689);
xor U21759 (N_21759,N_19770,N_19188);
nand U21760 (N_21760,N_18105,N_19392);
and U21761 (N_21761,N_19572,N_17505);
nand U21762 (N_21762,N_17782,N_18540);
or U21763 (N_21763,N_18804,N_19791);
xnor U21764 (N_21764,N_19434,N_19205);
and U21765 (N_21765,N_19905,N_17536);
xor U21766 (N_21766,N_18591,N_19489);
xor U21767 (N_21767,N_17917,N_18201);
nor U21768 (N_21768,N_19737,N_19743);
nor U21769 (N_21769,N_19182,N_17671);
xor U21770 (N_21770,N_19407,N_19587);
nor U21771 (N_21771,N_17773,N_18053);
and U21772 (N_21772,N_18704,N_19057);
and U21773 (N_21773,N_18471,N_18846);
nand U21774 (N_21774,N_18880,N_18010);
nand U21775 (N_21775,N_18490,N_18874);
or U21776 (N_21776,N_18748,N_18143);
or U21777 (N_21777,N_19515,N_18080);
and U21778 (N_21778,N_19340,N_19647);
and U21779 (N_21779,N_19059,N_18298);
or U21780 (N_21780,N_18343,N_17968);
and U21781 (N_21781,N_18836,N_19224);
or U21782 (N_21782,N_17695,N_19949);
nor U21783 (N_21783,N_18743,N_18489);
nand U21784 (N_21784,N_19217,N_17977);
nand U21785 (N_21785,N_19420,N_18724);
nand U21786 (N_21786,N_18615,N_19964);
or U21787 (N_21787,N_19707,N_17804);
or U21788 (N_21788,N_17966,N_18251);
or U21789 (N_21789,N_19903,N_19004);
xnor U21790 (N_21790,N_18276,N_18868);
nand U21791 (N_21791,N_17741,N_17580);
nand U21792 (N_21792,N_19166,N_17689);
xor U21793 (N_21793,N_17961,N_17579);
nand U21794 (N_21794,N_18174,N_19146);
and U21795 (N_21795,N_18983,N_18692);
nand U21796 (N_21796,N_19169,N_18225);
xor U21797 (N_21797,N_18045,N_19527);
xor U21798 (N_21798,N_18320,N_18017);
and U21799 (N_21799,N_18254,N_18033);
and U21800 (N_21800,N_19947,N_19234);
nand U21801 (N_21801,N_18602,N_19847);
nor U21802 (N_21802,N_19003,N_17629);
nor U21803 (N_21803,N_19942,N_17889);
xor U21804 (N_21804,N_19177,N_18430);
and U21805 (N_21805,N_19504,N_17613);
xor U21806 (N_21806,N_18536,N_19516);
xor U21807 (N_21807,N_18324,N_17982);
or U21808 (N_21808,N_17789,N_17532);
nand U21809 (N_21809,N_17635,N_19053);
nor U21810 (N_21810,N_19433,N_19504);
nor U21811 (N_21811,N_19337,N_19124);
xnor U21812 (N_21812,N_19511,N_18723);
or U21813 (N_21813,N_19757,N_17818);
nand U21814 (N_21814,N_19555,N_17753);
xnor U21815 (N_21815,N_17727,N_19260);
nand U21816 (N_21816,N_17844,N_18333);
xor U21817 (N_21817,N_18123,N_19439);
xnor U21818 (N_21818,N_18935,N_18495);
xnor U21819 (N_21819,N_19999,N_18857);
and U21820 (N_21820,N_19942,N_18528);
and U21821 (N_21821,N_17586,N_19747);
nor U21822 (N_21822,N_19565,N_18377);
xor U21823 (N_21823,N_18919,N_18353);
and U21824 (N_21824,N_18252,N_17681);
nand U21825 (N_21825,N_18657,N_17886);
nand U21826 (N_21826,N_18572,N_17857);
nor U21827 (N_21827,N_17966,N_18893);
nand U21828 (N_21828,N_18031,N_17840);
and U21829 (N_21829,N_19227,N_19074);
or U21830 (N_21830,N_18589,N_19749);
or U21831 (N_21831,N_19317,N_19844);
nor U21832 (N_21832,N_18400,N_18827);
and U21833 (N_21833,N_18881,N_18096);
xor U21834 (N_21834,N_17865,N_17750);
nor U21835 (N_21835,N_19253,N_18059);
xnor U21836 (N_21836,N_17923,N_19250);
xnor U21837 (N_21837,N_17858,N_18952);
and U21838 (N_21838,N_19428,N_18392);
and U21839 (N_21839,N_18860,N_18246);
or U21840 (N_21840,N_19561,N_19150);
nand U21841 (N_21841,N_18658,N_17867);
and U21842 (N_21842,N_18142,N_17526);
or U21843 (N_21843,N_19706,N_18409);
nand U21844 (N_21844,N_17870,N_18949);
or U21845 (N_21845,N_17598,N_17587);
nor U21846 (N_21846,N_18545,N_17968);
nand U21847 (N_21847,N_17508,N_18422);
nand U21848 (N_21848,N_19500,N_19119);
xor U21849 (N_21849,N_18935,N_19106);
nor U21850 (N_21850,N_18534,N_18652);
and U21851 (N_21851,N_18219,N_18050);
nor U21852 (N_21852,N_19392,N_19661);
nand U21853 (N_21853,N_19691,N_19982);
xnor U21854 (N_21854,N_18539,N_18919);
nand U21855 (N_21855,N_18089,N_19361);
or U21856 (N_21856,N_17583,N_18575);
xor U21857 (N_21857,N_19489,N_17861);
nand U21858 (N_21858,N_19313,N_18009);
xnor U21859 (N_21859,N_19828,N_18111);
xnor U21860 (N_21860,N_18547,N_19014);
nand U21861 (N_21861,N_19745,N_18712);
xnor U21862 (N_21862,N_19633,N_19510);
and U21863 (N_21863,N_18660,N_19642);
and U21864 (N_21864,N_18304,N_17782);
nand U21865 (N_21865,N_19057,N_18724);
or U21866 (N_21866,N_19681,N_18154);
xnor U21867 (N_21867,N_19594,N_19172);
nand U21868 (N_21868,N_18318,N_17936);
or U21869 (N_21869,N_19130,N_18404);
or U21870 (N_21870,N_19309,N_18775);
nand U21871 (N_21871,N_18177,N_18578);
nand U21872 (N_21872,N_19632,N_19865);
nor U21873 (N_21873,N_19271,N_19781);
nor U21874 (N_21874,N_19888,N_19234);
and U21875 (N_21875,N_19820,N_17754);
and U21876 (N_21876,N_19684,N_19506);
nand U21877 (N_21877,N_19190,N_18819);
or U21878 (N_21878,N_17700,N_18694);
xnor U21879 (N_21879,N_18329,N_17896);
or U21880 (N_21880,N_18350,N_18621);
and U21881 (N_21881,N_18111,N_19420);
nand U21882 (N_21882,N_19309,N_19615);
and U21883 (N_21883,N_19793,N_17849);
and U21884 (N_21884,N_17622,N_19602);
nor U21885 (N_21885,N_18780,N_18945);
nand U21886 (N_21886,N_19046,N_17674);
nor U21887 (N_21887,N_18555,N_18187);
and U21888 (N_21888,N_17697,N_18728);
nand U21889 (N_21889,N_17537,N_18788);
or U21890 (N_21890,N_18509,N_18988);
nor U21891 (N_21891,N_19221,N_19084);
nand U21892 (N_21892,N_19658,N_19153);
nand U21893 (N_21893,N_18235,N_17556);
nor U21894 (N_21894,N_19314,N_19143);
or U21895 (N_21895,N_17884,N_19450);
xnor U21896 (N_21896,N_18277,N_18141);
xor U21897 (N_21897,N_19185,N_17551);
nand U21898 (N_21898,N_18857,N_19731);
nand U21899 (N_21899,N_17929,N_19958);
and U21900 (N_21900,N_19788,N_19787);
nor U21901 (N_21901,N_19771,N_19431);
nor U21902 (N_21902,N_19161,N_19331);
nand U21903 (N_21903,N_19215,N_19235);
xor U21904 (N_21904,N_18320,N_19675);
nor U21905 (N_21905,N_17675,N_18929);
xor U21906 (N_21906,N_17566,N_17850);
nor U21907 (N_21907,N_19130,N_18322);
nor U21908 (N_21908,N_18471,N_19790);
nand U21909 (N_21909,N_17597,N_17500);
nor U21910 (N_21910,N_19982,N_19699);
or U21911 (N_21911,N_18385,N_19920);
xor U21912 (N_21912,N_19466,N_19358);
or U21913 (N_21913,N_18384,N_19795);
xnor U21914 (N_21914,N_18669,N_19707);
and U21915 (N_21915,N_19675,N_19264);
nand U21916 (N_21916,N_18267,N_18008);
nor U21917 (N_21917,N_18328,N_18326);
nor U21918 (N_21918,N_19168,N_17714);
or U21919 (N_21919,N_18406,N_17873);
nand U21920 (N_21920,N_18552,N_19907);
nand U21921 (N_21921,N_19449,N_18101);
or U21922 (N_21922,N_17595,N_18871);
nor U21923 (N_21923,N_19686,N_19320);
or U21924 (N_21924,N_18848,N_18495);
xor U21925 (N_21925,N_18107,N_18954);
and U21926 (N_21926,N_17601,N_18435);
nand U21927 (N_21927,N_19295,N_18601);
or U21928 (N_21928,N_18165,N_19939);
or U21929 (N_21929,N_19561,N_17856);
nand U21930 (N_21930,N_18763,N_18434);
nor U21931 (N_21931,N_17953,N_17635);
nand U21932 (N_21932,N_17694,N_18488);
or U21933 (N_21933,N_19953,N_17979);
and U21934 (N_21934,N_19434,N_19646);
nand U21935 (N_21935,N_18379,N_18277);
nor U21936 (N_21936,N_19735,N_18974);
nand U21937 (N_21937,N_18140,N_17991);
nor U21938 (N_21938,N_17808,N_18954);
or U21939 (N_21939,N_18305,N_19898);
nor U21940 (N_21940,N_19417,N_18147);
or U21941 (N_21941,N_18211,N_19576);
and U21942 (N_21942,N_19885,N_18456);
or U21943 (N_21943,N_17831,N_18534);
and U21944 (N_21944,N_18939,N_19924);
or U21945 (N_21945,N_17672,N_19223);
nand U21946 (N_21946,N_19403,N_19115);
nor U21947 (N_21947,N_19537,N_18547);
and U21948 (N_21948,N_19716,N_19660);
and U21949 (N_21949,N_17925,N_18677);
nor U21950 (N_21950,N_18953,N_19810);
nand U21951 (N_21951,N_17541,N_18519);
nor U21952 (N_21952,N_19111,N_19170);
nor U21953 (N_21953,N_18778,N_17552);
or U21954 (N_21954,N_17614,N_19768);
and U21955 (N_21955,N_19442,N_19733);
nor U21956 (N_21956,N_19450,N_17670);
and U21957 (N_21957,N_17920,N_19406);
nand U21958 (N_21958,N_19618,N_19992);
nand U21959 (N_21959,N_19182,N_18742);
nor U21960 (N_21960,N_19084,N_18771);
xnor U21961 (N_21961,N_18451,N_18843);
nor U21962 (N_21962,N_17621,N_19626);
nand U21963 (N_21963,N_17806,N_18200);
xor U21964 (N_21964,N_19761,N_17868);
nor U21965 (N_21965,N_17966,N_18444);
nor U21966 (N_21966,N_18475,N_17963);
nand U21967 (N_21967,N_18500,N_19038);
xor U21968 (N_21968,N_18127,N_18391);
nor U21969 (N_21969,N_19751,N_18404);
xnor U21970 (N_21970,N_17688,N_18038);
nand U21971 (N_21971,N_19582,N_19620);
nor U21972 (N_21972,N_17888,N_17708);
and U21973 (N_21973,N_19027,N_18178);
or U21974 (N_21974,N_18504,N_18680);
nand U21975 (N_21975,N_19600,N_17504);
nor U21976 (N_21976,N_18356,N_19857);
nor U21977 (N_21977,N_18173,N_19797);
nor U21978 (N_21978,N_17628,N_18063);
or U21979 (N_21979,N_18027,N_17936);
nand U21980 (N_21980,N_18855,N_19968);
xor U21981 (N_21981,N_19933,N_18749);
nand U21982 (N_21982,N_19621,N_17861);
and U21983 (N_21983,N_18629,N_18420);
nand U21984 (N_21984,N_17759,N_19589);
nor U21985 (N_21985,N_19155,N_18207);
xor U21986 (N_21986,N_19850,N_17787);
xor U21987 (N_21987,N_19652,N_17528);
or U21988 (N_21988,N_18034,N_17736);
and U21989 (N_21989,N_19549,N_18803);
or U21990 (N_21990,N_18135,N_18633);
xor U21991 (N_21991,N_18209,N_18132);
or U21992 (N_21992,N_17898,N_18357);
nand U21993 (N_21993,N_17794,N_19222);
nor U21994 (N_21994,N_19048,N_17913);
nand U21995 (N_21995,N_18596,N_18974);
nand U21996 (N_21996,N_18252,N_18225);
or U21997 (N_21997,N_17956,N_18496);
or U21998 (N_21998,N_17583,N_17835);
or U21999 (N_21999,N_18889,N_18968);
and U22000 (N_22000,N_18124,N_19733);
nand U22001 (N_22001,N_19361,N_17657);
nand U22002 (N_22002,N_18823,N_19842);
nand U22003 (N_22003,N_18421,N_19035);
nand U22004 (N_22004,N_18098,N_19004);
nor U22005 (N_22005,N_19001,N_19562);
and U22006 (N_22006,N_19740,N_18523);
nor U22007 (N_22007,N_18218,N_19273);
xnor U22008 (N_22008,N_19724,N_19003);
or U22009 (N_22009,N_19974,N_18135);
or U22010 (N_22010,N_18071,N_19181);
nand U22011 (N_22011,N_19331,N_18439);
nor U22012 (N_22012,N_19175,N_17886);
nor U22013 (N_22013,N_17839,N_18146);
and U22014 (N_22014,N_17801,N_19651);
xnor U22015 (N_22015,N_17979,N_19857);
nor U22016 (N_22016,N_19605,N_19739);
nor U22017 (N_22017,N_17555,N_19647);
or U22018 (N_22018,N_18408,N_17698);
nor U22019 (N_22019,N_19149,N_18761);
nand U22020 (N_22020,N_18803,N_18984);
and U22021 (N_22021,N_18901,N_18065);
and U22022 (N_22022,N_19799,N_17973);
or U22023 (N_22023,N_18445,N_19506);
nand U22024 (N_22024,N_19020,N_18849);
nand U22025 (N_22025,N_19174,N_18849);
xnor U22026 (N_22026,N_18530,N_18773);
or U22027 (N_22027,N_18700,N_17950);
and U22028 (N_22028,N_18247,N_18411);
nor U22029 (N_22029,N_18775,N_18659);
and U22030 (N_22030,N_19208,N_18109);
nor U22031 (N_22031,N_18117,N_19192);
or U22032 (N_22032,N_18858,N_17867);
and U22033 (N_22033,N_18687,N_18116);
xnor U22034 (N_22034,N_19840,N_17571);
nand U22035 (N_22035,N_17506,N_19949);
nand U22036 (N_22036,N_19717,N_18135);
xnor U22037 (N_22037,N_18685,N_18506);
or U22038 (N_22038,N_18921,N_18463);
or U22039 (N_22039,N_17897,N_17961);
or U22040 (N_22040,N_19178,N_18746);
nand U22041 (N_22041,N_18976,N_18578);
xnor U22042 (N_22042,N_19401,N_18453);
xor U22043 (N_22043,N_17668,N_19101);
and U22044 (N_22044,N_17949,N_19447);
nor U22045 (N_22045,N_18550,N_17927);
xor U22046 (N_22046,N_18949,N_19416);
xor U22047 (N_22047,N_19877,N_17907);
nand U22048 (N_22048,N_19389,N_19948);
and U22049 (N_22049,N_18151,N_19509);
nand U22050 (N_22050,N_19424,N_18228);
and U22051 (N_22051,N_19387,N_18938);
or U22052 (N_22052,N_18138,N_19254);
nand U22053 (N_22053,N_18175,N_17905);
or U22054 (N_22054,N_19661,N_18125);
nor U22055 (N_22055,N_18125,N_17842);
nand U22056 (N_22056,N_19200,N_19795);
nand U22057 (N_22057,N_17595,N_18803);
or U22058 (N_22058,N_19091,N_17568);
or U22059 (N_22059,N_18278,N_18896);
and U22060 (N_22060,N_18123,N_19286);
nor U22061 (N_22061,N_17698,N_18906);
or U22062 (N_22062,N_19244,N_19661);
or U22063 (N_22063,N_19922,N_18621);
nand U22064 (N_22064,N_17818,N_19016);
and U22065 (N_22065,N_17511,N_18124);
and U22066 (N_22066,N_19564,N_19098);
nor U22067 (N_22067,N_18552,N_19704);
or U22068 (N_22068,N_19882,N_19327);
nand U22069 (N_22069,N_17661,N_19984);
xnor U22070 (N_22070,N_19181,N_17545);
nand U22071 (N_22071,N_17545,N_17974);
and U22072 (N_22072,N_19668,N_19161);
and U22073 (N_22073,N_18411,N_18503);
nor U22074 (N_22074,N_18355,N_18463);
nor U22075 (N_22075,N_18581,N_17513);
nor U22076 (N_22076,N_19382,N_18445);
nor U22077 (N_22077,N_19286,N_18923);
or U22078 (N_22078,N_18740,N_18091);
xor U22079 (N_22079,N_19493,N_18241);
nor U22080 (N_22080,N_17889,N_18395);
and U22081 (N_22081,N_18364,N_19326);
or U22082 (N_22082,N_19553,N_18185);
and U22083 (N_22083,N_19662,N_18728);
nor U22084 (N_22084,N_18709,N_17923);
or U22085 (N_22085,N_19992,N_18462);
xnor U22086 (N_22086,N_18830,N_17796);
or U22087 (N_22087,N_19891,N_18390);
and U22088 (N_22088,N_17817,N_18055);
nand U22089 (N_22089,N_19432,N_18030);
or U22090 (N_22090,N_18937,N_19386);
nand U22091 (N_22091,N_18673,N_19397);
or U22092 (N_22092,N_19219,N_18186);
and U22093 (N_22093,N_18331,N_18233);
nand U22094 (N_22094,N_18167,N_19460);
nand U22095 (N_22095,N_19117,N_18235);
xnor U22096 (N_22096,N_19732,N_19444);
and U22097 (N_22097,N_18558,N_19936);
nand U22098 (N_22098,N_18572,N_18001);
nand U22099 (N_22099,N_19233,N_17709);
nand U22100 (N_22100,N_19070,N_18437);
xnor U22101 (N_22101,N_19654,N_18073);
nor U22102 (N_22102,N_19709,N_18238);
and U22103 (N_22103,N_19349,N_18629);
nor U22104 (N_22104,N_18957,N_17590);
nand U22105 (N_22105,N_19677,N_17757);
and U22106 (N_22106,N_19555,N_19877);
or U22107 (N_22107,N_19939,N_19154);
or U22108 (N_22108,N_19376,N_18612);
xor U22109 (N_22109,N_19172,N_17559);
nand U22110 (N_22110,N_18753,N_18074);
and U22111 (N_22111,N_18962,N_18324);
or U22112 (N_22112,N_19684,N_18780);
nand U22113 (N_22113,N_18863,N_18338);
nand U22114 (N_22114,N_18462,N_19665);
xnor U22115 (N_22115,N_19064,N_19113);
nand U22116 (N_22116,N_18262,N_19710);
and U22117 (N_22117,N_19653,N_17510);
xor U22118 (N_22118,N_19964,N_18631);
and U22119 (N_22119,N_18114,N_18605);
and U22120 (N_22120,N_19487,N_17892);
xnor U22121 (N_22121,N_17895,N_18028);
and U22122 (N_22122,N_19432,N_18067);
or U22123 (N_22123,N_19731,N_18502);
nor U22124 (N_22124,N_18507,N_19708);
nor U22125 (N_22125,N_19044,N_19090);
and U22126 (N_22126,N_18201,N_19122);
nand U22127 (N_22127,N_18232,N_19289);
nand U22128 (N_22128,N_19998,N_19253);
xnor U22129 (N_22129,N_18744,N_19291);
and U22130 (N_22130,N_17893,N_18191);
nor U22131 (N_22131,N_17620,N_19134);
xnor U22132 (N_22132,N_17639,N_19335);
xor U22133 (N_22133,N_19844,N_19882);
nand U22134 (N_22134,N_19523,N_19254);
nor U22135 (N_22135,N_19590,N_17720);
nand U22136 (N_22136,N_18489,N_18906);
and U22137 (N_22137,N_19368,N_18248);
xnor U22138 (N_22138,N_19390,N_17988);
nor U22139 (N_22139,N_19453,N_19517);
or U22140 (N_22140,N_18925,N_17764);
nor U22141 (N_22141,N_17672,N_18023);
and U22142 (N_22142,N_19289,N_18648);
nor U22143 (N_22143,N_18336,N_19368);
nor U22144 (N_22144,N_18542,N_18235);
nand U22145 (N_22145,N_18086,N_19274);
and U22146 (N_22146,N_19705,N_18889);
xor U22147 (N_22147,N_19659,N_19102);
nand U22148 (N_22148,N_19195,N_18285);
and U22149 (N_22149,N_17770,N_18977);
or U22150 (N_22150,N_18310,N_18514);
or U22151 (N_22151,N_19079,N_17993);
xor U22152 (N_22152,N_19590,N_18488);
nand U22153 (N_22153,N_17878,N_18001);
and U22154 (N_22154,N_17631,N_19339);
xor U22155 (N_22155,N_18009,N_18080);
or U22156 (N_22156,N_18021,N_19270);
nand U22157 (N_22157,N_18368,N_19294);
nand U22158 (N_22158,N_19854,N_18703);
or U22159 (N_22159,N_17890,N_19314);
and U22160 (N_22160,N_18645,N_18290);
or U22161 (N_22161,N_18906,N_19755);
nor U22162 (N_22162,N_18255,N_17569);
xor U22163 (N_22163,N_18164,N_19500);
and U22164 (N_22164,N_19074,N_19327);
or U22165 (N_22165,N_17657,N_17637);
or U22166 (N_22166,N_19903,N_19728);
and U22167 (N_22167,N_18399,N_19676);
xor U22168 (N_22168,N_19289,N_19031);
xor U22169 (N_22169,N_19248,N_18806);
nand U22170 (N_22170,N_17654,N_19257);
xnor U22171 (N_22171,N_18720,N_17655);
xor U22172 (N_22172,N_19885,N_17615);
xnor U22173 (N_22173,N_17504,N_18048);
or U22174 (N_22174,N_18610,N_19726);
nand U22175 (N_22175,N_18085,N_19354);
xnor U22176 (N_22176,N_17926,N_19612);
and U22177 (N_22177,N_19323,N_19314);
or U22178 (N_22178,N_18395,N_18886);
xnor U22179 (N_22179,N_19013,N_19408);
or U22180 (N_22180,N_18182,N_19013);
nor U22181 (N_22181,N_19704,N_19711);
or U22182 (N_22182,N_19052,N_18024);
or U22183 (N_22183,N_18427,N_19155);
or U22184 (N_22184,N_19850,N_18219);
nand U22185 (N_22185,N_17990,N_19233);
or U22186 (N_22186,N_19539,N_18738);
xor U22187 (N_22187,N_17992,N_19038);
nand U22188 (N_22188,N_17524,N_19528);
and U22189 (N_22189,N_19867,N_19936);
nor U22190 (N_22190,N_19708,N_17754);
nand U22191 (N_22191,N_19510,N_18104);
nor U22192 (N_22192,N_18857,N_18818);
nor U22193 (N_22193,N_19931,N_17844);
nor U22194 (N_22194,N_18731,N_19815);
and U22195 (N_22195,N_19413,N_19150);
xor U22196 (N_22196,N_17729,N_18697);
or U22197 (N_22197,N_18656,N_19482);
or U22198 (N_22198,N_17712,N_19632);
nand U22199 (N_22199,N_18445,N_18101);
nor U22200 (N_22200,N_19220,N_17715);
or U22201 (N_22201,N_18933,N_19770);
xnor U22202 (N_22202,N_19027,N_17851);
nand U22203 (N_22203,N_19361,N_19153);
and U22204 (N_22204,N_19672,N_18308);
nand U22205 (N_22205,N_19530,N_17621);
nor U22206 (N_22206,N_18663,N_18066);
nor U22207 (N_22207,N_19942,N_19017);
or U22208 (N_22208,N_19844,N_18978);
and U22209 (N_22209,N_18193,N_19860);
and U22210 (N_22210,N_17859,N_18148);
nand U22211 (N_22211,N_19239,N_19332);
or U22212 (N_22212,N_18637,N_18926);
or U22213 (N_22213,N_18388,N_19965);
xnor U22214 (N_22214,N_19208,N_18537);
xor U22215 (N_22215,N_17990,N_18622);
nor U22216 (N_22216,N_19518,N_19938);
xor U22217 (N_22217,N_18372,N_19415);
xnor U22218 (N_22218,N_18367,N_18314);
and U22219 (N_22219,N_19824,N_17607);
and U22220 (N_22220,N_19871,N_19165);
and U22221 (N_22221,N_18192,N_18348);
nor U22222 (N_22222,N_17798,N_19054);
or U22223 (N_22223,N_18462,N_19966);
nand U22224 (N_22224,N_19445,N_17861);
and U22225 (N_22225,N_19856,N_18352);
and U22226 (N_22226,N_18971,N_18325);
or U22227 (N_22227,N_18982,N_19439);
xnor U22228 (N_22228,N_17675,N_18549);
xor U22229 (N_22229,N_18227,N_19125);
and U22230 (N_22230,N_19803,N_19104);
or U22231 (N_22231,N_18471,N_19332);
nor U22232 (N_22232,N_18341,N_19661);
xnor U22233 (N_22233,N_17646,N_17811);
nand U22234 (N_22234,N_17655,N_17904);
nor U22235 (N_22235,N_18065,N_18152);
xnor U22236 (N_22236,N_17662,N_19241);
nand U22237 (N_22237,N_17670,N_18316);
nor U22238 (N_22238,N_19244,N_18252);
nand U22239 (N_22239,N_18651,N_19417);
xor U22240 (N_22240,N_18755,N_19089);
nand U22241 (N_22241,N_18849,N_19654);
and U22242 (N_22242,N_18646,N_18859);
nor U22243 (N_22243,N_17876,N_17735);
xor U22244 (N_22244,N_17574,N_19095);
nor U22245 (N_22245,N_18469,N_18189);
nand U22246 (N_22246,N_19418,N_17513);
nor U22247 (N_22247,N_17616,N_17545);
nor U22248 (N_22248,N_19998,N_18717);
xnor U22249 (N_22249,N_18533,N_19460);
nor U22250 (N_22250,N_17780,N_19163);
and U22251 (N_22251,N_19250,N_19102);
xor U22252 (N_22252,N_19917,N_17761);
and U22253 (N_22253,N_17918,N_19698);
and U22254 (N_22254,N_19429,N_18164);
xnor U22255 (N_22255,N_18421,N_18256);
nand U22256 (N_22256,N_17576,N_18660);
or U22257 (N_22257,N_18440,N_17641);
nor U22258 (N_22258,N_17943,N_18362);
or U22259 (N_22259,N_17780,N_18654);
or U22260 (N_22260,N_18058,N_18136);
xor U22261 (N_22261,N_18680,N_19193);
or U22262 (N_22262,N_17876,N_18738);
nor U22263 (N_22263,N_18283,N_17707);
nand U22264 (N_22264,N_19462,N_18644);
and U22265 (N_22265,N_17866,N_19111);
or U22266 (N_22266,N_18008,N_18330);
and U22267 (N_22267,N_17763,N_19231);
xor U22268 (N_22268,N_19313,N_19866);
nor U22269 (N_22269,N_19261,N_18457);
xnor U22270 (N_22270,N_18880,N_18263);
nand U22271 (N_22271,N_17970,N_18277);
nand U22272 (N_22272,N_17518,N_17678);
nand U22273 (N_22273,N_18554,N_18572);
xnor U22274 (N_22274,N_18303,N_19900);
nor U22275 (N_22275,N_19574,N_18091);
and U22276 (N_22276,N_19407,N_18754);
xnor U22277 (N_22277,N_19469,N_19785);
or U22278 (N_22278,N_18273,N_19841);
nand U22279 (N_22279,N_18910,N_18739);
xor U22280 (N_22280,N_19643,N_19855);
or U22281 (N_22281,N_19077,N_19469);
nor U22282 (N_22282,N_18731,N_18953);
and U22283 (N_22283,N_18165,N_18069);
nor U22284 (N_22284,N_18771,N_17751);
nor U22285 (N_22285,N_18316,N_19635);
and U22286 (N_22286,N_19383,N_18891);
and U22287 (N_22287,N_19787,N_18614);
and U22288 (N_22288,N_17900,N_18026);
xnor U22289 (N_22289,N_19020,N_18986);
or U22290 (N_22290,N_19669,N_19018);
and U22291 (N_22291,N_19453,N_17729);
and U22292 (N_22292,N_18472,N_17755);
or U22293 (N_22293,N_17877,N_19924);
or U22294 (N_22294,N_18768,N_18070);
nor U22295 (N_22295,N_19245,N_19968);
nor U22296 (N_22296,N_18280,N_19142);
nand U22297 (N_22297,N_17896,N_18229);
and U22298 (N_22298,N_19250,N_19473);
or U22299 (N_22299,N_18496,N_18672);
nand U22300 (N_22300,N_17715,N_19094);
or U22301 (N_22301,N_18606,N_18097);
or U22302 (N_22302,N_18444,N_19288);
and U22303 (N_22303,N_19588,N_18483);
nor U22304 (N_22304,N_19923,N_19599);
xnor U22305 (N_22305,N_17733,N_19195);
or U22306 (N_22306,N_18965,N_18861);
xnor U22307 (N_22307,N_18150,N_19327);
nor U22308 (N_22308,N_19127,N_17946);
and U22309 (N_22309,N_19269,N_17732);
xor U22310 (N_22310,N_18335,N_18173);
nor U22311 (N_22311,N_17799,N_18947);
xor U22312 (N_22312,N_18785,N_17658);
and U22313 (N_22313,N_18618,N_17875);
or U22314 (N_22314,N_19592,N_18701);
and U22315 (N_22315,N_19166,N_18264);
xor U22316 (N_22316,N_19036,N_19835);
or U22317 (N_22317,N_18106,N_19675);
or U22318 (N_22318,N_18189,N_18300);
nor U22319 (N_22319,N_17973,N_19416);
and U22320 (N_22320,N_17723,N_19222);
xor U22321 (N_22321,N_19543,N_19729);
nand U22322 (N_22322,N_18355,N_17526);
and U22323 (N_22323,N_17845,N_17519);
nand U22324 (N_22324,N_18547,N_17795);
nand U22325 (N_22325,N_18602,N_19407);
nor U22326 (N_22326,N_18436,N_19999);
or U22327 (N_22327,N_17715,N_19086);
nand U22328 (N_22328,N_19240,N_19120);
and U22329 (N_22329,N_18065,N_19362);
or U22330 (N_22330,N_17731,N_19456);
nor U22331 (N_22331,N_19068,N_19109);
nor U22332 (N_22332,N_18431,N_19102);
or U22333 (N_22333,N_19478,N_18592);
and U22334 (N_22334,N_19715,N_19903);
xor U22335 (N_22335,N_18211,N_17572);
nand U22336 (N_22336,N_19697,N_17668);
or U22337 (N_22337,N_19674,N_19279);
or U22338 (N_22338,N_19676,N_19339);
and U22339 (N_22339,N_19736,N_17624);
and U22340 (N_22340,N_19384,N_19770);
nor U22341 (N_22341,N_18292,N_18498);
nand U22342 (N_22342,N_18084,N_17886);
and U22343 (N_22343,N_18404,N_19067);
nor U22344 (N_22344,N_18933,N_17655);
nand U22345 (N_22345,N_19769,N_18896);
nand U22346 (N_22346,N_18442,N_18162);
xnor U22347 (N_22347,N_19705,N_19975);
or U22348 (N_22348,N_18265,N_18172);
or U22349 (N_22349,N_18282,N_18531);
nor U22350 (N_22350,N_18746,N_18433);
xnor U22351 (N_22351,N_19725,N_18285);
or U22352 (N_22352,N_18315,N_18536);
or U22353 (N_22353,N_19026,N_19078);
and U22354 (N_22354,N_19733,N_19685);
nand U22355 (N_22355,N_19056,N_18723);
nand U22356 (N_22356,N_17509,N_17918);
nand U22357 (N_22357,N_18738,N_17607);
or U22358 (N_22358,N_18506,N_18926);
nand U22359 (N_22359,N_17816,N_18534);
nand U22360 (N_22360,N_18886,N_18065);
nor U22361 (N_22361,N_19305,N_18334);
and U22362 (N_22362,N_18638,N_19149);
or U22363 (N_22363,N_19700,N_19955);
and U22364 (N_22364,N_19336,N_18709);
and U22365 (N_22365,N_19816,N_19043);
nand U22366 (N_22366,N_18625,N_18876);
nand U22367 (N_22367,N_17651,N_18877);
xor U22368 (N_22368,N_18366,N_19648);
xnor U22369 (N_22369,N_19636,N_17591);
xor U22370 (N_22370,N_19403,N_18929);
nor U22371 (N_22371,N_19354,N_19745);
and U22372 (N_22372,N_18279,N_17772);
and U22373 (N_22373,N_19781,N_17818);
or U22374 (N_22374,N_19693,N_18549);
nor U22375 (N_22375,N_19854,N_18386);
nand U22376 (N_22376,N_17794,N_19989);
xnor U22377 (N_22377,N_17532,N_18154);
nor U22378 (N_22378,N_18677,N_17857);
nor U22379 (N_22379,N_19818,N_17822);
nor U22380 (N_22380,N_19364,N_18737);
nand U22381 (N_22381,N_18620,N_19272);
and U22382 (N_22382,N_19264,N_18774);
nor U22383 (N_22383,N_18774,N_17926);
xor U22384 (N_22384,N_17791,N_19868);
or U22385 (N_22385,N_17790,N_19767);
xor U22386 (N_22386,N_17930,N_18320);
nand U22387 (N_22387,N_18409,N_17885);
xnor U22388 (N_22388,N_19642,N_17562);
nor U22389 (N_22389,N_19397,N_19101);
nor U22390 (N_22390,N_18898,N_19949);
xnor U22391 (N_22391,N_19927,N_18094);
nand U22392 (N_22392,N_19669,N_19399);
xnor U22393 (N_22393,N_19877,N_18969);
xnor U22394 (N_22394,N_18567,N_19181);
and U22395 (N_22395,N_18115,N_18269);
nor U22396 (N_22396,N_19943,N_19580);
and U22397 (N_22397,N_17707,N_18452);
xor U22398 (N_22398,N_18629,N_18401);
nand U22399 (N_22399,N_19149,N_17752);
xor U22400 (N_22400,N_19288,N_18083);
and U22401 (N_22401,N_19354,N_17761);
xor U22402 (N_22402,N_19458,N_18927);
nand U22403 (N_22403,N_18601,N_17625);
or U22404 (N_22404,N_19709,N_19312);
nor U22405 (N_22405,N_19656,N_19233);
and U22406 (N_22406,N_19538,N_18049);
nor U22407 (N_22407,N_17957,N_19328);
or U22408 (N_22408,N_18816,N_19206);
nor U22409 (N_22409,N_19712,N_18250);
or U22410 (N_22410,N_18881,N_17959);
nor U22411 (N_22411,N_17527,N_17929);
or U22412 (N_22412,N_18513,N_18191);
or U22413 (N_22413,N_18260,N_17669);
nor U22414 (N_22414,N_19460,N_18703);
or U22415 (N_22415,N_17664,N_19682);
nand U22416 (N_22416,N_17587,N_19652);
or U22417 (N_22417,N_19431,N_17584);
nor U22418 (N_22418,N_17852,N_18762);
xor U22419 (N_22419,N_17950,N_17616);
xnor U22420 (N_22420,N_19793,N_18448);
nor U22421 (N_22421,N_17944,N_19463);
nand U22422 (N_22422,N_19521,N_19649);
nor U22423 (N_22423,N_17546,N_17898);
nand U22424 (N_22424,N_17947,N_18804);
and U22425 (N_22425,N_17659,N_19171);
nand U22426 (N_22426,N_18226,N_19711);
nor U22427 (N_22427,N_18135,N_19778);
nor U22428 (N_22428,N_19980,N_19051);
or U22429 (N_22429,N_19053,N_18951);
nor U22430 (N_22430,N_18343,N_19814);
xor U22431 (N_22431,N_19099,N_19642);
and U22432 (N_22432,N_19538,N_17651);
xnor U22433 (N_22433,N_19597,N_18894);
or U22434 (N_22434,N_19793,N_19566);
and U22435 (N_22435,N_19293,N_18353);
and U22436 (N_22436,N_18132,N_17999);
nand U22437 (N_22437,N_18416,N_18166);
nand U22438 (N_22438,N_19014,N_19644);
and U22439 (N_22439,N_18083,N_17908);
xnor U22440 (N_22440,N_19293,N_19789);
nor U22441 (N_22441,N_19581,N_17770);
and U22442 (N_22442,N_17752,N_17941);
or U22443 (N_22443,N_18596,N_18693);
nor U22444 (N_22444,N_19314,N_19729);
xnor U22445 (N_22445,N_19683,N_17873);
nand U22446 (N_22446,N_19289,N_18999);
or U22447 (N_22447,N_19156,N_18657);
nand U22448 (N_22448,N_19239,N_17674);
xnor U22449 (N_22449,N_17512,N_19054);
nand U22450 (N_22450,N_19804,N_19463);
and U22451 (N_22451,N_18723,N_19375);
xnor U22452 (N_22452,N_18425,N_17502);
or U22453 (N_22453,N_17855,N_18867);
or U22454 (N_22454,N_17647,N_18776);
xor U22455 (N_22455,N_19919,N_17847);
or U22456 (N_22456,N_17678,N_19658);
and U22457 (N_22457,N_18118,N_18498);
nand U22458 (N_22458,N_17981,N_18014);
xor U22459 (N_22459,N_18942,N_18056);
and U22460 (N_22460,N_19729,N_17619);
and U22461 (N_22461,N_18531,N_17634);
nand U22462 (N_22462,N_19882,N_18725);
or U22463 (N_22463,N_18230,N_19448);
or U22464 (N_22464,N_17914,N_19142);
or U22465 (N_22465,N_17986,N_19022);
nand U22466 (N_22466,N_19763,N_19558);
and U22467 (N_22467,N_18689,N_18596);
nand U22468 (N_22468,N_18810,N_18011);
and U22469 (N_22469,N_18110,N_19155);
or U22470 (N_22470,N_19465,N_19440);
nand U22471 (N_22471,N_18628,N_19478);
nand U22472 (N_22472,N_19894,N_19768);
and U22473 (N_22473,N_19531,N_18107);
nand U22474 (N_22474,N_19862,N_19469);
nand U22475 (N_22475,N_19601,N_19317);
or U22476 (N_22476,N_17572,N_19694);
and U22477 (N_22477,N_19519,N_18934);
and U22478 (N_22478,N_17899,N_17596);
nand U22479 (N_22479,N_17976,N_18729);
and U22480 (N_22480,N_17544,N_19165);
and U22481 (N_22481,N_19011,N_19087);
and U22482 (N_22482,N_19165,N_19503);
and U22483 (N_22483,N_19104,N_19013);
or U22484 (N_22484,N_18327,N_19565);
or U22485 (N_22485,N_17966,N_19446);
xnor U22486 (N_22486,N_19937,N_18227);
and U22487 (N_22487,N_19999,N_19249);
and U22488 (N_22488,N_17543,N_18372);
and U22489 (N_22489,N_18416,N_19283);
nor U22490 (N_22490,N_17893,N_18330);
xor U22491 (N_22491,N_19342,N_18294);
nand U22492 (N_22492,N_19006,N_17750);
and U22493 (N_22493,N_18029,N_18662);
nand U22494 (N_22494,N_18813,N_18137);
nor U22495 (N_22495,N_17861,N_18886);
xor U22496 (N_22496,N_17815,N_19221);
or U22497 (N_22497,N_18746,N_19766);
xor U22498 (N_22498,N_17646,N_18761);
or U22499 (N_22499,N_19131,N_18772);
nand U22500 (N_22500,N_20107,N_21521);
xnor U22501 (N_22501,N_20279,N_21635);
or U22502 (N_22502,N_22271,N_21299);
xnor U22503 (N_22503,N_21801,N_20843);
nor U22504 (N_22504,N_20505,N_21633);
and U22505 (N_22505,N_20084,N_20424);
or U22506 (N_22506,N_20239,N_22300);
and U22507 (N_22507,N_22058,N_21509);
xnor U22508 (N_22508,N_20704,N_20834);
nand U22509 (N_22509,N_20861,N_21780);
nor U22510 (N_22510,N_20284,N_21857);
and U22511 (N_22511,N_20908,N_22257);
and U22512 (N_22512,N_20923,N_20484);
nor U22513 (N_22513,N_21649,N_20990);
nand U22514 (N_22514,N_20150,N_20082);
xor U22515 (N_22515,N_21277,N_21750);
or U22516 (N_22516,N_21420,N_22329);
or U22517 (N_22517,N_20862,N_20551);
and U22518 (N_22518,N_20492,N_21751);
and U22519 (N_22519,N_20606,N_20869);
and U22520 (N_22520,N_20522,N_22273);
and U22521 (N_22521,N_21659,N_21217);
nor U22522 (N_22522,N_22274,N_21760);
nand U22523 (N_22523,N_22135,N_20166);
and U22524 (N_22524,N_20087,N_20963);
nor U22525 (N_22525,N_22336,N_20197);
nand U22526 (N_22526,N_20219,N_21556);
nor U22527 (N_22527,N_20103,N_20318);
nor U22528 (N_22528,N_20732,N_21957);
nor U22529 (N_22529,N_22203,N_20675);
xnor U22530 (N_22530,N_21518,N_20609);
xor U22531 (N_22531,N_20473,N_20479);
or U22532 (N_22532,N_20196,N_21411);
xor U22533 (N_22533,N_20858,N_20835);
and U22534 (N_22534,N_20693,N_20199);
xnor U22535 (N_22535,N_21944,N_22068);
xnor U22536 (N_22536,N_21938,N_22441);
and U22537 (N_22537,N_22121,N_20477);
nor U22538 (N_22538,N_22376,N_20517);
and U22539 (N_22539,N_21579,N_20410);
nand U22540 (N_22540,N_21807,N_20458);
nor U22541 (N_22541,N_20626,N_20648);
xor U22542 (N_22542,N_20554,N_21464);
nor U22543 (N_22543,N_21990,N_20830);
and U22544 (N_22544,N_22155,N_21490);
and U22545 (N_22545,N_21914,N_21295);
nor U22546 (N_22546,N_21992,N_20922);
xnor U22547 (N_22547,N_21557,N_21113);
xor U22548 (N_22548,N_21347,N_21454);
and U22549 (N_22549,N_22287,N_22298);
or U22550 (N_22550,N_20428,N_20540);
xnor U22551 (N_22551,N_21993,N_22136);
or U22552 (N_22552,N_20478,N_21928);
xnor U22553 (N_22553,N_22031,N_21244);
and U22554 (N_22554,N_21466,N_20232);
nand U22555 (N_22555,N_21162,N_21543);
and U22556 (N_22556,N_20400,N_21772);
nand U22557 (N_22557,N_21744,N_20992);
or U22558 (N_22558,N_21813,N_20299);
xnor U22559 (N_22559,N_20737,N_20287);
xnor U22560 (N_22560,N_22333,N_21359);
xor U22561 (N_22561,N_20653,N_20720);
or U22562 (N_22562,N_21484,N_20759);
nand U22563 (N_22563,N_21125,N_21907);
nand U22564 (N_22564,N_20772,N_21200);
nor U22565 (N_22565,N_22045,N_20384);
and U22566 (N_22566,N_22489,N_22123);
or U22567 (N_22567,N_20355,N_22451);
or U22568 (N_22568,N_21191,N_21708);
or U22569 (N_22569,N_22067,N_20877);
nor U22570 (N_22570,N_21842,N_21847);
nand U22571 (N_22571,N_20128,N_21546);
xnor U22572 (N_22572,N_22106,N_20046);
nor U22573 (N_22573,N_21391,N_20102);
and U22574 (N_22574,N_20680,N_20707);
xnor U22575 (N_22575,N_22390,N_21048);
nand U22576 (N_22576,N_21925,N_21169);
nor U22577 (N_22577,N_21657,N_21201);
xor U22578 (N_22578,N_22127,N_21401);
xnor U22579 (N_22579,N_21565,N_21778);
xnor U22580 (N_22580,N_22150,N_20892);
nor U22581 (N_22581,N_20138,N_21493);
xor U22582 (N_22582,N_20174,N_20326);
or U22583 (N_22583,N_20701,N_21333);
nand U22584 (N_22584,N_20225,N_21810);
or U22585 (N_22585,N_20209,N_20577);
nor U22586 (N_22586,N_22404,N_20426);
and U22587 (N_22587,N_21133,N_21446);
xor U22588 (N_22588,N_20726,N_20635);
xnor U22589 (N_22589,N_22152,N_20984);
nand U22590 (N_22590,N_21507,N_20289);
or U22591 (N_22591,N_21770,N_21319);
nor U22592 (N_22592,N_20186,N_21260);
nand U22593 (N_22593,N_20934,N_22138);
xnor U22594 (N_22594,N_22165,N_22221);
nor U22595 (N_22595,N_20350,N_20709);
nor U22596 (N_22596,N_22284,N_20981);
xnor U22597 (N_22597,N_20555,N_20367);
xnor U22598 (N_22598,N_21423,N_21276);
or U22599 (N_22599,N_20283,N_22464);
nand U22600 (N_22600,N_20538,N_21433);
nor U22601 (N_22601,N_21603,N_21594);
xnor U22602 (N_22602,N_20987,N_21838);
xor U22603 (N_22603,N_20148,N_21562);
nor U22604 (N_22604,N_21432,N_21566);
nor U22605 (N_22605,N_20443,N_20574);
nor U22606 (N_22606,N_22264,N_21478);
nand U22607 (N_22607,N_20489,N_21979);
nand U22608 (N_22608,N_20749,N_22417);
and U22609 (N_22609,N_22492,N_20278);
xnor U22610 (N_22610,N_20831,N_22187);
or U22611 (N_22611,N_20151,N_22151);
nor U22612 (N_22612,N_20785,N_21101);
xor U22613 (N_22613,N_20994,N_22370);
nor U22614 (N_22614,N_20997,N_22076);
and U22615 (N_22615,N_22321,N_21088);
or U22616 (N_22616,N_21046,N_21430);
and U22617 (N_22617,N_21910,N_21749);
or U22618 (N_22618,N_22430,N_22447);
xnor U22619 (N_22619,N_22269,N_20180);
xor U22620 (N_22620,N_20684,N_20440);
xnor U22621 (N_22621,N_20565,N_22367);
xnor U22622 (N_22622,N_22178,N_21149);
xnor U22623 (N_22623,N_21077,N_22471);
nor U22624 (N_22624,N_21777,N_20114);
and U22625 (N_22625,N_21998,N_21026);
nor U22626 (N_22626,N_20872,N_21214);
nor U22627 (N_22627,N_22279,N_21577);
and U22628 (N_22628,N_21554,N_21398);
nand U22629 (N_22629,N_21251,N_21654);
nand U22630 (N_22630,N_21908,N_22019);
nor U22631 (N_22631,N_20634,N_21817);
xnor U22632 (N_22632,N_20343,N_20904);
and U22633 (N_22633,N_22387,N_21835);
nand U22634 (N_22634,N_21736,N_21177);
and U22635 (N_22635,N_21141,N_20322);
nor U22636 (N_22636,N_22224,N_21012);
and U22637 (N_22637,N_22063,N_21404);
xnor U22638 (N_22638,N_21374,N_20657);
or U22639 (N_22639,N_21618,N_21656);
and U22640 (N_22640,N_21519,N_21109);
xnor U22641 (N_22641,N_21589,N_22359);
nor U22642 (N_22642,N_21033,N_21245);
and U22643 (N_22643,N_20340,N_21799);
nor U22644 (N_22644,N_20051,N_22338);
nand U22645 (N_22645,N_20005,N_22236);
nor U22646 (N_22646,N_20569,N_20613);
nor U22647 (N_22647,N_21968,N_22427);
or U22648 (N_22648,N_21055,N_20757);
or U22649 (N_22649,N_22207,N_21246);
and U22650 (N_22650,N_21686,N_21087);
or U22651 (N_22651,N_21886,N_20253);
or U22652 (N_22652,N_20851,N_20794);
and U22653 (N_22653,N_22487,N_21131);
or U22654 (N_22654,N_21729,N_21114);
or U22655 (N_22655,N_20585,N_21505);
nand U22656 (N_22656,N_21892,N_20703);
or U22657 (N_22657,N_22073,N_21072);
and U22658 (N_22658,N_22107,N_22049);
nor U22659 (N_22659,N_20481,N_20805);
or U22660 (N_22660,N_20642,N_21850);
nor U22661 (N_22661,N_21220,N_21844);
nor U22662 (N_22662,N_20292,N_21210);
and U22663 (N_22663,N_20235,N_21935);
nand U22664 (N_22664,N_21642,N_21779);
xor U22665 (N_22665,N_20290,N_20752);
nand U22666 (N_22666,N_21877,N_21628);
or U22667 (N_22667,N_21984,N_20406);
nor U22668 (N_22668,N_20042,N_20931);
or U22669 (N_22669,N_21231,N_21624);
xor U22670 (N_22670,N_22122,N_20049);
and U22671 (N_22671,N_21690,N_20572);
or U22672 (N_22672,N_21467,N_21255);
and U22673 (N_22673,N_21631,N_20476);
or U22674 (N_22674,N_21038,N_21375);
nor U22675 (N_22675,N_22188,N_20695);
or U22676 (N_22676,N_22444,N_20860);
or U22677 (N_22677,N_20527,N_20890);
and U22678 (N_22678,N_20271,N_20390);
nor U22679 (N_22679,N_21314,N_21593);
nor U22680 (N_22680,N_20825,N_20142);
or U22681 (N_22681,N_22088,N_20706);
or U22682 (N_22682,N_20317,N_21897);
nand U22683 (N_22683,N_21045,N_20395);
xor U22684 (N_22684,N_21815,N_21717);
nand U22685 (N_22685,N_21014,N_21443);
nor U22686 (N_22686,N_20029,N_20467);
and U22687 (N_22687,N_22091,N_22109);
and U22688 (N_22688,N_21115,N_22498);
xor U22689 (N_22689,N_22086,N_21463);
xnor U22690 (N_22690,N_21158,N_21481);
and U22691 (N_22691,N_21684,N_20865);
and U22692 (N_22692,N_20070,N_21940);
nand U22693 (N_22693,N_22227,N_21735);
nor U22694 (N_22694,N_21117,N_21501);
nand U22695 (N_22695,N_22278,N_20829);
and U22696 (N_22696,N_22015,N_20113);
nand U22697 (N_22697,N_21187,N_20856);
and U22698 (N_22698,N_21873,N_20583);
nand U22699 (N_22699,N_20265,N_21473);
nor U22700 (N_22700,N_20779,N_22050);
or U22701 (N_22701,N_20533,N_20407);
nand U22702 (N_22702,N_21822,N_20286);
nor U22703 (N_22703,N_21915,N_22422);
or U22704 (N_22704,N_21899,N_21176);
nand U22705 (N_22705,N_21129,N_21243);
and U22706 (N_22706,N_21852,N_20991);
or U22707 (N_22707,N_22052,N_20535);
nor U22708 (N_22708,N_21737,N_20072);
or U22709 (N_22709,N_20466,N_20778);
and U22710 (N_22710,N_21261,N_20285);
and U22711 (N_22711,N_21235,N_20268);
nor U22712 (N_22712,N_22405,N_20414);
nand U22713 (N_22713,N_22162,N_22283);
nor U22714 (N_22714,N_20813,N_22199);
or U22715 (N_22715,N_20913,N_21880);
or U22716 (N_22716,N_20425,N_21067);
nor U22717 (N_22717,N_22130,N_22065);
or U22718 (N_22718,N_20347,N_20708);
xor U22719 (N_22719,N_22032,N_20669);
and U22720 (N_22720,N_21480,N_20746);
or U22721 (N_22721,N_22000,N_21174);
nor U22722 (N_22722,N_21280,N_21558);
or U22723 (N_22723,N_22411,N_21161);
and U22724 (N_22724,N_20625,N_21193);
or U22725 (N_22725,N_20989,N_21821);
or U22726 (N_22726,N_21641,N_20020);
nand U22727 (N_22727,N_21585,N_21450);
or U22728 (N_22728,N_22348,N_20777);
or U22729 (N_22729,N_22096,N_20526);
nand U22730 (N_22730,N_21494,N_21190);
xnor U22731 (N_22731,N_20611,N_21268);
nand U22732 (N_22732,N_21234,N_21078);
and U22733 (N_22733,N_20246,N_20823);
xnor U22734 (N_22734,N_20064,N_20628);
nand U22735 (N_22735,N_20164,N_20631);
nor U22736 (N_22736,N_21535,N_21582);
xnor U22737 (N_22737,N_21954,N_21284);
and U22738 (N_22738,N_22097,N_20584);
xnor U22739 (N_22739,N_21966,N_21932);
and U22740 (N_22740,N_21592,N_20968);
and U22741 (N_22741,N_21074,N_22239);
nor U22742 (N_22742,N_22228,N_21611);
xor U22743 (N_22743,N_22331,N_21977);
nand U22744 (N_22744,N_20621,N_22351);
and U22745 (N_22745,N_22077,N_20169);
or U22746 (N_22746,N_21983,N_22134);
nand U22747 (N_22747,N_22212,N_20422);
nand U22748 (N_22748,N_21459,N_20048);
nand U22749 (N_22749,N_22053,N_21264);
xnor U22750 (N_22750,N_22094,N_20755);
and U22751 (N_22751,N_20038,N_20412);
or U22752 (N_22752,N_22409,N_20172);
xnor U22753 (N_22753,N_21516,N_21016);
nand U22754 (N_22754,N_20610,N_21971);
nor U22755 (N_22755,N_20885,N_20773);
and U22756 (N_22756,N_20195,N_21923);
nor U22757 (N_22757,N_21901,N_20145);
nor U22758 (N_22758,N_21989,N_20076);
xnor U22759 (N_22759,N_20697,N_20000);
nor U22760 (N_22760,N_20506,N_20576);
xnor U22761 (N_22761,N_22243,N_21912);
or U22762 (N_22762,N_20089,N_21322);
nor U22763 (N_22763,N_22358,N_20348);
nand U22764 (N_22764,N_21706,N_20760);
and U22765 (N_22765,N_21279,N_20270);
nand U22766 (N_22766,N_21303,N_22310);
nand U22767 (N_22767,N_21053,N_21943);
and U22768 (N_22768,N_21597,N_20795);
xnor U22769 (N_22769,N_20266,N_21636);
nand U22770 (N_22770,N_21181,N_21561);
nor U22771 (N_22771,N_21685,N_21574);
or U22772 (N_22772,N_21816,N_20966);
and U22773 (N_22773,N_22491,N_20446);
nand U22774 (N_22774,N_21655,N_21147);
and U22775 (N_22775,N_20101,N_21236);
and U22776 (N_22776,N_20544,N_21694);
nand U22777 (N_22777,N_22379,N_20346);
xnor U22778 (N_22778,N_21394,N_20563);
and U22779 (N_22779,N_21027,N_21017);
nor U22780 (N_22780,N_21604,N_20105);
nand U22781 (N_22781,N_21136,N_21428);
or U22782 (N_22782,N_21044,N_21138);
xor U22783 (N_22783,N_20623,N_20601);
nand U22784 (N_22784,N_20809,N_20294);
nand U22785 (N_22785,N_20252,N_20342);
or U22786 (N_22786,N_22197,N_20911);
xnor U22787 (N_22787,N_20881,N_20824);
and U22788 (N_22788,N_20470,N_22309);
nor U22789 (N_22789,N_21005,N_20821);
nand U22790 (N_22790,N_21792,N_21447);
and U22791 (N_22791,N_22114,N_22128);
and U22792 (N_22792,N_22173,N_20345);
nor U22793 (N_22793,N_21682,N_20028);
xor U22794 (N_22794,N_20335,N_21793);
nor U22795 (N_22795,N_20850,N_20220);
nand U22796 (N_22796,N_22395,N_21922);
nand U22797 (N_22797,N_20661,N_20297);
and U22798 (N_22798,N_20887,N_21457);
or U22799 (N_22799,N_20321,N_20808);
nor U22800 (N_22800,N_21440,N_22182);
nor U22801 (N_22801,N_20723,N_21228);
xnor U22802 (N_22802,N_21036,N_22011);
nand U22803 (N_22803,N_21195,N_21542);
xor U22804 (N_22804,N_20663,N_20144);
nand U22805 (N_22805,N_20358,N_22057);
and U22806 (N_22806,N_21878,N_20036);
or U22807 (N_22807,N_22026,N_22434);
nor U22808 (N_22808,N_22323,N_20275);
or U22809 (N_22809,N_20421,N_22380);
and U22810 (N_22810,N_21933,N_21049);
xor U22811 (N_22811,N_21080,N_20387);
or U22812 (N_22812,N_20907,N_20498);
or U22813 (N_22813,N_21084,N_21266);
nor U22814 (N_22814,N_21950,N_20534);
xor U22815 (N_22815,N_22147,N_21119);
xnor U22816 (N_22816,N_21757,N_21165);
xnor U22817 (N_22817,N_20462,N_21728);
nand U22818 (N_22818,N_20351,N_21258);
nand U22819 (N_22819,N_21569,N_21707);
xor U22820 (N_22820,N_20868,N_22347);
nand U22821 (N_22821,N_20403,N_20231);
or U22822 (N_22822,N_22392,N_21959);
or U22823 (N_22823,N_21834,N_20018);
nor U22824 (N_22824,N_20328,N_20692);
or U22825 (N_22825,N_20641,N_20378);
nor U22826 (N_22826,N_22215,N_22341);
or U22827 (N_22827,N_21904,N_20796);
nand U22828 (N_22828,N_20874,N_22252);
or U22829 (N_22829,N_20415,N_22368);
and U22830 (N_22830,N_20152,N_21667);
nor U22831 (N_22831,N_21894,N_20333);
or U22832 (N_22832,N_20614,N_20799);
or U22833 (N_22833,N_21032,N_21610);
or U22834 (N_22834,N_21293,N_22175);
nand U22835 (N_22835,N_21285,N_21202);
nor U22836 (N_22836,N_20127,N_21924);
xor U22837 (N_22837,N_21126,N_21326);
xor U22838 (N_22838,N_21462,N_22126);
and U22839 (N_22839,N_20839,N_20095);
or U22840 (N_22840,N_21071,N_21124);
nor U22841 (N_22841,N_20735,N_20662);
or U22842 (N_22842,N_20451,N_21424);
or U22843 (N_22843,N_21584,N_21328);
nand U22844 (N_22844,N_22476,N_21881);
and U22845 (N_22845,N_22081,N_21186);
and U22846 (N_22846,N_20909,N_21302);
and U22847 (N_22847,N_21586,N_20916);
xnor U22848 (N_22848,N_22132,N_22457);
or U22849 (N_22849,N_20019,N_21468);
xor U22850 (N_22850,N_22322,N_21092);
nand U22851 (N_22851,N_22435,N_21313);
nor U22852 (N_22852,N_22270,N_20818);
nand U22853 (N_22853,N_20305,N_20588);
or U22854 (N_22854,N_20023,N_21762);
nor U22855 (N_22855,N_20817,N_22399);
nand U22856 (N_22856,N_21290,N_20147);
nor U22857 (N_22857,N_21864,N_22332);
xor U22858 (N_22858,N_22095,N_20007);
nand U22859 (N_22859,N_21547,N_20959);
or U22860 (N_22860,N_21363,N_22148);
nor U22861 (N_22861,N_22033,N_21184);
nand U22862 (N_22862,N_20591,N_20394);
or U22863 (N_22863,N_22013,N_21354);
nand U22864 (N_22864,N_20254,N_21068);
nor U22865 (N_22865,N_21112,N_21890);
or U22866 (N_22866,N_21796,N_21931);
nor U22867 (N_22867,N_20003,N_21323);
or U22868 (N_22868,N_21309,N_22497);
nor U22869 (N_22869,N_21645,N_20770);
or U22870 (N_22870,N_20359,N_22198);
nor U22871 (N_22871,N_22385,N_20941);
nand U22872 (N_22872,N_20751,N_22056);
nand U22873 (N_22873,N_20957,N_22048);
xor U22874 (N_22874,N_21221,N_20397);
xnor U22875 (N_22875,N_20867,N_22115);
and U22876 (N_22876,N_22458,N_22041);
xor U22877 (N_22877,N_21937,N_21608);
xor U22878 (N_22878,N_20699,N_20999);
xnor U22879 (N_22879,N_21951,N_22116);
or U22880 (N_22880,N_21035,N_21942);
nor U22881 (N_22881,N_22429,N_20607);
nor U22882 (N_22882,N_21709,N_20250);
nand U22883 (N_22883,N_21100,N_22070);
or U22884 (N_22884,N_20983,N_20686);
nor U22885 (N_22885,N_21142,N_20883);
nor U22886 (N_22886,N_20181,N_20579);
nand U22887 (N_22887,N_21360,N_22064);
and U22888 (N_22888,N_20120,N_21598);
nand U22889 (N_22889,N_20814,N_20083);
nor U22890 (N_22890,N_21758,N_20753);
nor U22891 (N_22891,N_21576,N_20188);
nand U22892 (N_22892,N_20832,N_20846);
and U22893 (N_22893,N_21530,N_20501);
nor U22894 (N_22894,N_22223,N_20810);
and U22895 (N_22895,N_20902,N_21389);
or U22896 (N_22896,N_22371,N_22245);
nor U22897 (N_22897,N_21564,N_21110);
nor U22898 (N_22898,N_20622,N_21339);
and U22899 (N_22899,N_20603,N_22410);
and U22900 (N_22900,N_21862,N_20047);
nor U22901 (N_22901,N_21687,N_20488);
nand U22902 (N_22902,N_22075,N_21330);
xor U22903 (N_22903,N_21733,N_21712);
and U22904 (N_22904,N_20004,N_20391);
and U22905 (N_22905,N_21437,N_21726);
xor U22906 (N_22906,N_22205,N_20500);
and U22907 (N_22907,N_20323,N_21015);
nand U22908 (N_22908,N_21525,N_20100);
and U22909 (N_22909,N_21056,N_21194);
or U22910 (N_22910,N_22299,N_21705);
and U22911 (N_22911,N_21668,N_20721);
or U22912 (N_22912,N_20092,N_20056);
or U22913 (N_22913,N_20096,N_22432);
nor U22914 (N_22914,N_21300,N_20034);
nand U22915 (N_22915,N_22420,N_21975);
or U22916 (N_22916,N_22060,N_22216);
nand U22917 (N_22917,N_21102,N_22484);
nor U22918 (N_22918,N_21541,N_20217);
and U22919 (N_22919,N_20205,N_20401);
nor U22920 (N_22920,N_21412,N_21622);
xnor U22921 (N_22921,N_20496,N_21527);
nor U22922 (N_22922,N_20936,N_20898);
nor U22923 (N_22923,N_20894,N_20947);
xnor U22924 (N_22924,N_21745,N_22112);
nand U22925 (N_22925,N_20893,N_21647);
xnor U22926 (N_22926,N_21306,N_22294);
nand U22927 (N_22927,N_21452,N_21637);
xnor U22928 (N_22928,N_20605,N_21572);
and U22929 (N_22929,N_20800,N_20025);
or U22930 (N_22930,N_21680,N_21583);
and U22931 (N_22931,N_21742,N_21601);
nor U22932 (N_22932,N_20929,N_21054);
xor U22933 (N_22933,N_20192,N_20393);
xnor U22934 (N_22934,N_20306,N_21848);
nor U22935 (N_22935,N_20719,N_21116);
and U22936 (N_22936,N_20198,N_22483);
nor U22937 (N_22937,N_22423,N_20943);
xor U22938 (N_22938,N_20654,N_20949);
nor U22939 (N_22939,N_21106,N_21781);
or U22940 (N_22940,N_20320,N_21639);
nand U22941 (N_22941,N_20903,N_21192);
and U22942 (N_22942,N_20967,N_20982);
and U22943 (N_22943,N_21765,N_21876);
and U22944 (N_22944,N_20149,N_20878);
and U22945 (N_22945,N_21427,N_21902);
or U22946 (N_22946,N_20153,N_22046);
or U22947 (N_22947,N_20157,N_20932);
nand U22948 (N_22948,N_22449,N_20889);
nor U22949 (N_22949,N_22494,N_21551);
and U22950 (N_22950,N_21338,N_21520);
nand U22951 (N_22951,N_20612,N_20691);
and U22952 (N_22952,N_20261,N_20132);
nor U22953 (N_22953,N_20389,N_21723);
and U22954 (N_22954,N_21840,N_20876);
nor U22955 (N_22955,N_22235,N_20314);
nand U22956 (N_22956,N_20366,N_21458);
nand U22957 (N_22957,N_20739,N_22231);
and U22958 (N_22958,N_22185,N_21063);
and U22959 (N_22959,N_21976,N_22098);
nor U22960 (N_22960,N_21486,N_22470);
nor U22961 (N_22961,N_20396,N_20357);
nand U22962 (N_22962,N_21963,N_20134);
and U22963 (N_22963,N_21416,N_22225);
xnor U22964 (N_22964,N_22263,N_20556);
nand U22965 (N_22965,N_20870,N_20586);
nand U22966 (N_22966,N_21410,N_21640);
and U22967 (N_22967,N_21393,N_20093);
and U22968 (N_22968,N_22397,N_21858);
and U22969 (N_22969,N_22232,N_20679);
nor U22970 (N_22970,N_21383,N_21934);
nor U22971 (N_22971,N_21230,N_20660);
nand U22972 (N_22972,N_20079,N_21075);
or U22973 (N_22973,N_22438,N_21528);
xor U22974 (N_22974,N_20125,N_20895);
xnor U22975 (N_22975,N_20696,N_22428);
nor U22976 (N_22976,N_21365,N_20081);
or U22977 (N_22977,N_21444,N_20175);
xor U22978 (N_22978,N_21345,N_22177);
nand U22979 (N_22979,N_20244,N_21948);
xor U22980 (N_22980,N_20578,N_22490);
and U22981 (N_22981,N_20480,N_20154);
nand U22982 (N_22982,N_20670,N_21034);
nand U22983 (N_22983,N_21698,N_22194);
xnor U22984 (N_22984,N_20986,N_20897);
xor U22985 (N_22985,N_20840,N_21414);
nor U22986 (N_22986,N_21377,N_20027);
xor U22987 (N_22987,N_21679,N_22149);
nand U22988 (N_22988,N_21089,N_22025);
xnor U22989 (N_22989,N_22102,N_21920);
nand U22990 (N_22990,N_20596,N_20449);
and U22991 (N_22991,N_22377,N_20155);
and U22992 (N_22992,N_21121,N_20536);
nor U22993 (N_22993,N_21238,N_20065);
nor U22994 (N_22994,N_21538,N_20854);
and U22995 (N_22995,N_22043,N_20516);
xnor U22996 (N_22996,N_22454,N_22030);
and U22997 (N_22997,N_20781,N_22036);
nor U22998 (N_22998,N_20274,N_21417);
nor U22999 (N_22999,N_21316,N_21178);
xor U23000 (N_23000,N_22266,N_22140);
and U23001 (N_23001,N_21638,N_20106);
nor U23002 (N_23002,N_21590,N_20515);
xnor U23003 (N_23003,N_21057,N_21134);
nor U23004 (N_23004,N_21919,N_20059);
or U23005 (N_23005,N_20728,N_20822);
nor U23006 (N_23006,N_20381,N_21241);
or U23007 (N_23007,N_21843,N_20216);
and U23008 (N_23008,N_20456,N_21956);
nor U23009 (N_23009,N_21491,N_21146);
or U23010 (N_23010,N_22373,N_21826);
nor U23011 (N_23011,N_20549,N_21421);
and U23012 (N_23012,N_22424,N_20423);
nand U23013 (N_23013,N_21903,N_21537);
xor U23014 (N_23014,N_21615,N_21160);
nand U23015 (N_23015,N_21725,N_21312);
and U23016 (N_23016,N_20671,N_20330);
nor U23017 (N_23017,N_22110,N_22414);
xor U23018 (N_23018,N_22349,N_20802);
or U23019 (N_23019,N_21581,N_20140);
and U23020 (N_23020,N_21946,N_20067);
and U23021 (N_23021,N_21820,N_21349);
or U23022 (N_23022,N_20530,N_20882);
or U23023 (N_23023,N_21171,N_20429);
or U23024 (N_23024,N_21855,N_20159);
nor U23025 (N_23025,N_20906,N_21732);
nand U23026 (N_23026,N_21665,N_22253);
nor U23027 (N_23027,N_21763,N_21105);
and U23028 (N_23028,N_21399,N_21651);
or U23029 (N_23029,N_22291,N_21434);
or U23030 (N_23030,N_21856,N_22211);
and U23031 (N_23031,N_21958,N_21371);
nand U23032 (N_23032,N_21104,N_21062);
or U23033 (N_23033,N_21381,N_22327);
nand U23034 (N_23034,N_21870,N_21508);
nand U23035 (N_23035,N_20380,N_20315);
or U23036 (N_23036,N_21213,N_21607);
nand U23037 (N_23037,N_20071,N_20228);
nor U23038 (N_23038,N_21691,N_22244);
nand U23039 (N_23039,N_22229,N_21692);
xnor U23040 (N_23040,N_21011,N_21866);
and U23041 (N_23041,N_22084,N_21634);
nand U23042 (N_23042,N_20630,N_22014);
xnor U23043 (N_23043,N_20838,N_20559);
nor U23044 (N_23044,N_22038,N_22002);
or U23045 (N_23045,N_20645,N_21941);
xnor U23046 (N_23046,N_22167,N_20420);
nor U23047 (N_23047,N_20097,N_21361);
or U23048 (N_23048,N_20765,N_20483);
or U23049 (N_23049,N_21311,N_22445);
and U23050 (N_23050,N_21091,N_20112);
or U23051 (N_23051,N_22394,N_22328);
and U23052 (N_23052,N_22054,N_21321);
nand U23053 (N_23053,N_20191,N_21419);
xnor U23054 (N_23054,N_20633,N_22452);
and U23055 (N_23055,N_22103,N_22442);
and U23056 (N_23056,N_20013,N_20363);
nand U23057 (N_23057,N_20873,N_20915);
and U23058 (N_23058,N_20589,N_21324);
or U23059 (N_23059,N_20465,N_21677);
or U23060 (N_23060,N_22201,N_21152);
nand U23061 (N_23061,N_22415,N_21836);
or U23062 (N_23062,N_20043,N_21713);
and U23063 (N_23063,N_22413,N_20667);
nor U23064 (N_23064,N_20638,N_20532);
and U23065 (N_23065,N_21079,N_21352);
nand U23066 (N_23066,N_20694,N_20241);
nor U23067 (N_23067,N_20190,N_20365);
or U23068 (N_23068,N_21663,N_22391);
nor U23069 (N_23069,N_20319,N_20441);
or U23070 (N_23070,N_20119,N_21672);
and U23071 (N_23071,N_21259,N_22383);
nand U23072 (N_23072,N_20541,N_20672);
and U23073 (N_23073,N_21402,N_20560);
nor U23074 (N_23074,N_21180,N_20958);
nand U23075 (N_23075,N_20828,N_21678);
nand U23076 (N_23076,N_20267,N_20552);
nor U23077 (N_23077,N_21719,N_20183);
nor U23078 (N_23078,N_21052,N_20940);
and U23079 (N_23079,N_21372,N_20845);
xor U23080 (N_23080,N_21753,N_21043);
or U23081 (N_23081,N_20313,N_20998);
and U23082 (N_23082,N_21747,N_20954);
xnor U23083 (N_23083,N_21553,N_21004);
and U23084 (N_23084,N_21872,N_21776);
or U23085 (N_23085,N_20702,N_21693);
and U23086 (N_23086,N_20309,N_21408);
nor U23087 (N_23087,N_21327,N_20689);
or U23088 (N_23088,N_20080,N_20411);
nand U23089 (N_23089,N_20417,N_21288);
nand U23090 (N_23090,N_20201,N_21827);
or U23091 (N_23091,N_20073,N_21369);
and U23092 (N_23092,N_21301,N_21442);
and U23093 (N_23093,N_22374,N_21911);
nand U23094 (N_23094,N_21814,N_21529);
nor U23095 (N_23095,N_21823,N_20497);
and U23096 (N_23096,N_21097,N_21479);
nor U23097 (N_23097,N_22164,N_22183);
xor U23098 (N_23098,N_21967,N_21185);
nand U23099 (N_23099,N_22354,N_20039);
and U23100 (N_23100,N_22499,N_20644);
and U23101 (N_23101,N_21504,N_21289);
nor U23102 (N_23102,N_20006,N_21451);
nor U23103 (N_23103,N_20581,N_21083);
or U23104 (N_23104,N_22143,N_20762);
xnor U23105 (N_23105,N_21580,N_20964);
and U23106 (N_23106,N_21155,N_20754);
xor U23107 (N_23107,N_21273,N_20859);
and U23108 (N_23108,N_22093,N_21829);
xnor U23109 (N_23109,N_21175,N_20117);
and U23110 (N_23110,N_21804,N_22007);
xnor U23111 (N_23111,N_21661,N_20063);
and U23112 (N_23112,N_21851,N_20260);
nor U23113 (N_23113,N_20126,N_22133);
and U23114 (N_23114,N_22277,N_20924);
nor U23115 (N_23115,N_20944,N_21346);
and U23116 (N_23116,N_22469,N_21304);
nor U23117 (N_23117,N_21837,N_20041);
nand U23118 (N_23118,N_22467,N_20058);
xor U23119 (N_23119,N_20742,N_20222);
xnor U23120 (N_23120,N_20602,N_21379);
and U23121 (N_23121,N_20372,N_20568);
nand U23122 (N_23122,N_22472,N_22010);
and U23123 (N_23123,N_20194,N_22171);
nand U23124 (N_23124,N_22267,N_20237);
and U23125 (N_23125,N_21341,N_21426);
and U23126 (N_23126,N_20637,N_20632);
xnor U23127 (N_23127,N_20062,N_21960);
and U23128 (N_23128,N_21358,N_20727);
nor U23129 (N_23129,N_20567,N_21620);
and U23130 (N_23130,N_22440,N_22190);
or U23131 (N_23131,N_22419,N_21673);
xor U23132 (N_23132,N_21150,N_21513);
nand U23133 (N_23133,N_21415,N_20961);
xnor U23134 (N_23134,N_20337,N_20598);
nor U23135 (N_23135,N_20160,N_20135);
nand U23136 (N_23136,N_21222,N_21031);
nor U23137 (N_23137,N_21800,N_22265);
nand U23138 (N_23138,N_21144,N_21845);
and U23139 (N_23139,N_21536,N_21961);
nand U23140 (N_23140,N_22308,N_21643);
nor U23141 (N_23141,N_20281,N_21489);
and U23142 (N_23142,N_20548,N_22035);
or U23143 (N_23143,N_22272,N_22268);
xnor U23144 (N_23144,N_21986,N_20111);
nor U23145 (N_23145,N_21107,N_21795);
and U23146 (N_23146,N_22478,N_22193);
or U23147 (N_23147,N_21335,N_21867);
or U23148 (N_23148,N_21808,N_20764);
nand U23149 (N_23149,N_22319,N_22393);
nor U23150 (N_23150,N_21145,N_21949);
nand U23151 (N_23151,N_21973,N_21179);
nand U23152 (N_23152,N_21108,N_21215);
and U23153 (N_23153,N_20690,N_21969);
xor U23154 (N_23154,N_20938,N_21738);
and U23155 (N_23155,N_22008,N_20121);
and U23156 (N_23156,N_20733,N_20833);
and U23157 (N_23157,N_20408,N_21283);
and U23158 (N_23158,N_21127,N_20055);
or U23159 (N_23159,N_20061,N_21006);
nor U23160 (N_23160,N_22131,N_21061);
and U23161 (N_23161,N_20768,N_22021);
nand U23162 (N_23162,N_20993,N_20826);
or U23163 (N_23163,N_22479,N_22255);
nor U23164 (N_23164,N_22456,N_20213);
and U23165 (N_23165,N_20539,N_20942);
nand U23166 (N_23166,N_20156,N_20431);
xor U23167 (N_23167,N_20507,N_21570);
xnor U23168 (N_23168,N_20187,N_21721);
nand U23169 (N_23169,N_22326,N_20341);
nand U23170 (N_23170,N_21522,N_20597);
or U23171 (N_23171,N_21588,N_20016);
xor U23172 (N_23172,N_21128,N_21094);
nand U23173 (N_23173,N_20077,N_20091);
nand U23174 (N_23174,N_20946,N_20962);
xor U23175 (N_23175,N_20710,N_21167);
nand U23176 (N_23176,N_20978,N_21240);
or U23177 (N_23177,N_20088,N_20837);
or U23178 (N_23178,N_21809,N_20439);
xor U23179 (N_23179,N_22468,N_20980);
nor U23180 (N_23180,N_20248,N_21010);
xor U23181 (N_23181,N_22023,N_21157);
nor U23182 (N_23182,N_22344,N_21366);
and U23183 (N_23183,N_21252,N_22361);
nand U23184 (N_23184,N_22408,N_21153);
and U23185 (N_23185,N_20469,N_20053);
and U23186 (N_23186,N_20774,N_21761);
nor U23187 (N_23187,N_20618,N_21906);
nand U23188 (N_23188,N_20383,N_21096);
or U23189 (N_23189,N_21270,N_21025);
nor U23190 (N_23190,N_21882,N_22184);
or U23191 (N_23191,N_20386,N_21249);
nor U23192 (N_23192,N_20951,N_21086);
nand U23193 (N_23193,N_20471,N_21343);
nor U23194 (N_23194,N_22485,N_20399);
and U23195 (N_23195,N_20339,N_20740);
nor U23196 (N_23196,N_22219,N_21515);
nand U23197 (N_23197,N_20976,N_20438);
nor U23198 (N_23198,N_22425,N_20712);
xor U23199 (N_23199,N_21262,N_21197);
nand U23200 (N_23200,N_20293,N_21342);
or U23201 (N_23201,N_20482,N_22364);
nand U23202 (N_23202,N_21492,N_20455);
nand U23203 (N_23203,N_21909,N_20952);
or U23204 (N_23204,N_20842,N_21898);
or U23205 (N_23205,N_20123,N_22317);
nor U23206 (N_23206,N_20879,N_22463);
nor U23207 (N_23207,N_20717,N_20173);
nand U23208 (N_23208,N_21787,N_21567);
or U23209 (N_23209,N_20171,N_20224);
xnor U23210 (N_23210,N_21759,N_21884);
xor U23211 (N_23211,N_21790,N_21991);
nand U23212 (N_23212,N_22433,N_21418);
xor U23213 (N_23213,N_22401,N_21429);
xor U23214 (N_23214,N_21103,N_20891);
and U23215 (N_23215,N_20705,N_20747);
or U23216 (N_23216,N_22181,N_20935);
nand U23217 (N_23217,N_20474,N_20599);
nor U23218 (N_23218,N_20682,N_21123);
nor U23219 (N_23219,N_21797,N_20259);
nor U23220 (N_23220,N_21495,N_20002);
nor U23221 (N_23221,N_22087,N_20948);
or U23222 (N_23222,N_22313,N_20640);
nor U23223 (N_23223,N_20880,N_21734);
nor U23224 (N_23224,N_22343,N_21839);
xor U23225 (N_23225,N_21517,N_22362);
or U23226 (N_23226,N_21090,N_22137);
or U23227 (N_23227,N_22249,N_22142);
or U23228 (N_23228,N_22139,N_21775);
xor U23229 (N_23229,N_20032,N_21198);
xnor U23230 (N_23230,N_22186,N_22486);
nor U23231 (N_23231,N_20398,N_21506);
nor U23232 (N_23232,N_22355,N_21545);
nand U23233 (N_23233,N_22386,N_21085);
xor U23234 (N_23234,N_20722,N_20888);
and U23235 (N_23235,N_21294,N_20143);
xnor U23236 (N_23236,N_21390,N_22493);
xnor U23237 (N_23237,N_22360,N_21019);
and U23238 (N_23238,N_21226,N_20900);
or U23239 (N_23239,N_21095,N_22431);
xor U23240 (N_23240,N_20793,N_21018);
nand U23241 (N_23241,N_21465,N_20026);
nor U23242 (N_23242,N_21436,N_21987);
nor U23243 (N_23243,N_20078,N_21784);
and U23244 (N_23244,N_22312,N_21344);
or U23245 (N_23245,N_20620,N_21664);
and U23246 (N_23246,N_21599,N_21703);
xnor U23247 (N_23247,N_20985,N_21207);
nand U23248 (N_23248,N_21806,N_20525);
and U23249 (N_23249,N_20238,N_20262);
nor U23250 (N_23250,N_20131,N_20937);
xor U23251 (N_23251,N_20230,N_20405);
nand U23252 (N_23252,N_22465,N_22311);
nor U23253 (N_23253,N_21563,N_20212);
and U23254 (N_23254,N_22295,N_21503);
and U23255 (N_23255,N_21253,N_21617);
xor U23256 (N_23256,N_21549,N_22350);
xnor U23257 (N_23257,N_21189,N_20687);
nand U23258 (N_23258,N_20184,N_22426);
xnor U23259 (N_23259,N_20256,N_20452);
xor U23260 (N_23260,N_20571,N_20109);
and U23261 (N_23261,N_21887,N_22237);
xor U23262 (N_23262,N_21970,N_21785);
nand U23263 (N_23263,N_20221,N_22448);
nor U23264 (N_23264,N_21208,N_20853);
and U23265 (N_23265,N_20057,N_22439);
and U23266 (N_23266,N_20307,N_21548);
nor U23267 (N_23267,N_21470,N_20920);
and U23268 (N_23268,N_20050,N_20519);
nor U23269 (N_23269,N_20334,N_21889);
nand U23270 (N_23270,N_20756,N_21472);
xnor U23271 (N_23271,N_21982,N_22259);
or U23272 (N_23272,N_20338,N_20996);
xor U23273 (N_23273,N_20282,N_21082);
nand U23274 (N_23274,N_22159,N_22018);
or U23275 (N_23275,N_21318,N_22117);
and U23276 (N_23276,N_21305,N_21774);
and U23277 (N_23277,N_21510,N_21929);
nand U23278 (N_23278,N_20214,N_20402);
and U23279 (N_23279,N_21168,N_21385);
nand U23280 (N_23280,N_21916,N_20392);
nand U23281 (N_23281,N_22466,N_20666);
and U23282 (N_23282,N_21456,N_20110);
xnor U23283 (N_23283,N_20730,N_22125);
xor U23284 (N_23284,N_22316,N_21298);
nand U23285 (N_23285,N_20910,N_20115);
nand U23286 (N_23286,N_21868,N_22334);
and U23287 (N_23287,N_21274,N_20528);
or U23288 (N_23288,N_21746,N_20362);
and U23289 (N_23289,N_20464,N_22337);
or U23290 (N_23290,N_20553,N_21502);
nor U23291 (N_23291,N_20863,N_20014);
nand U23292 (N_23292,N_20921,N_20901);
nor U23293 (N_23293,N_21605,N_20639);
and U23294 (N_23294,N_22482,N_20683);
xor U23295 (N_23295,N_21275,N_20457);
and U23296 (N_23296,N_22153,N_22378);
or U23297 (N_23297,N_21803,N_21353);
or U23298 (N_23298,N_22488,N_22495);
and U23299 (N_23299,N_20035,N_22302);
or U23300 (N_23300,N_21225,N_21482);
nor U23301 (N_23301,N_21137,N_20988);
and U23302 (N_23302,N_21209,N_21786);
nor U23303 (N_23303,N_21173,N_20247);
nand U23304 (N_23304,N_20529,N_20308);
and U23305 (N_23305,N_20801,N_21674);
and U23306 (N_23306,N_20673,N_20771);
xor U23307 (N_23307,N_21571,N_22475);
or U23308 (N_23308,N_20744,N_20665);
and U23309 (N_23309,N_21568,N_21865);
nor U23310 (N_23310,N_21683,N_22290);
and U23311 (N_23311,N_21888,N_20364);
and U23312 (N_23312,N_20060,N_20493);
xnor U23313 (N_23313,N_21040,N_20033);
nor U23314 (N_23314,N_20045,N_22218);
nor U23315 (N_23315,N_20734,N_20783);
or U23316 (N_23316,N_20448,N_21704);
xor U23317 (N_23317,N_21741,N_20327);
xor U23318 (N_23318,N_22398,N_22230);
nand U23319 (N_23319,N_20804,N_21699);
nor U23320 (N_23320,N_21575,N_20445);
nand U23321 (N_23321,N_21955,N_21256);
and U23322 (N_23322,N_21614,N_22192);
nor U23323 (N_23323,N_20463,N_21257);
and U23324 (N_23324,N_22174,N_20504);
nand U23325 (N_23325,N_20136,N_20509);
nor U23326 (N_23326,N_22047,N_21540);
nor U23327 (N_23327,N_22260,N_21695);
xor U23328 (N_23328,N_22365,N_21658);
nand U23329 (N_23329,N_21681,N_20647);
and U23330 (N_23330,N_21748,N_20788);
nand U23331 (N_23331,N_22403,N_21368);
and U23332 (N_23332,N_20273,N_21860);
or U23333 (N_23333,N_20356,N_20736);
xnor U23334 (N_23334,N_21060,N_20437);
nor U23335 (N_23335,N_22204,N_21170);
xor U23336 (N_23336,N_20798,N_22168);
nor U23337 (N_23337,N_20761,N_20316);
nor U23338 (N_23338,N_20382,N_21964);
or U23339 (N_23339,N_20566,N_20502);
nor U23340 (N_23340,N_20031,N_20022);
or U23341 (N_23341,N_22166,N_21697);
and U23342 (N_23342,N_22455,N_21205);
and U23343 (N_23343,N_21297,N_22242);
nor U23344 (N_23344,N_20668,N_21263);
nor U23345 (N_23345,N_22039,N_22017);
or U23346 (N_23346,N_22450,N_21475);
nand U23347 (N_23347,N_22208,N_20970);
xor U23348 (N_23348,N_21028,N_22330);
or U23349 (N_23349,N_21676,N_22388);
or U23350 (N_23350,N_21487,N_20514);
and U23351 (N_23351,N_21242,N_20510);
and U23352 (N_23352,N_20758,N_21320);
or U23353 (N_23353,N_20547,N_21849);
and U23354 (N_23354,N_20090,N_21559);
nand U23355 (N_23355,N_21250,N_20272);
nor U23356 (N_23356,N_21965,N_20236);
nand U23357 (N_23357,N_22460,N_22092);
and U23358 (N_23358,N_20812,N_20255);
or U23359 (N_23359,N_20664,N_22020);
or U23360 (N_23360,N_22037,N_21355);
and U23361 (N_23361,N_21766,N_20269);
xnor U23362 (N_23362,N_20775,N_21182);
nand U23363 (N_23363,N_21183,N_20674);
xnor U23364 (N_23364,N_21578,N_22078);
or U23365 (N_23365,N_22293,N_20745);
and U23366 (N_23366,N_22305,N_20914);
xnor U23367 (N_23367,N_20258,N_20459);
nand U23368 (N_23368,N_22157,N_21405);
or U23369 (N_23369,N_22069,N_20627);
or U23370 (N_23370,N_20218,N_21832);
nand U23371 (N_23371,N_21098,N_21794);
xor U23372 (N_23372,N_20896,N_22366);
nand U23373 (N_23373,N_21438,N_20130);
nand U23374 (N_23374,N_20688,N_20899);
nor U23375 (N_23375,N_20332,N_22004);
nand U23376 (N_23376,N_22461,N_20537);
nor U23377 (N_23377,N_20950,N_20168);
and U23378 (N_23378,N_20447,N_21609);
and U23379 (N_23379,N_22261,N_20678);
xor U23380 (N_23380,N_21172,N_20658);
and U23381 (N_23381,N_21833,N_21526);
xor U23382 (N_23382,N_21791,N_21523);
nor U23383 (N_23383,N_21051,N_21003);
or U23384 (N_23384,N_20587,N_22363);
nand U23385 (N_23385,N_21022,N_20543);
or U23386 (N_23386,N_20434,N_20167);
and U23387 (N_23387,N_20251,N_21913);
xnor U23388 (N_23388,N_22335,N_20763);
nand U23389 (N_23389,N_21895,N_20074);
nor U23390 (N_23390,N_21789,N_20017);
or U23391 (N_23391,N_21769,N_21893);
nand U23392 (N_23392,N_21921,N_20475);
and U23393 (N_23393,N_21981,N_21469);
nand U23394 (N_23394,N_21613,N_22104);
nor U23395 (N_23395,N_20349,N_21625);
or U23396 (N_23396,N_21700,N_20945);
nand U23397 (N_23397,N_22072,N_21818);
nand U23398 (N_23398,N_22144,N_21930);
nand U23399 (N_23399,N_21166,N_21653);
nand U23400 (N_23400,N_20617,N_22353);
nand U23401 (N_23401,N_21600,N_21151);
nand U23402 (N_23402,N_20223,N_22124);
and U23403 (N_23403,N_21666,N_22156);
nor U23404 (N_23404,N_20956,N_22453);
nand U23405 (N_23405,N_22301,N_20263);
nor U23406 (N_23406,N_20590,N_20416);
or U23407 (N_23407,N_20139,N_20979);
or U23408 (N_23408,N_21743,N_21223);
xor U23409 (N_23409,N_21148,N_20486);
nand U23410 (N_23410,N_22180,N_21539);
and U23411 (N_23411,N_21370,N_22089);
nor U23412 (N_23412,N_21500,N_21139);
nand U23413 (N_23413,N_21644,N_21453);
nand U23414 (N_23414,N_20331,N_22145);
nor U23415 (N_23415,N_21367,N_20354);
nand U23416 (N_23416,N_22281,N_21310);
or U23417 (N_23417,N_20200,N_20652);
xnor U23418 (N_23418,N_22044,N_20037);
or U23419 (N_23419,N_21771,N_21380);
nand U23420 (N_23420,N_20518,N_20054);
xnor U23421 (N_23421,N_20884,N_22028);
nor U23422 (N_23422,N_20304,N_20933);
nand U23423 (N_23423,N_20141,N_21224);
xnor U23424 (N_23424,N_20075,N_21927);
nor U23425 (N_23425,N_20158,N_21396);
nor U23426 (N_23426,N_21099,N_20729);
nand U23427 (N_23427,N_22246,N_20520);
nand U23428 (N_23428,N_21718,N_20177);
nor U23429 (N_23429,N_21831,N_22120);
or U23430 (N_23430,N_21945,N_20960);
or U23431 (N_23431,N_20508,N_21702);
nor U23432 (N_23432,N_20573,N_20276);
or U23433 (N_23433,N_20782,N_21066);
nor U23434 (N_23434,N_21292,N_20841);
and U23435 (N_23435,N_20816,N_21782);
xor U23436 (N_23436,N_22085,N_21212);
or U23437 (N_23437,N_21023,N_21271);
nor U23438 (N_23438,N_21863,N_20008);
or U23439 (N_23439,N_21514,N_22240);
or U23440 (N_23440,N_21560,N_21248);
xnor U23441 (N_23441,N_20524,N_21896);
nand U23442 (N_23442,N_22111,N_20178);
nor U23443 (N_23443,N_20094,N_20010);
xor U23444 (N_23444,N_20659,N_21626);
nand U23445 (N_23445,N_20953,N_21041);
nor U23446 (N_23446,N_21118,N_22352);
nor U23447 (N_23447,N_21247,N_22304);
and U23448 (N_23448,N_22241,N_20592);
or U23449 (N_23449,N_22129,N_22079);
nor U23450 (N_23450,N_21533,N_20249);
or U23451 (N_23451,N_22480,N_22324);
or U23452 (N_23452,N_20202,N_20124);
nor U23453 (N_23453,N_22357,N_20786);
and U23454 (N_23454,N_20624,N_21988);
nor U23455 (N_23455,N_20352,N_20928);
or U23456 (N_23456,N_20600,N_20616);
xnor U23457 (N_23457,N_20685,N_21461);
nor U23458 (N_23458,N_22416,N_20468);
nor U23459 (N_23459,N_20368,N_21819);
nand U23460 (N_23460,N_20651,N_21805);
xor U23461 (N_23461,N_20724,N_22382);
xor U23462 (N_23462,N_20646,N_21156);
nand U23463 (N_23463,N_20738,N_20234);
and U23464 (N_23464,N_21752,N_22315);
nor U23465 (N_23465,N_21999,N_20827);
xor U23466 (N_23466,N_21828,N_21841);
and U23467 (N_23467,N_20129,N_22108);
xnor U23468 (N_23468,N_20855,N_20681);
nand U23469 (N_23469,N_22282,N_20162);
nand U23470 (N_23470,N_20137,N_20848);
nor U23471 (N_23471,N_22055,N_20371);
xnor U23472 (N_23472,N_21332,N_21885);
nand U23473 (N_23473,N_20161,N_22473);
nor U23474 (N_23474,N_21474,N_20790);
nand U23475 (N_23475,N_21064,N_21013);
or U23476 (N_23476,N_20324,N_20965);
nand U23477 (N_23477,N_20542,N_20104);
nor U23478 (N_23478,N_21065,N_20494);
or U23479 (N_23479,N_22001,N_20791);
and U23480 (N_23480,N_21154,N_21632);
or U23481 (N_23481,N_20711,N_20972);
nor U23482 (N_23482,N_22407,N_20435);
and U23483 (N_23483,N_20301,N_21203);
xor U23484 (N_23484,N_21497,N_22320);
nor U23485 (N_23485,N_21824,N_21496);
or U23486 (N_23486,N_21739,N_22105);
nand U23487 (N_23487,N_20021,N_21286);
and U23488 (N_23488,N_20099,N_22176);
and U23489 (N_23489,N_21788,N_22034);
nand U23490 (N_23490,N_22325,N_20649);
or U23491 (N_23491,N_21196,N_21413);
nor U23492 (N_23492,N_20203,N_22303);
and U23493 (N_23493,N_21532,N_20955);
nand U23494 (N_23494,N_22066,N_20204);
nand U23495 (N_23495,N_22254,N_22381);
nor U23496 (N_23496,N_20163,N_20226);
nor U23497 (N_23497,N_21291,N_21859);
nand U23498 (N_23498,N_22003,N_21020);
or U23499 (N_23499,N_21953,N_21387);
xnor U23500 (N_23500,N_21364,N_21039);
and U23501 (N_23501,N_20713,N_21329);
xor U23502 (N_23502,N_20280,N_21853);
or U23503 (N_23503,N_21485,N_20844);
or U23504 (N_23504,N_21939,N_20925);
nor U23505 (N_23505,N_22226,N_21524);
xor U23506 (N_23506,N_20927,N_20849);
or U23507 (N_23507,N_20373,N_22082);
and U23508 (N_23508,N_21058,N_20460);
or U23509 (N_23509,N_21232,N_21406);
nand U23510 (N_23510,N_21455,N_21811);
xnor U23511 (N_23511,N_21802,N_21382);
nor U23512 (N_23512,N_20360,N_21740);
and U23513 (N_23513,N_21357,N_21477);
and U23514 (N_23514,N_20792,N_20011);
and U23515 (N_23515,N_20546,N_20977);
or U23516 (N_23516,N_20575,N_21730);
nand U23517 (N_23517,N_22051,N_21315);
xnor U23518 (N_23518,N_21648,N_20806);
nor U23519 (N_23519,N_21962,N_20836);
nand U23520 (N_23520,N_20491,N_21199);
nor U23521 (N_23521,N_20418,N_20939);
nor U23522 (N_23522,N_20595,N_20419);
xnor U23523 (N_23523,N_21307,N_21689);
nand U23524 (N_23524,N_20655,N_22275);
or U23525 (N_23525,N_22029,N_20550);
or U23526 (N_23526,N_20085,N_20030);
nor U23527 (N_23527,N_21386,N_21325);
nand U23528 (N_23528,N_21587,N_20310);
or U23529 (N_23529,N_22248,N_22074);
xor U23530 (N_23530,N_22009,N_21996);
or U23531 (N_23531,N_21047,N_21511);
or U23532 (N_23532,N_20444,N_21435);
nand U23533 (N_23533,N_22146,N_20743);
xnor U23534 (N_23534,N_21573,N_20677);
nor U23535 (N_23535,N_21431,N_20847);
or U23536 (N_23536,N_21267,N_22099);
nand U23537 (N_23537,N_22220,N_22384);
nor U23538 (N_23538,N_21952,N_22496);
xor U23539 (N_23539,N_20561,N_20643);
nand U23540 (N_23540,N_20608,N_20636);
and U23541 (N_23541,N_20442,N_22189);
nor U23542 (N_23542,N_21317,N_22356);
and U23543 (N_23543,N_20165,N_20629);
xor U23544 (N_23544,N_21544,N_21710);
nor U23545 (N_23545,N_20523,N_21926);
or U23546 (N_23546,N_20009,N_20302);
nor U23547 (N_23547,N_20377,N_21308);
nand U23548 (N_23548,N_20512,N_21534);
nand U23549 (N_23549,N_20185,N_20240);
or U23550 (N_23550,N_21350,N_20495);
nand U23551 (N_23551,N_21846,N_20044);
nand U23552 (N_23552,N_20108,N_22222);
nor U23553 (N_23553,N_20875,N_21448);
nor U23554 (N_23554,N_20871,N_21093);
or U23555 (N_23555,N_20066,N_21237);
or U23556 (N_23556,N_22286,N_20436);
nor U23557 (N_23557,N_21218,N_21591);
or U23558 (N_23558,N_22256,N_21650);
nand U23559 (N_23559,N_21720,N_20767);
and U23560 (N_23560,N_21351,N_22200);
or U23561 (N_23561,N_20303,N_20206);
or U23562 (N_23562,N_22083,N_20511);
nor U23563 (N_23563,N_21336,N_20503);
nor U23564 (N_23564,N_21008,N_22161);
nand U23565 (N_23565,N_21869,N_22345);
or U23566 (N_23566,N_20698,N_20570);
nor U23567 (N_23567,N_21675,N_21037);
nor U23568 (N_23568,N_20453,N_21001);
nor U23569 (N_23569,N_21555,N_21073);
or U23570 (N_23570,N_20182,N_20969);
or U23571 (N_23571,N_22169,N_22396);
nor U23572 (N_23572,N_22172,N_21348);
and U23573 (N_23573,N_20715,N_20919);
xnor U23574 (N_23574,N_21606,N_21163);
nor U23575 (N_23575,N_22196,N_21727);
nor U23576 (N_23576,N_21595,N_20995);
xnor U23577 (N_23577,N_20864,N_22369);
xnor U23578 (N_23578,N_20815,N_20015);
or U23579 (N_23579,N_22163,N_22005);
nor U23580 (N_23580,N_21715,N_22389);
or U23581 (N_23581,N_20766,N_20656);
or U23582 (N_23582,N_21334,N_21445);
or U23583 (N_23583,N_22214,N_20336);
nand U23584 (N_23584,N_21029,N_21120);
xor U23585 (N_23585,N_20619,N_20024);
nor U23586 (N_23586,N_21550,N_21985);
and U23587 (N_23587,N_21621,N_20545);
or U23588 (N_23588,N_22346,N_21227);
nor U23589 (N_23589,N_21879,N_20454);
nor U23590 (N_23590,N_22071,N_20472);
xor U23591 (N_23591,N_22285,N_20886);
xnor U23592 (N_23592,N_20325,N_20803);
or U23593 (N_23593,N_21030,N_21272);
and U23594 (N_23594,N_20811,N_21407);
xor U23595 (N_23595,N_22061,N_22418);
nor U23596 (N_23596,N_22024,N_21296);
nor U23597 (N_23597,N_21974,N_21397);
nor U23598 (N_23598,N_20700,N_20650);
xor U23599 (N_23599,N_21978,N_21754);
nand U23600 (N_23600,N_20344,N_22247);
xor U23601 (N_23601,N_20298,N_22446);
nor U23602 (N_23602,N_20564,N_22372);
nor U23603 (N_23603,N_21696,N_22339);
and U23604 (N_23604,N_21711,N_21995);
or U23605 (N_23605,N_21619,N_20208);
nor U23606 (N_23606,N_21627,N_21531);
nor U23607 (N_23607,N_20370,N_20784);
and U23608 (N_23608,N_20118,N_21356);
xor U23609 (N_23609,N_21936,N_21069);
nor U23610 (N_23610,N_20353,N_21211);
and U23611 (N_23611,N_22119,N_21652);
xor U23612 (N_23612,N_20716,N_21422);
or U23613 (N_23613,N_21441,N_20385);
or U23614 (N_23614,N_21756,N_20098);
and U23615 (N_23615,N_20971,N_20430);
nand U23616 (N_23616,N_21825,N_20300);
or U23617 (N_23617,N_20379,N_21376);
and U23618 (N_23618,N_21331,N_21042);
xnor U23619 (N_23619,N_22289,N_21768);
xnor U23620 (N_23620,N_21111,N_22276);
and U23621 (N_23621,N_20069,N_22400);
xor U23622 (N_23622,N_20189,N_20918);
and U23623 (N_23623,N_21233,N_20593);
nand U23624 (N_23624,N_22233,N_22296);
xnor U23625 (N_23625,N_20866,N_20376);
nand U23626 (N_23626,N_22101,N_21861);
or U23627 (N_23627,N_21714,N_20594);
xnor U23628 (N_23628,N_22297,N_21731);
nor U23629 (N_23629,N_22421,N_20257);
nand U23630 (N_23630,N_21830,N_22209);
and U23631 (N_23631,N_22022,N_21362);
nor U23632 (N_23632,N_20912,N_20487);
nor U23633 (N_23633,N_20312,N_21488);
and U23634 (N_23634,N_20780,N_21660);
and U23635 (N_23635,N_22154,N_21512);
nand U23636 (N_23636,N_20116,N_20714);
and U23637 (N_23637,N_20490,N_22234);
or U23638 (N_23638,N_20789,N_20291);
and U23639 (N_23639,N_21130,N_22016);
nor U23640 (N_23640,N_22006,N_20776);
or U23641 (N_23641,N_20857,N_20558);
xnor U23642 (N_23642,N_20748,N_20718);
nand U23643 (N_23643,N_20296,N_20604);
nor U23644 (N_23644,N_21716,N_22118);
nand U23645 (N_23645,N_21024,N_20388);
nand U23646 (N_23646,N_20133,N_22141);
or U23647 (N_23647,N_22195,N_21917);
nor U23648 (N_23648,N_22042,N_22318);
nor U23649 (N_23649,N_22258,N_21340);
nor U23650 (N_23650,N_22213,N_21403);
and U23651 (N_23651,N_21206,N_20427);
nor U23652 (N_23652,N_21409,N_22443);
nor U23653 (N_23653,N_22437,N_21281);
nor U23654 (N_23654,N_21000,N_20404);
and U23655 (N_23655,N_20207,N_20615);
nor U23656 (N_23656,N_21612,N_22100);
nand U23657 (N_23657,N_21460,N_21471);
nor U23658 (N_23658,N_20179,N_22288);
or U23659 (N_23659,N_20930,N_21602);
xor U23660 (N_23660,N_22217,N_21798);
nor U23661 (N_23661,N_21254,N_21671);
nand U23662 (N_23662,N_21439,N_20820);
xnor U23663 (N_23663,N_20513,N_20012);
or U23664 (N_23664,N_21388,N_21216);
xnor U23665 (N_23665,N_21009,N_20926);
xnor U23666 (N_23666,N_21425,N_20040);
or U23667 (N_23667,N_21997,N_21767);
and U23668 (N_23668,N_22210,N_22436);
nand U23669 (N_23669,N_22306,N_22251);
xor U23670 (N_23670,N_20676,N_21722);
nand U23671 (N_23671,N_20086,N_21269);
nand U23672 (N_23672,N_20052,N_21701);
nor U23673 (N_23673,N_20193,N_21278);
nand U23674 (N_23674,N_20001,N_20852);
nor U23675 (N_23675,N_20211,N_21629);
and U23676 (N_23676,N_21229,N_20311);
nor U23677 (N_23677,N_21132,N_20210);
and U23678 (N_23678,N_20557,N_21265);
or U23679 (N_23679,N_22412,N_20973);
nand U23680 (N_23680,N_21384,N_21688);
or U23681 (N_23681,N_21616,N_20215);
nor U23682 (N_23682,N_22481,N_20413);
or U23683 (N_23683,N_20582,N_20369);
xnor U23684 (N_23684,N_21499,N_21994);
nand U23685 (N_23685,N_22250,N_21980);
and U23686 (N_23686,N_20264,N_21854);
nor U23687 (N_23687,N_20450,N_22459);
xnor U23688 (N_23688,N_20797,N_22160);
nand U23689 (N_23689,N_21002,N_22191);
or U23690 (N_23690,N_21164,N_22202);
or U23691 (N_23691,N_20461,N_20170);
or U23692 (N_23692,N_20233,N_21395);
xor U23693 (N_23693,N_21662,N_22080);
nand U23694 (N_23694,N_22206,N_21476);
or U23695 (N_23695,N_21874,N_22059);
nor U23696 (N_23696,N_20485,N_21239);
nor U23697 (N_23697,N_21287,N_21081);
nand U23698 (N_23698,N_22113,N_21059);
or U23699 (N_23699,N_21623,N_21007);
or U23700 (N_23700,N_20361,N_21764);
nand U23701 (N_23701,N_21021,N_20068);
nand U23702 (N_23702,N_21143,N_20787);
or U23703 (N_23703,N_20329,N_21337);
xor U23704 (N_23704,N_22307,N_20432);
xor U23705 (N_23705,N_21670,N_20769);
nand U23706 (N_23706,N_20433,N_20288);
nand U23707 (N_23707,N_21378,N_20229);
xor U23708 (N_23708,N_20146,N_20295);
nand U23709 (N_23709,N_22179,N_20819);
nor U23710 (N_23710,N_21050,N_20227);
or U23711 (N_23711,N_21871,N_21483);
nand U23712 (N_23712,N_21392,N_20917);
and U23713 (N_23713,N_21373,N_21449);
and U23714 (N_23714,N_21755,N_22238);
xor U23715 (N_23715,N_20277,N_22158);
nor U23716 (N_23716,N_21159,N_20580);
xor U23717 (N_23717,N_20375,N_21204);
nand U23718 (N_23718,N_21400,N_20975);
or U23719 (N_23719,N_20374,N_21972);
nor U23720 (N_23720,N_22375,N_21905);
nor U23721 (N_23721,N_20807,N_21188);
and U23722 (N_23722,N_21282,N_21630);
and U23723 (N_23723,N_20521,N_22170);
nand U23724 (N_23724,N_21076,N_20562);
xnor U23725 (N_23725,N_20725,N_21883);
nor U23726 (N_23726,N_21596,N_21724);
xnor U23727 (N_23727,N_22474,N_22262);
nor U23728 (N_23728,N_22402,N_21947);
or U23729 (N_23729,N_21135,N_20242);
or U23730 (N_23730,N_20905,N_22292);
and U23731 (N_23731,N_22280,N_20741);
xor U23732 (N_23732,N_20409,N_21900);
xnor U23733 (N_23733,N_22314,N_21812);
nor U23734 (N_23734,N_22040,N_21552);
or U23735 (N_23735,N_21219,N_22462);
nand U23736 (N_23736,N_22027,N_21070);
nor U23737 (N_23737,N_22090,N_21773);
nand U23738 (N_23738,N_20750,N_21875);
nor U23739 (N_23739,N_22406,N_21669);
xor U23740 (N_23740,N_20243,N_22340);
xnor U23741 (N_23741,N_21891,N_22012);
and U23742 (N_23742,N_20122,N_21498);
nor U23743 (N_23743,N_22062,N_21122);
and U23744 (N_23744,N_20531,N_22342);
and U23745 (N_23745,N_20245,N_20974);
xor U23746 (N_23746,N_21918,N_21646);
or U23747 (N_23747,N_21783,N_21140);
nor U23748 (N_23748,N_22477,N_20499);
and U23749 (N_23749,N_20176,N_20731);
nand U23750 (N_23750,N_22168,N_20398);
or U23751 (N_23751,N_22480,N_21575);
xnor U23752 (N_23752,N_21094,N_21283);
nor U23753 (N_23753,N_20466,N_22348);
and U23754 (N_23754,N_21371,N_22178);
xnor U23755 (N_23755,N_22291,N_21783);
nor U23756 (N_23756,N_20863,N_21468);
and U23757 (N_23757,N_22169,N_21581);
or U23758 (N_23758,N_20786,N_21394);
xor U23759 (N_23759,N_20455,N_20196);
or U23760 (N_23760,N_22166,N_22317);
nor U23761 (N_23761,N_21953,N_20443);
xnor U23762 (N_23762,N_21259,N_21422);
and U23763 (N_23763,N_21991,N_22361);
or U23764 (N_23764,N_20561,N_21387);
xnor U23765 (N_23765,N_21181,N_20230);
xor U23766 (N_23766,N_21044,N_21744);
and U23767 (N_23767,N_20304,N_22245);
or U23768 (N_23768,N_21172,N_20638);
and U23769 (N_23769,N_21132,N_20288);
or U23770 (N_23770,N_21358,N_22203);
nor U23771 (N_23771,N_21369,N_22150);
nor U23772 (N_23772,N_21566,N_20582);
and U23773 (N_23773,N_22308,N_21891);
nor U23774 (N_23774,N_20177,N_22326);
xor U23775 (N_23775,N_21248,N_21087);
nor U23776 (N_23776,N_20303,N_20562);
xor U23777 (N_23777,N_20696,N_22078);
nand U23778 (N_23778,N_20096,N_20637);
and U23779 (N_23779,N_20082,N_21324);
nand U23780 (N_23780,N_20589,N_20389);
nor U23781 (N_23781,N_21882,N_22334);
xnor U23782 (N_23782,N_20040,N_21225);
nand U23783 (N_23783,N_21543,N_21844);
nor U23784 (N_23784,N_21218,N_20805);
xnor U23785 (N_23785,N_20280,N_20101);
xnor U23786 (N_23786,N_20443,N_21276);
or U23787 (N_23787,N_21146,N_21452);
xor U23788 (N_23788,N_22129,N_20255);
xor U23789 (N_23789,N_20046,N_21049);
nand U23790 (N_23790,N_20581,N_21716);
or U23791 (N_23791,N_21160,N_21233);
xor U23792 (N_23792,N_20086,N_21956);
xor U23793 (N_23793,N_20655,N_22381);
nand U23794 (N_23794,N_20848,N_20326);
nor U23795 (N_23795,N_20744,N_20520);
nor U23796 (N_23796,N_20587,N_21463);
xnor U23797 (N_23797,N_22450,N_22329);
or U23798 (N_23798,N_20616,N_20707);
nand U23799 (N_23799,N_22172,N_22217);
and U23800 (N_23800,N_20447,N_20186);
nor U23801 (N_23801,N_21035,N_21062);
xor U23802 (N_23802,N_21409,N_21429);
nor U23803 (N_23803,N_21990,N_21213);
and U23804 (N_23804,N_21420,N_21701);
nor U23805 (N_23805,N_20029,N_21416);
or U23806 (N_23806,N_20624,N_20449);
nand U23807 (N_23807,N_22353,N_20087);
xnor U23808 (N_23808,N_21503,N_20658);
nor U23809 (N_23809,N_21075,N_22221);
and U23810 (N_23810,N_20011,N_21315);
xor U23811 (N_23811,N_22487,N_21086);
nand U23812 (N_23812,N_22056,N_21180);
and U23813 (N_23813,N_20448,N_21900);
or U23814 (N_23814,N_22129,N_20150);
or U23815 (N_23815,N_21925,N_20630);
nor U23816 (N_23816,N_22192,N_20711);
and U23817 (N_23817,N_21021,N_21242);
nor U23818 (N_23818,N_21567,N_22273);
nand U23819 (N_23819,N_21635,N_20559);
and U23820 (N_23820,N_21358,N_22014);
nand U23821 (N_23821,N_20484,N_21521);
and U23822 (N_23822,N_20455,N_21085);
nor U23823 (N_23823,N_20858,N_21580);
xnor U23824 (N_23824,N_20619,N_20635);
or U23825 (N_23825,N_22262,N_21735);
nor U23826 (N_23826,N_22249,N_21897);
or U23827 (N_23827,N_21488,N_20769);
xor U23828 (N_23828,N_20473,N_21514);
nor U23829 (N_23829,N_20029,N_21191);
and U23830 (N_23830,N_21089,N_20900);
or U23831 (N_23831,N_20339,N_21041);
and U23832 (N_23832,N_21119,N_20957);
xor U23833 (N_23833,N_20275,N_20486);
nor U23834 (N_23834,N_21219,N_22233);
or U23835 (N_23835,N_21200,N_22251);
nand U23836 (N_23836,N_20671,N_20454);
or U23837 (N_23837,N_22178,N_20638);
xnor U23838 (N_23838,N_21213,N_20266);
or U23839 (N_23839,N_20518,N_22201);
xor U23840 (N_23840,N_20618,N_20255);
and U23841 (N_23841,N_20264,N_21563);
xnor U23842 (N_23842,N_22127,N_21610);
nand U23843 (N_23843,N_20621,N_21709);
xor U23844 (N_23844,N_22491,N_20154);
nor U23845 (N_23845,N_20633,N_21787);
nor U23846 (N_23846,N_20782,N_21906);
or U23847 (N_23847,N_21253,N_21129);
and U23848 (N_23848,N_20424,N_20763);
xor U23849 (N_23849,N_20590,N_21741);
xnor U23850 (N_23850,N_22194,N_20468);
nand U23851 (N_23851,N_21107,N_22036);
xor U23852 (N_23852,N_20737,N_21468);
or U23853 (N_23853,N_21118,N_20510);
or U23854 (N_23854,N_22342,N_21154);
nor U23855 (N_23855,N_20929,N_21123);
nor U23856 (N_23856,N_22206,N_20407);
and U23857 (N_23857,N_20553,N_20754);
nand U23858 (N_23858,N_20252,N_21140);
xor U23859 (N_23859,N_21516,N_20676);
nor U23860 (N_23860,N_20744,N_21510);
and U23861 (N_23861,N_21152,N_20706);
xor U23862 (N_23862,N_21487,N_20627);
or U23863 (N_23863,N_20646,N_20805);
xnor U23864 (N_23864,N_21260,N_20437);
nor U23865 (N_23865,N_22437,N_22278);
xnor U23866 (N_23866,N_22422,N_21001);
xnor U23867 (N_23867,N_20518,N_21279);
and U23868 (N_23868,N_21941,N_22396);
xor U23869 (N_23869,N_21357,N_21368);
nand U23870 (N_23870,N_20879,N_21237);
nand U23871 (N_23871,N_21528,N_20909);
and U23872 (N_23872,N_22488,N_20277);
or U23873 (N_23873,N_22415,N_20006);
nand U23874 (N_23874,N_22086,N_20817);
xor U23875 (N_23875,N_21566,N_22066);
xor U23876 (N_23876,N_21289,N_21244);
xor U23877 (N_23877,N_20750,N_21670);
xor U23878 (N_23878,N_22217,N_21989);
or U23879 (N_23879,N_20711,N_21490);
and U23880 (N_23880,N_21400,N_21551);
and U23881 (N_23881,N_21524,N_21903);
xnor U23882 (N_23882,N_20047,N_22207);
and U23883 (N_23883,N_21029,N_20889);
and U23884 (N_23884,N_21019,N_20190);
xor U23885 (N_23885,N_21028,N_20758);
nand U23886 (N_23886,N_21389,N_20251);
nand U23887 (N_23887,N_20599,N_21392);
and U23888 (N_23888,N_21149,N_22390);
nand U23889 (N_23889,N_20733,N_20112);
nand U23890 (N_23890,N_21724,N_20190);
and U23891 (N_23891,N_20163,N_21728);
nor U23892 (N_23892,N_21673,N_20719);
nand U23893 (N_23893,N_21882,N_20823);
and U23894 (N_23894,N_20050,N_22126);
nor U23895 (N_23895,N_20199,N_21786);
nand U23896 (N_23896,N_22332,N_22229);
nand U23897 (N_23897,N_21762,N_20055);
and U23898 (N_23898,N_21431,N_20668);
and U23899 (N_23899,N_20817,N_20291);
nor U23900 (N_23900,N_22464,N_22255);
nor U23901 (N_23901,N_22113,N_22380);
or U23902 (N_23902,N_20381,N_21140);
xor U23903 (N_23903,N_21266,N_22293);
nor U23904 (N_23904,N_20374,N_20476);
nor U23905 (N_23905,N_21119,N_21081);
or U23906 (N_23906,N_20281,N_21082);
or U23907 (N_23907,N_21234,N_21553);
xor U23908 (N_23908,N_20491,N_22477);
and U23909 (N_23909,N_21204,N_21863);
or U23910 (N_23910,N_20541,N_20187);
or U23911 (N_23911,N_21966,N_20219);
xnor U23912 (N_23912,N_20186,N_20689);
nand U23913 (N_23913,N_22129,N_20764);
or U23914 (N_23914,N_21702,N_20349);
nand U23915 (N_23915,N_21262,N_20617);
xnor U23916 (N_23916,N_20350,N_20648);
nor U23917 (N_23917,N_21391,N_20479);
nor U23918 (N_23918,N_21358,N_21457);
nor U23919 (N_23919,N_20265,N_21782);
or U23920 (N_23920,N_20264,N_20125);
nor U23921 (N_23921,N_22333,N_22176);
nor U23922 (N_23922,N_20737,N_21870);
and U23923 (N_23923,N_21035,N_22127);
and U23924 (N_23924,N_21632,N_20947);
nor U23925 (N_23925,N_21606,N_20462);
nand U23926 (N_23926,N_20798,N_20347);
nand U23927 (N_23927,N_20290,N_20684);
or U23928 (N_23928,N_20682,N_20416);
and U23929 (N_23929,N_21785,N_22346);
nand U23930 (N_23930,N_21790,N_21472);
or U23931 (N_23931,N_21751,N_21479);
nand U23932 (N_23932,N_22472,N_20630);
and U23933 (N_23933,N_22076,N_21852);
nor U23934 (N_23934,N_22301,N_20931);
and U23935 (N_23935,N_21908,N_21512);
and U23936 (N_23936,N_20069,N_21225);
or U23937 (N_23937,N_22292,N_21051);
nand U23938 (N_23938,N_21859,N_22385);
and U23939 (N_23939,N_20183,N_20804);
nand U23940 (N_23940,N_20337,N_20948);
or U23941 (N_23941,N_21983,N_22344);
or U23942 (N_23942,N_21490,N_20861);
nor U23943 (N_23943,N_22167,N_21901);
and U23944 (N_23944,N_22263,N_21594);
xor U23945 (N_23945,N_21783,N_21465);
or U23946 (N_23946,N_21185,N_21830);
nand U23947 (N_23947,N_20007,N_22363);
or U23948 (N_23948,N_21898,N_21350);
or U23949 (N_23949,N_20946,N_20358);
or U23950 (N_23950,N_20148,N_21962);
nor U23951 (N_23951,N_20679,N_22080);
nand U23952 (N_23952,N_22380,N_20874);
nor U23953 (N_23953,N_22065,N_20178);
and U23954 (N_23954,N_22495,N_20908);
and U23955 (N_23955,N_20838,N_20138);
xor U23956 (N_23956,N_22213,N_20425);
and U23957 (N_23957,N_20768,N_20586);
xnor U23958 (N_23958,N_20259,N_20114);
and U23959 (N_23959,N_20362,N_20998);
xnor U23960 (N_23960,N_21965,N_20181);
xnor U23961 (N_23961,N_20051,N_21023);
or U23962 (N_23962,N_21571,N_20992);
nor U23963 (N_23963,N_21609,N_20728);
nand U23964 (N_23964,N_21343,N_22248);
and U23965 (N_23965,N_22332,N_20759);
or U23966 (N_23966,N_22490,N_21659);
nand U23967 (N_23967,N_20422,N_22040);
nor U23968 (N_23968,N_21533,N_21191);
nor U23969 (N_23969,N_21326,N_21484);
and U23970 (N_23970,N_22044,N_20974);
and U23971 (N_23971,N_20079,N_21628);
nor U23972 (N_23972,N_22357,N_20401);
nor U23973 (N_23973,N_20960,N_21498);
xnor U23974 (N_23974,N_22496,N_21735);
xor U23975 (N_23975,N_20168,N_21796);
or U23976 (N_23976,N_22305,N_21733);
xnor U23977 (N_23977,N_20439,N_20697);
xnor U23978 (N_23978,N_20852,N_20944);
nand U23979 (N_23979,N_20989,N_21276);
and U23980 (N_23980,N_22177,N_21792);
or U23981 (N_23981,N_21267,N_22126);
nor U23982 (N_23982,N_21218,N_21354);
nor U23983 (N_23983,N_22218,N_21013);
or U23984 (N_23984,N_20052,N_20966);
and U23985 (N_23985,N_22460,N_22061);
and U23986 (N_23986,N_21416,N_21482);
nand U23987 (N_23987,N_21499,N_20239);
nand U23988 (N_23988,N_22233,N_21687);
nor U23989 (N_23989,N_21364,N_20169);
or U23990 (N_23990,N_21530,N_21381);
nor U23991 (N_23991,N_22057,N_20021);
xor U23992 (N_23992,N_20015,N_22488);
and U23993 (N_23993,N_20922,N_21252);
nor U23994 (N_23994,N_21621,N_22475);
nor U23995 (N_23995,N_22121,N_21409);
nand U23996 (N_23996,N_22196,N_21897);
and U23997 (N_23997,N_21199,N_21963);
xor U23998 (N_23998,N_20500,N_21301);
or U23999 (N_23999,N_21341,N_20566);
and U24000 (N_24000,N_21297,N_22483);
xnor U24001 (N_24001,N_20815,N_21492);
nor U24002 (N_24002,N_21235,N_21918);
and U24003 (N_24003,N_20233,N_21942);
or U24004 (N_24004,N_22269,N_20005);
nand U24005 (N_24005,N_21636,N_22497);
nor U24006 (N_24006,N_21776,N_22023);
nand U24007 (N_24007,N_21289,N_21456);
or U24008 (N_24008,N_22479,N_20861);
or U24009 (N_24009,N_21018,N_20015);
xor U24010 (N_24010,N_20776,N_20657);
or U24011 (N_24011,N_20136,N_21044);
nand U24012 (N_24012,N_20070,N_20469);
nand U24013 (N_24013,N_20513,N_20849);
nand U24014 (N_24014,N_21728,N_20475);
or U24015 (N_24015,N_21545,N_20130);
xnor U24016 (N_24016,N_21968,N_20410);
xor U24017 (N_24017,N_22474,N_21929);
and U24018 (N_24018,N_21622,N_20587);
nor U24019 (N_24019,N_20957,N_21956);
xnor U24020 (N_24020,N_21916,N_22452);
or U24021 (N_24021,N_20709,N_20249);
or U24022 (N_24022,N_20398,N_20970);
and U24023 (N_24023,N_21231,N_21395);
nor U24024 (N_24024,N_21519,N_22220);
and U24025 (N_24025,N_20069,N_21695);
nand U24026 (N_24026,N_20769,N_21904);
nand U24027 (N_24027,N_21901,N_21303);
xor U24028 (N_24028,N_21826,N_21895);
or U24029 (N_24029,N_20970,N_21059);
nor U24030 (N_24030,N_21067,N_20129);
xnor U24031 (N_24031,N_20617,N_20739);
xor U24032 (N_24032,N_20145,N_20103);
and U24033 (N_24033,N_22078,N_20491);
and U24034 (N_24034,N_20269,N_20503);
and U24035 (N_24035,N_21903,N_22119);
and U24036 (N_24036,N_21475,N_20415);
nor U24037 (N_24037,N_21465,N_21676);
xnor U24038 (N_24038,N_20838,N_20417);
or U24039 (N_24039,N_21635,N_22246);
or U24040 (N_24040,N_21354,N_21471);
nand U24041 (N_24041,N_22479,N_21226);
or U24042 (N_24042,N_22065,N_20026);
nor U24043 (N_24043,N_21666,N_21256);
or U24044 (N_24044,N_20240,N_21126);
nor U24045 (N_24045,N_21873,N_20186);
nand U24046 (N_24046,N_21101,N_20283);
nor U24047 (N_24047,N_21211,N_20645);
nor U24048 (N_24048,N_20643,N_20963);
nand U24049 (N_24049,N_21334,N_21238);
and U24050 (N_24050,N_22383,N_20457);
nand U24051 (N_24051,N_21103,N_21713);
xor U24052 (N_24052,N_22287,N_20193);
nand U24053 (N_24053,N_20374,N_21991);
and U24054 (N_24054,N_21146,N_21933);
and U24055 (N_24055,N_20516,N_21489);
and U24056 (N_24056,N_21088,N_20222);
nand U24057 (N_24057,N_20686,N_21813);
or U24058 (N_24058,N_20495,N_21259);
or U24059 (N_24059,N_21185,N_21763);
or U24060 (N_24060,N_21138,N_20817);
xnor U24061 (N_24061,N_20653,N_21850);
and U24062 (N_24062,N_22220,N_20105);
xnor U24063 (N_24063,N_20870,N_20066);
nand U24064 (N_24064,N_21436,N_21801);
nand U24065 (N_24065,N_21077,N_21400);
or U24066 (N_24066,N_20604,N_20645);
nor U24067 (N_24067,N_20679,N_20417);
and U24068 (N_24068,N_20334,N_21228);
and U24069 (N_24069,N_21974,N_20631);
nor U24070 (N_24070,N_20597,N_21328);
xnor U24071 (N_24071,N_20665,N_20670);
nand U24072 (N_24072,N_21516,N_20934);
nand U24073 (N_24073,N_20620,N_21338);
nand U24074 (N_24074,N_20801,N_22374);
nand U24075 (N_24075,N_21125,N_20698);
xnor U24076 (N_24076,N_21465,N_21018);
xnor U24077 (N_24077,N_21317,N_22210);
nand U24078 (N_24078,N_21767,N_20871);
or U24079 (N_24079,N_20515,N_22382);
nand U24080 (N_24080,N_22316,N_20720);
nor U24081 (N_24081,N_22431,N_22409);
nor U24082 (N_24082,N_22255,N_21357);
nor U24083 (N_24083,N_21407,N_22463);
nor U24084 (N_24084,N_20173,N_21679);
nand U24085 (N_24085,N_20538,N_22486);
and U24086 (N_24086,N_21103,N_21487);
nand U24087 (N_24087,N_22356,N_20622);
or U24088 (N_24088,N_21083,N_20042);
and U24089 (N_24089,N_20289,N_21181);
and U24090 (N_24090,N_20954,N_20896);
and U24091 (N_24091,N_20169,N_21901);
xor U24092 (N_24092,N_22237,N_20036);
and U24093 (N_24093,N_21936,N_21194);
or U24094 (N_24094,N_20595,N_22358);
nor U24095 (N_24095,N_20308,N_21695);
xnor U24096 (N_24096,N_20296,N_21510);
xnor U24097 (N_24097,N_20272,N_20739);
nor U24098 (N_24098,N_20209,N_20846);
nor U24099 (N_24099,N_21681,N_20303);
nor U24100 (N_24100,N_22328,N_22447);
nand U24101 (N_24101,N_20794,N_20999);
nor U24102 (N_24102,N_20933,N_22036);
nand U24103 (N_24103,N_20309,N_20056);
nand U24104 (N_24104,N_20564,N_21999);
nand U24105 (N_24105,N_21023,N_21549);
nor U24106 (N_24106,N_20187,N_20397);
or U24107 (N_24107,N_20919,N_22412);
xnor U24108 (N_24108,N_21104,N_20445);
nand U24109 (N_24109,N_20107,N_20482);
xnor U24110 (N_24110,N_21755,N_22073);
xnor U24111 (N_24111,N_22377,N_20549);
nor U24112 (N_24112,N_20015,N_20762);
and U24113 (N_24113,N_21150,N_21442);
xnor U24114 (N_24114,N_21867,N_20325);
nor U24115 (N_24115,N_20844,N_20826);
nand U24116 (N_24116,N_21670,N_22375);
or U24117 (N_24117,N_20670,N_20822);
and U24118 (N_24118,N_21013,N_21173);
nand U24119 (N_24119,N_22419,N_20065);
or U24120 (N_24120,N_21002,N_21997);
or U24121 (N_24121,N_21627,N_20202);
or U24122 (N_24122,N_20376,N_21889);
nand U24123 (N_24123,N_21197,N_20407);
or U24124 (N_24124,N_22004,N_21141);
xnor U24125 (N_24125,N_20389,N_21999);
and U24126 (N_24126,N_22246,N_22421);
xor U24127 (N_24127,N_22349,N_22197);
nand U24128 (N_24128,N_21566,N_21634);
nand U24129 (N_24129,N_22446,N_21970);
nor U24130 (N_24130,N_20071,N_21165);
and U24131 (N_24131,N_20465,N_21266);
nand U24132 (N_24132,N_22038,N_21878);
or U24133 (N_24133,N_20269,N_20555);
nor U24134 (N_24134,N_20761,N_21537);
xor U24135 (N_24135,N_21534,N_21107);
or U24136 (N_24136,N_21762,N_22440);
xnor U24137 (N_24137,N_20228,N_20971);
nand U24138 (N_24138,N_20438,N_20409);
nand U24139 (N_24139,N_20286,N_21052);
or U24140 (N_24140,N_20903,N_20583);
and U24141 (N_24141,N_20167,N_20710);
nand U24142 (N_24142,N_21814,N_22399);
or U24143 (N_24143,N_21166,N_20279);
or U24144 (N_24144,N_21126,N_21532);
nand U24145 (N_24145,N_20523,N_20680);
xnor U24146 (N_24146,N_22191,N_22192);
nand U24147 (N_24147,N_20918,N_20331);
nand U24148 (N_24148,N_20835,N_21823);
xnor U24149 (N_24149,N_20218,N_20830);
xnor U24150 (N_24150,N_20368,N_20631);
or U24151 (N_24151,N_22150,N_22198);
or U24152 (N_24152,N_20943,N_22405);
nand U24153 (N_24153,N_21602,N_21435);
xor U24154 (N_24154,N_21016,N_20940);
xnor U24155 (N_24155,N_20180,N_20242);
nor U24156 (N_24156,N_21592,N_20352);
nor U24157 (N_24157,N_20248,N_21913);
or U24158 (N_24158,N_21368,N_21801);
xnor U24159 (N_24159,N_21781,N_21883);
nor U24160 (N_24160,N_21643,N_21397);
nor U24161 (N_24161,N_20284,N_21988);
nand U24162 (N_24162,N_21425,N_22407);
and U24163 (N_24163,N_22379,N_20672);
nand U24164 (N_24164,N_20664,N_21141);
nor U24165 (N_24165,N_22214,N_21073);
or U24166 (N_24166,N_21212,N_20715);
nand U24167 (N_24167,N_21266,N_20415);
nor U24168 (N_24168,N_21276,N_20865);
and U24169 (N_24169,N_21169,N_21753);
and U24170 (N_24170,N_21349,N_21230);
xor U24171 (N_24171,N_21194,N_21074);
nand U24172 (N_24172,N_20593,N_20014);
nor U24173 (N_24173,N_20819,N_22039);
nor U24174 (N_24174,N_21681,N_21745);
nand U24175 (N_24175,N_21485,N_20375);
and U24176 (N_24176,N_20791,N_20519);
and U24177 (N_24177,N_20747,N_21148);
nand U24178 (N_24178,N_20094,N_21630);
or U24179 (N_24179,N_20082,N_20901);
nor U24180 (N_24180,N_22456,N_20475);
nor U24181 (N_24181,N_21770,N_20152);
or U24182 (N_24182,N_22114,N_21353);
nand U24183 (N_24183,N_20909,N_21548);
or U24184 (N_24184,N_20522,N_20654);
nand U24185 (N_24185,N_20716,N_21317);
or U24186 (N_24186,N_21756,N_21240);
or U24187 (N_24187,N_20082,N_21329);
xor U24188 (N_24188,N_21247,N_21950);
xnor U24189 (N_24189,N_20663,N_21616);
nand U24190 (N_24190,N_21641,N_22182);
or U24191 (N_24191,N_22188,N_20708);
nor U24192 (N_24192,N_20021,N_22310);
and U24193 (N_24193,N_20757,N_20029);
xor U24194 (N_24194,N_20728,N_21878);
nor U24195 (N_24195,N_20112,N_20869);
nor U24196 (N_24196,N_21356,N_20791);
nor U24197 (N_24197,N_21485,N_20084);
and U24198 (N_24198,N_20015,N_21338);
and U24199 (N_24199,N_20626,N_20794);
nor U24200 (N_24200,N_21632,N_22135);
or U24201 (N_24201,N_21982,N_22392);
or U24202 (N_24202,N_21371,N_22456);
nand U24203 (N_24203,N_21987,N_22482);
or U24204 (N_24204,N_21784,N_20803);
xnor U24205 (N_24205,N_21069,N_21616);
or U24206 (N_24206,N_22156,N_21502);
and U24207 (N_24207,N_20169,N_21875);
nand U24208 (N_24208,N_21920,N_22393);
nor U24209 (N_24209,N_22169,N_21463);
and U24210 (N_24210,N_20723,N_20520);
nand U24211 (N_24211,N_20529,N_21734);
or U24212 (N_24212,N_22167,N_20452);
or U24213 (N_24213,N_20994,N_20843);
and U24214 (N_24214,N_21485,N_20684);
nand U24215 (N_24215,N_20696,N_20602);
xor U24216 (N_24216,N_22229,N_22267);
nor U24217 (N_24217,N_20444,N_20006);
nor U24218 (N_24218,N_20269,N_22280);
nand U24219 (N_24219,N_20996,N_21806);
nand U24220 (N_24220,N_21509,N_20654);
and U24221 (N_24221,N_21922,N_20774);
xnor U24222 (N_24222,N_22150,N_20877);
and U24223 (N_24223,N_22228,N_20066);
or U24224 (N_24224,N_22282,N_22473);
nor U24225 (N_24225,N_21319,N_22310);
and U24226 (N_24226,N_22234,N_21317);
or U24227 (N_24227,N_22462,N_20034);
xnor U24228 (N_24228,N_20452,N_20338);
and U24229 (N_24229,N_21649,N_20861);
nor U24230 (N_24230,N_22359,N_21606);
xor U24231 (N_24231,N_20243,N_21240);
and U24232 (N_24232,N_21222,N_22172);
xor U24233 (N_24233,N_22124,N_20211);
and U24234 (N_24234,N_20296,N_20343);
xor U24235 (N_24235,N_22107,N_21741);
or U24236 (N_24236,N_21389,N_20832);
and U24237 (N_24237,N_20434,N_21480);
nand U24238 (N_24238,N_20633,N_22435);
and U24239 (N_24239,N_21406,N_20935);
or U24240 (N_24240,N_21857,N_22053);
nor U24241 (N_24241,N_21069,N_21022);
nor U24242 (N_24242,N_22452,N_20810);
nor U24243 (N_24243,N_22179,N_22164);
xnor U24244 (N_24244,N_21928,N_20985);
or U24245 (N_24245,N_21873,N_20905);
xor U24246 (N_24246,N_22118,N_20405);
xor U24247 (N_24247,N_20776,N_21495);
nor U24248 (N_24248,N_21177,N_21415);
or U24249 (N_24249,N_22116,N_22066);
nor U24250 (N_24250,N_21623,N_20522);
and U24251 (N_24251,N_20745,N_21979);
and U24252 (N_24252,N_21414,N_20563);
nand U24253 (N_24253,N_20533,N_21194);
nor U24254 (N_24254,N_21748,N_22400);
nand U24255 (N_24255,N_20706,N_20850);
xnor U24256 (N_24256,N_21616,N_22114);
nand U24257 (N_24257,N_22298,N_20405);
nor U24258 (N_24258,N_22031,N_22000);
nand U24259 (N_24259,N_21322,N_20712);
nand U24260 (N_24260,N_21755,N_20921);
and U24261 (N_24261,N_21841,N_20886);
and U24262 (N_24262,N_22142,N_20342);
or U24263 (N_24263,N_20936,N_20848);
nand U24264 (N_24264,N_21130,N_20211);
nor U24265 (N_24265,N_21576,N_22190);
and U24266 (N_24266,N_21046,N_22427);
and U24267 (N_24267,N_21078,N_21172);
xnor U24268 (N_24268,N_20413,N_21604);
nand U24269 (N_24269,N_22209,N_20382);
or U24270 (N_24270,N_20035,N_20534);
or U24271 (N_24271,N_20027,N_21109);
nand U24272 (N_24272,N_20931,N_21306);
xor U24273 (N_24273,N_20375,N_20799);
nand U24274 (N_24274,N_21280,N_20826);
xnor U24275 (N_24275,N_20497,N_20366);
or U24276 (N_24276,N_21899,N_21013);
or U24277 (N_24277,N_22058,N_20026);
nand U24278 (N_24278,N_21192,N_22305);
or U24279 (N_24279,N_21455,N_22490);
or U24280 (N_24280,N_21161,N_21086);
or U24281 (N_24281,N_20529,N_22174);
or U24282 (N_24282,N_21913,N_21223);
nand U24283 (N_24283,N_22439,N_20642);
nor U24284 (N_24284,N_22442,N_22341);
nand U24285 (N_24285,N_20886,N_21288);
and U24286 (N_24286,N_20430,N_20106);
and U24287 (N_24287,N_22063,N_22311);
or U24288 (N_24288,N_22008,N_20203);
xnor U24289 (N_24289,N_22007,N_21661);
nor U24290 (N_24290,N_21084,N_22466);
and U24291 (N_24291,N_21275,N_22252);
xnor U24292 (N_24292,N_20121,N_20861);
or U24293 (N_24293,N_21943,N_20055);
xor U24294 (N_24294,N_22481,N_20696);
nand U24295 (N_24295,N_21096,N_20758);
xnor U24296 (N_24296,N_20982,N_20447);
or U24297 (N_24297,N_21750,N_22132);
nor U24298 (N_24298,N_21151,N_22220);
nand U24299 (N_24299,N_22389,N_21573);
nand U24300 (N_24300,N_21072,N_22189);
xor U24301 (N_24301,N_21664,N_20725);
nand U24302 (N_24302,N_21891,N_22071);
nand U24303 (N_24303,N_20805,N_21206);
nand U24304 (N_24304,N_22054,N_20795);
or U24305 (N_24305,N_21925,N_21704);
nand U24306 (N_24306,N_22332,N_20877);
or U24307 (N_24307,N_20381,N_21891);
or U24308 (N_24308,N_20446,N_21913);
xor U24309 (N_24309,N_20154,N_21471);
and U24310 (N_24310,N_20601,N_21218);
nor U24311 (N_24311,N_21727,N_21823);
or U24312 (N_24312,N_20879,N_22491);
nor U24313 (N_24313,N_20751,N_20806);
and U24314 (N_24314,N_22391,N_20652);
or U24315 (N_24315,N_22086,N_20599);
or U24316 (N_24316,N_20564,N_21716);
and U24317 (N_24317,N_22027,N_20067);
and U24318 (N_24318,N_22247,N_21882);
or U24319 (N_24319,N_20904,N_21234);
and U24320 (N_24320,N_20308,N_20825);
xnor U24321 (N_24321,N_20415,N_21667);
nor U24322 (N_24322,N_22017,N_21825);
xor U24323 (N_24323,N_20475,N_21741);
xor U24324 (N_24324,N_20953,N_20051);
or U24325 (N_24325,N_21798,N_20541);
nor U24326 (N_24326,N_20211,N_20123);
nand U24327 (N_24327,N_22202,N_20359);
and U24328 (N_24328,N_20179,N_21366);
or U24329 (N_24329,N_21689,N_22079);
xnor U24330 (N_24330,N_20670,N_20823);
or U24331 (N_24331,N_21010,N_21103);
and U24332 (N_24332,N_20936,N_22344);
nor U24333 (N_24333,N_20132,N_22186);
nand U24334 (N_24334,N_21332,N_20875);
and U24335 (N_24335,N_21165,N_20724);
and U24336 (N_24336,N_20259,N_21641);
nand U24337 (N_24337,N_21878,N_21247);
or U24338 (N_24338,N_21352,N_20808);
and U24339 (N_24339,N_20998,N_21556);
or U24340 (N_24340,N_21029,N_21468);
or U24341 (N_24341,N_21858,N_20706);
nor U24342 (N_24342,N_20527,N_22173);
nor U24343 (N_24343,N_21474,N_21668);
xnor U24344 (N_24344,N_21886,N_22160);
or U24345 (N_24345,N_20788,N_20342);
nand U24346 (N_24346,N_22222,N_22193);
nand U24347 (N_24347,N_20852,N_22181);
or U24348 (N_24348,N_21563,N_20772);
nor U24349 (N_24349,N_21141,N_22459);
or U24350 (N_24350,N_21062,N_20387);
and U24351 (N_24351,N_21312,N_20734);
xor U24352 (N_24352,N_21567,N_22389);
nor U24353 (N_24353,N_21644,N_20573);
and U24354 (N_24354,N_20402,N_20384);
nand U24355 (N_24355,N_21009,N_20645);
xnor U24356 (N_24356,N_21777,N_21697);
nor U24357 (N_24357,N_20169,N_21178);
nand U24358 (N_24358,N_21257,N_21815);
xor U24359 (N_24359,N_22416,N_21514);
or U24360 (N_24360,N_20350,N_22294);
and U24361 (N_24361,N_22020,N_21880);
and U24362 (N_24362,N_21066,N_20978);
nor U24363 (N_24363,N_21250,N_21944);
xor U24364 (N_24364,N_20109,N_20372);
or U24365 (N_24365,N_21842,N_20801);
xor U24366 (N_24366,N_20822,N_21050);
xor U24367 (N_24367,N_21380,N_21390);
xor U24368 (N_24368,N_21744,N_20512);
and U24369 (N_24369,N_20327,N_22111);
nand U24370 (N_24370,N_21525,N_21698);
xnor U24371 (N_24371,N_21386,N_20394);
nor U24372 (N_24372,N_21936,N_20481);
nand U24373 (N_24373,N_20745,N_20658);
nand U24374 (N_24374,N_21963,N_21435);
nor U24375 (N_24375,N_20858,N_22011);
nor U24376 (N_24376,N_20937,N_20930);
and U24377 (N_24377,N_20777,N_21789);
nor U24378 (N_24378,N_22033,N_22487);
and U24379 (N_24379,N_20207,N_21216);
xnor U24380 (N_24380,N_21761,N_20105);
xor U24381 (N_24381,N_22386,N_20199);
nand U24382 (N_24382,N_20511,N_22139);
and U24383 (N_24383,N_22091,N_20303);
xor U24384 (N_24384,N_20896,N_20685);
nor U24385 (N_24385,N_20518,N_21994);
or U24386 (N_24386,N_20247,N_20469);
or U24387 (N_24387,N_20625,N_20531);
nand U24388 (N_24388,N_20392,N_20022);
nand U24389 (N_24389,N_20683,N_20113);
xor U24390 (N_24390,N_20767,N_21231);
and U24391 (N_24391,N_22147,N_21827);
nor U24392 (N_24392,N_21130,N_20694);
nor U24393 (N_24393,N_21240,N_22157);
xor U24394 (N_24394,N_20478,N_21180);
nor U24395 (N_24395,N_21082,N_21093);
nor U24396 (N_24396,N_22448,N_21191);
and U24397 (N_24397,N_21092,N_20551);
nor U24398 (N_24398,N_20744,N_21619);
nand U24399 (N_24399,N_21640,N_22309);
nand U24400 (N_24400,N_21958,N_20375);
xor U24401 (N_24401,N_21127,N_21727);
nor U24402 (N_24402,N_21671,N_22009);
and U24403 (N_24403,N_21739,N_21997);
and U24404 (N_24404,N_21812,N_21977);
nand U24405 (N_24405,N_20706,N_20418);
nand U24406 (N_24406,N_21090,N_20495);
nand U24407 (N_24407,N_21721,N_20052);
and U24408 (N_24408,N_21620,N_21785);
or U24409 (N_24409,N_22235,N_20617);
nand U24410 (N_24410,N_20273,N_21096);
xor U24411 (N_24411,N_20784,N_21153);
nor U24412 (N_24412,N_21220,N_20410);
nor U24413 (N_24413,N_22463,N_22394);
xor U24414 (N_24414,N_22069,N_21563);
nor U24415 (N_24415,N_22356,N_20612);
xor U24416 (N_24416,N_20714,N_21034);
xnor U24417 (N_24417,N_22255,N_20685);
nand U24418 (N_24418,N_22478,N_20986);
and U24419 (N_24419,N_20924,N_21640);
or U24420 (N_24420,N_22195,N_20396);
nand U24421 (N_24421,N_20377,N_20484);
nand U24422 (N_24422,N_22304,N_20614);
and U24423 (N_24423,N_21757,N_20873);
nor U24424 (N_24424,N_22025,N_20252);
xnor U24425 (N_24425,N_22210,N_20863);
or U24426 (N_24426,N_20781,N_21338);
nand U24427 (N_24427,N_20703,N_21423);
nand U24428 (N_24428,N_20210,N_20212);
xor U24429 (N_24429,N_21468,N_21879);
xnor U24430 (N_24430,N_20724,N_20794);
nor U24431 (N_24431,N_22353,N_21481);
nor U24432 (N_24432,N_20047,N_20518);
xor U24433 (N_24433,N_20312,N_21156);
nor U24434 (N_24434,N_22243,N_22493);
or U24435 (N_24435,N_20222,N_21159);
nand U24436 (N_24436,N_21428,N_20771);
nand U24437 (N_24437,N_20882,N_22211);
nor U24438 (N_24438,N_22093,N_22023);
or U24439 (N_24439,N_21843,N_20197);
or U24440 (N_24440,N_20890,N_20403);
and U24441 (N_24441,N_20017,N_20937);
and U24442 (N_24442,N_21078,N_22204);
xor U24443 (N_24443,N_20541,N_20714);
nor U24444 (N_24444,N_20553,N_20761);
or U24445 (N_24445,N_20820,N_21306);
or U24446 (N_24446,N_20542,N_20842);
and U24447 (N_24447,N_21822,N_20579);
and U24448 (N_24448,N_22349,N_21275);
or U24449 (N_24449,N_21173,N_21538);
xor U24450 (N_24450,N_21734,N_22238);
xnor U24451 (N_24451,N_21902,N_21196);
xnor U24452 (N_24452,N_21360,N_21185);
or U24453 (N_24453,N_20986,N_21227);
xor U24454 (N_24454,N_22457,N_20319);
nand U24455 (N_24455,N_21206,N_22029);
xor U24456 (N_24456,N_20423,N_22335);
nand U24457 (N_24457,N_21726,N_20306);
nand U24458 (N_24458,N_22110,N_21985);
or U24459 (N_24459,N_21128,N_21959);
nand U24460 (N_24460,N_21526,N_21623);
xnor U24461 (N_24461,N_22035,N_21418);
and U24462 (N_24462,N_21684,N_21513);
and U24463 (N_24463,N_21135,N_20626);
nor U24464 (N_24464,N_22097,N_20310);
nand U24465 (N_24465,N_20538,N_20704);
xnor U24466 (N_24466,N_20440,N_21094);
or U24467 (N_24467,N_20661,N_21415);
or U24468 (N_24468,N_20745,N_22138);
xor U24469 (N_24469,N_21025,N_20665);
or U24470 (N_24470,N_21776,N_22139);
or U24471 (N_24471,N_22105,N_22021);
or U24472 (N_24472,N_22181,N_21883);
and U24473 (N_24473,N_20350,N_22029);
xor U24474 (N_24474,N_20401,N_20474);
or U24475 (N_24475,N_20989,N_20239);
nand U24476 (N_24476,N_21267,N_21507);
and U24477 (N_24477,N_22180,N_20285);
xnor U24478 (N_24478,N_20670,N_20304);
or U24479 (N_24479,N_21844,N_21644);
nand U24480 (N_24480,N_20867,N_21298);
nor U24481 (N_24481,N_21828,N_21013);
nor U24482 (N_24482,N_20262,N_21285);
nor U24483 (N_24483,N_20620,N_20575);
and U24484 (N_24484,N_21877,N_21866);
nor U24485 (N_24485,N_21406,N_22338);
nand U24486 (N_24486,N_20412,N_22463);
and U24487 (N_24487,N_21475,N_22178);
xor U24488 (N_24488,N_22454,N_20173);
or U24489 (N_24489,N_21586,N_20288);
xor U24490 (N_24490,N_21386,N_21290);
nand U24491 (N_24491,N_20295,N_20009);
xnor U24492 (N_24492,N_20076,N_20825);
xor U24493 (N_24493,N_20072,N_21247);
and U24494 (N_24494,N_21982,N_22115);
or U24495 (N_24495,N_21369,N_20255);
nor U24496 (N_24496,N_21787,N_22013);
and U24497 (N_24497,N_20924,N_21746);
or U24498 (N_24498,N_20080,N_21900);
nor U24499 (N_24499,N_21068,N_21400);
and U24500 (N_24500,N_20902,N_20557);
or U24501 (N_24501,N_20180,N_20392);
xor U24502 (N_24502,N_20698,N_22484);
xor U24503 (N_24503,N_20520,N_21198);
nand U24504 (N_24504,N_21885,N_20388);
and U24505 (N_24505,N_21394,N_20225);
nand U24506 (N_24506,N_21719,N_22116);
nor U24507 (N_24507,N_20513,N_21305);
xor U24508 (N_24508,N_21948,N_22206);
or U24509 (N_24509,N_20466,N_20897);
and U24510 (N_24510,N_20344,N_21898);
xnor U24511 (N_24511,N_20162,N_21856);
or U24512 (N_24512,N_20139,N_21469);
or U24513 (N_24513,N_20008,N_20373);
xor U24514 (N_24514,N_20385,N_21488);
or U24515 (N_24515,N_20536,N_22438);
nand U24516 (N_24516,N_21419,N_22440);
nor U24517 (N_24517,N_20807,N_20906);
nor U24518 (N_24518,N_20051,N_21201);
and U24519 (N_24519,N_20408,N_22384);
and U24520 (N_24520,N_21319,N_20664);
xor U24521 (N_24521,N_22438,N_21949);
nand U24522 (N_24522,N_22459,N_21159);
or U24523 (N_24523,N_22153,N_20425);
xnor U24524 (N_24524,N_21395,N_22036);
and U24525 (N_24525,N_21904,N_22446);
and U24526 (N_24526,N_20934,N_22480);
nand U24527 (N_24527,N_20524,N_20521);
and U24528 (N_24528,N_21988,N_22223);
nand U24529 (N_24529,N_22009,N_20015);
or U24530 (N_24530,N_20088,N_21305);
nand U24531 (N_24531,N_21904,N_20762);
nor U24532 (N_24532,N_21625,N_22174);
xor U24533 (N_24533,N_20008,N_21287);
nor U24534 (N_24534,N_20600,N_21437);
and U24535 (N_24535,N_20168,N_20172);
nand U24536 (N_24536,N_20870,N_20884);
and U24537 (N_24537,N_22179,N_20988);
or U24538 (N_24538,N_20276,N_22495);
nor U24539 (N_24539,N_20718,N_21083);
and U24540 (N_24540,N_22315,N_20615);
nand U24541 (N_24541,N_20822,N_20423);
nor U24542 (N_24542,N_22256,N_20593);
xnor U24543 (N_24543,N_20541,N_22245);
or U24544 (N_24544,N_20696,N_20113);
and U24545 (N_24545,N_20720,N_22356);
and U24546 (N_24546,N_22294,N_21587);
or U24547 (N_24547,N_20961,N_20452);
and U24548 (N_24548,N_22157,N_20467);
nand U24549 (N_24549,N_20912,N_22209);
nor U24550 (N_24550,N_20938,N_22257);
or U24551 (N_24551,N_20417,N_21411);
nor U24552 (N_24552,N_21762,N_22053);
or U24553 (N_24553,N_21357,N_22162);
nor U24554 (N_24554,N_21304,N_20907);
nand U24555 (N_24555,N_21016,N_20564);
xnor U24556 (N_24556,N_20762,N_21511);
or U24557 (N_24557,N_20184,N_21925);
and U24558 (N_24558,N_22419,N_22363);
xnor U24559 (N_24559,N_21266,N_21149);
and U24560 (N_24560,N_21207,N_20288);
or U24561 (N_24561,N_21426,N_21675);
xnor U24562 (N_24562,N_21480,N_20213);
nor U24563 (N_24563,N_20305,N_20643);
nand U24564 (N_24564,N_22432,N_22309);
or U24565 (N_24565,N_21112,N_21110);
or U24566 (N_24566,N_21103,N_20545);
or U24567 (N_24567,N_20377,N_21232);
or U24568 (N_24568,N_22160,N_21214);
nand U24569 (N_24569,N_20182,N_20189);
nand U24570 (N_24570,N_21181,N_20462);
nand U24571 (N_24571,N_20418,N_20197);
nand U24572 (N_24572,N_21040,N_21241);
and U24573 (N_24573,N_20082,N_22466);
xor U24574 (N_24574,N_20669,N_20209);
nand U24575 (N_24575,N_21118,N_22277);
nand U24576 (N_24576,N_20985,N_20442);
or U24577 (N_24577,N_22300,N_21761);
and U24578 (N_24578,N_21450,N_21503);
and U24579 (N_24579,N_20733,N_20209);
or U24580 (N_24580,N_22445,N_22388);
nand U24581 (N_24581,N_20218,N_20528);
xor U24582 (N_24582,N_20700,N_21254);
or U24583 (N_24583,N_21162,N_21090);
or U24584 (N_24584,N_21220,N_20062);
and U24585 (N_24585,N_22393,N_21867);
nand U24586 (N_24586,N_20297,N_21038);
nand U24587 (N_24587,N_21651,N_21592);
or U24588 (N_24588,N_20444,N_21520);
nand U24589 (N_24589,N_21543,N_21458);
nand U24590 (N_24590,N_22399,N_21802);
nor U24591 (N_24591,N_21727,N_20094);
or U24592 (N_24592,N_21403,N_21990);
nand U24593 (N_24593,N_20700,N_20746);
nand U24594 (N_24594,N_22235,N_20316);
nand U24595 (N_24595,N_21215,N_21576);
or U24596 (N_24596,N_21953,N_22268);
nor U24597 (N_24597,N_21309,N_20184);
nand U24598 (N_24598,N_20805,N_21331);
nor U24599 (N_24599,N_20788,N_20854);
nor U24600 (N_24600,N_20190,N_20560);
nor U24601 (N_24601,N_20850,N_22493);
xor U24602 (N_24602,N_22444,N_21780);
xnor U24603 (N_24603,N_20615,N_21569);
nor U24604 (N_24604,N_21060,N_20352);
nand U24605 (N_24605,N_20908,N_21404);
nor U24606 (N_24606,N_21956,N_22076);
or U24607 (N_24607,N_21353,N_20429);
xnor U24608 (N_24608,N_20145,N_21359);
nand U24609 (N_24609,N_20259,N_22231);
and U24610 (N_24610,N_20065,N_21104);
and U24611 (N_24611,N_20556,N_21189);
nand U24612 (N_24612,N_22474,N_20057);
or U24613 (N_24613,N_22253,N_20701);
xnor U24614 (N_24614,N_20566,N_20288);
and U24615 (N_24615,N_22244,N_20996);
xor U24616 (N_24616,N_20160,N_20313);
and U24617 (N_24617,N_21115,N_21597);
nor U24618 (N_24618,N_22037,N_21549);
xnor U24619 (N_24619,N_22134,N_21103);
xor U24620 (N_24620,N_21168,N_22410);
and U24621 (N_24621,N_21007,N_21667);
nand U24622 (N_24622,N_21670,N_21841);
and U24623 (N_24623,N_21317,N_20312);
and U24624 (N_24624,N_20488,N_20294);
nor U24625 (N_24625,N_21657,N_20716);
nor U24626 (N_24626,N_21381,N_20730);
nor U24627 (N_24627,N_20301,N_22352);
and U24628 (N_24628,N_22101,N_20279);
xnor U24629 (N_24629,N_20732,N_20932);
nand U24630 (N_24630,N_20278,N_21823);
nand U24631 (N_24631,N_20857,N_21751);
xnor U24632 (N_24632,N_22074,N_20839);
xnor U24633 (N_24633,N_20468,N_21261);
nand U24634 (N_24634,N_21505,N_20797);
and U24635 (N_24635,N_21311,N_22055);
nor U24636 (N_24636,N_21308,N_20225);
nand U24637 (N_24637,N_21049,N_20646);
and U24638 (N_24638,N_22012,N_22419);
nor U24639 (N_24639,N_20883,N_20811);
or U24640 (N_24640,N_21886,N_20514);
and U24641 (N_24641,N_21816,N_22183);
or U24642 (N_24642,N_20281,N_20630);
nand U24643 (N_24643,N_21189,N_21400);
xnor U24644 (N_24644,N_20979,N_21377);
nand U24645 (N_24645,N_21761,N_21736);
and U24646 (N_24646,N_21520,N_20283);
xor U24647 (N_24647,N_21422,N_22220);
and U24648 (N_24648,N_22458,N_20267);
nor U24649 (N_24649,N_21578,N_21180);
nand U24650 (N_24650,N_21595,N_21677);
xor U24651 (N_24651,N_20243,N_20805);
and U24652 (N_24652,N_20344,N_21963);
or U24653 (N_24653,N_21055,N_22150);
or U24654 (N_24654,N_21808,N_21771);
xor U24655 (N_24655,N_20092,N_21775);
or U24656 (N_24656,N_20123,N_20491);
nand U24657 (N_24657,N_21530,N_21638);
nand U24658 (N_24658,N_22409,N_20436);
and U24659 (N_24659,N_21305,N_21065);
or U24660 (N_24660,N_21861,N_20290);
or U24661 (N_24661,N_21965,N_20920);
nor U24662 (N_24662,N_20466,N_20974);
nor U24663 (N_24663,N_20069,N_20447);
and U24664 (N_24664,N_20173,N_20334);
xnor U24665 (N_24665,N_20731,N_20267);
xnor U24666 (N_24666,N_22449,N_20421);
nor U24667 (N_24667,N_21675,N_22300);
nor U24668 (N_24668,N_21680,N_21083);
nor U24669 (N_24669,N_20001,N_21885);
nor U24670 (N_24670,N_20705,N_20428);
nand U24671 (N_24671,N_21176,N_20178);
nand U24672 (N_24672,N_21660,N_22043);
xnor U24673 (N_24673,N_22008,N_20177);
nor U24674 (N_24674,N_22259,N_21273);
xor U24675 (N_24675,N_22443,N_22186);
or U24676 (N_24676,N_21890,N_22422);
nor U24677 (N_24677,N_22298,N_21285);
or U24678 (N_24678,N_20605,N_21697);
nor U24679 (N_24679,N_21771,N_20366);
xor U24680 (N_24680,N_21848,N_21366);
nor U24681 (N_24681,N_22093,N_21071);
nor U24682 (N_24682,N_22004,N_22048);
xor U24683 (N_24683,N_22096,N_21971);
xor U24684 (N_24684,N_21420,N_21454);
nand U24685 (N_24685,N_21770,N_21064);
and U24686 (N_24686,N_20647,N_21451);
nand U24687 (N_24687,N_22137,N_22407);
xnor U24688 (N_24688,N_21106,N_22054);
nor U24689 (N_24689,N_20065,N_21750);
xnor U24690 (N_24690,N_21692,N_22135);
xor U24691 (N_24691,N_21983,N_22319);
nor U24692 (N_24692,N_22184,N_21963);
nor U24693 (N_24693,N_20647,N_20617);
nor U24694 (N_24694,N_21351,N_20207);
nor U24695 (N_24695,N_22246,N_21125);
nor U24696 (N_24696,N_22152,N_22327);
nor U24697 (N_24697,N_20308,N_22365);
nor U24698 (N_24698,N_21822,N_20887);
nand U24699 (N_24699,N_20588,N_21143);
nor U24700 (N_24700,N_20835,N_21978);
or U24701 (N_24701,N_21800,N_21531);
or U24702 (N_24702,N_21681,N_22091);
nor U24703 (N_24703,N_20062,N_22322);
and U24704 (N_24704,N_22448,N_21660);
and U24705 (N_24705,N_21747,N_20405);
or U24706 (N_24706,N_21564,N_20217);
or U24707 (N_24707,N_21007,N_20025);
nor U24708 (N_24708,N_20286,N_21571);
or U24709 (N_24709,N_20775,N_21741);
and U24710 (N_24710,N_20532,N_22192);
and U24711 (N_24711,N_20904,N_20931);
or U24712 (N_24712,N_21828,N_21882);
xnor U24713 (N_24713,N_22088,N_20018);
nand U24714 (N_24714,N_20648,N_22348);
xnor U24715 (N_24715,N_21305,N_20391);
nand U24716 (N_24716,N_20580,N_21994);
nand U24717 (N_24717,N_22092,N_22433);
or U24718 (N_24718,N_22136,N_21273);
nand U24719 (N_24719,N_20866,N_22124);
nand U24720 (N_24720,N_22098,N_21245);
nor U24721 (N_24721,N_20724,N_21075);
xnor U24722 (N_24722,N_21747,N_21976);
and U24723 (N_24723,N_20365,N_20124);
and U24724 (N_24724,N_20859,N_22411);
nand U24725 (N_24725,N_20343,N_21695);
nand U24726 (N_24726,N_21368,N_20470);
and U24727 (N_24727,N_20692,N_20632);
xor U24728 (N_24728,N_22272,N_21869);
and U24729 (N_24729,N_20320,N_21679);
xor U24730 (N_24730,N_20618,N_21065);
nor U24731 (N_24731,N_22386,N_20374);
or U24732 (N_24732,N_21545,N_22055);
and U24733 (N_24733,N_22411,N_22460);
nand U24734 (N_24734,N_21894,N_22341);
nand U24735 (N_24735,N_22218,N_20901);
nand U24736 (N_24736,N_21534,N_22024);
nor U24737 (N_24737,N_21180,N_20406);
nor U24738 (N_24738,N_22057,N_20789);
nand U24739 (N_24739,N_20472,N_20967);
nor U24740 (N_24740,N_21563,N_22182);
and U24741 (N_24741,N_21288,N_21753);
and U24742 (N_24742,N_22465,N_20006);
or U24743 (N_24743,N_21141,N_21678);
nand U24744 (N_24744,N_22072,N_20274);
or U24745 (N_24745,N_21396,N_22439);
or U24746 (N_24746,N_21571,N_20022);
and U24747 (N_24747,N_20297,N_20320);
or U24748 (N_24748,N_20764,N_21389);
nor U24749 (N_24749,N_20941,N_20223);
nor U24750 (N_24750,N_20113,N_20549);
or U24751 (N_24751,N_20036,N_20407);
nor U24752 (N_24752,N_21606,N_20460);
and U24753 (N_24753,N_21930,N_22471);
xnor U24754 (N_24754,N_21693,N_21585);
xor U24755 (N_24755,N_21481,N_20641);
xor U24756 (N_24756,N_22053,N_22398);
nand U24757 (N_24757,N_20163,N_21761);
nand U24758 (N_24758,N_20585,N_20329);
or U24759 (N_24759,N_22471,N_21131);
xor U24760 (N_24760,N_22144,N_21994);
and U24761 (N_24761,N_21393,N_22328);
nor U24762 (N_24762,N_22024,N_20451);
nor U24763 (N_24763,N_21479,N_20431);
or U24764 (N_24764,N_22014,N_21372);
xnor U24765 (N_24765,N_22001,N_21622);
and U24766 (N_24766,N_21161,N_20382);
nand U24767 (N_24767,N_20273,N_20737);
or U24768 (N_24768,N_21524,N_20995);
xor U24769 (N_24769,N_20578,N_21191);
and U24770 (N_24770,N_21551,N_20685);
xor U24771 (N_24771,N_20458,N_21058);
nor U24772 (N_24772,N_22207,N_21977);
or U24773 (N_24773,N_22193,N_21684);
nor U24774 (N_24774,N_20095,N_21959);
nor U24775 (N_24775,N_22458,N_21691);
or U24776 (N_24776,N_22072,N_20169);
nand U24777 (N_24777,N_20312,N_20596);
or U24778 (N_24778,N_21055,N_22363);
and U24779 (N_24779,N_20630,N_21544);
nand U24780 (N_24780,N_22340,N_22420);
and U24781 (N_24781,N_20275,N_21250);
nand U24782 (N_24782,N_21759,N_22105);
and U24783 (N_24783,N_20313,N_21133);
nand U24784 (N_24784,N_21558,N_21302);
nand U24785 (N_24785,N_21853,N_20464);
xor U24786 (N_24786,N_21037,N_22421);
or U24787 (N_24787,N_21601,N_21410);
nand U24788 (N_24788,N_21708,N_21985);
or U24789 (N_24789,N_20048,N_22106);
and U24790 (N_24790,N_20768,N_22154);
xor U24791 (N_24791,N_20224,N_20016);
or U24792 (N_24792,N_20674,N_21214);
and U24793 (N_24793,N_22359,N_20277);
nand U24794 (N_24794,N_20327,N_20051);
and U24795 (N_24795,N_21928,N_20644);
or U24796 (N_24796,N_21875,N_20243);
or U24797 (N_24797,N_22234,N_21937);
and U24798 (N_24798,N_22190,N_22187);
and U24799 (N_24799,N_21457,N_21717);
nand U24800 (N_24800,N_20757,N_20335);
and U24801 (N_24801,N_20617,N_21603);
nand U24802 (N_24802,N_21155,N_21715);
or U24803 (N_24803,N_20061,N_21886);
xnor U24804 (N_24804,N_22039,N_20648);
nand U24805 (N_24805,N_20744,N_22429);
nand U24806 (N_24806,N_20177,N_21049);
nand U24807 (N_24807,N_22060,N_20546);
nand U24808 (N_24808,N_22300,N_22082);
nor U24809 (N_24809,N_22162,N_20343);
nand U24810 (N_24810,N_22068,N_22039);
xnor U24811 (N_24811,N_22416,N_20198);
and U24812 (N_24812,N_21648,N_21819);
nor U24813 (N_24813,N_20831,N_20905);
nand U24814 (N_24814,N_21368,N_22285);
nand U24815 (N_24815,N_20627,N_21239);
xnor U24816 (N_24816,N_20568,N_20376);
nand U24817 (N_24817,N_20271,N_21501);
xnor U24818 (N_24818,N_21399,N_22372);
nand U24819 (N_24819,N_22117,N_20637);
nand U24820 (N_24820,N_21729,N_21531);
nand U24821 (N_24821,N_22465,N_21287);
nand U24822 (N_24822,N_22099,N_21729);
nor U24823 (N_24823,N_21134,N_22108);
nand U24824 (N_24824,N_20464,N_21987);
nor U24825 (N_24825,N_20047,N_21593);
xnor U24826 (N_24826,N_20077,N_20378);
nor U24827 (N_24827,N_21026,N_21888);
nor U24828 (N_24828,N_21862,N_22189);
or U24829 (N_24829,N_20710,N_21261);
nor U24830 (N_24830,N_20361,N_22450);
nand U24831 (N_24831,N_22354,N_22342);
and U24832 (N_24832,N_21747,N_21643);
nor U24833 (N_24833,N_20521,N_22174);
xor U24834 (N_24834,N_20602,N_20131);
xnor U24835 (N_24835,N_22143,N_20436);
or U24836 (N_24836,N_21025,N_21116);
and U24837 (N_24837,N_22464,N_20955);
and U24838 (N_24838,N_21504,N_21382);
nand U24839 (N_24839,N_21346,N_21616);
xor U24840 (N_24840,N_22070,N_20398);
or U24841 (N_24841,N_22178,N_21421);
or U24842 (N_24842,N_21637,N_21376);
xnor U24843 (N_24843,N_20423,N_20781);
xnor U24844 (N_24844,N_21104,N_22236);
or U24845 (N_24845,N_22180,N_20552);
xor U24846 (N_24846,N_22131,N_20426);
and U24847 (N_24847,N_21520,N_20267);
nand U24848 (N_24848,N_22002,N_20779);
nor U24849 (N_24849,N_21284,N_20274);
nand U24850 (N_24850,N_21195,N_20816);
or U24851 (N_24851,N_20294,N_21996);
or U24852 (N_24852,N_22326,N_21092);
and U24853 (N_24853,N_21093,N_21088);
and U24854 (N_24854,N_22477,N_21763);
and U24855 (N_24855,N_20943,N_20928);
xnor U24856 (N_24856,N_20900,N_22026);
xor U24857 (N_24857,N_20356,N_21648);
nand U24858 (N_24858,N_20913,N_20262);
and U24859 (N_24859,N_22126,N_20635);
nor U24860 (N_24860,N_20831,N_21920);
xnor U24861 (N_24861,N_20475,N_20860);
and U24862 (N_24862,N_21830,N_22040);
nand U24863 (N_24863,N_21841,N_20965);
and U24864 (N_24864,N_21147,N_20051);
nor U24865 (N_24865,N_22395,N_20722);
nand U24866 (N_24866,N_20728,N_20721);
nand U24867 (N_24867,N_22347,N_20947);
and U24868 (N_24868,N_21233,N_21390);
nor U24869 (N_24869,N_22269,N_20858);
or U24870 (N_24870,N_20271,N_21553);
nand U24871 (N_24871,N_21088,N_20209);
or U24872 (N_24872,N_21926,N_21363);
or U24873 (N_24873,N_22126,N_21633);
nor U24874 (N_24874,N_20838,N_21696);
and U24875 (N_24875,N_21264,N_20094);
or U24876 (N_24876,N_20620,N_20917);
nand U24877 (N_24877,N_20034,N_21642);
and U24878 (N_24878,N_21523,N_21532);
nor U24879 (N_24879,N_20062,N_20218);
or U24880 (N_24880,N_22124,N_22098);
nand U24881 (N_24881,N_21776,N_20609);
nor U24882 (N_24882,N_20835,N_21906);
nand U24883 (N_24883,N_21579,N_20385);
and U24884 (N_24884,N_22148,N_21260);
nand U24885 (N_24885,N_20676,N_20356);
and U24886 (N_24886,N_21925,N_20591);
nand U24887 (N_24887,N_20723,N_21973);
xnor U24888 (N_24888,N_22099,N_21132);
nor U24889 (N_24889,N_22131,N_21347);
and U24890 (N_24890,N_20776,N_21175);
nor U24891 (N_24891,N_22010,N_22079);
or U24892 (N_24892,N_21035,N_20729);
nand U24893 (N_24893,N_20169,N_20330);
or U24894 (N_24894,N_21983,N_21338);
nor U24895 (N_24895,N_21139,N_20784);
nor U24896 (N_24896,N_21731,N_22376);
nand U24897 (N_24897,N_21020,N_22484);
nand U24898 (N_24898,N_21070,N_20553);
xor U24899 (N_24899,N_21573,N_22073);
and U24900 (N_24900,N_22497,N_21277);
nor U24901 (N_24901,N_21762,N_21068);
and U24902 (N_24902,N_20964,N_20939);
or U24903 (N_24903,N_20040,N_21954);
and U24904 (N_24904,N_22212,N_20463);
nor U24905 (N_24905,N_22338,N_20374);
nor U24906 (N_24906,N_21785,N_20233);
nand U24907 (N_24907,N_20738,N_21787);
nor U24908 (N_24908,N_21501,N_21304);
and U24909 (N_24909,N_20609,N_20775);
xor U24910 (N_24910,N_20703,N_21485);
or U24911 (N_24911,N_21523,N_21291);
and U24912 (N_24912,N_21425,N_20379);
or U24913 (N_24913,N_21345,N_20261);
xnor U24914 (N_24914,N_21556,N_20731);
or U24915 (N_24915,N_21909,N_22204);
or U24916 (N_24916,N_21812,N_22361);
or U24917 (N_24917,N_21335,N_22052);
nand U24918 (N_24918,N_22189,N_21713);
and U24919 (N_24919,N_20651,N_20258);
xor U24920 (N_24920,N_20681,N_20366);
or U24921 (N_24921,N_20491,N_21851);
or U24922 (N_24922,N_20776,N_21666);
or U24923 (N_24923,N_21357,N_22307);
or U24924 (N_24924,N_21574,N_21644);
or U24925 (N_24925,N_20056,N_22292);
and U24926 (N_24926,N_20507,N_22233);
xor U24927 (N_24927,N_20375,N_20844);
xnor U24928 (N_24928,N_21294,N_21404);
nand U24929 (N_24929,N_20500,N_22355);
nor U24930 (N_24930,N_22006,N_20142);
or U24931 (N_24931,N_20772,N_20511);
nand U24932 (N_24932,N_22206,N_20184);
and U24933 (N_24933,N_21253,N_21845);
xor U24934 (N_24934,N_21320,N_22284);
nand U24935 (N_24935,N_20224,N_21034);
or U24936 (N_24936,N_22200,N_20511);
nand U24937 (N_24937,N_21875,N_20503);
nor U24938 (N_24938,N_20530,N_20897);
and U24939 (N_24939,N_20016,N_21903);
nand U24940 (N_24940,N_20111,N_20403);
nand U24941 (N_24941,N_20116,N_21314);
or U24942 (N_24942,N_22222,N_21712);
or U24943 (N_24943,N_21031,N_22293);
xnor U24944 (N_24944,N_20389,N_21739);
nor U24945 (N_24945,N_20162,N_20155);
or U24946 (N_24946,N_22371,N_20158);
xor U24947 (N_24947,N_21916,N_20288);
and U24948 (N_24948,N_20138,N_21065);
nor U24949 (N_24949,N_20902,N_21719);
nor U24950 (N_24950,N_20759,N_20488);
nor U24951 (N_24951,N_21154,N_20152);
or U24952 (N_24952,N_22034,N_22288);
nor U24953 (N_24953,N_20745,N_21179);
nand U24954 (N_24954,N_20766,N_20089);
nand U24955 (N_24955,N_22488,N_22478);
or U24956 (N_24956,N_21483,N_21161);
or U24957 (N_24957,N_20649,N_22094);
xnor U24958 (N_24958,N_21449,N_20961);
xor U24959 (N_24959,N_21876,N_22306);
xnor U24960 (N_24960,N_20146,N_22473);
nor U24961 (N_24961,N_21313,N_22352);
nand U24962 (N_24962,N_20043,N_20176);
or U24963 (N_24963,N_20982,N_20772);
nand U24964 (N_24964,N_21254,N_21949);
nor U24965 (N_24965,N_21034,N_22027);
nor U24966 (N_24966,N_22080,N_20822);
nor U24967 (N_24967,N_20632,N_20081);
nand U24968 (N_24968,N_22283,N_22017);
nand U24969 (N_24969,N_20592,N_22026);
nor U24970 (N_24970,N_21994,N_21826);
nor U24971 (N_24971,N_20735,N_22422);
nand U24972 (N_24972,N_20566,N_20488);
xnor U24973 (N_24973,N_21940,N_21711);
xnor U24974 (N_24974,N_22438,N_21660);
nor U24975 (N_24975,N_21214,N_20475);
nor U24976 (N_24976,N_22319,N_21741);
and U24977 (N_24977,N_21260,N_22224);
and U24978 (N_24978,N_21370,N_21445);
xor U24979 (N_24979,N_21566,N_20920);
xor U24980 (N_24980,N_21101,N_20255);
or U24981 (N_24981,N_20060,N_22230);
nand U24982 (N_24982,N_21297,N_22001);
nor U24983 (N_24983,N_21040,N_22219);
and U24984 (N_24984,N_22228,N_22010);
nor U24985 (N_24985,N_20247,N_22047);
xor U24986 (N_24986,N_21083,N_22246);
and U24987 (N_24987,N_21726,N_20010);
nand U24988 (N_24988,N_21545,N_21811);
or U24989 (N_24989,N_21840,N_22169);
or U24990 (N_24990,N_22021,N_21779);
or U24991 (N_24991,N_20475,N_22019);
nor U24992 (N_24992,N_20818,N_20605);
xnor U24993 (N_24993,N_20611,N_21845);
nor U24994 (N_24994,N_22498,N_20544);
or U24995 (N_24995,N_21179,N_21712);
xor U24996 (N_24996,N_21351,N_22175);
and U24997 (N_24997,N_22341,N_20718);
and U24998 (N_24998,N_20285,N_20898);
or U24999 (N_24999,N_21508,N_21465);
and U25000 (N_25000,N_24191,N_22622);
xor U25001 (N_25001,N_23082,N_24462);
xnor U25002 (N_25002,N_23788,N_24030);
or U25003 (N_25003,N_22812,N_24338);
and U25004 (N_25004,N_22672,N_23341);
xnor U25005 (N_25005,N_23630,N_24696);
nand U25006 (N_25006,N_22788,N_23045);
xor U25007 (N_25007,N_24291,N_22720);
nor U25008 (N_25008,N_22693,N_23573);
nand U25009 (N_25009,N_23653,N_23142);
nor U25010 (N_25010,N_23842,N_24487);
nand U25011 (N_25011,N_22866,N_24852);
or U25012 (N_25012,N_24150,N_24471);
or U25013 (N_25013,N_23294,N_22536);
nand U25014 (N_25014,N_23518,N_24947);
and U25015 (N_25015,N_22774,N_24490);
and U25016 (N_25016,N_24472,N_22530);
xnor U25017 (N_25017,N_22817,N_24516);
and U25018 (N_25018,N_23137,N_24101);
nor U25019 (N_25019,N_24033,N_23458);
nor U25020 (N_25020,N_22845,N_24991);
or U25021 (N_25021,N_23544,N_23475);
nor U25022 (N_25022,N_23741,N_24697);
nor U25023 (N_25023,N_23574,N_24394);
or U25024 (N_25024,N_23049,N_23388);
xor U25025 (N_25025,N_24458,N_23827);
nand U25026 (N_25026,N_23925,N_24190);
and U25027 (N_25027,N_23107,N_23570);
nand U25028 (N_25028,N_22885,N_23516);
and U25029 (N_25029,N_23395,N_22811);
xnor U25030 (N_25030,N_24570,N_23365);
or U25031 (N_25031,N_23414,N_23227);
and U25032 (N_25032,N_24295,N_23742);
xnor U25033 (N_25033,N_23411,N_24773);
or U25034 (N_25034,N_24774,N_24066);
or U25035 (N_25035,N_23609,N_23638);
or U25036 (N_25036,N_23718,N_24767);
nor U25037 (N_25037,N_24715,N_22963);
xnor U25038 (N_25038,N_23121,N_23471);
xnor U25039 (N_25039,N_23891,N_24902);
nor U25040 (N_25040,N_22697,N_22784);
or U25041 (N_25041,N_24287,N_22907);
or U25042 (N_25042,N_22517,N_22971);
or U25043 (N_25043,N_24615,N_23831);
xor U25044 (N_25044,N_23649,N_23938);
and U25045 (N_25045,N_23571,N_23915);
or U25046 (N_25046,N_23992,N_24451);
and U25047 (N_25047,N_24638,N_23665);
nand U25048 (N_25048,N_24138,N_24561);
or U25049 (N_25049,N_23507,N_23093);
nand U25050 (N_25050,N_23729,N_24145);
nand U25051 (N_25051,N_24447,N_22991);
or U25052 (N_25052,N_23958,N_23246);
or U25053 (N_25053,N_22883,N_23619);
xor U25054 (N_25054,N_24165,N_23690);
nand U25055 (N_25055,N_23862,N_22700);
nor U25056 (N_25056,N_24370,N_23401);
nand U25057 (N_25057,N_23044,N_24569);
or U25058 (N_25058,N_23282,N_23855);
nor U25059 (N_25059,N_23375,N_24979);
xor U25060 (N_25060,N_24685,N_22712);
xor U25061 (N_25061,N_24061,N_23789);
nand U25062 (N_25062,N_23556,N_23013);
and U25063 (N_25063,N_22943,N_24804);
xor U25064 (N_25064,N_22834,N_23519);
xor U25065 (N_25065,N_23515,N_22641);
xnor U25066 (N_25066,N_23616,N_24015);
xnor U25067 (N_25067,N_24938,N_22704);
nor U25068 (N_25068,N_24851,N_24203);
xor U25069 (N_25069,N_24357,N_24987);
or U25070 (N_25070,N_24022,N_22540);
xnor U25071 (N_25071,N_23140,N_24481);
nand U25072 (N_25072,N_23034,N_24620);
nand U25073 (N_25073,N_23525,N_22962);
nand U25074 (N_25074,N_24379,N_24673);
xnor U25075 (N_25075,N_24726,N_23203);
xor U25076 (N_25076,N_23845,N_23770);
nand U25077 (N_25077,N_23380,N_24466);
nor U25078 (N_25078,N_23250,N_22630);
and U25079 (N_25079,N_23091,N_23153);
or U25080 (N_25080,N_23982,N_23627);
nand U25081 (N_25081,N_22793,N_22930);
or U25082 (N_25082,N_23979,N_23870);
or U25083 (N_25083,N_24442,N_24353);
or U25084 (N_25084,N_23578,N_24996);
nor U25085 (N_25085,N_24185,N_22768);
and U25086 (N_25086,N_22782,N_24328);
nor U25087 (N_25087,N_23366,N_22518);
nand U25088 (N_25088,N_23465,N_24812);
and U25089 (N_25089,N_24577,N_23782);
or U25090 (N_25090,N_23815,N_23933);
or U25091 (N_25091,N_22719,N_22875);
or U25092 (N_25092,N_23917,N_24843);
xnor U25093 (N_25093,N_24054,N_23432);
or U25094 (N_25094,N_24867,N_24565);
nor U25095 (N_25095,N_23807,N_23099);
nand U25096 (N_25096,N_23071,N_24688);
nand U25097 (N_25097,N_23408,N_23932);
xor U25098 (N_25098,N_23115,N_24563);
or U25099 (N_25099,N_23779,N_24588);
nand U25100 (N_25100,N_23248,N_24684);
nor U25101 (N_25101,N_22614,N_23368);
and U25102 (N_25102,N_24452,N_24963);
and U25103 (N_25103,N_24955,N_24722);
nor U25104 (N_25104,N_23311,N_24250);
or U25105 (N_25105,N_24656,N_23672);
nor U25106 (N_25106,N_23639,N_23670);
nand U25107 (N_25107,N_24690,N_24853);
or U25108 (N_25108,N_22915,N_23088);
or U25109 (N_25109,N_24470,N_24412);
nand U25110 (N_25110,N_24512,N_22769);
nand U25111 (N_25111,N_23101,N_22957);
nor U25112 (N_25112,N_22613,N_22571);
nand U25113 (N_25113,N_24085,N_24670);
xnor U25114 (N_25114,N_23547,N_23890);
nand U25115 (N_25115,N_22946,N_24854);
xnor U25116 (N_25116,N_22561,N_24074);
and U25117 (N_25117,N_24510,N_23269);
nor U25118 (N_25118,N_24971,N_24933);
nor U25119 (N_25119,N_23764,N_23846);
xnor U25120 (N_25120,N_24477,N_23675);
nor U25121 (N_25121,N_22678,N_24527);
nand U25122 (N_25122,N_24498,N_24855);
xnor U25123 (N_25123,N_24461,N_23355);
nand U25124 (N_25124,N_23505,N_23343);
and U25125 (N_25125,N_23572,N_24411);
nor U25126 (N_25126,N_23717,N_23620);
xnor U25127 (N_25127,N_23364,N_24278);
xnor U25128 (N_25128,N_22772,N_24021);
nor U25129 (N_25129,N_24446,N_23084);
or U25130 (N_25130,N_23874,N_24251);
nand U25131 (N_25131,N_24778,N_24305);
nor U25132 (N_25132,N_22878,N_22770);
xor U25133 (N_25133,N_24738,N_22773);
or U25134 (N_25134,N_24339,N_24678);
nor U25135 (N_25135,N_22526,N_23530);
xnor U25136 (N_25136,N_23751,N_24849);
or U25137 (N_25137,N_23967,N_24432);
nor U25138 (N_25138,N_23042,N_22699);
or U25139 (N_25139,N_23180,N_24292);
nor U25140 (N_25140,N_24247,N_23275);
nor U25141 (N_25141,N_23497,N_23976);
nor U25142 (N_25142,N_24395,N_24980);
nor U25143 (N_25143,N_22575,N_24886);
nand U25144 (N_25144,N_24671,N_23017);
nor U25145 (N_25145,N_23456,N_24386);
nor U25146 (N_25146,N_23126,N_22671);
or U25147 (N_25147,N_23305,N_23549);
or U25148 (N_25148,N_23299,N_24329);
nand U25149 (N_25149,N_22532,N_23687);
xnor U25150 (N_25150,N_23541,N_23236);
and U25151 (N_25151,N_23800,N_24589);
and U25152 (N_25152,N_23942,N_23469);
nand U25153 (N_25153,N_22795,N_24969);
nand U25154 (N_25154,N_23908,N_23217);
or U25155 (N_25155,N_23796,N_24239);
nand U25156 (N_25156,N_23724,N_23464);
xor U25157 (N_25157,N_24972,N_23132);
nor U25158 (N_25158,N_23256,N_23390);
xor U25159 (N_25159,N_23075,N_24916);
and U25160 (N_25160,N_23928,N_24616);
nor U25161 (N_25161,N_22757,N_24946);
xnor U25162 (N_25162,N_24923,N_23155);
nor U25163 (N_25163,N_24331,N_24230);
or U25164 (N_25164,N_24982,N_23445);
and U25165 (N_25165,N_23583,N_23715);
nor U25166 (N_25166,N_23266,N_23863);
xor U25167 (N_25167,N_22708,N_23416);
or U25168 (N_25168,N_23008,N_24374);
nand U25169 (N_25169,N_23241,N_22804);
nor U25170 (N_25170,N_23035,N_23479);
nand U25171 (N_25171,N_24376,N_22982);
and U25172 (N_25172,N_24023,N_24060);
or U25173 (N_25173,N_23960,N_24574);
nor U25174 (N_25174,N_24534,N_23524);
nor U25175 (N_25175,N_23146,N_24749);
nand U25176 (N_25176,N_23067,N_24123);
nor U25177 (N_25177,N_24856,N_23185);
and U25178 (N_25178,N_23777,N_23955);
and U25179 (N_25179,N_23667,N_22642);
xnor U25180 (N_25180,N_22574,N_24482);
or U25181 (N_25181,N_23454,N_23184);
and U25182 (N_25182,N_22789,N_22709);
nor U25183 (N_25183,N_24554,N_23655);
xor U25184 (N_25184,N_24485,N_23929);
xnor U25185 (N_25185,N_24739,N_22761);
xnor U25186 (N_25186,N_24467,N_24114);
and U25187 (N_25187,N_22625,N_23695);
nand U25188 (N_25188,N_24113,N_24007);
xnor U25189 (N_25189,N_22856,N_24084);
nor U25190 (N_25190,N_23950,N_23357);
or U25191 (N_25191,N_24349,N_24270);
or U25192 (N_25192,N_24235,N_23613);
nor U25193 (N_25193,N_23892,N_24202);
xor U25194 (N_25194,N_24961,N_23872);
xnor U25195 (N_25195,N_24273,N_23521);
nand U25196 (N_25196,N_24801,N_23405);
or U25197 (N_25197,N_24552,N_23755);
nand U25198 (N_25198,N_24909,N_23797);
nor U25199 (N_25199,N_24747,N_24325);
or U25200 (N_25200,N_24122,N_23597);
nor U25201 (N_25201,N_23252,N_23658);
and U25202 (N_25202,N_24197,N_24850);
nor U25203 (N_25203,N_23430,N_23174);
nand U25204 (N_25204,N_22758,N_23813);
xor U25205 (N_25205,N_22750,N_23888);
or U25206 (N_25206,N_23165,N_23385);
nor U25207 (N_25207,N_24795,N_23188);
nor U25208 (N_25208,N_22594,N_24936);
nand U25209 (N_25209,N_22872,N_24188);
or U25210 (N_25210,N_22889,N_22760);
xor U25211 (N_25211,N_22867,N_23199);
or U25212 (N_25212,N_22835,N_23809);
and U25213 (N_25213,N_23832,N_24222);
or U25214 (N_25214,N_23194,N_24931);
nand U25215 (N_25215,N_24364,N_23125);
or U25216 (N_25216,N_24241,N_23588);
nor U25217 (N_25217,N_23720,N_23429);
xnor U25218 (N_25218,N_24492,N_22911);
xor U25219 (N_25219,N_23060,N_23331);
or U25220 (N_25220,N_23859,N_23635);
nand U25221 (N_25221,N_23511,N_24284);
xnor U25222 (N_25222,N_23024,N_22777);
or U25223 (N_25223,N_23335,N_24881);
and U25224 (N_25224,N_23230,N_23632);
nand U25225 (N_25225,N_23555,N_23484);
xnor U25226 (N_25226,N_24429,N_23758);
or U25227 (N_25227,N_24324,N_23738);
or U25228 (N_25228,N_24264,N_23190);
or U25229 (N_25229,N_24934,N_23799);
and U25230 (N_25230,N_23163,N_22860);
nor U25231 (N_25231,N_24870,N_23098);
and U25232 (N_25232,N_24057,N_24887);
nor U25233 (N_25233,N_24956,N_23293);
xnor U25234 (N_25234,N_24562,N_22947);
or U25235 (N_25235,N_22895,N_22893);
xnor U25236 (N_25236,N_24160,N_24153);
and U25237 (N_25237,N_24392,N_22559);
and U25238 (N_25238,N_23659,N_24826);
and U25239 (N_25239,N_23914,N_24725);
or U25240 (N_25240,N_24905,N_23714);
nor U25241 (N_25241,N_23354,N_24419);
xnor U25242 (N_25242,N_24459,N_24187);
nand U25243 (N_25243,N_24425,N_24463);
and U25244 (N_25244,N_22545,N_24269);
or U25245 (N_25245,N_24166,N_22601);
or U25246 (N_25246,N_24137,N_24667);
or U25247 (N_25247,N_24152,N_24149);
nand U25248 (N_25248,N_24775,N_24402);
or U25249 (N_25249,N_23076,N_23240);
and U25250 (N_25250,N_24096,N_23784);
nor U25251 (N_25251,N_23503,N_23923);
nand U25252 (N_25252,N_23852,N_24694);
or U25253 (N_25253,N_23326,N_24848);
and U25254 (N_25254,N_24018,N_24316);
xor U25255 (N_25255,N_23730,N_24640);
or U25256 (N_25256,N_23993,N_23805);
nor U25257 (N_25257,N_22799,N_22808);
nand U25258 (N_25258,N_22595,N_23737);
xor U25259 (N_25259,N_23795,N_24474);
nor U25260 (N_25260,N_23766,N_24192);
xnor U25261 (N_25261,N_24128,N_24687);
nand U25262 (N_25262,N_22548,N_24530);
nand U25263 (N_25263,N_23025,N_23733);
or U25264 (N_25264,N_24479,N_22767);
and U25265 (N_25265,N_22562,N_24340);
xor U25266 (N_25266,N_22800,N_24026);
or U25267 (N_25267,N_23565,N_23297);
nor U25268 (N_25268,N_23333,N_22721);
or U25269 (N_25269,N_24960,N_24896);
and U25270 (N_25270,N_24922,N_24120);
nor U25271 (N_25271,N_23212,N_22729);
nor U25272 (N_25272,N_24103,N_24875);
nor U25273 (N_25273,N_24426,N_24653);
and U25274 (N_25274,N_22775,N_23791);
or U25275 (N_25275,N_22981,N_23587);
or U25276 (N_25276,N_23685,N_23569);
xor U25277 (N_25277,N_24205,N_24974);
xnor U25278 (N_25278,N_23889,N_24127);
xnor U25279 (N_25279,N_23397,N_22948);
nor U25280 (N_25280,N_24508,N_24857);
or U25281 (N_25281,N_23052,N_23666);
xnor U25282 (N_25282,N_23593,N_22612);
and U25283 (N_25283,N_24518,N_22778);
nand U25284 (N_25284,N_22522,N_24603);
nor U25285 (N_25285,N_23003,N_24031);
and U25286 (N_25286,N_23171,N_24825);
or U25287 (N_25287,N_23922,N_23911);
or U25288 (N_25288,N_24469,N_22810);
nor U25289 (N_25289,N_24377,N_24798);
and U25290 (N_25290,N_23356,N_22927);
nor U25291 (N_25291,N_23873,N_23498);
and U25292 (N_25292,N_24836,N_24448);
and U25293 (N_25293,N_24600,N_24617);
and U25294 (N_25294,N_24834,N_22986);
xnor U25295 (N_25295,N_24794,N_23073);
xnor U25296 (N_25296,N_23279,N_23509);
or U25297 (N_25297,N_23843,N_24124);
nand U25298 (N_25298,N_24267,N_23147);
nand U25299 (N_25299,N_24208,N_24303);
nor U25300 (N_25300,N_23886,N_22752);
nor U25301 (N_25301,N_23358,N_22728);
xor U25302 (N_25302,N_24871,N_22882);
or U25303 (N_25303,N_24069,N_23904);
and U25304 (N_25304,N_23441,N_23821);
xnor U25305 (N_25305,N_22565,N_24970);
or U25306 (N_25306,N_24999,N_23679);
xor U25307 (N_25307,N_24983,N_22869);
and U25308 (N_25308,N_23962,N_23550);
nand U25309 (N_25309,N_24657,N_23057);
xor U25310 (N_25310,N_22791,N_23192);
xor U25311 (N_25311,N_22572,N_23007);
and U25312 (N_25312,N_24913,N_24763);
nand U25313 (N_25313,N_24423,N_22838);
xor U25314 (N_25314,N_22711,N_24089);
xnor U25315 (N_25315,N_23696,N_22537);
nor U25316 (N_25316,N_22790,N_23642);
xor U25317 (N_25317,N_22636,N_23881);
nand U25318 (N_25318,N_23118,N_23273);
nor U25319 (N_25319,N_23531,N_24546);
and U25320 (N_25320,N_24175,N_23191);
and U25321 (N_25321,N_22951,N_23462);
nor U25322 (N_25322,N_23901,N_24951);
xor U25323 (N_25323,N_22906,N_24587);
nor U25324 (N_25324,N_22533,N_23491);
xnor U25325 (N_25325,N_23263,N_22714);
nand U25326 (N_25326,N_23924,N_22515);
nand U25327 (N_25327,N_23941,N_24141);
or U25328 (N_25328,N_24664,N_24396);
nand U25329 (N_25329,N_24584,N_24360);
nor U25330 (N_25330,N_24660,N_24373);
and U25331 (N_25331,N_24993,N_23810);
nor U25332 (N_25332,N_24520,N_24154);
nor U25333 (N_25333,N_24078,N_23444);
or U25334 (N_25334,N_23243,N_24680);
xnor U25335 (N_25335,N_23258,N_24874);
nor U25336 (N_25336,N_23480,N_23016);
xnor U25337 (N_25337,N_24381,N_23372);
nand U25338 (N_25338,N_23840,N_23334);
xor U25339 (N_25339,N_23736,N_22934);
and U25340 (N_25340,N_23999,N_22736);
and U25341 (N_25341,N_22753,N_22566);
and U25342 (N_25342,N_23568,N_23223);
xor U25343 (N_25343,N_23085,N_23272);
nand U25344 (N_25344,N_23161,N_24814);
nand U25345 (N_25345,N_23514,N_23548);
and U25346 (N_25346,N_22617,N_23400);
and U25347 (N_25347,N_23222,N_24217);
or U25348 (N_25348,N_23041,N_24254);
or U25349 (N_25349,N_23945,N_24212);
or U25350 (N_25350,N_24788,N_22843);
xor U25351 (N_25351,N_24371,N_22921);
xnor U25352 (N_25352,N_24206,N_23621);
or U25353 (N_25353,N_24008,N_22797);
or U25354 (N_25354,N_23473,N_23854);
and U25355 (N_25355,N_23399,N_24966);
and U25356 (N_25356,N_22820,N_23557);
and U25357 (N_25357,N_22632,N_22591);
and U25358 (N_25358,N_23213,N_23281);
and U25359 (N_25359,N_24585,N_22846);
nor U25360 (N_25360,N_23624,N_24862);
or U25361 (N_25361,N_22655,N_23195);
or U25362 (N_25362,N_23691,N_22637);
and U25363 (N_25363,N_23504,N_24476);
and U25364 (N_25364,N_23238,N_23037);
and U25365 (N_25365,N_22519,N_22501);
or U25366 (N_25366,N_23502,N_23526);
nand U25367 (N_25367,N_24596,N_24721);
or U25368 (N_25368,N_24255,N_24313);
and U25369 (N_25369,N_24178,N_24525);
nor U25370 (N_25370,N_24288,N_23551);
and U25371 (N_25371,N_24358,N_22598);
nor U25372 (N_25372,N_23181,N_23000);
nand U25373 (N_25373,N_22573,N_22504);
xor U25374 (N_25374,N_24714,N_24944);
or U25375 (N_25375,N_23461,N_24318);
xor U25376 (N_25376,N_23939,N_24215);
xor U25377 (N_25377,N_24837,N_23662);
nor U25378 (N_25378,N_24627,N_23319);
and U25379 (N_25379,N_24543,N_22953);
or U25380 (N_25380,N_24176,N_24783);
nor U25381 (N_25381,N_24681,N_23698);
or U25382 (N_25382,N_22684,N_23466);
nand U25383 (N_25383,N_23606,N_24575);
nor U25384 (N_25384,N_22675,N_24382);
nor U25385 (N_25385,N_24428,N_24362);
xnor U25386 (N_25386,N_23819,N_22739);
nor U25387 (N_25387,N_23612,N_24119);
xnor U25388 (N_25388,N_23776,N_23058);
nand U25389 (N_25389,N_24658,N_24894);
nor U25390 (N_25390,N_24702,N_23394);
and U25391 (N_25391,N_23274,N_23646);
xnor U25392 (N_25392,N_23338,N_23261);
and U25393 (N_25393,N_22706,N_23716);
xor U25394 (N_25394,N_23953,N_24491);
nand U25395 (N_25395,N_23833,N_24456);
xnor U25396 (N_25396,N_23794,N_23905);
nand U25397 (N_25397,N_22939,N_24401);
xnor U25398 (N_25398,N_24105,N_23637);
nor U25399 (N_25399,N_23706,N_24051);
nand U25400 (N_25400,N_24865,N_24024);
nor U25401 (N_25401,N_24918,N_23902);
and U25402 (N_25402,N_23267,N_24590);
nor U25403 (N_25403,N_22597,N_24117);
nand U25404 (N_25404,N_23972,N_22914);
or U25405 (N_25405,N_22604,N_23420);
xnor U25406 (N_25406,N_24302,N_24092);
and U25407 (N_25407,N_24258,N_23934);
xnor U25408 (N_25408,N_23887,N_24891);
nor U25409 (N_25409,N_23880,N_24583);
or U25410 (N_25410,N_22936,N_22917);
nand U25411 (N_25411,N_23750,N_23189);
nand U25412 (N_25412,N_23315,N_24935);
or U25413 (N_25413,N_22661,N_23291);
nand U25414 (N_25414,N_23585,N_22521);
or U25415 (N_25415,N_24285,N_24131);
or U25416 (N_25416,N_24743,N_22588);
xor U25417 (N_25417,N_22871,N_23749);
xnor U25418 (N_25418,N_24751,N_23773);
nand U25419 (N_25419,N_24252,N_24387);
xor U25420 (N_25420,N_24760,N_23158);
xnor U25421 (N_25421,N_24740,N_24319);
or U25422 (N_25422,N_22904,N_24514);
xor U25423 (N_25423,N_24296,N_23176);
nand U25424 (N_25424,N_23701,N_24689);
nand U25425 (N_25425,N_23292,N_24706);
nor U25426 (N_25426,N_22932,N_23242);
nor U25427 (N_25427,N_24771,N_23801);
or U25428 (N_25428,N_24659,N_22664);
xor U25429 (N_25429,N_23671,N_23753);
and U25430 (N_25430,N_23847,N_24977);
nor U25431 (N_25431,N_24607,N_24772);
nand U25432 (N_25432,N_23975,N_24785);
and U25433 (N_25433,N_24654,N_24967);
xor U25434 (N_25434,N_23981,N_23481);
and U25435 (N_25435,N_24496,N_24244);
xnor U25436 (N_25436,N_24139,N_23065);
or U25437 (N_25437,N_22512,N_23139);
xnor U25438 (N_25438,N_24637,N_23861);
nand U25439 (N_25439,N_23536,N_24676);
nand U25440 (N_25440,N_23131,N_23907);
nand U25441 (N_25441,N_23307,N_24758);
nand U25442 (N_25442,N_23496,N_23183);
and U25443 (N_25443,N_23079,N_24422);
or U25444 (N_25444,N_24790,N_22568);
or U25445 (N_25445,N_23965,N_23247);
or U25446 (N_25446,N_24953,N_24348);
or U25447 (N_25447,N_24489,N_22590);
xnor U25448 (N_25448,N_24614,N_23652);
or U25449 (N_25449,N_23792,N_24201);
nand U25450 (N_25450,N_24522,N_22987);
nand U25451 (N_25451,N_23362,N_22901);
xor U25452 (N_25452,N_24049,N_24326);
or U25453 (N_25453,N_23412,N_22765);
nor U25454 (N_25454,N_23170,N_23709);
nand U25455 (N_25455,N_22570,N_23560);
and U25456 (N_25456,N_23558,N_24723);
xor U25457 (N_25457,N_23943,N_24473);
and U25458 (N_25458,N_24962,N_22653);
nor U25459 (N_25459,N_23398,N_24440);
xnor U25460 (N_25460,N_23211,N_22896);
or U25461 (N_25461,N_24805,N_24196);
nor U25462 (N_25462,N_22696,N_24907);
nor U25463 (N_25463,N_24538,N_24777);
and U25464 (N_25464,N_24890,N_22621);
nand U25465 (N_25465,N_24332,N_23517);
and U25466 (N_25466,N_24151,N_23070);
nand U25467 (N_25467,N_23725,N_22756);
or U25468 (N_25468,N_22755,N_23734);
nand U25469 (N_25469,N_23692,N_23301);
and U25470 (N_25470,N_24355,N_23712);
nand U25471 (N_25471,N_24877,N_23601);
and U25472 (N_25472,N_23543,N_24892);
nor U25473 (N_25473,N_23327,N_23106);
nand U25474 (N_25474,N_24115,N_23012);
and U25475 (N_25475,N_22841,N_23564);
and U25476 (N_25476,N_24718,N_24417);
xnor U25477 (N_25477,N_23493,N_23022);
xor U25478 (N_25478,N_24304,N_24350);
nand U25479 (N_25479,N_24665,N_24356);
xnor U25480 (N_25480,N_24579,N_24056);
or U25481 (N_25481,N_24431,N_24879);
or U25482 (N_25482,N_24820,N_23650);
and U25483 (N_25483,N_23823,N_23721);
xor U25484 (N_25484,N_24949,N_22918);
xor U25485 (N_25485,N_24483,N_23231);
xnor U25486 (N_25486,N_22801,N_23997);
nand U25487 (N_25487,N_24793,N_23726);
and U25488 (N_25488,N_23244,N_22546);
or U25489 (N_25489,N_24162,N_23618);
nor U25490 (N_25490,N_23136,N_24634);
nor U25491 (N_25491,N_22610,N_23596);
or U25492 (N_25492,N_23451,N_24142);
nand U25493 (N_25493,N_22520,N_23677);
and U25494 (N_25494,N_23878,N_24321);
xor U25495 (N_25495,N_24744,N_24441);
or U25496 (N_25496,N_22746,N_24495);
and U25497 (N_25497,N_23144,N_23693);
nor U25498 (N_25498,N_22876,N_22967);
and U25499 (N_25499,N_22707,N_24502);
nand U25500 (N_25500,N_24073,N_24540);
nand U25501 (N_25501,N_24121,N_24911);
or U25502 (N_25502,N_22603,N_24271);
nor U25503 (N_25503,N_23875,N_24864);
or U25504 (N_25504,N_23903,N_24730);
and U25505 (N_25505,N_24047,N_24941);
or U25506 (N_25506,N_22989,N_23463);
and U25507 (N_25507,N_24352,N_23657);
nand U25508 (N_25508,N_23378,N_22759);
or U25509 (N_25509,N_22766,N_24833);
xnor U25510 (N_25510,N_23109,N_24389);
xnor U25511 (N_25511,N_23336,N_23255);
nor U25512 (N_25512,N_24034,N_22928);
nand U25513 (N_25513,N_23694,N_24578);
and U25514 (N_25514,N_23018,N_22500);
xnor U25515 (N_25515,N_24404,N_23913);
nor U25516 (N_25516,N_23961,N_22599);
xnor U25517 (N_25517,N_24802,N_22865);
xnor U25518 (N_25518,N_22887,N_23739);
nand U25519 (N_25519,N_23160,N_23537);
nor U25520 (N_25520,N_23330,N_24858);
nor U25521 (N_25521,N_22624,N_24573);
and U25522 (N_25522,N_24253,N_23916);
and U25523 (N_25523,N_22718,N_24301);
nand U25524 (N_25524,N_24365,N_22535);
and U25525 (N_25525,N_22674,N_23081);
nand U25526 (N_25526,N_22830,N_24475);
nor U25527 (N_25527,N_22949,N_23825);
and U25528 (N_25528,N_23628,N_23019);
nand U25529 (N_25529,N_24037,N_23234);
xor U25530 (N_25530,N_24182,N_23425);
xnor U25531 (N_25531,N_24869,N_23957);
nand U25532 (N_25532,N_24104,N_23539);
and U25533 (N_25533,N_24263,N_24385);
nand U25534 (N_25534,N_22958,N_22880);
xnor U25535 (N_25535,N_23450,N_24899);
or U25536 (N_25536,N_24560,N_23415);
and U25537 (N_25537,N_24405,N_24803);
nand U25538 (N_25538,N_23029,N_23651);
and U25539 (N_25539,N_24011,N_24630);
nand U25540 (N_25540,N_23756,N_22503);
or U25541 (N_25541,N_24580,N_22513);
nand U25542 (N_25542,N_22724,N_22861);
nand U25543 (N_25543,N_23681,N_24985);
xor U25544 (N_25544,N_22596,N_22669);
or U25545 (N_25545,N_24391,N_22993);
xnor U25546 (N_25546,N_24237,N_24409);
nor U25547 (N_25547,N_23439,N_22748);
or U25548 (N_25548,N_24866,N_22933);
and U25549 (N_25549,N_23178,N_22528);
or U25550 (N_25550,N_23968,N_24808);
or U25551 (N_25551,N_22997,N_23912);
and U25552 (N_25552,N_23457,N_24062);
xor U25553 (N_25553,N_24418,N_22960);
xnor U25554 (N_25554,N_23990,N_22740);
nor U25555 (N_25555,N_24861,N_23748);
or U25556 (N_25556,N_22805,N_23202);
xnor U25557 (N_25557,N_24091,N_24261);
or U25558 (N_25558,N_24298,N_24499);
xor U25559 (N_25559,N_22938,N_24286);
nand U25560 (N_25560,N_22681,N_22780);
or U25561 (N_25561,N_24082,N_22553);
or U25562 (N_25562,N_24832,N_23864);
nand U25563 (N_25563,N_23489,N_22980);
xor U25564 (N_25564,N_22821,N_23046);
xnor U25565 (N_25565,N_23542,N_24629);
xor U25566 (N_25566,N_23159,N_24184);
or U25567 (N_25567,N_24029,N_22550);
or U25568 (N_25568,N_24965,N_24240);
and U25569 (N_25569,N_23032,N_24524);
and U25570 (N_25570,N_24752,N_22502);
xor U25571 (N_25571,N_24478,N_23009);
and U25572 (N_25572,N_22909,N_24544);
nand U25573 (N_25573,N_24080,N_24888);
xnor U25574 (N_25574,N_24529,N_23452);
xor U25575 (N_25575,N_23604,N_22822);
xnor U25576 (N_25576,N_23232,N_24919);
or U25577 (N_25577,N_22839,N_22965);
and U25578 (N_25578,N_23237,N_22689);
nor U25579 (N_25579,N_23320,N_23446);
nor U25580 (N_25580,N_23152,N_22516);
and U25581 (N_25581,N_23296,N_23278);
nand U25582 (N_25582,N_24755,N_22639);
nor U25583 (N_25583,N_24842,N_23674);
or U25584 (N_25584,N_23954,N_23586);
xnor U25585 (N_25585,N_22648,N_23783);
and U25586 (N_25586,N_23533,N_24322);
nand U25587 (N_25587,N_23219,N_23063);
xor U25588 (N_25588,N_24500,N_23527);
nand U25589 (N_25589,N_24390,N_24077);
xnor U25590 (N_25590,N_23608,N_24821);
nor U25591 (N_25591,N_23221,N_23759);
nand U25592 (N_25592,N_24171,N_24236);
xor U25593 (N_25593,N_22995,N_23949);
nand U25594 (N_25594,N_23404,N_23200);
and U25595 (N_25595,N_24207,N_23808);
or U25596 (N_25596,N_24380,N_24939);
xnor U25597 (N_25597,N_22956,N_23918);
xnor U25598 (N_25598,N_24351,N_24148);
and U25599 (N_25599,N_24532,N_22623);
nand U25600 (N_25600,N_23249,N_23002);
or U25601 (N_25601,N_24968,N_24260);
or U25602 (N_25602,N_24734,N_22673);
or U25603 (N_25603,N_23468,N_24761);
and U25604 (N_25604,N_23253,N_24609);
and U25605 (N_25605,N_24827,N_24006);
xor U25606 (N_25606,N_24526,N_23952);
xor U25607 (N_25607,N_23595,N_24822);
nand U25608 (N_25608,N_22813,N_24219);
or U25609 (N_25609,N_24097,N_24564);
nand U25610 (N_25610,N_24238,N_23765);
or U25611 (N_25611,N_22905,N_24576);
xnor U25612 (N_25612,N_22920,N_24277);
and U25613 (N_25613,N_22552,N_22605);
or U25614 (N_25614,N_24581,N_24780);
and U25615 (N_25615,N_23111,N_23707);
and U25616 (N_25616,N_24354,N_23971);
or U25617 (N_25617,N_23359,N_22607);
and U25618 (N_25618,N_23006,N_23660);
and U25619 (N_25619,N_23494,N_24731);
xor U25620 (N_25620,N_24135,N_24547);
and U25621 (N_25621,N_24975,N_22735);
nor U25622 (N_25622,N_23844,N_22666);
xnor U25623 (N_25623,N_23014,N_22734);
and U25624 (N_25624,N_24159,N_23935);
xor U25625 (N_25625,N_24100,N_24845);
xnor U25626 (N_25626,N_24636,N_24943);
nor U25627 (N_25627,N_22716,N_22635);
and U25628 (N_25628,N_24551,N_24071);
xnor U25629 (N_25629,N_24306,N_22660);
nand U25630 (N_25630,N_24531,N_23561);
nand U25631 (N_25631,N_24052,N_23216);
or U25632 (N_25632,N_23103,N_24204);
nor U25633 (N_25633,N_22629,N_22923);
nor U25634 (N_25634,N_24792,N_22690);
xor U25635 (N_25635,N_22964,N_24199);
or U25636 (N_25636,N_24789,N_24335);
nand U25637 (N_25637,N_22640,N_23314);
or U25638 (N_25638,N_24523,N_24156);
nand U25639 (N_25639,N_24639,N_24186);
and U25640 (N_25640,N_22634,N_24180);
nor U25641 (N_25641,N_24901,N_23814);
nor U25642 (N_25642,N_23360,N_22705);
nor U25643 (N_25643,N_23043,N_24791);
nand U25644 (N_25644,N_24841,N_23811);
nor U25645 (N_25645,N_23337,N_23036);
nor U25646 (N_25646,N_23495,N_24797);
or U25647 (N_25647,N_22730,N_22606);
and U25648 (N_25648,N_24406,N_23686);
xor U25649 (N_25649,N_24484,N_24895);
and U25650 (N_25650,N_24311,N_22762);
nor U25651 (N_25651,N_24372,N_24509);
nand U25652 (N_25652,N_23309,N_24628);
nor U25653 (N_25653,N_24109,N_22754);
nor U25654 (N_25654,N_23731,N_24729);
or U25655 (N_25655,N_22683,N_23828);
or U25656 (N_25656,N_24612,N_23640);
or U25657 (N_25657,N_24602,N_23787);
xor U25658 (N_25658,N_23026,N_22833);
nand U25659 (N_25659,N_23930,N_23702);
and U25660 (N_25660,N_24809,N_24439);
or U25661 (N_25661,N_22798,N_23259);
nand U25662 (N_25662,N_22691,N_22983);
or U25663 (N_25663,N_24274,N_24558);
xor U25664 (N_25664,N_24548,N_24976);
or U25665 (N_25665,N_24289,N_24625);
nand U25666 (N_25666,N_23529,N_23944);
xnor U25667 (N_25667,N_22998,N_24606);
nand U25668 (N_25668,N_24921,N_24450);
and U25669 (N_25669,N_24415,N_22658);
and U25670 (N_25670,N_23317,N_24661);
xor U25671 (N_25671,N_22886,N_23853);
nand U25672 (N_25672,N_22514,N_23592);
nor U25673 (N_25673,N_22589,N_24028);
xor U25674 (N_25674,N_22955,N_24133);
or U25675 (N_25675,N_23027,N_24649);
xnor U25676 (N_25676,N_23102,N_23431);
nand U25677 (N_25677,N_24799,N_24420);
nand U25678 (N_25678,N_22628,N_24915);
or U25679 (N_25679,N_23321,N_22667);
and U25680 (N_25680,N_24621,N_24712);
nor U25681 (N_25681,N_24810,N_22643);
or U25682 (N_25682,N_23141,N_24668);
nand U25683 (N_25683,N_23781,N_23417);
or U25684 (N_25684,N_24282,N_22733);
or U25685 (N_25685,N_24908,N_23406);
and U25686 (N_25686,N_24177,N_23987);
xnor U25687 (N_25687,N_23407,N_23028);
xor U25688 (N_25688,N_22582,N_24880);
and U25689 (N_25689,N_24605,N_24672);
and U25690 (N_25690,N_23806,N_24727);
nand U25691 (N_25691,N_23678,N_24917);
nor U25692 (N_25692,N_23154,N_24193);
xor U25693 (N_25693,N_23798,N_22783);
nor U25694 (N_25694,N_23156,N_23838);
or U25695 (N_25695,N_23104,N_24161);
nor U25696 (N_25696,N_24710,N_23817);
or U25697 (N_25697,N_23442,N_23500);
or U25698 (N_25698,N_24806,N_23276);
nand U25699 (N_25699,N_24214,N_23713);
and U25700 (N_25700,N_24677,N_22881);
or U25701 (N_25701,N_24228,N_23193);
or U25702 (N_25702,N_23077,N_24598);
nor U25703 (N_25703,N_23704,N_24736);
or U25704 (N_25704,N_24198,N_23785);
and U25705 (N_25705,N_22903,N_24327);
and U25706 (N_25706,N_22609,N_22732);
and U25707 (N_25707,N_24599,N_22935);
nand U25708 (N_25708,N_24674,N_24597);
and U25709 (N_25709,N_22952,N_23963);
or U25710 (N_25710,N_24622,N_23994);
nor U25711 (N_25711,N_22557,N_24945);
and U25712 (N_25712,N_23054,N_23580);
xnor U25713 (N_25713,N_23689,N_24948);
and U25714 (N_25714,N_23927,N_24424);
nor U25715 (N_25715,N_23988,N_23906);
nand U25716 (N_25716,N_23804,N_24231);
nor U25717 (N_25717,N_23332,N_23850);
and U25718 (N_25718,N_23921,N_23270);
nor U25719 (N_25719,N_24618,N_23563);
and U25720 (N_25720,N_24663,N_24209);
nand U25721 (N_25721,N_24717,N_23123);
nand U25722 (N_25722,N_24754,N_22826);
nand U25723 (N_25723,N_23757,N_24984);
and U25724 (N_25724,N_22710,N_23841);
nor U25725 (N_25725,N_23470,N_24112);
nand U25726 (N_25726,N_24582,N_23680);
nand U25727 (N_25727,N_22832,N_23345);
nand U25728 (N_25728,N_23883,N_24724);
or U25729 (N_25729,N_24090,N_22563);
xnor U25730 (N_25730,N_24817,N_24566);
and U25731 (N_25731,N_22919,N_23708);
nor U25732 (N_25732,N_24695,N_23728);
nand U25733 (N_25733,N_23735,N_22857);
and U25734 (N_25734,N_24859,N_23617);
xnor U25735 (N_25735,N_22823,N_24025);
nor U25736 (N_25736,N_23984,N_24748);
and U25737 (N_25737,N_22898,N_22579);
nand U25738 (N_25738,N_22942,N_24505);
nor U25739 (N_25739,N_24644,N_22659);
nand U25740 (N_25740,N_24146,N_22985);
nand U25741 (N_25741,N_24604,N_23534);
nor U25742 (N_25742,N_23631,N_23786);
or U25743 (N_25743,N_23031,N_22644);
nor U25744 (N_25744,N_24086,N_22807);
nor U25745 (N_25745,N_24824,N_23262);
xnor U25746 (N_25746,N_22973,N_23508);
nor U25747 (N_25747,N_24067,N_24435);
xnor U25748 (N_25748,N_23867,N_22827);
or U25749 (N_25749,N_23204,N_24682);
and U25750 (N_25750,N_23030,N_22910);
nor U25751 (N_25751,N_24087,N_24705);
nand U25752 (N_25752,N_24537,N_24140);
xnor U25753 (N_25753,N_22968,N_24094);
or U25754 (N_25754,N_23047,N_24320);
nand U25755 (N_25755,N_24134,N_23520);
nor U25756 (N_25756,N_22633,N_24453);
nor U25757 (N_25757,N_23233,N_23422);
and U25758 (N_25758,N_23937,N_22694);
and U25759 (N_25759,N_23582,N_23664);
nor U25760 (N_25760,N_24796,N_23167);
nand U25761 (N_25761,N_22862,N_24130);
and U25762 (N_25762,N_24926,N_22852);
nor U25763 (N_25763,N_24698,N_23313);
nand U25764 (N_25764,N_24224,N_22567);
nand U25765 (N_25765,N_22558,N_23096);
xor U25766 (N_25766,N_24075,N_24517);
nor U25767 (N_25767,N_23129,N_24550);
or U25768 (N_25768,N_24129,N_23361);
or U25769 (N_25769,N_23478,N_24272);
xor U25770 (N_25770,N_24876,N_23207);
nor U25771 (N_25771,N_23829,N_24126);
nor U25772 (N_25772,N_24317,N_23615);
nor U25773 (N_25773,N_23866,N_22586);
nor U25774 (N_25774,N_24457,N_23166);
xor U25775 (N_25775,N_23501,N_24081);
xor U25776 (N_25776,N_22925,N_24013);
xnor U25777 (N_25777,N_24720,N_23289);
xnor U25778 (N_25778,N_23339,N_23251);
nand U25779 (N_25779,N_23705,N_24957);
and U25780 (N_25780,N_23623,N_22723);
or U25781 (N_25781,N_24713,N_23377);
nor U25782 (N_25782,N_23826,N_23512);
and U25783 (N_25783,N_23625,N_22627);
or U25784 (N_25784,N_23996,N_24375);
nor U25785 (N_25785,N_24163,N_24964);
and U25786 (N_25786,N_23438,N_24998);
or U25787 (N_25787,N_24737,N_23304);
xor U25788 (N_25788,N_22715,N_24992);
xnor U25789 (N_25789,N_23409,N_24940);
and U25790 (N_25790,N_22771,N_23931);
and U25791 (N_25791,N_24733,N_22650);
xor U25792 (N_25792,N_24623,N_23575);
or U25793 (N_25793,N_23072,N_23600);
xnor U25794 (N_25794,N_24035,N_22940);
xor U25795 (N_25795,N_24398,N_24571);
xor U25796 (N_25796,N_22619,N_24414);
or U25797 (N_25797,N_24692,N_22806);
xor U25798 (N_25798,N_24064,N_23856);
nand U25799 (N_25799,N_24281,N_23284);
xnor U25800 (N_25800,N_24268,N_22688);
xnor U25801 (N_25801,N_24044,N_24924);
and U25802 (N_25802,N_24040,N_23168);
nand U25803 (N_25803,N_24632,N_23893);
and U25804 (N_25804,N_24189,N_23062);
nor U25805 (N_25805,N_23396,N_24027);
nor U25806 (N_25806,N_23460,N_22631);
or U25807 (N_25807,N_24416,N_23956);
xnor U25808 (N_25808,N_22787,N_24882);
nor U25809 (N_25809,N_24242,N_24521);
nand U25810 (N_25810,N_23959,N_24883);
and U25811 (N_25811,N_24297,N_22970);
xnor U25812 (N_25812,N_24511,N_24732);
or U25813 (N_25813,N_24334,N_22908);
nor U25814 (N_25814,N_22929,N_24932);
nand U25815 (N_25815,N_24536,N_23021);
and U25816 (N_25816,N_22701,N_23641);
and U25817 (N_25817,N_23910,N_24050);
nand U25818 (N_25818,N_22816,N_24342);
nor U25819 (N_25819,N_23611,N_22577);
nor U25820 (N_25820,N_24002,N_22600);
or U25821 (N_25821,N_22877,N_24572);
nand U25822 (N_25822,N_24914,N_22864);
nor U25823 (N_25823,N_24378,N_24541);
nor U25824 (N_25824,N_23419,N_24686);
nand U25825 (N_25825,N_23381,N_23577);
and U25826 (N_25826,N_24703,N_22850);
nor U25827 (N_25827,N_24225,N_22560);
or U25828 (N_25828,N_23347,N_23124);
nand U25829 (N_25829,N_24642,N_23120);
nand U25830 (N_25830,N_22680,N_23745);
and U25831 (N_25831,N_22966,N_24746);
xnor U25832 (N_25832,N_23837,N_24800);
and U25833 (N_25833,N_24245,N_22616);
nor U25834 (N_25834,N_22916,N_24157);
nand U25835 (N_25835,N_23353,N_24098);
xnor U25836 (N_25836,N_22972,N_24647);
or U25837 (N_25837,N_23522,N_22615);
nand U25838 (N_25838,N_22538,N_24344);
and U25839 (N_25839,N_23023,N_22645);
xor U25840 (N_25840,N_24211,N_22863);
nor U25841 (N_25841,N_23506,N_22763);
and U25842 (N_25842,N_22581,N_22541);
or U25843 (N_25843,N_24904,N_24635);
and U25844 (N_25844,N_23428,N_22979);
xnor U25845 (N_25845,N_24294,N_23435);
nand U25846 (N_25846,N_24181,N_24144);
nor U25847 (N_25847,N_22890,N_23218);
xor U25848 (N_25848,N_23834,N_23771);
nand U25849 (N_25849,N_23896,N_22764);
nand U25850 (N_25850,N_22555,N_24183);
xnor U25851 (N_25851,N_22779,N_23898);
xor U25852 (N_25852,N_22879,N_23114);
xnor U25853 (N_25853,N_23769,N_23727);
and U25854 (N_25854,N_24400,N_23351);
xnor U25855 (N_25855,N_22587,N_23768);
or U25856 (N_25856,N_24000,N_24643);
and U25857 (N_25857,N_24055,N_24168);
nand U25858 (N_25858,N_23567,N_24952);
nand U25859 (N_25859,N_24910,N_23117);
nand U25860 (N_25860,N_22990,N_23562);
or U25861 (N_25861,N_24010,N_23590);
nor U25862 (N_25862,N_22819,N_22853);
xor U25863 (N_25863,N_24611,N_24937);
xor U25864 (N_25864,N_23644,N_24045);
and U25865 (N_25865,N_23040,N_23350);
or U25866 (N_25866,N_23780,N_24515);
nor U25867 (N_25867,N_22510,N_22902);
and U25868 (N_25868,N_23926,N_23048);
and U25869 (N_25869,N_22663,N_24107);
or U25870 (N_25870,N_23089,N_24093);
xor U25871 (N_25871,N_23605,N_23352);
or U25872 (N_25872,N_23492,N_22662);
xor U25873 (N_25873,N_23647,N_24226);
nand U25874 (N_25874,N_24393,N_24675);
nand U25875 (N_25875,N_23064,N_24567);
and U25876 (N_25876,N_24897,N_24700);
nor U25877 (N_25877,N_24345,N_23410);
nand U25878 (N_25878,N_23775,N_24170);
nor U25879 (N_25879,N_23105,N_23818);
xnor U25880 (N_25880,N_23328,N_23349);
xnor U25881 (N_25881,N_23426,N_23271);
xor U25882 (N_25882,N_23162,N_23602);
and U25883 (N_25883,N_24004,N_24701);
and U25884 (N_25884,N_22961,N_23835);
and U25885 (N_25885,N_22695,N_24449);
and U25886 (N_25886,N_23039,N_24079);
nor U25887 (N_25887,N_23969,N_23148);
xor U25888 (N_25888,N_24807,N_24844);
nand U25889 (N_25889,N_22749,N_24594);
xor U25890 (N_25890,N_24383,N_24195);
nand U25891 (N_25891,N_24262,N_24835);
xor U25892 (N_25892,N_24336,N_23225);
and U25893 (N_25893,N_24601,N_24959);
xnor U25894 (N_25894,N_22894,N_22945);
nand U25895 (N_25895,N_23329,N_23983);
nor U25896 (N_25896,N_24549,N_24179);
xor U25897 (N_25897,N_24781,N_24735);
nand U25898 (N_25898,N_23340,N_22569);
xor U25899 (N_25899,N_23214,N_24981);
and U25900 (N_25900,N_22969,N_23760);
xor U25901 (N_25901,N_24408,N_22551);
nand U25902 (N_25902,N_23487,N_24503);
and U25903 (N_25903,N_23599,N_24454);
nand U25904 (N_25904,N_23820,N_23220);
xor U25905 (N_25905,N_24929,N_23711);
nand U25906 (N_25906,N_24645,N_24847);
nor U25907 (N_25907,N_23732,N_23055);
or U25908 (N_25908,N_23387,N_23286);
and U25909 (N_25909,N_24480,N_23895);
and U25910 (N_25910,N_24828,N_23703);
and U25911 (N_25911,N_24756,N_23175);
nor U25912 (N_25912,N_23839,N_23483);
nand U25913 (N_25913,N_23566,N_23803);
and U25914 (N_25914,N_24762,N_23363);
or U25915 (N_25915,N_23239,N_24693);
and U25916 (N_25916,N_24369,N_22897);
or U25917 (N_25917,N_24994,N_22682);
nand U25918 (N_25918,N_24065,N_22542);
xor U25919 (N_25919,N_23298,N_22988);
nand U25920 (N_25920,N_22786,N_23951);
xnor U25921 (N_25921,N_23157,N_24003);
and U25922 (N_25922,N_23633,N_24072);
xnor U25923 (N_25923,N_24058,N_24266);
and U25924 (N_25924,N_23964,N_22737);
and U25925 (N_25925,N_24276,N_24669);
nand U25926 (N_25926,N_22725,N_23177);
or U25927 (N_25927,N_22847,N_24246);
xor U25928 (N_25928,N_24779,N_23245);
or U25929 (N_25929,N_23970,N_23589);
nand U25930 (N_25930,N_23164,N_24046);
nor U25931 (N_25931,N_24586,N_22868);
nand U25932 (N_25932,N_23851,N_23122);
and U25933 (N_25933,N_22676,N_24893);
nand U25934 (N_25934,N_22618,N_22668);
and U25935 (N_25935,N_22829,N_23443);
and U25936 (N_25936,N_23061,N_24885);
and U25937 (N_25937,N_22525,N_24545);
or U25938 (N_25938,N_22529,N_24315);
and U25939 (N_25939,N_24059,N_23802);
nor U25940 (N_25940,N_24819,N_22564);
xnor U25941 (N_25941,N_24265,N_22527);
nor U25942 (N_25942,N_24218,N_22745);
and U25943 (N_25943,N_23205,N_24155);
nor U25944 (N_25944,N_23486,N_22999);
nand U25945 (N_25945,N_24333,N_23308);
or U25946 (N_25946,N_24243,N_23090);
nand U25947 (N_25947,N_23145,N_24118);
nand U25948 (N_25948,N_23312,N_22738);
xor U25949 (N_25949,N_23290,N_24314);
nor U25950 (N_25950,N_22554,N_24053);
or U25951 (N_25951,N_22854,N_23068);
xnor U25952 (N_25952,N_24036,N_23778);
and U25953 (N_25953,N_23318,N_22656);
xor U25954 (N_25954,N_22647,N_22509);
xnor U25955 (N_25955,N_24978,N_23143);
or U25956 (N_25956,N_24257,N_23812);
nor U25957 (N_25957,N_22803,N_23433);
and U25958 (N_25958,N_23697,N_23598);
nor U25959 (N_25959,N_24591,N_23661);
or U25960 (N_25960,N_24839,N_23283);
nor U25961 (N_25961,N_23112,N_23909);
xor U25962 (N_25962,N_24210,N_24468);
nor U25963 (N_25963,N_22505,N_24816);
xor U25964 (N_25964,N_24384,N_23858);
and U25965 (N_25965,N_24770,N_22922);
nor U25966 (N_25966,N_22549,N_24070);
nor U25967 (N_25967,N_24290,N_24308);
nand U25968 (N_25968,N_24460,N_22620);
and U25969 (N_25969,N_24493,N_24213);
and U25970 (N_25970,N_24111,N_22994);
nand U25971 (N_25971,N_24346,N_23300);
xor U25972 (N_25972,N_23172,N_24147);
or U25973 (N_25973,N_23523,N_24641);
and U25974 (N_25974,N_23346,N_23824);
nor U25975 (N_25975,N_22828,N_24279);
nor U25976 (N_25976,N_24403,N_24465);
or U25977 (N_25977,N_22698,N_23447);
xnor U25978 (N_25978,N_24132,N_22900);
nand U25979 (N_25979,N_23919,N_24811);
or U25980 (N_25980,N_23116,N_24742);
nand U25981 (N_25981,N_23374,N_22507);
xnor U25982 (N_25982,N_22731,N_24519);
or U25983 (N_25983,N_23643,N_23226);
nand U25984 (N_25984,N_24997,N_24652);
nand U25985 (N_25985,N_22976,N_24259);
or U25986 (N_25986,N_23488,N_23306);
or U25987 (N_25987,N_24019,N_22802);
and U25988 (N_25988,N_22702,N_22792);
xnor U25989 (N_25989,N_22844,N_24221);
nor U25990 (N_25990,N_24076,N_23966);
and U25991 (N_25991,N_24136,N_22851);
and U25992 (N_25992,N_23719,N_23389);
nor U25993 (N_25993,N_24906,N_24216);
nand U25994 (N_25994,N_24776,N_22576);
or U25995 (N_25995,N_24248,N_22837);
or U25996 (N_25996,N_23684,N_24359);
and U25997 (N_25997,N_23538,N_24535);
nor U25998 (N_25998,N_23885,N_24172);
or U25999 (N_25999,N_23295,N_23010);
or U26000 (N_26000,N_22544,N_23173);
nor U26001 (N_26001,N_23848,N_24095);
nand U26002 (N_26002,N_23545,N_22840);
or U26003 (N_26003,N_23379,N_23449);
xor U26004 (N_26004,N_23663,N_23392);
or U26005 (N_26005,N_24988,N_23594);
and U26006 (N_26006,N_24283,N_22592);
and U26007 (N_26007,N_23130,N_24341);
nand U26008 (N_26008,N_23087,N_24872);
or U26009 (N_26009,N_24728,N_23700);
nand U26010 (N_26010,N_23138,N_24173);
nor U26011 (N_26011,N_24068,N_24041);
xor U26012 (N_26012,N_22611,N_22626);
nor U26013 (N_26013,N_24220,N_24624);
nor U26014 (N_26014,N_24555,N_23150);
nand U26015 (N_26015,N_24662,N_24430);
nor U26016 (N_26016,N_23051,N_23038);
and U26017 (N_26017,N_24707,N_23467);
nand U26018 (N_26018,N_24108,N_24950);
and U26019 (N_26019,N_23197,N_23083);
nand U26020 (N_26020,N_23206,N_23553);
nor U26021 (N_26021,N_23857,N_23059);
and U26022 (N_26022,N_24765,N_22679);
xnor U26023 (N_26023,N_24299,N_23424);
or U26024 (N_26024,N_24164,N_23869);
or U26025 (N_26025,N_24631,N_24223);
xnor U26026 (N_26026,N_23722,N_24759);
nor U26027 (N_26027,N_24928,N_22531);
nand U26028 (N_26028,N_24256,N_24513);
or U26029 (N_26029,N_23614,N_24610);
or U26030 (N_26030,N_23455,N_24741);
and U26031 (N_26031,N_23762,N_23936);
and U26032 (N_26032,N_24438,N_24504);
and U26033 (N_26033,N_23229,N_23656);
and U26034 (N_26034,N_22722,N_23302);
or U26035 (N_26035,N_23584,N_24307);
nor U26036 (N_26036,N_23532,N_23897);
or U26037 (N_26037,N_23187,N_24437);
xor U26038 (N_26038,N_24413,N_22543);
xnor U26039 (N_26039,N_23393,N_23050);
or U26040 (N_26040,N_24958,N_23752);
xnor U26041 (N_26041,N_23285,N_22873);
nand U26042 (N_26042,N_24200,N_22888);
and U26043 (N_26043,N_23636,N_24388);
nand U26044 (N_26044,N_23369,N_24249);
nor U26045 (N_26045,N_23790,N_23228);
nor U26046 (N_26046,N_23603,N_24039);
and U26047 (N_26047,N_23215,N_24232);
or U26048 (N_26048,N_24234,N_24568);
xnor U26049 (N_26049,N_22815,N_23472);
nand U26050 (N_26050,N_24407,N_24898);
xor U26051 (N_26051,N_22975,N_23436);
nand U26052 (N_26052,N_23427,N_24830);
xor U26053 (N_26053,N_24542,N_23134);
nand U26054 (N_26054,N_24497,N_23499);
and U26055 (N_26055,N_23980,N_23260);
xor U26056 (N_26056,N_23280,N_24410);
or U26057 (N_26057,N_23978,N_23303);
or U26058 (N_26058,N_22524,N_23413);
or U26059 (N_26059,N_24020,N_22742);
xnor U26060 (N_26060,N_24063,N_23287);
nor U26061 (N_26061,N_24032,N_24716);
or U26062 (N_26062,N_22511,N_23900);
nor U26063 (N_26063,N_23591,N_23421);
or U26064 (N_26064,N_23940,N_22992);
nor U26065 (N_26065,N_22580,N_24995);
or U26066 (N_26066,N_23482,N_24648);
and U26067 (N_26067,N_24347,N_24048);
nor U26068 (N_26068,N_23179,N_22785);
and U26069 (N_26069,N_23877,N_24900);
or U26070 (N_26070,N_23201,N_22859);
xor U26071 (N_26071,N_24275,N_24427);
and U26072 (N_26072,N_22954,N_22899);
nand U26073 (N_26073,N_23344,N_22687);
nor U26074 (N_26074,N_23973,N_24361);
xor U26075 (N_26075,N_24507,N_22824);
nor U26076 (N_26076,N_22654,N_22818);
nand U26077 (N_26077,N_23376,N_23384);
or U26078 (N_26078,N_23186,N_23348);
xnor U26079 (N_26079,N_23836,N_23699);
and U26080 (N_26080,N_23322,N_24330);
and U26081 (N_26081,N_24227,N_24533);
xnor U26082 (N_26082,N_24293,N_23868);
nor U26083 (N_26083,N_23948,N_23894);
xnor U26084 (N_26084,N_24709,N_23474);
nor U26085 (N_26085,N_23610,N_24954);
xnor U26086 (N_26086,N_23133,N_22585);
and U26087 (N_26087,N_24884,N_23011);
xnor U26088 (N_26088,N_24421,N_24501);
nand U26089 (N_26089,N_23989,N_22713);
and U26090 (N_26090,N_23277,N_22593);
or U26091 (N_26091,N_22638,N_23654);
xor U26092 (N_26092,N_24651,N_22870);
xnor U26093 (N_26093,N_24973,N_22849);
xnor U26094 (N_26094,N_23437,N_22959);
xor U26095 (N_26095,N_24745,N_22814);
or U26096 (N_26096,N_24930,N_23876);
or U26097 (N_26097,N_24691,N_23793);
or U26098 (N_26098,N_23946,N_23367);
nand U26099 (N_26099,N_22913,N_22556);
nand U26100 (N_26100,N_24167,N_23066);
or U26101 (N_26101,N_24655,N_23710);
nor U26102 (N_26102,N_24143,N_24436);
nor U26103 (N_26103,N_23078,N_24556);
and U26104 (N_26104,N_23559,N_24633);
or U26105 (N_26105,N_23985,N_24106);
nand U26106 (N_26106,N_23740,N_23402);
nor U26107 (N_26107,N_24903,N_23264);
nand U26108 (N_26108,N_24559,N_22858);
xnor U26109 (N_26109,N_22741,N_22794);
nor U26110 (N_26110,N_24595,N_23579);
nand U26111 (N_26111,N_22984,N_23774);
xnor U26112 (N_26112,N_22977,N_23510);
and U26113 (N_26113,N_22912,N_23899);
or U26114 (N_26114,N_23182,N_23634);
xor U26115 (N_26115,N_23257,N_24650);
nand U26116 (N_26116,N_24366,N_24766);
or U26117 (N_26117,N_24557,N_24646);
xor U26118 (N_26118,N_22583,N_23554);
and U26119 (N_26119,N_23746,N_24038);
nand U26120 (N_26120,N_24757,N_24838);
nand U26121 (N_26121,N_23198,N_24704);
nor U26122 (N_26122,N_22996,N_22848);
or U26123 (N_26123,N_23386,N_24434);
xnor U26124 (N_26124,N_24001,N_24989);
or U26125 (N_26125,N_23476,N_23453);
xor U26126 (N_26126,N_22978,N_22747);
xnor U26127 (N_26127,N_24626,N_22842);
nor U26128 (N_26128,N_22944,N_24666);
and U26129 (N_26129,N_23092,N_23224);
xor U26130 (N_26130,N_23119,N_24363);
nor U26131 (N_26131,N_22665,N_23772);
and U26132 (N_26132,N_23540,N_24831);
xnor U26133 (N_26133,N_24592,N_22652);
nor U26134 (N_26134,N_24813,N_23669);
nand U26135 (N_26135,N_23015,N_24494);
or U26136 (N_26136,N_24829,N_24309);
xor U26137 (N_26137,N_23513,N_24863);
or U26138 (N_26138,N_23723,N_24005);
or U26139 (N_26139,N_24506,N_24110);
or U26140 (N_26140,N_24455,N_24399);
and U26141 (N_26141,N_23629,N_24125);
nand U26142 (N_26142,N_23645,N_23004);
nor U26143 (N_26143,N_22891,N_24116);
xor U26144 (N_26144,N_23822,N_24769);
or U26145 (N_26145,N_23676,N_24042);
nand U26146 (N_26146,N_22831,N_24750);
or U26147 (N_26147,N_22685,N_23325);
nand U26148 (N_26148,N_23477,N_23403);
and U26149 (N_26149,N_23094,N_22651);
or U26150 (N_26150,N_23434,N_23576);
nor U26151 (N_26151,N_23743,N_24016);
or U26152 (N_26152,N_23020,N_24619);
nor U26153 (N_26153,N_23830,N_23001);
xor U26154 (N_26154,N_22534,N_23080);
or U26155 (N_26155,N_22602,N_24158);
or U26156 (N_26156,N_23816,N_24699);
nor U26157 (N_26157,N_22584,N_23974);
and U26158 (N_26158,N_24860,N_23235);
xnor U26159 (N_26159,N_23947,N_22809);
nor U26160 (N_26160,N_22776,N_24679);
or U26161 (N_26161,N_24784,N_23688);
nor U26162 (N_26162,N_22717,N_22646);
xor U26163 (N_26163,N_23423,N_23053);
xor U26164 (N_26164,N_24719,N_24878);
and U26165 (N_26165,N_24229,N_24343);
xnor U26166 (N_26166,N_23998,N_23767);
nor U26167 (N_26167,N_24300,N_22937);
xnor U26168 (N_26168,N_23074,N_24539);
or U26169 (N_26169,N_23086,N_24986);
nor U26170 (N_26170,N_23622,N_22931);
or U26171 (N_26171,N_23418,N_22657);
nand U26172 (N_26172,N_24043,N_23324);
and U26173 (N_26173,N_24768,N_23005);
nor U26174 (N_26174,N_23860,N_23683);
nor U26175 (N_26175,N_24613,N_23208);
nand U26176 (N_26176,N_23865,N_22825);
xnor U26177 (N_26177,N_24099,N_22751);
nand U26178 (N_26178,N_23871,N_23151);
nand U26179 (N_26179,N_22892,N_22796);
nor U26180 (N_26180,N_24169,N_22649);
or U26181 (N_26181,N_23552,N_24014);
nor U26182 (N_26182,N_24593,N_23288);
nor U26183 (N_26183,N_22539,N_24868);
nand U26184 (N_26184,N_23108,N_24174);
nand U26185 (N_26185,N_23391,N_23323);
xor U26186 (N_26186,N_23135,N_24920);
xor U26187 (N_26187,N_24017,N_23268);
and U26188 (N_26188,N_23342,N_24815);
nand U26189 (N_26189,N_22744,N_22855);
nand U26190 (N_26190,N_22686,N_23448);
xnor U26191 (N_26191,N_24233,N_22578);
nor U26192 (N_26192,N_23626,N_22692);
or U26193 (N_26193,N_22884,N_23995);
nor U26194 (N_26194,N_24927,N_23882);
xnor U26195 (N_26195,N_24818,N_24873);
nor U26196 (N_26196,N_22506,N_23754);
xor U26197 (N_26197,N_23440,N_23265);
nand U26198 (N_26198,N_24444,N_23316);
nor U26199 (N_26199,N_24912,N_24312);
nor U26200 (N_26200,N_23884,N_23100);
and U26201 (N_26201,N_24009,N_24528);
nor U26202 (N_26202,N_23459,N_22781);
and U26203 (N_26203,N_23879,N_23196);
nor U26204 (N_26204,N_24368,N_24846);
nand U26205 (N_26205,N_24782,N_24823);
nor U26206 (N_26206,N_24367,N_23113);
or U26207 (N_26207,N_23607,N_23382);
or U26208 (N_26208,N_23986,N_23485);
nor U26209 (N_26209,N_23991,N_22677);
xor U26210 (N_26210,N_24443,N_23490);
or U26211 (N_26211,N_24764,N_23373);
xor U26212 (N_26212,N_22508,N_24786);
or U26213 (N_26213,N_23069,N_22726);
or U26214 (N_26214,N_24990,N_24486);
or U26215 (N_26215,N_23744,N_23546);
or U26216 (N_26216,N_23920,N_24753);
xnor U26217 (N_26217,N_23535,N_24464);
xnor U26218 (N_26218,N_22941,N_22670);
nand U26219 (N_26219,N_23761,N_23383);
and U26220 (N_26220,N_24433,N_24194);
and U26221 (N_26221,N_23763,N_22836);
nand U26222 (N_26222,N_23110,N_22926);
xnor U26223 (N_26223,N_24012,N_24088);
or U26224 (N_26224,N_23095,N_24711);
nand U26225 (N_26225,N_22974,N_23169);
and U26226 (N_26226,N_23254,N_22547);
and U26227 (N_26227,N_23149,N_24787);
and U26228 (N_26228,N_24840,N_23210);
and U26229 (N_26229,N_23747,N_23668);
or U26230 (N_26230,N_23209,N_23528);
or U26231 (N_26231,N_23977,N_24280);
nand U26232 (N_26232,N_23033,N_24310);
xnor U26233 (N_26233,N_24102,N_24553);
nor U26234 (N_26234,N_22727,N_23127);
xnor U26235 (N_26235,N_22608,N_23648);
xor U26236 (N_26236,N_23682,N_23310);
or U26237 (N_26237,N_22924,N_24942);
nand U26238 (N_26238,N_24337,N_23056);
nor U26239 (N_26239,N_24488,N_22743);
or U26240 (N_26240,N_23128,N_24445);
nor U26241 (N_26241,N_24397,N_23371);
xor U26242 (N_26242,N_24925,N_22523);
xor U26243 (N_26243,N_24608,N_24323);
nand U26244 (N_26244,N_22950,N_23581);
nor U26245 (N_26245,N_23849,N_23370);
nor U26246 (N_26246,N_24083,N_24683);
xor U26247 (N_26247,N_24889,N_22874);
xor U26248 (N_26248,N_24708,N_22703);
nor U26249 (N_26249,N_23673,N_23097);
and U26250 (N_26250,N_23102,N_24214);
xnor U26251 (N_26251,N_23913,N_23494);
xor U26252 (N_26252,N_23705,N_23939);
and U26253 (N_26253,N_24146,N_24588);
and U26254 (N_26254,N_24731,N_24972);
and U26255 (N_26255,N_23005,N_23372);
and U26256 (N_26256,N_24186,N_24450);
and U26257 (N_26257,N_23670,N_23632);
or U26258 (N_26258,N_23998,N_22788);
or U26259 (N_26259,N_24699,N_23932);
nor U26260 (N_26260,N_24284,N_24133);
xnor U26261 (N_26261,N_23833,N_23583);
and U26262 (N_26262,N_22617,N_24891);
nand U26263 (N_26263,N_23992,N_23026);
nand U26264 (N_26264,N_22707,N_22893);
nand U26265 (N_26265,N_24442,N_24489);
or U26266 (N_26266,N_23491,N_22650);
and U26267 (N_26267,N_24258,N_23394);
and U26268 (N_26268,N_24601,N_24021);
and U26269 (N_26269,N_23787,N_22838);
or U26270 (N_26270,N_23376,N_23545);
nor U26271 (N_26271,N_23009,N_24445);
and U26272 (N_26272,N_22633,N_23007);
and U26273 (N_26273,N_23638,N_24156);
nand U26274 (N_26274,N_23419,N_24784);
xnor U26275 (N_26275,N_24959,N_22724);
nor U26276 (N_26276,N_24887,N_22571);
or U26277 (N_26277,N_23088,N_23175);
and U26278 (N_26278,N_23069,N_23094);
nor U26279 (N_26279,N_24075,N_24107);
nor U26280 (N_26280,N_23133,N_24762);
or U26281 (N_26281,N_24535,N_24534);
nand U26282 (N_26282,N_22856,N_24630);
xnor U26283 (N_26283,N_23276,N_24054);
nand U26284 (N_26284,N_24235,N_24443);
or U26285 (N_26285,N_23655,N_24163);
or U26286 (N_26286,N_22960,N_23903);
nand U26287 (N_26287,N_22641,N_24684);
nor U26288 (N_26288,N_23233,N_22668);
nand U26289 (N_26289,N_24080,N_24328);
nor U26290 (N_26290,N_24665,N_23122);
or U26291 (N_26291,N_23520,N_23203);
and U26292 (N_26292,N_22970,N_24430);
and U26293 (N_26293,N_23442,N_22749);
nand U26294 (N_26294,N_24996,N_23040);
and U26295 (N_26295,N_22840,N_23108);
nor U26296 (N_26296,N_24882,N_24035);
nand U26297 (N_26297,N_24578,N_23027);
nand U26298 (N_26298,N_22773,N_24557);
nor U26299 (N_26299,N_23265,N_22951);
xor U26300 (N_26300,N_22658,N_23141);
or U26301 (N_26301,N_24276,N_24105);
xor U26302 (N_26302,N_23240,N_23685);
xnor U26303 (N_26303,N_24796,N_23666);
nand U26304 (N_26304,N_23745,N_24349);
xnor U26305 (N_26305,N_24520,N_23585);
nand U26306 (N_26306,N_23380,N_23186);
nand U26307 (N_26307,N_24887,N_24169);
xnor U26308 (N_26308,N_22519,N_23880);
xor U26309 (N_26309,N_23479,N_24620);
xnor U26310 (N_26310,N_22881,N_24520);
nor U26311 (N_26311,N_22587,N_24316);
or U26312 (N_26312,N_24095,N_23501);
nor U26313 (N_26313,N_24131,N_22843);
nand U26314 (N_26314,N_23554,N_23758);
xnor U26315 (N_26315,N_22984,N_22916);
or U26316 (N_26316,N_23772,N_23667);
and U26317 (N_26317,N_24754,N_23078);
or U26318 (N_26318,N_23919,N_24671);
xor U26319 (N_26319,N_24142,N_23793);
nor U26320 (N_26320,N_23220,N_23029);
and U26321 (N_26321,N_24880,N_24615);
nand U26322 (N_26322,N_24046,N_22950);
nand U26323 (N_26323,N_23180,N_24891);
xor U26324 (N_26324,N_23352,N_24796);
nor U26325 (N_26325,N_24929,N_22519);
nor U26326 (N_26326,N_24458,N_22710);
nor U26327 (N_26327,N_22523,N_24530);
nor U26328 (N_26328,N_24065,N_24948);
nand U26329 (N_26329,N_24079,N_22720);
and U26330 (N_26330,N_23319,N_24310);
nand U26331 (N_26331,N_23386,N_23960);
nor U26332 (N_26332,N_23696,N_23987);
or U26333 (N_26333,N_23226,N_24132);
nor U26334 (N_26334,N_23192,N_23381);
nand U26335 (N_26335,N_22975,N_24220);
and U26336 (N_26336,N_24600,N_23996);
nand U26337 (N_26337,N_23027,N_23179);
or U26338 (N_26338,N_23139,N_22636);
or U26339 (N_26339,N_23372,N_23157);
nand U26340 (N_26340,N_23003,N_23514);
or U26341 (N_26341,N_24591,N_23910);
nand U26342 (N_26342,N_22564,N_24837);
or U26343 (N_26343,N_23992,N_24412);
and U26344 (N_26344,N_24767,N_23117);
nor U26345 (N_26345,N_24487,N_24894);
xnor U26346 (N_26346,N_24453,N_22895);
xor U26347 (N_26347,N_22926,N_24336);
or U26348 (N_26348,N_23675,N_24586);
and U26349 (N_26349,N_22858,N_24113);
nor U26350 (N_26350,N_22836,N_22965);
nand U26351 (N_26351,N_24354,N_24472);
xor U26352 (N_26352,N_24873,N_24122);
nand U26353 (N_26353,N_23584,N_23877);
xor U26354 (N_26354,N_23085,N_24638);
xor U26355 (N_26355,N_22751,N_23035);
or U26356 (N_26356,N_22550,N_23179);
xnor U26357 (N_26357,N_22998,N_24891);
and U26358 (N_26358,N_22947,N_23937);
xnor U26359 (N_26359,N_23319,N_23124);
nand U26360 (N_26360,N_22548,N_22762);
or U26361 (N_26361,N_22506,N_23348);
or U26362 (N_26362,N_23849,N_23336);
xor U26363 (N_26363,N_22715,N_23228);
nand U26364 (N_26364,N_24883,N_23203);
nor U26365 (N_26365,N_24212,N_24651);
and U26366 (N_26366,N_22919,N_22822);
nand U26367 (N_26367,N_23125,N_24683);
or U26368 (N_26368,N_24630,N_24134);
nor U26369 (N_26369,N_24848,N_22743);
or U26370 (N_26370,N_24950,N_24490);
or U26371 (N_26371,N_24606,N_23220);
nor U26372 (N_26372,N_24881,N_23894);
or U26373 (N_26373,N_23083,N_23855);
and U26374 (N_26374,N_24603,N_24206);
and U26375 (N_26375,N_24935,N_22765);
or U26376 (N_26376,N_24628,N_23211);
nor U26377 (N_26377,N_22852,N_24632);
xnor U26378 (N_26378,N_23266,N_23355);
nand U26379 (N_26379,N_24271,N_22946);
and U26380 (N_26380,N_24074,N_24909);
or U26381 (N_26381,N_23699,N_22825);
nand U26382 (N_26382,N_23708,N_23979);
xnor U26383 (N_26383,N_24429,N_24262);
nand U26384 (N_26384,N_23445,N_23215);
nor U26385 (N_26385,N_23409,N_23495);
and U26386 (N_26386,N_23352,N_23253);
and U26387 (N_26387,N_23317,N_22963);
xnor U26388 (N_26388,N_23931,N_24101);
nor U26389 (N_26389,N_24252,N_24235);
and U26390 (N_26390,N_23484,N_23805);
xnor U26391 (N_26391,N_24129,N_24102);
nand U26392 (N_26392,N_23844,N_23530);
and U26393 (N_26393,N_23869,N_24196);
xor U26394 (N_26394,N_23640,N_22765);
and U26395 (N_26395,N_23132,N_22927);
or U26396 (N_26396,N_23423,N_23618);
xor U26397 (N_26397,N_24097,N_24028);
xnor U26398 (N_26398,N_23374,N_22706);
or U26399 (N_26399,N_24564,N_23151);
nand U26400 (N_26400,N_23109,N_24650);
xor U26401 (N_26401,N_23391,N_24249);
nor U26402 (N_26402,N_23536,N_22755);
nand U26403 (N_26403,N_23618,N_22689);
xor U26404 (N_26404,N_22576,N_23700);
xor U26405 (N_26405,N_23626,N_22843);
xnor U26406 (N_26406,N_23384,N_22505);
and U26407 (N_26407,N_23097,N_22936);
nor U26408 (N_26408,N_23964,N_22566);
and U26409 (N_26409,N_23262,N_24022);
xor U26410 (N_26410,N_23339,N_23752);
nand U26411 (N_26411,N_23276,N_23270);
xor U26412 (N_26412,N_24679,N_23581);
nor U26413 (N_26413,N_23828,N_24184);
or U26414 (N_26414,N_22657,N_24552);
nand U26415 (N_26415,N_23373,N_22561);
nor U26416 (N_26416,N_23478,N_23229);
nand U26417 (N_26417,N_24573,N_24822);
and U26418 (N_26418,N_22802,N_22903);
xor U26419 (N_26419,N_24028,N_23025);
xor U26420 (N_26420,N_23792,N_23244);
xor U26421 (N_26421,N_24514,N_22606);
or U26422 (N_26422,N_23417,N_23023);
nor U26423 (N_26423,N_23588,N_23323);
and U26424 (N_26424,N_23083,N_22834);
or U26425 (N_26425,N_24513,N_22871);
nand U26426 (N_26426,N_22556,N_24770);
xnor U26427 (N_26427,N_24095,N_23470);
nand U26428 (N_26428,N_23370,N_23774);
or U26429 (N_26429,N_24952,N_24674);
nor U26430 (N_26430,N_22751,N_23550);
nor U26431 (N_26431,N_24156,N_23676);
and U26432 (N_26432,N_22661,N_23664);
and U26433 (N_26433,N_24319,N_24637);
xnor U26434 (N_26434,N_24818,N_24214);
xnor U26435 (N_26435,N_22537,N_24276);
xor U26436 (N_26436,N_24140,N_24918);
or U26437 (N_26437,N_22906,N_23728);
or U26438 (N_26438,N_22956,N_22845);
and U26439 (N_26439,N_24820,N_23532);
nand U26440 (N_26440,N_23419,N_24435);
or U26441 (N_26441,N_23266,N_24270);
nand U26442 (N_26442,N_23341,N_23330);
or U26443 (N_26443,N_23943,N_24595);
nand U26444 (N_26444,N_23130,N_23435);
xnor U26445 (N_26445,N_23177,N_23438);
nand U26446 (N_26446,N_22509,N_23001);
xnor U26447 (N_26447,N_22513,N_23776);
xnor U26448 (N_26448,N_23302,N_23155);
or U26449 (N_26449,N_23706,N_24033);
nand U26450 (N_26450,N_24274,N_22917);
and U26451 (N_26451,N_23556,N_23642);
xor U26452 (N_26452,N_23309,N_22702);
xnor U26453 (N_26453,N_23446,N_22860);
or U26454 (N_26454,N_22599,N_23914);
xnor U26455 (N_26455,N_23725,N_22520);
and U26456 (N_26456,N_23023,N_22880);
or U26457 (N_26457,N_23142,N_24220);
xor U26458 (N_26458,N_24031,N_23216);
or U26459 (N_26459,N_23338,N_22644);
or U26460 (N_26460,N_23132,N_23846);
or U26461 (N_26461,N_24169,N_24861);
or U26462 (N_26462,N_22935,N_23996);
xor U26463 (N_26463,N_23492,N_23956);
nand U26464 (N_26464,N_24610,N_23176);
and U26465 (N_26465,N_23143,N_23851);
nor U26466 (N_26466,N_23200,N_22651);
and U26467 (N_26467,N_24004,N_22764);
xnor U26468 (N_26468,N_24402,N_23302);
or U26469 (N_26469,N_23694,N_23732);
xor U26470 (N_26470,N_23056,N_23096);
xor U26471 (N_26471,N_24736,N_22874);
nor U26472 (N_26472,N_24481,N_24125);
nor U26473 (N_26473,N_23498,N_23793);
nor U26474 (N_26474,N_24714,N_24523);
nand U26475 (N_26475,N_24765,N_22759);
and U26476 (N_26476,N_24510,N_22707);
nand U26477 (N_26477,N_22614,N_23529);
nand U26478 (N_26478,N_24382,N_24129);
xor U26479 (N_26479,N_24059,N_23142);
nor U26480 (N_26480,N_23938,N_23719);
or U26481 (N_26481,N_24440,N_24457);
nand U26482 (N_26482,N_24189,N_24209);
and U26483 (N_26483,N_24447,N_24454);
xnor U26484 (N_26484,N_24917,N_24446);
xor U26485 (N_26485,N_22642,N_23095);
and U26486 (N_26486,N_23264,N_24756);
nor U26487 (N_26487,N_24196,N_24128);
nand U26488 (N_26488,N_23186,N_24683);
nand U26489 (N_26489,N_23336,N_24235);
nor U26490 (N_26490,N_23892,N_24320);
and U26491 (N_26491,N_22884,N_22870);
nand U26492 (N_26492,N_22586,N_23759);
nand U26493 (N_26493,N_23482,N_23267);
nor U26494 (N_26494,N_22726,N_23462);
or U26495 (N_26495,N_23172,N_23572);
or U26496 (N_26496,N_23356,N_22559);
and U26497 (N_26497,N_24389,N_24203);
or U26498 (N_26498,N_22927,N_22868);
nor U26499 (N_26499,N_23728,N_22505);
and U26500 (N_26500,N_23590,N_22660);
or U26501 (N_26501,N_23570,N_24098);
xor U26502 (N_26502,N_22564,N_24910);
and U26503 (N_26503,N_24510,N_22763);
nor U26504 (N_26504,N_23664,N_23456);
nand U26505 (N_26505,N_24326,N_23375);
and U26506 (N_26506,N_23930,N_23791);
xor U26507 (N_26507,N_22990,N_23959);
xor U26508 (N_26508,N_23855,N_23553);
nor U26509 (N_26509,N_24750,N_24768);
and U26510 (N_26510,N_22910,N_24450);
nor U26511 (N_26511,N_24163,N_24584);
and U26512 (N_26512,N_23507,N_24903);
xor U26513 (N_26513,N_23265,N_22986);
xor U26514 (N_26514,N_24745,N_23885);
xor U26515 (N_26515,N_24102,N_23375);
and U26516 (N_26516,N_22941,N_24843);
xor U26517 (N_26517,N_22501,N_24242);
and U26518 (N_26518,N_23996,N_24880);
nor U26519 (N_26519,N_23174,N_24183);
nor U26520 (N_26520,N_23685,N_23067);
nor U26521 (N_26521,N_24491,N_23084);
or U26522 (N_26522,N_24232,N_24226);
and U26523 (N_26523,N_22810,N_22617);
nor U26524 (N_26524,N_24095,N_22696);
or U26525 (N_26525,N_24449,N_23853);
nand U26526 (N_26526,N_24737,N_22885);
xnor U26527 (N_26527,N_23733,N_23797);
xor U26528 (N_26528,N_24457,N_24637);
or U26529 (N_26529,N_23381,N_22840);
or U26530 (N_26530,N_24482,N_23901);
and U26531 (N_26531,N_22988,N_22682);
and U26532 (N_26532,N_23682,N_24853);
xor U26533 (N_26533,N_23037,N_22685);
xnor U26534 (N_26534,N_23047,N_24712);
nor U26535 (N_26535,N_23099,N_22839);
or U26536 (N_26536,N_24491,N_23150);
or U26537 (N_26537,N_23486,N_24455);
and U26538 (N_26538,N_22770,N_23843);
and U26539 (N_26539,N_24151,N_23604);
nand U26540 (N_26540,N_24250,N_23411);
nand U26541 (N_26541,N_24766,N_24412);
xor U26542 (N_26542,N_23215,N_24584);
nor U26543 (N_26543,N_24189,N_24945);
nand U26544 (N_26544,N_24680,N_23828);
nor U26545 (N_26545,N_22847,N_23895);
and U26546 (N_26546,N_24725,N_24143);
and U26547 (N_26547,N_24936,N_23232);
or U26548 (N_26548,N_23218,N_22542);
xnor U26549 (N_26549,N_22972,N_24281);
nand U26550 (N_26550,N_23941,N_23497);
xnor U26551 (N_26551,N_22666,N_24630);
nand U26552 (N_26552,N_22608,N_24864);
or U26553 (N_26553,N_23993,N_23703);
nor U26554 (N_26554,N_22541,N_23636);
xnor U26555 (N_26555,N_24550,N_23544);
and U26556 (N_26556,N_23525,N_23715);
and U26557 (N_26557,N_23401,N_24691);
or U26558 (N_26558,N_24562,N_23701);
nor U26559 (N_26559,N_24610,N_24507);
or U26560 (N_26560,N_23475,N_23853);
or U26561 (N_26561,N_24944,N_23082);
xnor U26562 (N_26562,N_24171,N_22606);
nand U26563 (N_26563,N_23797,N_24059);
or U26564 (N_26564,N_22798,N_23891);
xnor U26565 (N_26565,N_23369,N_24051);
xor U26566 (N_26566,N_24069,N_23494);
or U26567 (N_26567,N_24989,N_22897);
and U26568 (N_26568,N_24863,N_22729);
and U26569 (N_26569,N_24911,N_23649);
xnor U26570 (N_26570,N_23534,N_23942);
and U26571 (N_26571,N_24048,N_24463);
xnor U26572 (N_26572,N_24960,N_24349);
and U26573 (N_26573,N_22824,N_24817);
xnor U26574 (N_26574,N_23364,N_24273);
nor U26575 (N_26575,N_24862,N_24300);
xnor U26576 (N_26576,N_24038,N_23917);
xor U26577 (N_26577,N_22673,N_23617);
nor U26578 (N_26578,N_23181,N_24126);
xnor U26579 (N_26579,N_24208,N_23177);
xor U26580 (N_26580,N_23224,N_23089);
and U26581 (N_26581,N_24489,N_24719);
nor U26582 (N_26582,N_23754,N_24436);
nor U26583 (N_26583,N_24614,N_23671);
and U26584 (N_26584,N_22711,N_24647);
nand U26585 (N_26585,N_24350,N_22764);
nand U26586 (N_26586,N_24925,N_24964);
xor U26587 (N_26587,N_22887,N_24017);
xnor U26588 (N_26588,N_24121,N_24827);
and U26589 (N_26589,N_24551,N_23020);
nor U26590 (N_26590,N_22955,N_23683);
nor U26591 (N_26591,N_23851,N_24445);
nand U26592 (N_26592,N_23235,N_24278);
nand U26593 (N_26593,N_22536,N_23590);
nand U26594 (N_26594,N_24407,N_22674);
nor U26595 (N_26595,N_22636,N_24865);
nor U26596 (N_26596,N_24227,N_22975);
nor U26597 (N_26597,N_23913,N_24417);
xnor U26598 (N_26598,N_23491,N_23215);
or U26599 (N_26599,N_24188,N_24717);
or U26600 (N_26600,N_24226,N_23086);
xnor U26601 (N_26601,N_23018,N_23446);
nor U26602 (N_26602,N_24538,N_24688);
nor U26603 (N_26603,N_24747,N_24987);
and U26604 (N_26604,N_24326,N_22519);
xnor U26605 (N_26605,N_23193,N_24182);
or U26606 (N_26606,N_24206,N_22767);
nor U26607 (N_26607,N_23735,N_22691);
nand U26608 (N_26608,N_22999,N_22729);
xnor U26609 (N_26609,N_23339,N_24222);
or U26610 (N_26610,N_24699,N_24057);
and U26611 (N_26611,N_24154,N_23436);
nor U26612 (N_26612,N_23108,N_23748);
nor U26613 (N_26613,N_23040,N_24934);
or U26614 (N_26614,N_24206,N_23657);
xnor U26615 (N_26615,N_23510,N_22512);
xor U26616 (N_26616,N_24622,N_23006);
or U26617 (N_26617,N_24660,N_23260);
or U26618 (N_26618,N_23018,N_23348);
and U26619 (N_26619,N_24576,N_22620);
nor U26620 (N_26620,N_24818,N_24420);
xor U26621 (N_26621,N_24447,N_24155);
nand U26622 (N_26622,N_22544,N_23276);
nand U26623 (N_26623,N_24744,N_24299);
xor U26624 (N_26624,N_22517,N_23891);
or U26625 (N_26625,N_23683,N_23702);
or U26626 (N_26626,N_23611,N_24292);
nor U26627 (N_26627,N_23921,N_23229);
or U26628 (N_26628,N_22707,N_23172);
xor U26629 (N_26629,N_23546,N_23781);
and U26630 (N_26630,N_24338,N_23159);
and U26631 (N_26631,N_23081,N_22720);
xnor U26632 (N_26632,N_24771,N_23987);
or U26633 (N_26633,N_22566,N_23389);
nand U26634 (N_26634,N_23188,N_24194);
nor U26635 (N_26635,N_22925,N_23865);
nor U26636 (N_26636,N_24795,N_23721);
xnor U26637 (N_26637,N_22677,N_23249);
nor U26638 (N_26638,N_23572,N_24768);
or U26639 (N_26639,N_23399,N_22840);
and U26640 (N_26640,N_23747,N_24863);
xor U26641 (N_26641,N_24070,N_23372);
or U26642 (N_26642,N_23900,N_22968);
nor U26643 (N_26643,N_23622,N_24678);
and U26644 (N_26644,N_24514,N_22925);
nand U26645 (N_26645,N_23001,N_23969);
xor U26646 (N_26646,N_23823,N_22924);
or U26647 (N_26647,N_22729,N_24657);
xnor U26648 (N_26648,N_23549,N_23805);
and U26649 (N_26649,N_24161,N_22853);
and U26650 (N_26650,N_23898,N_23978);
and U26651 (N_26651,N_22808,N_23979);
nand U26652 (N_26652,N_22968,N_24274);
nor U26653 (N_26653,N_24948,N_24127);
nor U26654 (N_26654,N_23513,N_22843);
and U26655 (N_26655,N_23156,N_23947);
nand U26656 (N_26656,N_24633,N_23590);
xnor U26657 (N_26657,N_22888,N_24017);
xor U26658 (N_26658,N_24132,N_23010);
xnor U26659 (N_26659,N_23494,N_22892);
xnor U26660 (N_26660,N_23467,N_23602);
xnor U26661 (N_26661,N_23121,N_23774);
nand U26662 (N_26662,N_24678,N_22501);
and U26663 (N_26663,N_23600,N_24088);
or U26664 (N_26664,N_23981,N_23458);
xor U26665 (N_26665,N_24398,N_22780);
nand U26666 (N_26666,N_23889,N_24757);
nor U26667 (N_26667,N_24370,N_24058);
or U26668 (N_26668,N_23523,N_22520);
nor U26669 (N_26669,N_24403,N_24657);
xor U26670 (N_26670,N_23072,N_24086);
or U26671 (N_26671,N_24489,N_22701);
xor U26672 (N_26672,N_24613,N_24788);
nand U26673 (N_26673,N_23740,N_24285);
and U26674 (N_26674,N_22900,N_23346);
nor U26675 (N_26675,N_24640,N_24247);
nor U26676 (N_26676,N_24586,N_24595);
and U26677 (N_26677,N_24064,N_24451);
nor U26678 (N_26678,N_24274,N_23535);
nand U26679 (N_26679,N_23977,N_24225);
xor U26680 (N_26680,N_24402,N_23425);
nand U26681 (N_26681,N_23872,N_22693);
and U26682 (N_26682,N_24610,N_22929);
nor U26683 (N_26683,N_23844,N_24670);
nand U26684 (N_26684,N_22926,N_23919);
or U26685 (N_26685,N_23818,N_24017);
xnor U26686 (N_26686,N_22999,N_24980);
and U26687 (N_26687,N_24656,N_24521);
nand U26688 (N_26688,N_22594,N_23062);
or U26689 (N_26689,N_23700,N_23296);
and U26690 (N_26690,N_24302,N_24305);
or U26691 (N_26691,N_23517,N_22560);
nor U26692 (N_26692,N_22864,N_23371);
nor U26693 (N_26693,N_22868,N_24954);
and U26694 (N_26694,N_22951,N_24586);
nand U26695 (N_26695,N_23955,N_22716);
xor U26696 (N_26696,N_24105,N_24726);
and U26697 (N_26697,N_23272,N_24436);
nor U26698 (N_26698,N_24062,N_23349);
and U26699 (N_26699,N_22688,N_23800);
or U26700 (N_26700,N_24463,N_24974);
nor U26701 (N_26701,N_23894,N_22677);
nand U26702 (N_26702,N_23660,N_23704);
and U26703 (N_26703,N_23511,N_22585);
nor U26704 (N_26704,N_22973,N_23846);
nor U26705 (N_26705,N_24178,N_24203);
xnor U26706 (N_26706,N_22908,N_24351);
nand U26707 (N_26707,N_23465,N_24502);
xor U26708 (N_26708,N_23908,N_22640);
and U26709 (N_26709,N_24952,N_24155);
nand U26710 (N_26710,N_24099,N_22782);
nand U26711 (N_26711,N_23220,N_22503);
or U26712 (N_26712,N_22815,N_23587);
xnor U26713 (N_26713,N_22754,N_24136);
nand U26714 (N_26714,N_24188,N_24567);
nand U26715 (N_26715,N_23430,N_23172);
xnor U26716 (N_26716,N_23194,N_24371);
and U26717 (N_26717,N_23008,N_22614);
xor U26718 (N_26718,N_23679,N_24691);
or U26719 (N_26719,N_23760,N_23587);
or U26720 (N_26720,N_24569,N_22631);
and U26721 (N_26721,N_24430,N_23645);
xor U26722 (N_26722,N_24518,N_24210);
nand U26723 (N_26723,N_24354,N_23040);
nor U26724 (N_26724,N_23151,N_23614);
or U26725 (N_26725,N_24438,N_24442);
nand U26726 (N_26726,N_22594,N_22580);
or U26727 (N_26727,N_24702,N_24618);
or U26728 (N_26728,N_24053,N_23356);
or U26729 (N_26729,N_24264,N_23860);
and U26730 (N_26730,N_23740,N_24661);
and U26731 (N_26731,N_24563,N_24941);
nor U26732 (N_26732,N_24606,N_22912);
nand U26733 (N_26733,N_24640,N_23527);
nand U26734 (N_26734,N_22781,N_22789);
or U26735 (N_26735,N_22840,N_23371);
xnor U26736 (N_26736,N_23633,N_23875);
xnor U26737 (N_26737,N_23278,N_23790);
or U26738 (N_26738,N_23456,N_24856);
xor U26739 (N_26739,N_23469,N_23281);
and U26740 (N_26740,N_24069,N_24672);
nor U26741 (N_26741,N_23759,N_23825);
and U26742 (N_26742,N_23087,N_24471);
and U26743 (N_26743,N_24789,N_23065);
nand U26744 (N_26744,N_23065,N_23156);
and U26745 (N_26745,N_23612,N_22739);
xnor U26746 (N_26746,N_22700,N_22515);
or U26747 (N_26747,N_24614,N_24341);
nand U26748 (N_26748,N_22561,N_23254);
and U26749 (N_26749,N_24723,N_24602);
or U26750 (N_26750,N_23836,N_23742);
xor U26751 (N_26751,N_22509,N_24523);
xor U26752 (N_26752,N_24160,N_23863);
and U26753 (N_26753,N_22524,N_23635);
nor U26754 (N_26754,N_23934,N_22775);
or U26755 (N_26755,N_23006,N_23154);
nand U26756 (N_26756,N_23770,N_24455);
or U26757 (N_26757,N_24804,N_24500);
and U26758 (N_26758,N_24562,N_23475);
or U26759 (N_26759,N_22532,N_24416);
xor U26760 (N_26760,N_22943,N_23789);
or U26761 (N_26761,N_23915,N_23614);
xor U26762 (N_26762,N_24290,N_23425);
and U26763 (N_26763,N_24441,N_22926);
nor U26764 (N_26764,N_23132,N_24246);
nand U26765 (N_26765,N_23591,N_23086);
nand U26766 (N_26766,N_24692,N_23109);
or U26767 (N_26767,N_22582,N_23344);
or U26768 (N_26768,N_23702,N_24136);
xnor U26769 (N_26769,N_23175,N_24326);
xnor U26770 (N_26770,N_23751,N_24524);
and U26771 (N_26771,N_23565,N_23623);
nor U26772 (N_26772,N_24522,N_24646);
and U26773 (N_26773,N_24556,N_22844);
nor U26774 (N_26774,N_22612,N_22611);
nand U26775 (N_26775,N_22651,N_23907);
or U26776 (N_26776,N_22574,N_23600);
nand U26777 (N_26777,N_22593,N_23733);
xor U26778 (N_26778,N_24056,N_24455);
xnor U26779 (N_26779,N_24139,N_24088);
and U26780 (N_26780,N_24447,N_23767);
or U26781 (N_26781,N_24640,N_23782);
and U26782 (N_26782,N_24738,N_22607);
or U26783 (N_26783,N_22583,N_23604);
or U26784 (N_26784,N_24705,N_24230);
and U26785 (N_26785,N_23369,N_24871);
xnor U26786 (N_26786,N_23094,N_24462);
nand U26787 (N_26787,N_22769,N_24188);
and U26788 (N_26788,N_23694,N_24311);
xnor U26789 (N_26789,N_23404,N_23707);
nand U26790 (N_26790,N_22515,N_24915);
or U26791 (N_26791,N_23973,N_23649);
xor U26792 (N_26792,N_24440,N_23018);
nand U26793 (N_26793,N_24780,N_24362);
or U26794 (N_26794,N_24376,N_24985);
xor U26795 (N_26795,N_22555,N_23834);
nor U26796 (N_26796,N_23480,N_23477);
and U26797 (N_26797,N_24655,N_24269);
and U26798 (N_26798,N_23645,N_24847);
xor U26799 (N_26799,N_23975,N_23607);
or U26800 (N_26800,N_23358,N_23988);
or U26801 (N_26801,N_24716,N_22637);
or U26802 (N_26802,N_22662,N_24471);
xnor U26803 (N_26803,N_22531,N_24046);
and U26804 (N_26804,N_23169,N_23021);
xor U26805 (N_26805,N_23666,N_24444);
nand U26806 (N_26806,N_23770,N_23199);
xor U26807 (N_26807,N_24909,N_23621);
nand U26808 (N_26808,N_24503,N_23164);
or U26809 (N_26809,N_24500,N_23093);
xnor U26810 (N_26810,N_23674,N_24573);
xor U26811 (N_26811,N_24385,N_24080);
nand U26812 (N_26812,N_24538,N_24786);
nand U26813 (N_26813,N_23643,N_24948);
or U26814 (N_26814,N_23649,N_23735);
and U26815 (N_26815,N_24229,N_23567);
xnor U26816 (N_26816,N_24186,N_23049);
nand U26817 (N_26817,N_24211,N_22615);
or U26818 (N_26818,N_24771,N_24845);
nand U26819 (N_26819,N_24674,N_24266);
nand U26820 (N_26820,N_23828,N_24942);
xor U26821 (N_26821,N_23250,N_23500);
nor U26822 (N_26822,N_24760,N_22849);
nand U26823 (N_26823,N_23182,N_24315);
or U26824 (N_26824,N_23729,N_24047);
nand U26825 (N_26825,N_24465,N_23739);
xor U26826 (N_26826,N_24991,N_24943);
and U26827 (N_26827,N_24277,N_23266);
and U26828 (N_26828,N_24848,N_24280);
or U26829 (N_26829,N_23479,N_23968);
nand U26830 (N_26830,N_23138,N_23179);
xnor U26831 (N_26831,N_22556,N_23409);
nand U26832 (N_26832,N_24813,N_23067);
nor U26833 (N_26833,N_24762,N_24284);
xor U26834 (N_26834,N_22671,N_23659);
xnor U26835 (N_26835,N_23796,N_22944);
and U26836 (N_26836,N_24782,N_23893);
xnor U26837 (N_26837,N_23473,N_22644);
nor U26838 (N_26838,N_23056,N_22677);
and U26839 (N_26839,N_24055,N_23510);
or U26840 (N_26840,N_24198,N_23598);
nand U26841 (N_26841,N_23570,N_24838);
or U26842 (N_26842,N_24661,N_23342);
nor U26843 (N_26843,N_23227,N_24978);
and U26844 (N_26844,N_22859,N_24741);
nor U26845 (N_26845,N_23339,N_22616);
nor U26846 (N_26846,N_23216,N_23157);
and U26847 (N_26847,N_23703,N_22684);
nand U26848 (N_26848,N_23910,N_24191);
xor U26849 (N_26849,N_24811,N_23921);
nor U26850 (N_26850,N_23452,N_22610);
or U26851 (N_26851,N_23596,N_23526);
or U26852 (N_26852,N_22826,N_22503);
or U26853 (N_26853,N_24059,N_22650);
xor U26854 (N_26854,N_23855,N_22774);
nand U26855 (N_26855,N_24387,N_22791);
xnor U26856 (N_26856,N_23006,N_24998);
and U26857 (N_26857,N_24782,N_24514);
nand U26858 (N_26858,N_23020,N_24785);
nand U26859 (N_26859,N_24388,N_23381);
xnor U26860 (N_26860,N_23167,N_24086);
or U26861 (N_26861,N_22765,N_23180);
nor U26862 (N_26862,N_23653,N_24421);
nor U26863 (N_26863,N_24948,N_23867);
nand U26864 (N_26864,N_24152,N_23272);
xnor U26865 (N_26865,N_23418,N_24352);
or U26866 (N_26866,N_24849,N_22992);
nand U26867 (N_26867,N_24568,N_22794);
nor U26868 (N_26868,N_23533,N_24707);
xor U26869 (N_26869,N_23674,N_23369);
and U26870 (N_26870,N_23712,N_23794);
nor U26871 (N_26871,N_23847,N_23205);
xor U26872 (N_26872,N_24544,N_22779);
xor U26873 (N_26873,N_22722,N_23256);
and U26874 (N_26874,N_23422,N_23251);
and U26875 (N_26875,N_24730,N_24939);
or U26876 (N_26876,N_23432,N_24633);
or U26877 (N_26877,N_24864,N_23022);
nor U26878 (N_26878,N_24792,N_24768);
nor U26879 (N_26879,N_22891,N_23479);
nand U26880 (N_26880,N_22815,N_24296);
nor U26881 (N_26881,N_24382,N_24977);
and U26882 (N_26882,N_24094,N_24713);
and U26883 (N_26883,N_24428,N_23378);
or U26884 (N_26884,N_24194,N_24405);
nand U26885 (N_26885,N_22678,N_23126);
xor U26886 (N_26886,N_23036,N_22566);
or U26887 (N_26887,N_23350,N_23227);
and U26888 (N_26888,N_23513,N_24086);
nand U26889 (N_26889,N_23000,N_23430);
nand U26890 (N_26890,N_22906,N_22718);
or U26891 (N_26891,N_24684,N_23602);
or U26892 (N_26892,N_23481,N_22832);
and U26893 (N_26893,N_23342,N_24239);
nand U26894 (N_26894,N_22728,N_23730);
or U26895 (N_26895,N_24985,N_23001);
nor U26896 (N_26896,N_22685,N_24742);
xnor U26897 (N_26897,N_24486,N_23502);
nand U26898 (N_26898,N_22576,N_24186);
nand U26899 (N_26899,N_23401,N_22566);
nand U26900 (N_26900,N_23110,N_22886);
or U26901 (N_26901,N_22989,N_23674);
xor U26902 (N_26902,N_24111,N_22889);
xor U26903 (N_26903,N_24020,N_23961);
and U26904 (N_26904,N_22956,N_23280);
xnor U26905 (N_26905,N_23054,N_23373);
and U26906 (N_26906,N_23415,N_24306);
xnor U26907 (N_26907,N_24977,N_23881);
nand U26908 (N_26908,N_23148,N_24550);
nor U26909 (N_26909,N_23295,N_22939);
or U26910 (N_26910,N_23503,N_22633);
and U26911 (N_26911,N_23483,N_23228);
and U26912 (N_26912,N_24662,N_22563);
nor U26913 (N_26913,N_22919,N_24442);
and U26914 (N_26914,N_23398,N_23133);
or U26915 (N_26915,N_23739,N_24069);
xnor U26916 (N_26916,N_24616,N_23119);
and U26917 (N_26917,N_22813,N_22615);
nor U26918 (N_26918,N_22870,N_23932);
nor U26919 (N_26919,N_24325,N_22632);
nand U26920 (N_26920,N_24720,N_23648);
and U26921 (N_26921,N_24696,N_24311);
or U26922 (N_26922,N_24267,N_23464);
and U26923 (N_26923,N_24078,N_22878);
nor U26924 (N_26924,N_22524,N_23012);
nand U26925 (N_26925,N_23951,N_23921);
nor U26926 (N_26926,N_24735,N_23546);
nand U26927 (N_26927,N_22761,N_23674);
nor U26928 (N_26928,N_24962,N_23486);
nand U26929 (N_26929,N_23806,N_23340);
xnor U26930 (N_26930,N_23791,N_24810);
xor U26931 (N_26931,N_23028,N_23677);
nand U26932 (N_26932,N_23662,N_23933);
nor U26933 (N_26933,N_23284,N_24078);
xnor U26934 (N_26934,N_23010,N_22652);
nand U26935 (N_26935,N_23505,N_24518);
and U26936 (N_26936,N_24326,N_23738);
nor U26937 (N_26937,N_22919,N_24432);
nor U26938 (N_26938,N_24866,N_23338);
and U26939 (N_26939,N_22621,N_23397);
nand U26940 (N_26940,N_24206,N_23551);
or U26941 (N_26941,N_24520,N_23281);
nand U26942 (N_26942,N_22595,N_22956);
nand U26943 (N_26943,N_24597,N_23122);
and U26944 (N_26944,N_24563,N_24304);
or U26945 (N_26945,N_22554,N_23116);
nor U26946 (N_26946,N_24322,N_24470);
nand U26947 (N_26947,N_22535,N_22955);
xor U26948 (N_26948,N_24499,N_23102);
or U26949 (N_26949,N_22824,N_22880);
and U26950 (N_26950,N_23446,N_23234);
xnor U26951 (N_26951,N_23724,N_22754);
and U26952 (N_26952,N_24377,N_23565);
nand U26953 (N_26953,N_23332,N_24713);
nor U26954 (N_26954,N_22935,N_22852);
nor U26955 (N_26955,N_22819,N_23459);
and U26956 (N_26956,N_24220,N_22812);
xnor U26957 (N_26957,N_23162,N_24880);
nor U26958 (N_26958,N_24364,N_23320);
and U26959 (N_26959,N_23179,N_24455);
xor U26960 (N_26960,N_24451,N_24038);
nand U26961 (N_26961,N_23299,N_24697);
nor U26962 (N_26962,N_24947,N_24862);
and U26963 (N_26963,N_22912,N_24951);
and U26964 (N_26964,N_22667,N_24318);
nor U26965 (N_26965,N_24642,N_22929);
or U26966 (N_26966,N_23533,N_23143);
and U26967 (N_26967,N_22624,N_22723);
or U26968 (N_26968,N_24110,N_24374);
xor U26969 (N_26969,N_23470,N_22635);
nor U26970 (N_26970,N_23566,N_22656);
xnor U26971 (N_26971,N_23750,N_24358);
or U26972 (N_26972,N_24786,N_24258);
nand U26973 (N_26973,N_24138,N_22820);
xnor U26974 (N_26974,N_23851,N_24211);
or U26975 (N_26975,N_24669,N_23556);
nand U26976 (N_26976,N_23136,N_23911);
nand U26977 (N_26977,N_24250,N_23290);
and U26978 (N_26978,N_24460,N_23482);
xnor U26979 (N_26979,N_24458,N_23831);
xor U26980 (N_26980,N_22546,N_24632);
or U26981 (N_26981,N_22900,N_22550);
or U26982 (N_26982,N_22996,N_23571);
nor U26983 (N_26983,N_23602,N_24669);
or U26984 (N_26984,N_23567,N_23304);
and U26985 (N_26985,N_23548,N_23481);
xor U26986 (N_26986,N_24565,N_24212);
nor U26987 (N_26987,N_23803,N_24426);
and U26988 (N_26988,N_22952,N_23587);
or U26989 (N_26989,N_24894,N_24660);
xor U26990 (N_26990,N_22767,N_24632);
nand U26991 (N_26991,N_24512,N_23842);
xor U26992 (N_26992,N_23760,N_24538);
and U26993 (N_26993,N_24729,N_22908);
nand U26994 (N_26994,N_23114,N_23975);
xnor U26995 (N_26995,N_23249,N_24230);
nor U26996 (N_26996,N_24008,N_23931);
nand U26997 (N_26997,N_22529,N_22631);
or U26998 (N_26998,N_24070,N_23253);
and U26999 (N_26999,N_24522,N_24432);
and U27000 (N_27000,N_24342,N_22714);
nand U27001 (N_27001,N_23101,N_24776);
nor U27002 (N_27002,N_22745,N_24414);
nor U27003 (N_27003,N_23900,N_24170);
nor U27004 (N_27004,N_23653,N_23852);
or U27005 (N_27005,N_23926,N_24700);
nor U27006 (N_27006,N_22739,N_24346);
or U27007 (N_27007,N_23502,N_24687);
and U27008 (N_27008,N_24390,N_23163);
or U27009 (N_27009,N_22629,N_24161);
xor U27010 (N_27010,N_22512,N_23660);
and U27011 (N_27011,N_23330,N_23997);
and U27012 (N_27012,N_23695,N_24607);
nand U27013 (N_27013,N_23657,N_23586);
and U27014 (N_27014,N_22523,N_23943);
or U27015 (N_27015,N_24890,N_23066);
xnor U27016 (N_27016,N_22854,N_22597);
or U27017 (N_27017,N_24621,N_23832);
xnor U27018 (N_27018,N_23633,N_23486);
nor U27019 (N_27019,N_24731,N_22550);
or U27020 (N_27020,N_23831,N_24139);
xnor U27021 (N_27021,N_24881,N_24014);
and U27022 (N_27022,N_23184,N_24084);
and U27023 (N_27023,N_22643,N_22699);
xnor U27024 (N_27024,N_23254,N_24326);
xnor U27025 (N_27025,N_24389,N_23546);
and U27026 (N_27026,N_23537,N_24093);
and U27027 (N_27027,N_22930,N_23176);
nor U27028 (N_27028,N_24819,N_24755);
or U27029 (N_27029,N_23022,N_24744);
or U27030 (N_27030,N_22834,N_23242);
or U27031 (N_27031,N_23150,N_23697);
nor U27032 (N_27032,N_24169,N_23537);
nor U27033 (N_27033,N_24152,N_22996);
nand U27034 (N_27034,N_23729,N_23159);
xor U27035 (N_27035,N_23982,N_22722);
and U27036 (N_27036,N_23597,N_24935);
xor U27037 (N_27037,N_23249,N_23522);
nand U27038 (N_27038,N_22767,N_22703);
nand U27039 (N_27039,N_22585,N_24731);
nor U27040 (N_27040,N_24890,N_23692);
nand U27041 (N_27041,N_23561,N_24896);
or U27042 (N_27042,N_22538,N_24542);
nor U27043 (N_27043,N_23674,N_24155);
xor U27044 (N_27044,N_22927,N_22820);
nor U27045 (N_27045,N_23149,N_23046);
nor U27046 (N_27046,N_24933,N_24411);
xnor U27047 (N_27047,N_22708,N_23199);
and U27048 (N_27048,N_24980,N_24198);
xnor U27049 (N_27049,N_24771,N_23298);
or U27050 (N_27050,N_22731,N_22811);
and U27051 (N_27051,N_24462,N_23113);
and U27052 (N_27052,N_23883,N_24578);
nand U27053 (N_27053,N_23841,N_22683);
or U27054 (N_27054,N_23109,N_23715);
or U27055 (N_27055,N_23107,N_22653);
nor U27056 (N_27056,N_23054,N_24000);
and U27057 (N_27057,N_22567,N_23337);
xor U27058 (N_27058,N_24667,N_23206);
nor U27059 (N_27059,N_24215,N_24598);
or U27060 (N_27060,N_23896,N_22703);
nor U27061 (N_27061,N_22502,N_23956);
nor U27062 (N_27062,N_22806,N_23946);
and U27063 (N_27063,N_23188,N_23197);
nor U27064 (N_27064,N_23138,N_23441);
xor U27065 (N_27065,N_23886,N_24747);
xor U27066 (N_27066,N_22887,N_24336);
and U27067 (N_27067,N_23145,N_23808);
xor U27068 (N_27068,N_24865,N_22991);
and U27069 (N_27069,N_23555,N_23498);
nand U27070 (N_27070,N_23009,N_23628);
and U27071 (N_27071,N_24040,N_23876);
xor U27072 (N_27072,N_24208,N_22904);
nor U27073 (N_27073,N_24385,N_24253);
xor U27074 (N_27074,N_23034,N_22509);
and U27075 (N_27075,N_24487,N_23114);
and U27076 (N_27076,N_24659,N_24407);
xnor U27077 (N_27077,N_23931,N_22944);
and U27078 (N_27078,N_23630,N_24248);
nand U27079 (N_27079,N_22852,N_23020);
and U27080 (N_27080,N_23766,N_24750);
and U27081 (N_27081,N_22915,N_23673);
nor U27082 (N_27082,N_24397,N_22891);
or U27083 (N_27083,N_24669,N_24826);
and U27084 (N_27084,N_24160,N_23532);
nand U27085 (N_27085,N_24063,N_24791);
or U27086 (N_27086,N_24680,N_22870);
or U27087 (N_27087,N_24347,N_23840);
nor U27088 (N_27088,N_22545,N_23577);
and U27089 (N_27089,N_22716,N_23945);
or U27090 (N_27090,N_22643,N_22636);
and U27091 (N_27091,N_24753,N_23065);
nor U27092 (N_27092,N_24676,N_23950);
nand U27093 (N_27093,N_22877,N_24736);
or U27094 (N_27094,N_24969,N_23148);
nand U27095 (N_27095,N_24578,N_23190);
nor U27096 (N_27096,N_24131,N_24083);
nand U27097 (N_27097,N_23104,N_24155);
xor U27098 (N_27098,N_24542,N_23813);
xnor U27099 (N_27099,N_23439,N_22783);
nor U27100 (N_27100,N_23031,N_23006);
nand U27101 (N_27101,N_24203,N_23085);
nand U27102 (N_27102,N_23853,N_24622);
xnor U27103 (N_27103,N_23069,N_22585);
nand U27104 (N_27104,N_24927,N_24415);
nand U27105 (N_27105,N_22779,N_23239);
and U27106 (N_27106,N_24371,N_24091);
or U27107 (N_27107,N_23345,N_24921);
or U27108 (N_27108,N_24532,N_24583);
nand U27109 (N_27109,N_23744,N_23009);
or U27110 (N_27110,N_24587,N_24020);
nand U27111 (N_27111,N_24821,N_22762);
xnor U27112 (N_27112,N_23321,N_22755);
and U27113 (N_27113,N_23728,N_24254);
nor U27114 (N_27114,N_23810,N_23873);
nand U27115 (N_27115,N_23331,N_23811);
or U27116 (N_27116,N_23050,N_23179);
and U27117 (N_27117,N_23120,N_24719);
nor U27118 (N_27118,N_24295,N_24185);
xor U27119 (N_27119,N_24721,N_24779);
xor U27120 (N_27120,N_24333,N_22627);
or U27121 (N_27121,N_23281,N_24517);
nand U27122 (N_27122,N_23311,N_23497);
xnor U27123 (N_27123,N_24492,N_23786);
and U27124 (N_27124,N_23852,N_24408);
nand U27125 (N_27125,N_22914,N_23171);
nand U27126 (N_27126,N_22507,N_22838);
and U27127 (N_27127,N_24584,N_22981);
xor U27128 (N_27128,N_24814,N_22917);
or U27129 (N_27129,N_23550,N_24479);
nor U27130 (N_27130,N_24277,N_23176);
or U27131 (N_27131,N_23926,N_24301);
or U27132 (N_27132,N_22530,N_23286);
nor U27133 (N_27133,N_24647,N_24726);
and U27134 (N_27134,N_23622,N_24538);
or U27135 (N_27135,N_24070,N_22587);
nand U27136 (N_27136,N_22926,N_24149);
nand U27137 (N_27137,N_22818,N_23405);
or U27138 (N_27138,N_23510,N_23273);
nor U27139 (N_27139,N_24948,N_22949);
and U27140 (N_27140,N_24081,N_22618);
or U27141 (N_27141,N_24793,N_24593);
xor U27142 (N_27142,N_24479,N_23098);
and U27143 (N_27143,N_23237,N_24609);
nand U27144 (N_27144,N_23082,N_23112);
xnor U27145 (N_27145,N_24713,N_22840);
nand U27146 (N_27146,N_24808,N_23644);
or U27147 (N_27147,N_24193,N_23838);
xor U27148 (N_27148,N_23572,N_23471);
nand U27149 (N_27149,N_24393,N_23007);
and U27150 (N_27150,N_23007,N_23694);
nand U27151 (N_27151,N_23756,N_23717);
or U27152 (N_27152,N_24165,N_23470);
nand U27153 (N_27153,N_23261,N_24599);
or U27154 (N_27154,N_23116,N_23547);
xor U27155 (N_27155,N_22935,N_24073);
nor U27156 (N_27156,N_24085,N_24354);
nand U27157 (N_27157,N_24327,N_23654);
nor U27158 (N_27158,N_24364,N_22744);
and U27159 (N_27159,N_23264,N_24785);
and U27160 (N_27160,N_24329,N_24394);
nand U27161 (N_27161,N_22906,N_24127);
nand U27162 (N_27162,N_24591,N_24095);
and U27163 (N_27163,N_22885,N_23065);
nand U27164 (N_27164,N_22882,N_23574);
nand U27165 (N_27165,N_24741,N_23943);
nand U27166 (N_27166,N_22761,N_23965);
and U27167 (N_27167,N_22520,N_22605);
xor U27168 (N_27168,N_23922,N_23322);
and U27169 (N_27169,N_24954,N_23480);
nor U27170 (N_27170,N_24562,N_22726);
or U27171 (N_27171,N_24750,N_24948);
nand U27172 (N_27172,N_24293,N_22517);
nand U27173 (N_27173,N_24839,N_24157);
and U27174 (N_27174,N_23558,N_23652);
and U27175 (N_27175,N_24109,N_22863);
or U27176 (N_27176,N_24306,N_23933);
nand U27177 (N_27177,N_22795,N_24199);
nor U27178 (N_27178,N_23802,N_23844);
and U27179 (N_27179,N_23127,N_24041);
xnor U27180 (N_27180,N_22553,N_23342);
and U27181 (N_27181,N_24877,N_24526);
xnor U27182 (N_27182,N_24353,N_24113);
or U27183 (N_27183,N_24077,N_22604);
xor U27184 (N_27184,N_23096,N_23851);
or U27185 (N_27185,N_23577,N_22606);
and U27186 (N_27186,N_24355,N_23901);
nor U27187 (N_27187,N_23996,N_22630);
xnor U27188 (N_27188,N_22982,N_23243);
or U27189 (N_27189,N_23983,N_23556);
xor U27190 (N_27190,N_24473,N_24690);
and U27191 (N_27191,N_24301,N_23304);
nor U27192 (N_27192,N_24734,N_22637);
or U27193 (N_27193,N_22529,N_23162);
nand U27194 (N_27194,N_23377,N_24189);
xor U27195 (N_27195,N_23997,N_23928);
nand U27196 (N_27196,N_22627,N_24668);
or U27197 (N_27197,N_24417,N_23129);
and U27198 (N_27198,N_24299,N_22554);
or U27199 (N_27199,N_24180,N_24789);
xor U27200 (N_27200,N_24853,N_24324);
and U27201 (N_27201,N_24217,N_22745);
nand U27202 (N_27202,N_23443,N_24944);
or U27203 (N_27203,N_22632,N_24407);
and U27204 (N_27204,N_22753,N_24020);
or U27205 (N_27205,N_23426,N_24881);
nand U27206 (N_27206,N_22572,N_23492);
and U27207 (N_27207,N_23686,N_22638);
nor U27208 (N_27208,N_24906,N_24004);
nor U27209 (N_27209,N_24456,N_24732);
and U27210 (N_27210,N_22623,N_22928);
xnor U27211 (N_27211,N_22521,N_23730);
and U27212 (N_27212,N_22743,N_22695);
nor U27213 (N_27213,N_24530,N_24464);
nand U27214 (N_27214,N_24054,N_22570);
and U27215 (N_27215,N_23677,N_23916);
xor U27216 (N_27216,N_23744,N_23276);
xnor U27217 (N_27217,N_23546,N_22617);
and U27218 (N_27218,N_23652,N_22686);
nor U27219 (N_27219,N_24337,N_24494);
nand U27220 (N_27220,N_23043,N_22589);
nand U27221 (N_27221,N_23429,N_24155);
nand U27222 (N_27222,N_22845,N_24811);
nor U27223 (N_27223,N_22602,N_24747);
nand U27224 (N_27224,N_22859,N_24131);
nand U27225 (N_27225,N_23013,N_24638);
nand U27226 (N_27226,N_23579,N_23157);
or U27227 (N_27227,N_23160,N_23808);
xor U27228 (N_27228,N_23353,N_24097);
and U27229 (N_27229,N_23505,N_23371);
or U27230 (N_27230,N_22543,N_24983);
or U27231 (N_27231,N_24178,N_23949);
or U27232 (N_27232,N_23815,N_24143);
nand U27233 (N_27233,N_23047,N_24710);
and U27234 (N_27234,N_22618,N_23304);
nor U27235 (N_27235,N_24347,N_22721);
xnor U27236 (N_27236,N_23057,N_24687);
and U27237 (N_27237,N_23138,N_23956);
nor U27238 (N_27238,N_23311,N_23426);
or U27239 (N_27239,N_23436,N_22891);
nor U27240 (N_27240,N_24885,N_24757);
nand U27241 (N_27241,N_23574,N_23568);
xnor U27242 (N_27242,N_23657,N_22818);
nand U27243 (N_27243,N_24428,N_24812);
and U27244 (N_27244,N_24440,N_22554);
and U27245 (N_27245,N_23895,N_24385);
and U27246 (N_27246,N_24008,N_22840);
nand U27247 (N_27247,N_24524,N_22687);
nor U27248 (N_27248,N_24031,N_22803);
xnor U27249 (N_27249,N_22855,N_24029);
nor U27250 (N_27250,N_24436,N_24423);
xor U27251 (N_27251,N_24601,N_22918);
or U27252 (N_27252,N_22849,N_23444);
or U27253 (N_27253,N_22820,N_24183);
or U27254 (N_27254,N_24568,N_23658);
and U27255 (N_27255,N_23856,N_24748);
nor U27256 (N_27256,N_22500,N_24735);
or U27257 (N_27257,N_23998,N_23427);
or U27258 (N_27258,N_22942,N_24300);
and U27259 (N_27259,N_24536,N_24883);
or U27260 (N_27260,N_22801,N_23189);
nor U27261 (N_27261,N_24980,N_23457);
xor U27262 (N_27262,N_23894,N_23017);
and U27263 (N_27263,N_24283,N_23289);
nor U27264 (N_27264,N_24945,N_24307);
nor U27265 (N_27265,N_24882,N_23417);
or U27266 (N_27266,N_22999,N_24598);
nand U27267 (N_27267,N_22976,N_22977);
xnor U27268 (N_27268,N_23170,N_24350);
xnor U27269 (N_27269,N_23733,N_24047);
nor U27270 (N_27270,N_23467,N_24029);
or U27271 (N_27271,N_23972,N_22957);
nand U27272 (N_27272,N_22647,N_22772);
nand U27273 (N_27273,N_23939,N_24838);
nor U27274 (N_27274,N_22733,N_23505);
nor U27275 (N_27275,N_23653,N_23954);
nor U27276 (N_27276,N_23445,N_22574);
nand U27277 (N_27277,N_23318,N_22522);
nor U27278 (N_27278,N_24298,N_24626);
or U27279 (N_27279,N_23362,N_24453);
xnor U27280 (N_27280,N_24998,N_24414);
nor U27281 (N_27281,N_24178,N_23167);
and U27282 (N_27282,N_24263,N_22912);
and U27283 (N_27283,N_22616,N_24477);
nand U27284 (N_27284,N_23568,N_24415);
and U27285 (N_27285,N_23980,N_24243);
nand U27286 (N_27286,N_24416,N_24991);
and U27287 (N_27287,N_24396,N_24087);
nand U27288 (N_27288,N_24758,N_23418);
nand U27289 (N_27289,N_24027,N_22808);
and U27290 (N_27290,N_24287,N_23256);
nor U27291 (N_27291,N_24158,N_23836);
xor U27292 (N_27292,N_23229,N_23728);
nand U27293 (N_27293,N_24496,N_24719);
xnor U27294 (N_27294,N_22766,N_22570);
and U27295 (N_27295,N_24398,N_22514);
or U27296 (N_27296,N_22700,N_23452);
and U27297 (N_27297,N_24005,N_23553);
nand U27298 (N_27298,N_22985,N_23694);
or U27299 (N_27299,N_24710,N_23848);
nor U27300 (N_27300,N_23978,N_23246);
xnor U27301 (N_27301,N_24994,N_24775);
nand U27302 (N_27302,N_23765,N_23481);
or U27303 (N_27303,N_23260,N_22757);
nand U27304 (N_27304,N_24134,N_22919);
nor U27305 (N_27305,N_22945,N_23246);
nand U27306 (N_27306,N_23955,N_24052);
or U27307 (N_27307,N_24661,N_23172);
xor U27308 (N_27308,N_23965,N_23648);
nand U27309 (N_27309,N_23191,N_24686);
nand U27310 (N_27310,N_24988,N_22942);
nor U27311 (N_27311,N_23671,N_24490);
nand U27312 (N_27312,N_23402,N_23000);
and U27313 (N_27313,N_24727,N_23560);
nor U27314 (N_27314,N_24351,N_22734);
xor U27315 (N_27315,N_24009,N_23098);
xnor U27316 (N_27316,N_24032,N_24007);
xor U27317 (N_27317,N_24917,N_24818);
xnor U27318 (N_27318,N_23179,N_23107);
nor U27319 (N_27319,N_24450,N_24242);
nand U27320 (N_27320,N_23772,N_22629);
and U27321 (N_27321,N_23847,N_24531);
and U27322 (N_27322,N_23176,N_24392);
xnor U27323 (N_27323,N_24564,N_23291);
nand U27324 (N_27324,N_23546,N_22860);
or U27325 (N_27325,N_23433,N_24162);
or U27326 (N_27326,N_23442,N_23045);
or U27327 (N_27327,N_23535,N_23892);
or U27328 (N_27328,N_23877,N_23092);
nand U27329 (N_27329,N_23843,N_24165);
nand U27330 (N_27330,N_22707,N_24383);
nand U27331 (N_27331,N_23248,N_22628);
nand U27332 (N_27332,N_23325,N_22725);
xnor U27333 (N_27333,N_24081,N_24209);
or U27334 (N_27334,N_24114,N_23863);
xnor U27335 (N_27335,N_23877,N_24993);
xor U27336 (N_27336,N_24621,N_22671);
and U27337 (N_27337,N_22878,N_23681);
and U27338 (N_27338,N_24073,N_23029);
and U27339 (N_27339,N_23014,N_23617);
xor U27340 (N_27340,N_22958,N_23486);
or U27341 (N_27341,N_24909,N_22996);
nor U27342 (N_27342,N_22852,N_23824);
and U27343 (N_27343,N_23077,N_24739);
nor U27344 (N_27344,N_24093,N_24574);
or U27345 (N_27345,N_24989,N_24749);
and U27346 (N_27346,N_23377,N_24891);
xnor U27347 (N_27347,N_22725,N_24452);
nor U27348 (N_27348,N_24736,N_24878);
or U27349 (N_27349,N_23998,N_23215);
and U27350 (N_27350,N_24891,N_22906);
nand U27351 (N_27351,N_24645,N_24519);
xnor U27352 (N_27352,N_22746,N_24303);
or U27353 (N_27353,N_24236,N_24026);
and U27354 (N_27354,N_24531,N_24755);
nand U27355 (N_27355,N_24166,N_23731);
nor U27356 (N_27356,N_24837,N_23643);
nor U27357 (N_27357,N_23155,N_23893);
and U27358 (N_27358,N_24729,N_24306);
xnor U27359 (N_27359,N_22724,N_22977);
or U27360 (N_27360,N_24835,N_24270);
and U27361 (N_27361,N_23022,N_24000);
nand U27362 (N_27362,N_23452,N_23954);
and U27363 (N_27363,N_22601,N_24484);
xor U27364 (N_27364,N_22752,N_23682);
or U27365 (N_27365,N_23627,N_24745);
or U27366 (N_27366,N_24662,N_23660);
and U27367 (N_27367,N_23248,N_22509);
or U27368 (N_27368,N_24566,N_23809);
and U27369 (N_27369,N_24237,N_23911);
xnor U27370 (N_27370,N_23860,N_24409);
or U27371 (N_27371,N_24886,N_24233);
nand U27372 (N_27372,N_22803,N_23089);
and U27373 (N_27373,N_23750,N_23217);
nor U27374 (N_27374,N_23874,N_23840);
and U27375 (N_27375,N_22965,N_23456);
xor U27376 (N_27376,N_23188,N_24977);
nor U27377 (N_27377,N_24571,N_24454);
xor U27378 (N_27378,N_22945,N_24289);
nor U27379 (N_27379,N_23503,N_22680);
xor U27380 (N_27380,N_22791,N_23702);
xnor U27381 (N_27381,N_23023,N_24315);
nor U27382 (N_27382,N_23917,N_23599);
or U27383 (N_27383,N_22666,N_24308);
or U27384 (N_27384,N_24725,N_22930);
nor U27385 (N_27385,N_24838,N_23564);
xnor U27386 (N_27386,N_23599,N_22628);
xor U27387 (N_27387,N_24817,N_23819);
and U27388 (N_27388,N_23562,N_22771);
nand U27389 (N_27389,N_23602,N_24347);
and U27390 (N_27390,N_24455,N_24651);
nor U27391 (N_27391,N_22931,N_24876);
or U27392 (N_27392,N_24076,N_23498);
xor U27393 (N_27393,N_22603,N_24056);
nand U27394 (N_27394,N_24205,N_23197);
or U27395 (N_27395,N_24177,N_24881);
xor U27396 (N_27396,N_24311,N_23426);
xor U27397 (N_27397,N_24544,N_23344);
nand U27398 (N_27398,N_24354,N_23871);
nor U27399 (N_27399,N_24873,N_23328);
and U27400 (N_27400,N_22912,N_23300);
or U27401 (N_27401,N_24771,N_24336);
and U27402 (N_27402,N_22545,N_22651);
nor U27403 (N_27403,N_23827,N_23742);
nand U27404 (N_27404,N_23885,N_22581);
nor U27405 (N_27405,N_24824,N_24158);
or U27406 (N_27406,N_22607,N_22902);
xnor U27407 (N_27407,N_23079,N_22959);
nand U27408 (N_27408,N_24998,N_22765);
nand U27409 (N_27409,N_23133,N_23697);
nand U27410 (N_27410,N_23449,N_24328);
or U27411 (N_27411,N_23231,N_23400);
or U27412 (N_27412,N_24038,N_24302);
xor U27413 (N_27413,N_23440,N_24378);
or U27414 (N_27414,N_22927,N_24583);
or U27415 (N_27415,N_22889,N_22532);
and U27416 (N_27416,N_23987,N_23746);
nor U27417 (N_27417,N_22684,N_22967);
nand U27418 (N_27418,N_24080,N_24440);
or U27419 (N_27419,N_22986,N_24534);
or U27420 (N_27420,N_24266,N_24855);
nor U27421 (N_27421,N_23566,N_23319);
xor U27422 (N_27422,N_22725,N_23062);
xnor U27423 (N_27423,N_23108,N_23771);
nand U27424 (N_27424,N_24962,N_24943);
nand U27425 (N_27425,N_24756,N_24382);
xnor U27426 (N_27426,N_23863,N_24484);
or U27427 (N_27427,N_22755,N_22850);
nor U27428 (N_27428,N_24857,N_24027);
or U27429 (N_27429,N_22753,N_23563);
nor U27430 (N_27430,N_24505,N_22726);
and U27431 (N_27431,N_22518,N_24745);
or U27432 (N_27432,N_24383,N_23680);
nand U27433 (N_27433,N_24352,N_23902);
nand U27434 (N_27434,N_24317,N_22953);
nor U27435 (N_27435,N_24413,N_22678);
nor U27436 (N_27436,N_24472,N_22508);
nor U27437 (N_27437,N_22683,N_22526);
or U27438 (N_27438,N_24907,N_23667);
or U27439 (N_27439,N_23449,N_22784);
and U27440 (N_27440,N_24500,N_24761);
nor U27441 (N_27441,N_24488,N_22847);
nor U27442 (N_27442,N_24782,N_23972);
xor U27443 (N_27443,N_24206,N_24970);
nor U27444 (N_27444,N_24645,N_23732);
or U27445 (N_27445,N_23544,N_23275);
xor U27446 (N_27446,N_22549,N_24089);
or U27447 (N_27447,N_23907,N_24086);
xnor U27448 (N_27448,N_23851,N_23212);
and U27449 (N_27449,N_24885,N_24331);
nand U27450 (N_27450,N_24220,N_24514);
xor U27451 (N_27451,N_23108,N_22962);
and U27452 (N_27452,N_24550,N_23168);
nor U27453 (N_27453,N_22600,N_22795);
xor U27454 (N_27454,N_22627,N_23652);
nand U27455 (N_27455,N_23463,N_24886);
and U27456 (N_27456,N_23183,N_24414);
nand U27457 (N_27457,N_23776,N_24477);
xor U27458 (N_27458,N_24140,N_22769);
and U27459 (N_27459,N_23628,N_23473);
nor U27460 (N_27460,N_24999,N_22541);
xor U27461 (N_27461,N_23870,N_24490);
and U27462 (N_27462,N_22974,N_23452);
nor U27463 (N_27463,N_22959,N_24454);
and U27464 (N_27464,N_24366,N_22827);
or U27465 (N_27465,N_23276,N_24619);
xor U27466 (N_27466,N_24026,N_23667);
nand U27467 (N_27467,N_23978,N_23488);
nand U27468 (N_27468,N_24582,N_24480);
xor U27469 (N_27469,N_22650,N_23062);
xor U27470 (N_27470,N_24351,N_22586);
xor U27471 (N_27471,N_24566,N_23877);
nand U27472 (N_27472,N_23783,N_23844);
nand U27473 (N_27473,N_24168,N_22979);
xor U27474 (N_27474,N_24787,N_24811);
nand U27475 (N_27475,N_23591,N_22506);
nand U27476 (N_27476,N_24944,N_24864);
xor U27477 (N_27477,N_24236,N_22823);
or U27478 (N_27478,N_24305,N_22755);
xnor U27479 (N_27479,N_22729,N_23704);
or U27480 (N_27480,N_22866,N_23247);
nor U27481 (N_27481,N_24613,N_24412);
nand U27482 (N_27482,N_22585,N_23026);
and U27483 (N_27483,N_22561,N_22691);
nor U27484 (N_27484,N_24635,N_22554);
nand U27485 (N_27485,N_24954,N_23170);
nand U27486 (N_27486,N_22825,N_24439);
nor U27487 (N_27487,N_22589,N_23878);
nand U27488 (N_27488,N_24267,N_22838);
and U27489 (N_27489,N_22540,N_24172);
xor U27490 (N_27490,N_24958,N_24266);
and U27491 (N_27491,N_22549,N_23918);
and U27492 (N_27492,N_23797,N_23414);
nand U27493 (N_27493,N_23656,N_24401);
nand U27494 (N_27494,N_24677,N_22588);
and U27495 (N_27495,N_23148,N_23610);
and U27496 (N_27496,N_24414,N_23666);
and U27497 (N_27497,N_24262,N_22616);
nand U27498 (N_27498,N_24043,N_24379);
nor U27499 (N_27499,N_24591,N_22866);
nor U27500 (N_27500,N_25487,N_25771);
and U27501 (N_27501,N_25926,N_26181);
nor U27502 (N_27502,N_27244,N_27181);
xnor U27503 (N_27503,N_27391,N_25269);
and U27504 (N_27504,N_25683,N_26375);
or U27505 (N_27505,N_26255,N_26742);
nor U27506 (N_27506,N_27130,N_27192);
nand U27507 (N_27507,N_25428,N_27371);
or U27508 (N_27508,N_26735,N_26118);
nand U27509 (N_27509,N_27396,N_27322);
xor U27510 (N_27510,N_26387,N_25472);
or U27511 (N_27511,N_27302,N_26248);
nor U27512 (N_27512,N_25271,N_26270);
or U27513 (N_27513,N_25152,N_26922);
xnor U27514 (N_27514,N_26697,N_27333);
and U27515 (N_27515,N_27126,N_25214);
xor U27516 (N_27516,N_27451,N_25609);
nand U27517 (N_27517,N_26228,N_26763);
nor U27518 (N_27518,N_25542,N_25333);
nand U27519 (N_27519,N_25827,N_26772);
xnor U27520 (N_27520,N_25565,N_26744);
nor U27521 (N_27521,N_26075,N_26645);
nand U27522 (N_27522,N_26594,N_27384);
xnor U27523 (N_27523,N_26409,N_26995);
and U27524 (N_27524,N_25492,N_25929);
nand U27525 (N_27525,N_27463,N_26837);
nand U27526 (N_27526,N_26258,N_27061);
nand U27527 (N_27527,N_26700,N_26084);
nor U27528 (N_27528,N_27057,N_26470);
nor U27529 (N_27529,N_26465,N_27088);
xor U27530 (N_27530,N_25276,N_26058);
nand U27531 (N_27531,N_25007,N_25281);
and U27532 (N_27532,N_26866,N_27430);
or U27533 (N_27533,N_25006,N_26687);
xnor U27534 (N_27534,N_25248,N_25120);
xnor U27535 (N_27535,N_25033,N_25256);
nor U27536 (N_27536,N_25113,N_26278);
nand U27537 (N_27537,N_25088,N_27195);
nor U27538 (N_27538,N_26684,N_25694);
nor U27539 (N_27539,N_26405,N_25317);
nand U27540 (N_27540,N_27102,N_26968);
or U27541 (N_27541,N_27415,N_25455);
or U27542 (N_27542,N_25510,N_25580);
and U27543 (N_27543,N_26741,N_25201);
or U27544 (N_27544,N_26949,N_25785);
nand U27545 (N_27545,N_26044,N_26189);
and U27546 (N_27546,N_26456,N_27316);
or U27547 (N_27547,N_26948,N_26434);
xnor U27548 (N_27548,N_25945,N_27053);
and U27549 (N_27549,N_26033,N_27291);
nand U27550 (N_27550,N_27264,N_25810);
nor U27551 (N_27551,N_26757,N_26670);
xnor U27552 (N_27552,N_25849,N_26726);
or U27553 (N_27553,N_26595,N_26091);
nand U27554 (N_27554,N_26624,N_25679);
or U27555 (N_27555,N_27434,N_26144);
nor U27556 (N_27556,N_25224,N_25636);
and U27557 (N_27557,N_27447,N_25767);
xnor U27558 (N_27558,N_26206,N_26857);
nor U27559 (N_27559,N_26392,N_26141);
or U27560 (N_27560,N_27213,N_27094);
nor U27561 (N_27561,N_26355,N_25350);
and U27562 (N_27562,N_27035,N_25812);
or U27563 (N_27563,N_27338,N_26219);
or U27564 (N_27564,N_26923,N_26107);
and U27565 (N_27565,N_26378,N_25588);
xnor U27566 (N_27566,N_25336,N_26719);
or U27567 (N_27567,N_25844,N_25040);
nand U27568 (N_27568,N_27107,N_25342);
or U27569 (N_27569,N_26856,N_26888);
nor U27570 (N_27570,N_25501,N_25024);
nor U27571 (N_27571,N_25950,N_26362);
xnor U27572 (N_27572,N_25092,N_26108);
xor U27573 (N_27573,N_27393,N_27177);
nor U27574 (N_27574,N_26109,N_27127);
and U27575 (N_27575,N_26022,N_25441);
and U27576 (N_27576,N_26785,N_25131);
nor U27577 (N_27577,N_25548,N_26492);
nor U27578 (N_27578,N_26993,N_25703);
or U27579 (N_27579,N_27077,N_26399);
xor U27580 (N_27580,N_25523,N_25124);
nand U27581 (N_27581,N_26782,N_27394);
nor U27582 (N_27582,N_26926,N_27199);
and U27583 (N_27583,N_26243,N_26501);
or U27584 (N_27584,N_27267,N_26983);
and U27585 (N_27585,N_25118,N_27113);
and U27586 (N_27586,N_27301,N_25566);
and U27587 (N_27587,N_27014,N_25458);
nand U27588 (N_27588,N_26938,N_25035);
nand U27589 (N_27589,N_25520,N_27037);
nor U27590 (N_27590,N_26724,N_26579);
xor U27591 (N_27591,N_25559,N_25864);
xnor U27592 (N_27592,N_25747,N_25625);
and U27593 (N_27593,N_27168,N_25901);
nand U27594 (N_27594,N_25757,N_25315);
xor U27595 (N_27595,N_26667,N_25569);
xnor U27596 (N_27596,N_25323,N_25474);
or U27597 (N_27597,N_26304,N_25973);
xor U27598 (N_27598,N_25010,N_26069);
or U27599 (N_27599,N_25439,N_27040);
xor U27600 (N_27600,N_25257,N_25401);
and U27601 (N_27601,N_26650,N_27071);
xnor U27602 (N_27602,N_26202,N_27481);
nand U27603 (N_27603,N_25989,N_27445);
nor U27604 (N_27604,N_26641,N_26083);
xnor U27605 (N_27605,N_26070,N_25642);
nand U27606 (N_27606,N_25788,N_27066);
and U27607 (N_27607,N_26804,N_27253);
xnor U27608 (N_27608,N_25185,N_25195);
nor U27609 (N_27609,N_25652,N_26442);
nor U27610 (N_27610,N_26997,N_27188);
nor U27611 (N_27611,N_25225,N_25285);
nor U27612 (N_27612,N_26485,N_26244);
nor U27613 (N_27613,N_26261,N_26854);
nor U27614 (N_27614,N_27050,N_25452);
nand U27615 (N_27615,N_27157,N_26572);
and U27616 (N_27616,N_26281,N_25602);
xnor U27617 (N_27617,N_26256,N_25138);
or U27618 (N_27618,N_26575,N_27047);
and U27619 (N_27619,N_27399,N_27266);
and U27620 (N_27620,N_25662,N_27201);
nor U27621 (N_27621,N_27386,N_26191);
xor U27622 (N_27622,N_27004,N_27010);
or U27623 (N_27623,N_27361,N_25453);
or U27624 (N_27624,N_25050,N_26389);
and U27625 (N_27625,N_27209,N_25084);
and U27626 (N_27626,N_26495,N_27326);
or U27627 (N_27627,N_25199,N_27373);
nor U27628 (N_27628,N_25431,N_26630);
nand U27629 (N_27629,N_27474,N_26077);
nand U27630 (N_27630,N_26774,N_25255);
or U27631 (N_27631,N_27225,N_25066);
nor U27632 (N_27632,N_26010,N_26941);
xor U27633 (N_27633,N_27388,N_26373);
xor U27634 (N_27634,N_25895,N_26746);
and U27635 (N_27635,N_26009,N_25707);
or U27636 (N_27636,N_27365,N_25465);
and U27637 (N_27637,N_26336,N_26499);
or U27638 (N_27638,N_25831,N_25669);
and U27639 (N_27639,N_25615,N_26863);
nor U27640 (N_27640,N_27214,N_26388);
or U27641 (N_27641,N_25300,N_25110);
nand U27642 (N_27642,N_25970,N_26482);
and U27643 (N_27643,N_26306,N_26099);
and U27644 (N_27644,N_26566,N_25109);
nand U27645 (N_27645,N_26316,N_26357);
nand U27646 (N_27646,N_25292,N_26159);
nand U27647 (N_27647,N_25903,N_27364);
nor U27648 (N_27648,N_25412,N_27479);
nand U27649 (N_27649,N_26376,N_26066);
and U27650 (N_27650,N_25394,N_25598);
xnor U27651 (N_27651,N_26655,N_25606);
xnor U27652 (N_27652,N_27406,N_25979);
xor U27653 (N_27653,N_25801,N_25198);
xnor U27654 (N_27654,N_27086,N_25784);
or U27655 (N_27655,N_27016,N_26062);
xor U27656 (N_27656,N_26221,N_26800);
xor U27657 (N_27657,N_25427,N_25820);
nand U27658 (N_27658,N_26751,N_25127);
and U27659 (N_27659,N_27346,N_27330);
xor U27660 (N_27660,N_26418,N_25994);
xnor U27661 (N_27661,N_25765,N_26640);
nor U27662 (N_27662,N_25797,N_26691);
and U27663 (N_27663,N_25197,N_26155);
and U27664 (N_27664,N_26454,N_25561);
nor U27665 (N_27665,N_26262,N_25909);
or U27666 (N_27666,N_26733,N_26975);
and U27667 (N_27667,N_27369,N_27011);
nor U27668 (N_27668,N_25957,N_26209);
xor U27669 (N_27669,N_27460,N_27172);
or U27670 (N_27670,N_26750,N_25689);
nand U27671 (N_27671,N_25511,N_26550);
nor U27672 (N_27672,N_25599,N_27072);
xor U27673 (N_27673,N_27295,N_26048);
nand U27674 (N_27674,N_25880,N_26193);
xnor U27675 (N_27675,N_26540,N_25987);
nor U27676 (N_27676,N_26198,N_27429);
and U27677 (N_27677,N_25769,N_27424);
or U27678 (N_27678,N_26942,N_25090);
and U27679 (N_27679,N_25376,N_26130);
or U27680 (N_27680,N_25772,N_26266);
and U27681 (N_27681,N_26783,N_25532);
xnor U27682 (N_27682,N_26416,N_25644);
and U27683 (N_27683,N_26176,N_25943);
nor U27684 (N_27684,N_26711,N_25435);
or U27685 (N_27685,N_25639,N_27404);
nand U27686 (N_27686,N_26977,N_27262);
nor U27687 (N_27687,N_26528,N_27392);
and U27688 (N_27688,N_27411,N_27256);
nand U27689 (N_27689,N_25675,N_26623);
and U27690 (N_27690,N_27117,N_26531);
xor U27691 (N_27691,N_25912,N_26424);
xnor U27692 (N_27692,N_26690,N_26057);
xor U27693 (N_27693,N_25729,N_27490);
nor U27694 (N_27694,N_26521,N_25166);
nor U27695 (N_27695,N_27018,N_27417);
nand U27696 (N_27696,N_25605,N_27332);
nor U27697 (N_27697,N_25026,N_25478);
nor U27698 (N_27698,N_26541,N_26188);
nand U27699 (N_27699,N_25776,N_25388);
xnor U27700 (N_27700,N_26115,N_25251);
nor U27701 (N_27701,N_26639,N_27347);
xnor U27702 (N_27702,N_26950,N_26583);
or U27703 (N_27703,N_26829,N_26564);
or U27704 (N_27704,N_26601,N_25136);
nor U27705 (N_27705,N_25930,N_27198);
nor U27706 (N_27706,N_25868,N_26335);
nor U27707 (N_27707,N_26343,N_25732);
nand U27708 (N_27708,N_26469,N_25305);
nand U27709 (N_27709,N_25661,N_25444);
and U27710 (N_27710,N_25028,N_27249);
nand U27711 (N_27711,N_25437,N_27313);
nor U27712 (N_27712,N_26615,N_26161);
nand U27713 (N_27713,N_27390,N_25287);
or U27714 (N_27714,N_27111,N_25250);
and U27715 (N_27715,N_27208,N_25621);
nand U27716 (N_27716,N_26245,N_25204);
xor U27717 (N_27717,N_25823,N_25803);
xnor U27718 (N_27718,N_25706,N_25061);
or U27719 (N_27719,N_25175,N_25809);
xnor U27720 (N_27720,N_27320,N_26535);
and U27721 (N_27721,N_25894,N_27427);
nor U27722 (N_27722,N_26860,N_27397);
and U27723 (N_27723,N_25378,N_26821);
or U27724 (N_27724,N_25725,N_27207);
xor U27725 (N_27725,N_27165,N_25572);
and U27726 (N_27726,N_26151,N_25904);
nand U27727 (N_27727,N_26391,N_26769);
xor U27728 (N_27728,N_25701,N_25527);
xor U27729 (N_27729,N_25731,N_25573);
xor U27730 (N_27730,N_25074,N_27233);
nor U27731 (N_27731,N_25282,N_26849);
xor U27732 (N_27732,N_25881,N_25167);
or U27733 (N_27733,N_26139,N_25782);
or U27734 (N_27734,N_27410,N_25964);
or U27735 (N_27735,N_25991,N_25211);
or U27736 (N_27736,N_25237,N_26078);
and U27737 (N_27737,N_26101,N_25371);
nor U27738 (N_27738,N_26920,N_25633);
nand U27739 (N_27739,N_27005,N_26511);
xnor U27740 (N_27740,N_26167,N_26567);
and U27741 (N_27741,N_25303,N_25815);
nand U27742 (N_27742,N_25089,N_27211);
nor U27743 (N_27743,N_27138,N_25948);
and U27744 (N_27744,N_26530,N_26771);
nor U27745 (N_27745,N_25736,N_25314);
xnor U27746 (N_27746,N_25181,N_25860);
or U27747 (N_27747,N_27166,N_25663);
and U27748 (N_27748,N_25783,N_26710);
nor U27749 (N_27749,N_26621,N_26914);
and U27750 (N_27750,N_27452,N_27203);
and U27751 (N_27751,N_26584,N_26525);
or U27752 (N_27752,N_25746,N_26395);
nand U27753 (N_27753,N_25922,N_25684);
nand U27754 (N_27754,N_25162,N_27043);
and U27755 (N_27755,N_26036,N_25877);
nand U27756 (N_27756,N_26859,N_26321);
and U27757 (N_27757,N_26073,N_25958);
or U27758 (N_27758,N_26215,N_25519);
nor U27759 (N_27759,N_26738,N_26874);
xor U27760 (N_27760,N_26756,N_25846);
nor U27761 (N_27761,N_26397,N_26802);
xnor U27762 (N_27762,N_26199,N_27377);
and U27763 (N_27763,N_26590,N_25470);
or U27764 (N_27764,N_26127,N_26298);
and U27765 (N_27765,N_25210,N_27380);
nor U27766 (N_27766,N_26097,N_26008);
nand U27767 (N_27767,N_26678,N_25941);
and U27768 (N_27768,N_26398,N_25666);
nand U27769 (N_27769,N_25424,N_25751);
nor U27770 (N_27770,N_25862,N_25221);
and U27771 (N_27771,N_26940,N_25245);
nor U27772 (N_27772,N_25219,N_25130);
nor U27773 (N_27773,N_25889,N_25299);
nand U27774 (N_27774,N_26897,N_27095);
or U27775 (N_27775,N_25500,N_27067);
xor U27776 (N_27776,N_26094,N_26049);
xnor U27777 (N_27777,N_25536,N_26648);
nor U27778 (N_27778,N_26384,N_26162);
or U27779 (N_27779,N_26663,N_25539);
or U27780 (N_27780,N_26720,N_27248);
nand U27781 (N_27781,N_27265,N_25349);
and U27782 (N_27782,N_26573,N_25337);
nor U27783 (N_27783,N_26140,N_26096);
xnor U27784 (N_27784,N_25828,N_25900);
nor U27785 (N_27785,N_25921,N_25589);
and U27786 (N_27786,N_26156,N_26707);
xor U27787 (N_27787,N_26435,N_26116);
xnor U27788 (N_27788,N_25591,N_26458);
nand U27789 (N_27789,N_25592,N_27217);
xor U27790 (N_27790,N_26329,N_26027);
xnor U27791 (N_27791,N_26822,N_25253);
xor U27792 (N_27792,N_25231,N_26104);
nand U27793 (N_27793,N_25220,N_27036);
or U27794 (N_27794,N_25170,N_27023);
nand U27795 (N_27795,N_27308,N_26784);
nand U27796 (N_27796,N_25398,N_26381);
nand U27797 (N_27797,N_26227,N_26893);
nor U27798 (N_27798,N_26136,N_26658);
and U27799 (N_27799,N_25230,N_27475);
xor U27800 (N_27800,N_25792,N_26168);
or U27801 (N_27801,N_27079,N_25467);
or U27802 (N_27802,N_25284,N_26537);
nor U27803 (N_27803,N_26869,N_25522);
or U27804 (N_27804,N_25372,N_25976);
xor U27805 (N_27805,N_25992,N_25920);
nand U27806 (N_27806,N_27028,N_26249);
and U27807 (N_27807,N_26235,N_26134);
xnor U27808 (N_27808,N_25272,N_25132);
xnor U27809 (N_27809,N_25296,N_26277);
or U27810 (N_27810,N_26295,N_26423);
xor U27811 (N_27811,N_27008,N_25872);
xor U27812 (N_27812,N_26000,N_25270);
or U27813 (N_27813,N_27241,N_25242);
xor U27814 (N_27814,N_25916,N_26301);
xor U27815 (N_27815,N_25114,N_26150);
and U27816 (N_27816,N_27112,N_26432);
xnor U27817 (N_27817,N_25086,N_25787);
nor U27818 (N_27818,N_25884,N_26587);
or U27819 (N_27819,N_26106,N_25311);
nor U27820 (N_27820,N_25046,N_27432);
nor U27821 (N_27821,N_25631,N_25854);
xnor U27822 (N_27822,N_26732,N_27342);
nand U27823 (N_27823,N_25188,N_26239);
nand U27824 (N_27824,N_26504,N_27465);
xor U27825 (N_27825,N_25791,N_26200);
nor U27826 (N_27826,N_26740,N_27306);
xor U27827 (N_27827,N_26544,N_26135);
and U27828 (N_27828,N_27351,N_27292);
and U27829 (N_27829,N_25843,N_25355);
or U27830 (N_27830,N_26280,N_27194);
nand U27831 (N_27831,N_25538,N_27414);
nor U27832 (N_27832,N_26425,N_26138);
or U27833 (N_27833,N_25603,N_26481);
and U27834 (N_27834,N_27356,N_25168);
nand U27835 (N_27835,N_26994,N_25544);
or U27836 (N_27836,N_26734,N_25687);
xnor U27837 (N_27837,N_25325,N_25883);
or U27838 (N_27838,N_26050,N_26089);
and U27839 (N_27839,N_27012,N_27403);
or U27840 (N_27840,N_25475,N_26322);
xnor U27841 (N_27841,N_27285,N_27343);
and U27842 (N_27842,N_26196,N_25720);
xnor U27843 (N_27843,N_26591,N_26713);
and U27844 (N_27844,N_25381,N_26833);
and U27845 (N_27845,N_25807,N_26124);
nor U27846 (N_27846,N_26024,N_27484);
xor U27847 (N_27847,N_26317,N_27024);
and U27848 (N_27848,N_25658,N_26081);
xor U27849 (N_27849,N_25507,N_26194);
nor U27850 (N_27850,N_25585,N_26716);
nor U27851 (N_27851,N_25345,N_27362);
or U27852 (N_27852,N_26131,N_25575);
xnor U27853 (N_27853,N_27176,N_26468);
nor U27854 (N_27854,N_26001,N_25485);
and U27855 (N_27855,N_25202,N_27060);
xnor U27856 (N_27856,N_27270,N_26160);
nand U27857 (N_27857,N_26467,N_25052);
or U27858 (N_27858,N_27137,N_26493);
nor U27859 (N_27859,N_25865,N_25838);
and U27860 (N_27860,N_26892,N_26925);
nor U27861 (N_27861,N_25626,N_26788);
nor U27862 (N_27862,N_26533,N_25288);
or U27863 (N_27863,N_27064,N_25885);
and U27864 (N_27864,N_25917,N_25614);
and U27865 (N_27865,N_26017,N_26755);
or U27866 (N_27866,N_27026,N_26618);
nor U27867 (N_27867,N_25360,N_25223);
or U27868 (N_27868,N_25962,N_27161);
or U27869 (N_27869,N_25705,N_26045);
nand U27870 (N_27870,N_26065,N_25552);
and U27871 (N_27871,N_27379,N_26273);
xnor U27872 (N_27872,N_26413,N_25268);
xor U27873 (N_27873,N_26717,N_27297);
nand U27874 (N_27874,N_27142,N_25906);
nand U27875 (N_27875,N_27467,N_26582);
or U27876 (N_27876,N_26886,N_25554);
nand U27877 (N_27877,N_25334,N_25058);
or U27878 (N_27878,N_27085,N_26931);
or U27879 (N_27879,N_25359,N_26466);
and U27880 (N_27880,N_27228,N_25463);
or U27881 (N_27881,N_26832,N_25399);
or U27882 (N_27882,N_27435,N_25344);
nand U27883 (N_27883,N_27476,N_25260);
or U27884 (N_27884,N_26477,N_25149);
or U27885 (N_27885,N_26806,N_25456);
nand U27886 (N_27886,N_25674,N_25307);
nand U27887 (N_27887,N_26676,N_25209);
nor U27888 (N_27888,N_25739,N_25429);
or U27889 (N_27889,N_27280,N_25172);
xor U27890 (N_27890,N_26471,N_26709);
and U27891 (N_27891,N_26747,N_25932);
nor U27892 (N_27892,N_27464,N_25207);
nor U27893 (N_27893,N_26986,N_26129);
nand U27894 (N_27894,N_26170,N_26163);
xor U27895 (N_27895,N_26723,N_27020);
nor U27896 (N_27896,N_27068,N_26332);
and U27897 (N_27897,N_25668,N_25145);
and U27898 (N_27898,N_25102,N_26444);
nor U27899 (N_27899,N_25933,N_27129);
xnor U27900 (N_27900,N_27093,N_26282);
or U27901 (N_27901,N_25949,N_26440);
nand U27902 (N_27902,N_25280,N_27056);
xnor U27903 (N_27903,N_26921,N_26727);
nor U27904 (N_27904,N_26007,N_25002);
xor U27905 (N_27905,N_27335,N_26452);
or U27906 (N_27906,N_26169,N_26463);
and U27907 (N_27907,N_25630,N_27473);
and U27908 (N_27908,N_25190,N_27175);
or U27909 (N_27909,N_26218,N_26792);
nor U27910 (N_27910,N_26677,N_26984);
xnor U27911 (N_27911,N_27100,N_26040);
or U27912 (N_27912,N_26207,N_26339);
xor U27913 (N_27913,N_25648,N_25514);
xor U27914 (N_27914,N_25693,N_25959);
nand U27915 (N_27915,N_26636,N_25254);
nor U27916 (N_27916,N_26421,N_27013);
nand U27917 (N_27917,N_26900,N_25034);
xnor U27918 (N_27918,N_25714,N_26119);
xnor U27919 (N_27919,N_26480,N_25512);
and U27920 (N_27920,N_25274,N_26177);
nand U27921 (N_27921,N_25710,N_26128);
nor U27922 (N_27922,N_25407,N_25721);
nand U27923 (N_27923,N_25200,N_25400);
nand U27924 (N_27924,N_25076,N_25745);
nand U27925 (N_27925,N_26674,N_27132);
or U27926 (N_27926,N_26538,N_27183);
and U27927 (N_27927,N_25135,N_25899);
nand U27928 (N_27928,N_27075,N_25117);
xor U27929 (N_27929,N_26029,N_27259);
nor U27930 (N_27930,N_25859,N_26403);
nand U27931 (N_27931,N_25806,N_25306);
and U27932 (N_27932,N_26363,N_25396);
nand U27933 (N_27933,N_25908,N_26289);
nor U27934 (N_27934,N_27499,N_26743);
and U27935 (N_27935,N_25696,N_27196);
nand U27936 (N_27936,N_25704,N_27469);
xnor U27937 (N_27937,N_26345,N_25688);
nor U27938 (N_27938,N_26872,N_25163);
nor U27939 (N_27939,N_26730,N_26342);
nor U27940 (N_27940,N_25795,N_25940);
xnor U27941 (N_27941,N_25418,N_27096);
and U27942 (N_27942,N_27300,N_25331);
or U27943 (N_27943,N_26523,N_25983);
or U27944 (N_27944,N_25645,N_25030);
xnor U27945 (N_27945,N_26505,N_25414);
xnor U27946 (N_27946,N_26086,N_25780);
nand U27947 (N_27947,N_25003,N_25808);
xor U27948 (N_27948,N_25386,N_25081);
nand U27949 (N_27949,N_26323,N_27378);
or U27950 (N_27950,N_26402,N_25001);
nand U27951 (N_27951,N_25097,N_25196);
or U27952 (N_27952,N_27030,N_27443);
or U27953 (N_27953,N_25871,N_26944);
nor U27954 (N_27954,N_26148,N_25036);
nor U27955 (N_27955,N_27349,N_25981);
and U27956 (N_27956,N_27257,N_26149);
nor U27957 (N_27957,N_26915,N_27450);
xnor U27958 (N_27958,N_27099,N_25878);
nand U27959 (N_27959,N_25064,N_27059);
nor U27960 (N_27960,N_25169,N_25087);
xnor U27961 (N_27961,N_26913,N_25758);
nor U27962 (N_27962,N_26246,N_25643);
xor U27963 (N_27963,N_26310,N_25029);
nor U27964 (N_27964,N_27092,N_27219);
nand U27965 (N_27965,N_26074,N_25419);
nand U27966 (N_27966,N_25116,N_26222);
nand U27967 (N_27967,N_25586,N_25310);
and U27968 (N_27968,N_25655,N_27345);
xnor U27969 (N_27969,N_26928,N_27027);
nand U27970 (N_27970,N_27167,N_25761);
xor U27971 (N_27971,N_25121,N_26616);
and U27972 (N_27972,N_26241,N_25489);
or U27973 (N_27973,N_26093,N_27163);
nor U27974 (N_27974,N_25499,N_27131);
nand U27975 (N_27975,N_27368,N_26839);
nand U27976 (N_27976,N_25839,N_25157);
nor U27977 (N_27977,N_27105,N_25763);
nor U27978 (N_27978,N_26608,N_26887);
or U27979 (N_27979,N_26059,N_26642);
nand U27980 (N_27980,N_26229,N_25447);
xnor U27981 (N_27981,N_26197,N_25583);
and U27982 (N_27982,N_25380,N_25283);
nor U27983 (N_27983,N_25907,N_27054);
or U27984 (N_27984,N_26385,N_26905);
and U27985 (N_27985,N_25411,N_25953);
nor U27986 (N_27986,N_25265,N_27402);
and U27987 (N_27987,N_25252,N_26341);
xnor U27988 (N_27988,N_25647,N_27455);
nor U27989 (N_27989,N_25752,N_27472);
nand U27990 (N_27990,N_27210,N_25576);
nor U27991 (N_27991,N_26380,N_27303);
and U27992 (N_27992,N_27389,N_26520);
nor U27993 (N_27993,N_25829,N_26333);
nor U27994 (N_27994,N_27304,N_25484);
or U27995 (N_27995,N_26878,N_25309);
nand U27996 (N_27996,N_27318,N_27359);
nor U27997 (N_27997,N_27152,N_26396);
or U27998 (N_27998,N_26154,N_25348);
xor U27999 (N_27999,N_27405,N_26653);
or U28000 (N_28000,N_25890,N_27287);
nand U28001 (N_28001,N_26698,N_26060);
nand U28002 (N_28002,N_25497,N_27206);
nand U28003 (N_28003,N_27245,N_26754);
xnor U28004 (N_28004,N_26401,N_25461);
xnor U28005 (N_28005,N_27492,N_26693);
xor U28006 (N_28006,N_25343,N_25887);
and U28007 (N_28007,N_26367,N_25770);
nor U28008 (N_28008,N_26419,N_26996);
nor U28009 (N_28009,N_25753,N_26637);
xor U28010 (N_28010,N_25328,N_26314);
xor U28011 (N_28011,N_25613,N_26216);
nor U28012 (N_28012,N_26908,N_25678);
or U28013 (N_28013,N_26682,N_26517);
nor U28014 (N_28014,N_26880,N_25619);
nand U28015 (N_28015,N_25570,N_26665);
xor U28016 (N_28016,N_25213,N_25154);
nand U28017 (N_28017,N_25518,N_25147);
xnor U28018 (N_28018,N_25390,N_27216);
and U28019 (N_28019,N_26669,N_27136);
nor U28020 (N_28020,N_25711,N_26588);
nor U28021 (N_28021,N_25960,N_26371);
nand U28022 (N_28022,N_25476,N_26805);
xor U28023 (N_28023,N_25733,N_25841);
and U28024 (N_28024,N_26361,N_26267);
nand U28025 (N_28025,N_27232,N_25366);
or U28026 (N_28026,N_27276,N_26153);
or U28027 (N_28027,N_26808,N_27007);
nand U28028 (N_28028,N_26250,N_26386);
nor U28029 (N_28029,N_27202,N_25161);
nand U28030 (N_28030,N_27261,N_26120);
xor U28031 (N_28031,N_26230,N_25016);
nand U28032 (N_28032,N_26491,N_25897);
or U28033 (N_28033,N_25356,N_25931);
nand U28034 (N_28034,N_26930,N_25620);
or U28035 (N_28035,N_27252,N_25082);
xor U28036 (N_28036,N_26820,N_25316);
or U28037 (N_28037,N_26909,N_25212);
nor U28038 (N_28038,N_26354,N_25850);
nor U28039 (N_28039,N_25954,N_25071);
and U28040 (N_28040,N_25238,N_25395);
and U28041 (N_28041,N_25143,N_25672);
nor U28042 (N_28042,N_27323,N_26999);
and U28043 (N_28043,N_25448,N_27083);
nor U28044 (N_28044,N_26943,N_26980);
nand U28045 (N_28045,N_26415,N_26753);
and U28046 (N_28046,N_25649,N_25208);
and U28047 (N_28047,N_25697,N_25724);
nand U28048 (N_28048,N_26546,N_26761);
xnor U28049 (N_28049,N_25150,N_27423);
xor U28050 (N_28050,N_25261,N_26217);
xor U28051 (N_28051,N_26276,N_25443);
xnor U28052 (N_28052,N_27065,N_25851);
nand U28053 (N_28053,N_26502,N_25234);
xor U28054 (N_28054,N_25557,N_25290);
nor U28055 (N_28055,N_26843,N_27051);
and U28056 (N_28056,N_27352,N_25335);
xnor U28057 (N_28057,N_26848,N_26411);
and U28058 (N_28058,N_27029,N_25302);
nor U28059 (N_28059,N_26935,N_25653);
nor U28060 (N_28060,N_26319,N_25955);
xnor U28061 (N_28061,N_26064,N_25618);
or U28062 (N_28062,N_27310,N_25070);
nand U28063 (N_28063,N_26870,N_26126);
nor U28064 (N_28064,N_27184,N_25529);
xor U28065 (N_28065,N_27109,N_27220);
or U28066 (N_28066,N_25743,N_27296);
xnor U28067 (N_28067,N_27062,N_25821);
and U28068 (N_28068,N_26494,N_26646);
nor U28069 (N_28069,N_27491,N_25875);
nor U28070 (N_28070,N_25660,N_27258);
xor U28071 (N_28071,N_27477,N_27048);
nand U28072 (N_28072,N_26801,N_26509);
nand U28073 (N_28073,N_25873,N_25560);
nor U28074 (N_28074,N_27003,N_25413);
xor U28075 (N_28075,N_26003,N_25000);
nand U28076 (N_28076,N_26021,N_26302);
nand U28077 (N_28077,N_27186,N_26831);
nand U28078 (N_28078,N_25651,N_25085);
nand U28079 (N_28079,N_25737,N_27034);
or U28080 (N_28080,N_25490,N_25055);
nor U28081 (N_28081,N_26764,N_26692);
or U28082 (N_28082,N_27237,N_25579);
or U28083 (N_28083,N_25768,N_26946);
xnor U28084 (N_28084,N_26703,N_25641);
and U28085 (N_28085,N_27145,N_25189);
nor U28086 (N_28086,N_26779,N_26516);
and U28087 (N_28087,N_26146,N_26840);
xnor U28088 (N_28088,N_25158,N_27074);
nor U28089 (N_28089,N_25151,N_25818);
nor U28090 (N_28090,N_25847,N_26842);
or U28091 (N_28091,N_27250,N_25845);
nand U28092 (N_28092,N_25246,N_27178);
xnor U28093 (N_28093,N_25805,N_25927);
and U28094 (N_28094,N_25075,N_25879);
and U28095 (N_28095,N_25528,N_27339);
xor U28096 (N_28096,N_25100,N_26475);
nor U28097 (N_28097,N_25129,N_27153);
nand U28098 (N_28098,N_26180,N_25650);
nand U28099 (N_28099,N_25377,N_27084);
nand U28100 (N_28100,N_25415,N_27033);
xnor U28101 (N_28101,N_26457,N_25365);
nand U28102 (N_28102,N_26026,N_27459);
xor U28103 (N_28103,N_25867,N_25556);
nand U28104 (N_28104,N_25664,N_26079);
and U28105 (N_28105,N_27360,N_25623);
xor U28106 (N_28106,N_25910,N_26962);
xor U28107 (N_28107,N_27017,N_27089);
or U28108 (N_28108,N_25794,N_25496);
or U28109 (N_28109,N_25341,N_26661);
xor U28110 (N_28110,N_25346,N_26807);
xnor U28111 (N_28111,N_25186,N_26752);
nor U28112 (N_28112,N_25382,N_26791);
and U28113 (N_28113,N_26953,N_25919);
and U28114 (N_28114,N_25298,N_25712);
and U28115 (N_28115,N_27147,N_25543);
or U28116 (N_28116,N_26417,N_27324);
nor U28117 (N_28117,N_26688,N_25263);
and U28118 (N_28118,N_25133,N_27421);
xor U28119 (N_28119,N_25480,N_26088);
or U28120 (N_28120,N_26508,N_27236);
nor U28121 (N_28121,N_25057,N_25027);
nand U28122 (N_28122,N_26011,N_25708);
and U28123 (N_28123,N_25194,N_27282);
nor U28124 (N_28124,N_26173,N_25009);
xnor U28125 (N_28125,N_26054,N_26643);
nand U28126 (N_28126,N_26577,N_25819);
or U28127 (N_28127,N_26850,N_25079);
nand U28128 (N_28128,N_26513,N_26279);
and U28129 (N_28129,N_26609,N_27321);
or U28130 (N_28130,N_25893,N_26344);
nor U28131 (N_28131,N_27144,N_25673);
nand U28132 (N_28132,N_25468,N_25164);
and U28133 (N_28133,N_26702,N_25442);
nor U28134 (N_28134,N_26496,N_27069);
xor U28135 (N_28135,N_26632,N_25627);
or U28136 (N_28136,N_26208,N_26865);
nor U28137 (N_28137,N_27187,N_27021);
and U28138 (N_28138,N_26296,N_26350);
xnor U28139 (N_28139,N_26631,N_26325);
nor U28140 (N_28140,N_27382,N_25184);
and U28141 (N_28141,N_27180,N_26911);
and U28142 (N_28142,N_25312,N_26768);
nand U28143 (N_28143,N_27260,N_25692);
xnor U28144 (N_28144,N_26600,N_25773);
nor U28145 (N_28145,N_26890,N_27407);
or U28146 (N_28146,N_25977,N_25562);
and U28147 (N_28147,N_25938,N_26759);
xor U28148 (N_28148,N_26959,N_26916);
xnor U28149 (N_28149,N_27272,N_27334);
and U28150 (N_28150,N_26773,N_26318);
xor U28151 (N_28151,N_27418,N_25587);
nand U28152 (N_28152,N_26453,N_27073);
nand U28153 (N_28153,N_26014,N_25059);
nor U28154 (N_28154,N_27081,N_25713);
nor U28155 (N_28155,N_26681,N_26826);
nand U28156 (N_28156,N_25266,N_25279);
nand U28157 (N_28157,N_27193,N_26647);
nand U28158 (N_28158,N_26006,N_25956);
nand U28159 (N_28159,N_26778,N_27354);
or U28160 (N_28160,N_26777,N_26795);
or U28161 (N_28161,N_26718,N_25065);
or U28162 (N_28162,N_25896,N_27271);
nor U28163 (N_28163,N_26596,N_27169);
and U28164 (N_28164,N_26899,N_25393);
and U28165 (N_28165,N_25134,N_25993);
and U28166 (N_28166,N_26225,N_26627);
xor U28167 (N_28167,N_26599,N_26654);
and U28168 (N_28168,N_25798,N_25142);
or U28169 (N_28169,N_25313,N_26861);
and U28170 (N_28170,N_26668,N_26272);
nand U28171 (N_28171,N_26234,N_26474);
xnor U28172 (N_28172,N_25551,N_26972);
nor U28173 (N_28173,N_26087,N_25239);
nand U28174 (N_28174,N_27456,N_26657);
and U28175 (N_28175,N_26428,N_27239);
or U28176 (N_28176,N_26903,N_25123);
xor U28177 (N_28177,N_25358,N_26534);
nor U28178 (N_28178,N_27370,N_25032);
or U28179 (N_28179,N_25362,N_27348);
xnor U28180 (N_28180,N_26490,N_26560);
nand U28181 (N_28181,N_26845,N_25426);
and U28182 (N_28182,N_25493,N_26610);
or U28183 (N_28183,N_25037,N_25462);
nor U28184 (N_28184,N_25856,N_27190);
nor U28185 (N_28185,N_26519,N_26041);
and U28186 (N_28186,N_25324,N_26247);
nor U28187 (N_28187,N_25436,N_25837);
nor U28188 (N_28188,N_25165,N_26451);
and U28189 (N_28189,N_27243,N_25217);
xnor U28190 (N_28190,N_25546,N_26512);
nor U28191 (N_28191,N_26090,N_25469);
and U28192 (N_28192,N_27289,N_26110);
nor U28193 (N_28193,N_25374,N_25218);
nand U28194 (N_28194,N_27224,N_27438);
nor U28195 (N_28195,N_27387,N_26358);
xnor U28196 (N_28196,N_26137,N_25596);
and U28197 (N_28197,N_26547,N_26563);
or U28198 (N_28198,N_26503,N_26793);
nor U28199 (N_28199,N_25275,N_26963);
or U28200 (N_28200,N_25892,N_26383);
and U28201 (N_28201,N_26443,N_26896);
xor U28202 (N_28202,N_27022,N_25425);
or U28203 (N_28203,N_26855,N_25486);
xnor U28204 (N_28204,N_26815,N_26192);
nor U28205 (N_28205,N_25781,N_27114);
or U28206 (N_28206,N_26351,N_25963);
nor U28207 (N_28207,N_26448,N_26379);
and U28208 (N_28208,N_27269,N_25822);
and U28209 (N_28209,N_26557,N_27274);
or U28210 (N_28210,N_25568,N_26299);
xor U28211 (N_28211,N_25637,N_25495);
nand U28212 (N_28212,N_26284,N_26543);
nand U28213 (N_28213,N_27140,N_25549);
nand U28214 (N_28214,N_26092,N_25698);
xnor U28215 (N_28215,N_26420,N_26377);
nor U28216 (N_28216,N_25691,N_25640);
or U28217 (N_28217,N_25700,N_26775);
nand U28218 (N_28218,N_25481,N_26252);
nor U28219 (N_28219,N_27281,N_26257);
nor U28220 (N_28220,N_26500,N_26240);
and U28221 (N_28221,N_25205,N_25939);
and U28222 (N_28222,N_26955,N_27185);
nand U28223 (N_28223,N_25813,N_27277);
xnor U28224 (N_28224,N_27444,N_26326);
nor U28225 (N_28225,N_25686,N_27284);
nand U28226 (N_28226,N_27383,N_26725);
and U28227 (N_28227,N_26067,N_25777);
and U28228 (N_28228,N_26028,N_25183);
nand U28229 (N_28229,N_27468,N_26565);
nor U28230 (N_28230,N_26214,N_26739);
xnor U28231 (N_28231,N_25728,N_27409);
and U28232 (N_28232,N_26125,N_27489);
and U28233 (N_28233,N_25319,N_27433);
xor U28234 (N_28234,N_26998,N_26945);
xnor U28235 (N_28235,N_26548,N_27097);
xor U28236 (N_28236,N_26597,N_25975);
or U28237 (N_28237,N_25604,N_27376);
nand U28238 (N_28238,N_26731,N_26598);
or U28239 (N_28239,N_27355,N_26864);
nand U28240 (N_28240,N_26568,N_25391);
and U28241 (N_28241,N_25293,N_25054);
or U28242 (N_28242,N_25584,N_25545);
and U28243 (N_28243,N_26300,N_26796);
xnor U28244 (N_28244,N_26924,N_25073);
or U28245 (N_28245,N_25715,N_26365);
nand U28246 (N_28246,N_27408,N_26527);
or U28247 (N_28247,N_26827,N_25445);
or U28248 (N_28248,N_25322,N_25128);
nand U28249 (N_28249,N_25327,N_27426);
nand U28250 (N_28250,N_25582,N_27374);
xnor U28251 (N_28251,N_27098,N_25363);
and U28252 (N_28252,N_25352,N_26545);
xnor U28253 (N_28253,N_25774,N_25607);
or U28254 (N_28254,N_25126,N_27212);
or U28255 (N_28255,N_27428,N_25137);
xnor U28256 (N_28256,N_27437,N_25612);
or U28257 (N_28257,N_25379,N_25364);
or U28258 (N_28258,N_26030,N_26918);
and U28259 (N_28259,N_25051,N_25244);
xor U28260 (N_28260,N_27118,N_26617);
and U28261 (N_28261,N_27416,N_25454);
or U28262 (N_28262,N_27159,N_27340);
nand U28263 (N_28263,N_26910,N_25778);
and U28264 (N_28264,N_25329,N_26407);
nand U28265 (N_28265,N_25056,N_26714);
nor U28266 (N_28266,N_25508,N_25115);
and U28267 (N_28267,N_27133,N_27204);
xnor U28268 (N_28268,N_25722,N_25567);
nor U28269 (N_28269,N_26290,N_25600);
nand U28270 (N_28270,N_26076,N_27135);
or U28271 (N_28271,N_26012,N_27120);
or U28272 (N_28272,N_25905,N_25759);
or U28273 (N_28273,N_26797,N_25531);
and U28274 (N_28274,N_25503,N_26112);
or U28275 (N_28275,N_25332,N_25719);
nor U28276 (N_28276,N_25451,N_25180);
or U28277 (N_28277,N_26607,N_26238);
nand U28278 (N_28278,N_25734,N_27466);
and U28279 (N_28279,N_26459,N_26708);
xnor U28280 (N_28280,N_25339,N_26659);
nor U28281 (N_28281,N_25417,N_27160);
nor U28282 (N_28282,N_26844,N_26408);
nor U28283 (N_28283,N_26901,N_25654);
nand U28284 (N_28284,N_26576,N_25748);
or U28285 (N_28285,N_25656,N_25835);
nor U28286 (N_28286,N_27197,N_25775);
or U28287 (N_28287,N_26514,N_26780);
nand U28288 (N_28288,N_25923,N_26695);
and U28289 (N_28289,N_26589,N_26551);
or U28290 (N_28290,N_25853,N_25972);
nand U28291 (N_28291,N_27336,N_25646);
and U28292 (N_28292,N_25833,N_25083);
nand U28293 (N_28293,N_25825,N_25915);
or U28294 (N_28294,N_26737,N_25942);
and U28295 (N_28295,N_27251,N_26460);
nor U28296 (N_28296,N_26331,N_25537);
or U28297 (N_28297,N_26271,N_25318);
or U28298 (N_28298,N_27319,N_25155);
or U28299 (N_28299,N_26231,N_26085);
or U28300 (N_28300,N_26187,N_27311);
or U28301 (N_28301,N_27357,N_27317);
or U28302 (N_28302,N_25671,N_26671);
nor U28303 (N_28303,N_25968,N_26364);
xor U28304 (N_28304,N_26781,N_26004);
or U28305 (N_28305,N_27229,N_25804);
or U28306 (N_28306,N_26510,N_25961);
or U28307 (N_28307,N_26895,N_26578);
xor U28308 (N_28308,N_26293,N_25353);
xor U28309 (N_28309,N_25232,N_25577);
or U28310 (N_28310,N_25375,N_27122);
or U28311 (N_28311,N_26823,N_25243);
and U28312 (N_28312,N_26410,N_25148);
nor U28313 (N_28313,N_25440,N_26063);
nand U28314 (N_28314,N_27441,N_26429);
nand U28315 (N_28315,N_26786,N_27156);
and U28316 (N_28316,N_27448,N_25980);
xnor U28317 (N_28317,N_27009,N_27148);
nand U28318 (N_28318,N_25521,N_25944);
nand U28319 (N_28319,N_25354,N_25038);
nand U28320 (N_28320,N_25861,N_27487);
nor U28321 (N_28321,N_26035,N_26696);
xor U28322 (N_28322,N_26013,N_25125);
xnor U28323 (N_28323,N_25294,N_25842);
or U28324 (N_28324,N_26794,N_26152);
nor U28325 (N_28325,N_26664,N_25525);
nand U28326 (N_28326,N_26883,N_27255);
or U28327 (N_28327,N_26515,N_26952);
xnor U28328 (N_28328,N_26729,N_26360);
xnor U28329 (N_28329,N_26539,N_25067);
nor U28330 (N_28330,N_27182,N_26626);
and U28331 (N_28331,N_27246,N_25988);
xor U28332 (N_28332,N_26369,N_25515);
xnor U28333 (N_28333,N_26982,N_26461);
or U28334 (N_28334,N_26876,N_26052);
and U28335 (N_28335,N_26330,N_26171);
or U28336 (N_28336,N_25473,N_25095);
or U28337 (N_28337,N_26558,N_26478);
nand U28338 (N_28338,N_27449,N_26721);
and U28339 (N_28339,N_26016,N_25432);
or U28340 (N_28340,N_25141,N_25924);
and U28341 (N_28341,N_26603,N_25574);
nor U28342 (N_28342,N_27025,N_25869);
or U28343 (N_28343,N_27478,N_27412);
and U28344 (N_28344,N_25855,N_25624);
nand U28345 (N_28345,N_26812,N_26974);
and U28346 (N_28346,N_25999,N_25995);
or U28347 (N_28347,N_27200,N_27278);
or U28348 (N_28348,N_26745,N_27366);
or U28349 (N_28349,N_25119,N_26929);
or U28350 (N_28350,N_26991,N_25421);
xnor U28351 (N_28351,N_26205,N_25937);
and U28352 (N_28352,N_25227,N_26285);
and U28353 (N_28353,N_27453,N_26305);
or U28354 (N_28354,N_26536,N_26937);
nand U28355 (N_28355,N_25558,N_27128);
nor U28356 (N_28356,N_27226,N_25581);
and U28357 (N_28357,N_25068,N_27171);
nor U28358 (N_28358,N_25397,N_26912);
nand U28359 (N_28359,N_26989,N_25043);
and U28360 (N_28360,N_26018,N_26988);
and U28361 (N_28361,N_25509,N_27116);
nand U28362 (N_28362,N_27002,N_26532);
xnor U28363 (N_28363,N_25913,N_25601);
nand U28364 (N_28364,N_25048,N_26473);
nand U28365 (N_28365,N_25477,N_25041);
and U28366 (N_28366,N_26479,N_25947);
nand U28367 (N_28367,N_27385,N_25685);
nand U28368 (N_28368,N_25802,N_25498);
or U28369 (N_28369,N_25021,N_26370);
and U28370 (N_28370,N_26656,N_25247);
xnor U28371 (N_28371,N_26133,N_26570);
and U28372 (N_28372,N_26286,N_27143);
xor U28373 (N_28373,N_26762,N_27141);
and U28374 (N_28374,N_26613,N_27038);
nor U28375 (N_28375,N_26680,N_26212);
nor U28376 (N_28376,N_27315,N_26633);
or U28377 (N_28377,N_26851,N_25695);
or U28378 (N_28378,N_26486,N_27486);
nand U28379 (N_28379,N_25383,N_27493);
and U28380 (N_28380,N_25361,N_26704);
xor U28381 (N_28381,N_25547,N_25796);
and U28382 (N_28382,N_26967,N_25741);
or U28383 (N_28383,N_26080,N_25540);
and U28384 (N_28384,N_26056,N_25044);
xnor U28385 (N_28385,N_25505,N_26185);
nand U28386 (N_28386,N_27337,N_26303);
nand U28387 (N_28387,N_26809,N_26265);
and U28388 (N_28388,N_26635,N_25965);
and U28389 (N_28389,N_27125,N_27019);
nand U28390 (N_28390,N_25667,N_26122);
xnor U28391 (N_28391,N_27327,N_26082);
nor U28392 (N_28392,N_25347,N_25098);
nand U28393 (N_28393,N_25289,N_25982);
nand U28394 (N_28394,N_27222,N_27358);
xnor U28395 (N_28395,N_25320,N_26447);
or U28396 (N_28396,N_25762,N_26061);
nand U28397 (N_28397,N_26437,N_25216);
and U28398 (N_28398,N_25022,N_25277);
nor U28399 (N_28399,N_25608,N_26906);
or U28400 (N_28400,N_25182,N_25139);
nand U28401 (N_28401,N_25422,N_26705);
nor U28402 (N_28402,N_26957,N_26414);
nor U28403 (N_28403,N_25094,N_26356);
and U28404 (N_28404,N_25308,N_26694);
nor U28405 (N_28405,N_27480,N_26581);
xor U28406 (N_28406,N_26552,N_27328);
or U28407 (N_28407,N_26366,N_26102);
nand U28408 (N_28408,N_25106,N_26683);
or U28409 (N_28409,N_27325,N_26830);
xor U28410 (N_28410,N_26835,N_25446);
nand U28411 (N_28411,N_26347,N_27275);
or U28412 (N_28412,N_25998,N_27082);
and U28413 (N_28413,N_26592,N_26158);
and U28414 (N_28414,N_25450,N_25101);
and U28415 (N_28415,N_26799,N_25952);
nand U28416 (N_28416,N_27044,N_26877);
and U28417 (N_28417,N_27055,N_26736);
nor U28418 (N_28418,N_27495,N_26340);
nor U28419 (N_28419,N_26232,N_26472);
nor U28420 (N_28420,N_25590,N_27058);
or U28421 (N_28421,N_27121,N_25008);
and U28422 (N_28422,N_26195,N_25832);
and U28423 (N_28423,N_25676,N_26614);
or U28424 (N_28424,N_25482,N_26554);
or U28425 (N_28425,N_26334,N_26580);
and U28426 (N_28426,N_26891,N_27279);
nand U28427 (N_28427,N_27179,N_27032);
nor U28428 (N_28428,N_25717,N_26749);
nor U28429 (N_28429,N_26183,N_26629);
xor U28430 (N_28430,N_26605,N_25793);
or U28431 (N_28431,N_26072,N_27151);
and U28432 (N_28432,N_25273,N_25249);
and U28433 (N_28433,N_25814,N_26970);
nand U28434 (N_28434,N_25483,N_25014);
or U28435 (N_28435,N_27052,N_25925);
nand U28436 (N_28436,N_27344,N_25104);
nor U28437 (N_28437,N_26939,N_27041);
and U28438 (N_28438,N_26147,N_26651);
nor U28439 (N_28439,N_25502,N_27119);
or U28440 (N_28440,N_25659,N_25726);
nand U28441 (N_28441,N_25742,N_25857);
nor U28442 (N_28442,N_26561,N_25258);
xor U28443 (N_28443,N_25078,N_26619);
or U28444 (N_28444,N_27309,N_27091);
nor U28445 (N_28445,N_25790,N_25632);
and U28446 (N_28446,N_26174,N_25053);
and U28447 (N_28447,N_27149,N_27442);
nor U28448 (N_28448,N_26881,N_25107);
xor U28449 (N_28449,N_27305,N_26917);
nor U28450 (N_28450,N_25914,N_25786);
or U28451 (N_28451,N_25176,N_26445);
and U28452 (N_28452,N_26025,N_25727);
or U28453 (N_28453,N_27247,N_26224);
nand U28454 (N_28454,N_27070,N_25766);
nor U28455 (N_28455,N_26105,N_25338);
xnor U28456 (N_28456,N_26113,N_25019);
nor U28457 (N_28457,N_26593,N_25215);
nand U28458 (N_28458,N_27263,N_26433);
xnor U28459 (N_28459,N_26497,N_26489);
and U28460 (N_28460,N_25330,N_27312);
nand U28461 (N_28461,N_27006,N_26838);
xor U28462 (N_28462,N_26868,N_25526);
nor U28463 (N_28463,N_25433,N_25384);
nor U28464 (N_28464,N_26051,N_26098);
nand U28465 (N_28465,N_26312,N_26766);
xor U28466 (N_28466,N_25863,N_27381);
or U28467 (N_28467,N_26611,N_27283);
or U28468 (N_28468,N_25122,N_26157);
xnor U28469 (N_28469,N_26254,N_27401);
or U28470 (N_28470,N_26846,N_25852);
and U28471 (N_28471,N_26522,N_25262);
xor U28472 (N_28472,N_26042,N_26053);
or U28473 (N_28473,N_25978,N_26237);
nor U28474 (N_28474,N_26706,N_25241);
nand U28475 (N_28475,N_26034,N_25236);
or U28476 (N_28476,N_27294,N_27049);
nand U28477 (N_28477,N_26374,N_27440);
nor U28478 (N_28478,N_25171,N_25013);
and U28479 (N_28479,N_27436,N_25351);
xnor U28480 (N_28480,N_25888,N_26166);
nand U28481 (N_28481,N_25156,N_27076);
nor U28482 (N_28482,N_26288,N_26172);
nor U28483 (N_28483,N_26043,N_25011);
nand U28484 (N_28484,N_25764,N_27400);
nor U28485 (N_28485,N_25235,N_26349);
and U28486 (N_28486,N_26606,N_26602);
or U28487 (N_28487,N_25096,N_27189);
nor U28488 (N_28488,N_25749,N_26039);
or U28489 (N_28489,N_26853,N_26660);
xnor U28490 (N_28490,N_26455,N_27494);
nor U28491 (N_28491,N_27425,N_25681);
and U28492 (N_28492,N_25410,N_26979);
nand U28493 (N_28493,N_25740,N_25834);
or U28494 (N_28494,N_26987,N_27235);
nor U28495 (N_28495,N_25012,N_27483);
nor U28496 (N_28496,N_26662,N_25513);
and U28497 (N_28497,N_26862,N_26142);
xnor U28498 (N_28498,N_26644,N_26292);
nor U28499 (N_28499,N_27498,N_25321);
or U28500 (N_28500,N_25902,N_27363);
nand U28501 (N_28501,N_27286,N_26524);
nand U28502 (N_28502,N_26211,N_26203);
nand U28503 (N_28503,N_25634,N_25635);
nand U28504 (N_28504,N_26518,N_26858);
xor U28505 (N_28505,N_26223,N_26894);
and U28506 (N_28506,N_26346,N_25858);
and U28507 (N_28507,N_25459,N_25610);
or U28508 (N_28508,N_25146,N_25039);
or U28509 (N_28509,N_25430,N_26390);
xnor U28510 (N_28510,N_25760,N_25240);
nor U28511 (N_28511,N_27238,N_27162);
nor U28512 (N_28512,N_25326,N_25826);
or U28513 (N_28513,N_26353,N_25228);
nand U28514 (N_28514,N_25951,N_26038);
xnor U28515 (N_28515,N_27331,N_25799);
xnor U28516 (N_28516,N_26841,N_27314);
nor U28517 (N_28517,N_25203,N_26020);
nand U28518 (N_28518,N_26111,N_25286);
nor U28519 (N_28519,N_26046,N_25840);
nand U28520 (N_28520,N_27158,N_26123);
and U28521 (N_28521,N_25144,N_26143);
and U28522 (N_28522,N_25817,N_25996);
xnor U28523 (N_28523,N_25191,N_27273);
or U28524 (N_28524,N_25986,N_27398);
xnor U28525 (N_28525,N_26005,N_26032);
nand U28526 (N_28526,N_26372,N_26852);
xor U28527 (N_28527,N_26649,N_26268);
nand U28528 (N_28528,N_25504,N_26884);
nor U28529 (N_28529,N_27139,N_25779);
xor U28530 (N_28530,N_26612,N_25882);
nor U28531 (N_28531,N_25063,N_25665);
nand U28532 (N_28532,N_26978,N_27170);
nor U28533 (N_28533,N_27293,N_26932);
nor U28534 (N_28534,N_25045,N_25471);
and U28535 (N_28535,N_25077,N_26165);
xor U28536 (N_28536,N_26348,N_27307);
nor U28537 (N_28537,N_26604,N_25023);
xnor U28538 (N_28538,N_27078,N_26338);
nand U28539 (N_28539,N_27015,N_26828);
or U28540 (N_28540,N_26847,N_26585);
or U28541 (N_28541,N_27080,N_26526);
nor U28542 (N_28542,N_26438,N_26562);
or U28543 (N_28543,N_26055,N_26569);
xnor U28544 (N_28544,N_26758,N_25744);
and U28545 (N_28545,N_25594,N_26352);
nor U28546 (N_28546,N_26464,N_26699);
or U28547 (N_28547,N_26586,N_26095);
or U28548 (N_28548,N_26186,N_26023);
xnor U28549 (N_28549,N_25340,N_26311);
nand U28550 (N_28550,N_25578,N_26770);
xor U28551 (N_28551,N_27350,N_25229);
nand U28552 (N_28552,N_25990,N_27288);
and U28553 (N_28553,N_25080,N_27497);
nor U28554 (N_28554,N_26117,N_27174);
or U28555 (N_28555,N_26824,N_25616);
or U28556 (N_28556,N_26259,N_26969);
nand U28557 (N_28557,N_26919,N_26446);
nor U28558 (N_28558,N_26439,N_25404);
nor U28559 (N_28559,N_25099,N_25680);
and U28560 (N_28560,N_27000,N_25494);
and U28561 (N_28561,N_27372,N_26686);
nor U28562 (N_28562,N_26961,N_27218);
or U28563 (N_28563,N_27462,N_27164);
or U28564 (N_28564,N_27205,N_26190);
and U28565 (N_28565,N_27101,N_26260);
or U28566 (N_28566,N_25259,N_25226);
nand U28567 (N_28567,N_27496,N_26819);
nand U28568 (N_28568,N_25369,N_25304);
nand U28569 (N_28569,N_25800,N_27329);
nand U28570 (N_28570,N_27146,N_25563);
or U28571 (N_28571,N_25541,N_25530);
nand U28572 (N_28572,N_26422,N_25756);
or U28573 (N_28573,N_25392,N_27230);
nor U28574 (N_28574,N_27042,N_26936);
nand U28575 (N_28575,N_26767,N_26816);
nand U28576 (N_28576,N_26889,N_26068);
nor U28577 (N_28577,N_26487,N_25179);
or U28578 (N_28578,N_26427,N_25571);
nor U28579 (N_28579,N_25206,N_27461);
nand U28580 (N_28580,N_25984,N_26818);
nand U28581 (N_28581,N_26242,N_26406);
nor U28582 (N_28582,N_25534,N_25457);
and U28583 (N_28583,N_27124,N_26748);
xor U28584 (N_28584,N_27154,N_27103);
nor U28585 (N_28585,N_26549,N_26450);
and U28586 (N_28586,N_26182,N_26675);
nor U28587 (N_28587,N_25091,N_25153);
nor U28588 (N_28588,N_27446,N_26506);
or U28589 (N_28589,N_26294,N_25677);
xnor U28590 (N_28590,N_26834,N_25434);
xor U28591 (N_28591,N_25140,N_27470);
or U28592 (N_28592,N_26313,N_25611);
nand U28593 (N_28593,N_25222,N_26882);
xor U28594 (N_28594,N_26927,N_27150);
and U28595 (N_28595,N_25911,N_25716);
and U28596 (N_28596,N_25449,N_25368);
nand U28597 (N_28597,N_27482,N_25370);
nand U28598 (N_28598,N_27375,N_26426);
xor U28599 (N_28599,N_25886,N_25173);
and U28600 (N_28600,N_26287,N_27439);
nand U28601 (N_28601,N_25971,N_26103);
xor U28602 (N_28602,N_26556,N_25406);
nand U28603 (N_28603,N_25967,N_27395);
nor U28604 (N_28604,N_25874,N_25373);
nand U28605 (N_28605,N_26879,N_26790);
xnor U28606 (N_28606,N_26971,N_27242);
and U28607 (N_28607,N_26571,N_26201);
or U28608 (N_28608,N_26673,N_25017);
and U28609 (N_28609,N_27234,N_25093);
xor U28610 (N_28610,N_25108,N_26269);
or U28611 (N_28611,N_27046,N_25160);
xnor U28612 (N_28612,N_26400,N_27299);
or U28613 (N_28613,N_25898,N_27367);
and U28614 (N_28614,N_25866,N_25985);
nor U28615 (N_28615,N_25709,N_25389);
nand U28616 (N_28616,N_27173,N_25295);
nor U28617 (N_28617,N_26798,N_27227);
and U28618 (N_28618,N_26715,N_26393);
nand U28619 (N_28619,N_25622,N_27106);
nor U28620 (N_28620,N_27290,N_26291);
nor U28621 (N_28621,N_26015,N_26542);
nor U28622 (N_28622,N_25966,N_25177);
or U28623 (N_28623,N_25750,N_25718);
nand U28624 (N_28624,N_26652,N_27087);
nand U28625 (N_28625,N_26867,N_25848);
nor U28626 (N_28626,N_27454,N_27031);
nor U28627 (N_28627,N_27240,N_25730);
nand U28628 (N_28628,N_25702,N_26620);
nor U28629 (N_28629,N_26071,N_25617);
or U28630 (N_28630,N_25464,N_26638);
nor U28631 (N_28631,N_26836,N_26803);
or U28632 (N_28632,N_26382,N_25755);
and U28633 (N_28633,N_25025,N_26484);
or U28634 (N_28634,N_25178,N_27108);
nand U28635 (N_28635,N_27419,N_25187);
and U28636 (N_28636,N_25555,N_26810);
nand U28637 (N_28637,N_27104,N_25997);
nor U28638 (N_28638,N_27123,N_26811);
nand U28639 (N_28639,N_26907,N_25811);
or U28640 (N_28640,N_26436,N_26404);
nor U28641 (N_28641,N_25103,N_26327);
or U28642 (N_28642,N_25946,N_26990);
and U28643 (N_28643,N_25524,N_26825);
nand U28644 (N_28644,N_26965,N_25004);
nor U28645 (N_28645,N_25387,N_25060);
and U28646 (N_28646,N_25174,N_26555);
or U28647 (N_28647,N_25420,N_25491);
xor U28648 (N_28648,N_26476,N_25682);
or U28649 (N_28649,N_26871,N_27420);
nand U28650 (N_28650,N_26274,N_25105);
or U28651 (N_28651,N_26488,N_26947);
and U28652 (N_28652,N_25015,N_26253);
nor U28653 (N_28653,N_26431,N_27488);
and U28654 (N_28654,N_25629,N_25408);
nor U28655 (N_28655,N_25233,N_27458);
xor U28656 (N_28656,N_26787,N_26324);
nor U28657 (N_28657,N_25409,N_26985);
and U28658 (N_28658,N_26430,N_25479);
and U28659 (N_28659,N_25533,N_26498);
nor U28660 (N_28660,N_26902,N_26898);
xnor U28661 (N_28661,N_26981,N_26712);
and U28662 (N_28662,N_25193,N_26814);
and U28663 (N_28663,N_25264,N_25405);
or U28664 (N_28664,N_26184,N_25062);
nor U28665 (N_28665,N_26976,N_25918);
and U28666 (N_28666,N_25934,N_27231);
xor U28667 (N_28667,N_26047,N_26685);
or U28668 (N_28668,N_26958,N_25738);
nor U28669 (N_28669,N_26875,N_26559);
and U28670 (N_28670,N_26297,N_26634);
or U28671 (N_28671,N_26359,N_27223);
nor U28672 (N_28672,N_26622,N_27039);
and U28673 (N_28673,N_27045,N_26019);
or U28674 (N_28674,N_25403,N_26309);
nor U28675 (N_28675,N_26765,N_25657);
xnor U28676 (N_28676,N_25735,N_25357);
xor U28677 (N_28677,N_26164,N_25423);
nor U28678 (N_28678,N_26368,N_26933);
xor U28679 (N_28679,N_25699,N_26789);
xnor U28680 (N_28680,N_25553,N_25595);
nor U28681 (N_28681,N_25466,N_26210);
and U28682 (N_28682,N_25005,N_26956);
and U28683 (N_28683,N_25416,N_27298);
nand U28684 (N_28684,N_25297,N_25112);
or U28685 (N_28685,N_25974,N_26701);
and U28686 (N_28686,N_25928,N_26100);
or U28687 (N_28687,N_26529,N_26394);
and U28688 (N_28688,N_27001,N_25460);
nor U28689 (N_28689,N_27268,N_26722);
nor U28690 (N_28690,N_26283,N_25069);
and U28691 (N_28691,N_25670,N_26002);
xor U28692 (N_28692,N_26308,N_26817);
nor U28693 (N_28693,N_25936,N_26263);
or U28694 (N_28694,N_27115,N_25891);
nand U28695 (N_28695,N_27090,N_27457);
nand U28696 (N_28696,N_26679,N_25192);
or U28697 (N_28697,N_27191,N_25402);
or U28698 (N_28698,N_26179,N_25047);
nor U28699 (N_28699,N_26031,N_26412);
nor U28700 (N_28700,N_26462,N_25628);
nand U28701 (N_28701,N_25597,N_25564);
nand U28702 (N_28702,N_27485,N_25690);
xnor U28703 (N_28703,N_26483,N_26441);
and U28704 (N_28704,N_25438,N_25789);
nand U28705 (N_28705,N_26307,N_25072);
or U28706 (N_28706,N_25488,N_25018);
and U28707 (N_28707,N_25830,N_26574);
nor U28708 (N_28708,N_25638,N_27063);
nor U28709 (N_28709,N_26251,N_26553);
xor U28710 (N_28710,N_27155,N_26760);
nor U28711 (N_28711,N_26320,N_26121);
nand U28712 (N_28712,N_27471,N_26813);
or U28713 (N_28713,N_25301,N_25031);
or U28714 (N_28714,N_26275,N_26960);
or U28715 (N_28715,N_25516,N_27422);
nor U28716 (N_28716,N_26233,N_26337);
nor U28717 (N_28717,N_26954,N_26689);
nor U28718 (N_28718,N_26666,N_27353);
xor U28719 (N_28719,N_25020,N_26145);
nor U28720 (N_28720,N_25870,N_26885);
xor U28721 (N_28721,N_26264,N_25278);
xnor U28722 (N_28722,N_27215,N_25385);
nand U28723 (N_28723,N_25267,N_25836);
nand U28724 (N_28724,N_27254,N_26114);
and U28725 (N_28725,N_25754,N_25049);
and U28726 (N_28726,N_25593,N_26934);
xnor U28727 (N_28727,N_26220,N_26992);
xor U28728 (N_28728,N_25111,N_26449);
nor U28729 (N_28729,N_26672,N_26951);
and U28730 (N_28730,N_25506,N_26204);
nor U28731 (N_28731,N_26966,N_25824);
and U28732 (N_28732,N_26132,N_27221);
nor U28733 (N_28733,N_26625,N_25816);
or U28734 (N_28734,N_26973,N_25969);
nor U28735 (N_28735,N_27431,N_26776);
and U28736 (N_28736,N_27134,N_26964);
or U28737 (N_28737,N_26213,N_26175);
nand U28738 (N_28738,N_26507,N_27341);
or U28739 (N_28739,N_26904,N_25550);
xnor U28740 (N_28740,N_26328,N_26873);
or U28741 (N_28741,N_26037,N_26628);
xor U28742 (N_28742,N_25723,N_26226);
and U28743 (N_28743,N_26178,N_26236);
xnor U28744 (N_28744,N_25517,N_25367);
nand U28745 (N_28745,N_25291,N_26315);
xor U28746 (N_28746,N_27413,N_25535);
and U28747 (N_28747,N_25935,N_27110);
nor U28748 (N_28748,N_25876,N_25159);
or U28749 (N_28749,N_26728,N_25042);
xnor U28750 (N_28750,N_27365,N_27415);
or U28751 (N_28751,N_26457,N_27373);
nand U28752 (N_28752,N_27303,N_27405);
nand U28753 (N_28753,N_26548,N_25660);
and U28754 (N_28754,N_25130,N_26739);
or U28755 (N_28755,N_26041,N_26333);
or U28756 (N_28756,N_25015,N_25721);
xnor U28757 (N_28757,N_26833,N_26254);
and U28758 (N_28758,N_26303,N_25312);
and U28759 (N_28759,N_26352,N_27341);
xnor U28760 (N_28760,N_26071,N_27396);
xor U28761 (N_28761,N_26565,N_25585);
nor U28762 (N_28762,N_25630,N_26481);
or U28763 (N_28763,N_26149,N_26414);
and U28764 (N_28764,N_25630,N_25344);
or U28765 (N_28765,N_27419,N_26080);
xor U28766 (N_28766,N_26885,N_25851);
nand U28767 (N_28767,N_25790,N_26913);
or U28768 (N_28768,N_25793,N_25972);
nand U28769 (N_28769,N_26157,N_25489);
xor U28770 (N_28770,N_27339,N_25944);
and U28771 (N_28771,N_26579,N_26441);
and U28772 (N_28772,N_26852,N_25925);
nand U28773 (N_28773,N_26143,N_25639);
nand U28774 (N_28774,N_25716,N_26702);
and U28775 (N_28775,N_26801,N_26301);
or U28776 (N_28776,N_27091,N_27351);
nand U28777 (N_28777,N_27215,N_25837);
or U28778 (N_28778,N_25125,N_27077);
nor U28779 (N_28779,N_25644,N_25107);
nand U28780 (N_28780,N_25929,N_26372);
and U28781 (N_28781,N_25622,N_27346);
and U28782 (N_28782,N_26939,N_27428);
nor U28783 (N_28783,N_26728,N_25010);
or U28784 (N_28784,N_25972,N_25175);
xor U28785 (N_28785,N_27348,N_27324);
and U28786 (N_28786,N_27462,N_26748);
nand U28787 (N_28787,N_26648,N_26633);
nand U28788 (N_28788,N_26703,N_25814);
or U28789 (N_28789,N_25764,N_25153);
and U28790 (N_28790,N_27280,N_26123);
and U28791 (N_28791,N_26466,N_25466);
xor U28792 (N_28792,N_26779,N_26382);
and U28793 (N_28793,N_26242,N_27402);
and U28794 (N_28794,N_26786,N_26219);
nand U28795 (N_28795,N_26807,N_26680);
nand U28796 (N_28796,N_27373,N_26396);
xor U28797 (N_28797,N_27063,N_27073);
and U28798 (N_28798,N_25388,N_25163);
or U28799 (N_28799,N_26854,N_25240);
nand U28800 (N_28800,N_25196,N_25328);
or U28801 (N_28801,N_26357,N_27039);
or U28802 (N_28802,N_25387,N_25438);
xor U28803 (N_28803,N_26480,N_26332);
and U28804 (N_28804,N_26197,N_25011);
xor U28805 (N_28805,N_25720,N_27454);
xnor U28806 (N_28806,N_25517,N_26821);
nand U28807 (N_28807,N_27448,N_25441);
or U28808 (N_28808,N_25430,N_25438);
or U28809 (N_28809,N_26467,N_25433);
and U28810 (N_28810,N_25301,N_26735);
or U28811 (N_28811,N_25780,N_26155);
nor U28812 (N_28812,N_25155,N_27171);
nand U28813 (N_28813,N_25072,N_26318);
nand U28814 (N_28814,N_25586,N_26738);
nand U28815 (N_28815,N_25705,N_26291);
xnor U28816 (N_28816,N_27189,N_27132);
nand U28817 (N_28817,N_25394,N_25294);
and U28818 (N_28818,N_27011,N_25158);
or U28819 (N_28819,N_25658,N_25340);
or U28820 (N_28820,N_26599,N_26935);
or U28821 (N_28821,N_26887,N_25088);
and U28822 (N_28822,N_26124,N_27198);
nor U28823 (N_28823,N_26475,N_25476);
or U28824 (N_28824,N_25148,N_26073);
and U28825 (N_28825,N_25864,N_26453);
nor U28826 (N_28826,N_27236,N_26081);
and U28827 (N_28827,N_27111,N_26437);
and U28828 (N_28828,N_25947,N_27361);
or U28829 (N_28829,N_25118,N_26939);
nand U28830 (N_28830,N_27079,N_27142);
nor U28831 (N_28831,N_26165,N_26146);
nor U28832 (N_28832,N_27074,N_26965);
nand U28833 (N_28833,N_26863,N_26809);
or U28834 (N_28834,N_26116,N_25625);
nor U28835 (N_28835,N_25824,N_26178);
or U28836 (N_28836,N_27222,N_26016);
and U28837 (N_28837,N_27379,N_27144);
nand U28838 (N_28838,N_25288,N_25209);
and U28839 (N_28839,N_26820,N_26819);
or U28840 (N_28840,N_27252,N_27387);
nor U28841 (N_28841,N_26711,N_27312);
nand U28842 (N_28842,N_26015,N_25784);
nor U28843 (N_28843,N_27169,N_26704);
and U28844 (N_28844,N_25147,N_26875);
and U28845 (N_28845,N_27440,N_25096);
xnor U28846 (N_28846,N_26118,N_26588);
xnor U28847 (N_28847,N_26039,N_25616);
and U28848 (N_28848,N_25618,N_26322);
xnor U28849 (N_28849,N_27305,N_25151);
and U28850 (N_28850,N_25894,N_27132);
xnor U28851 (N_28851,N_26723,N_26523);
or U28852 (N_28852,N_26512,N_25555);
nand U28853 (N_28853,N_25835,N_26483);
nand U28854 (N_28854,N_25880,N_25895);
nand U28855 (N_28855,N_26157,N_27308);
nand U28856 (N_28856,N_25042,N_26876);
xor U28857 (N_28857,N_27323,N_26942);
or U28858 (N_28858,N_25526,N_26757);
and U28859 (N_28859,N_27066,N_27012);
nor U28860 (N_28860,N_26069,N_26477);
and U28861 (N_28861,N_25883,N_25620);
or U28862 (N_28862,N_27094,N_27199);
xnor U28863 (N_28863,N_25578,N_27223);
nand U28864 (N_28864,N_27025,N_25595);
nand U28865 (N_28865,N_26858,N_25888);
or U28866 (N_28866,N_27391,N_26154);
or U28867 (N_28867,N_27113,N_25941);
xnor U28868 (N_28868,N_26627,N_26714);
nand U28869 (N_28869,N_26400,N_25967);
nand U28870 (N_28870,N_27450,N_27396);
xor U28871 (N_28871,N_26995,N_25582);
and U28872 (N_28872,N_27283,N_25595);
nand U28873 (N_28873,N_26428,N_26435);
and U28874 (N_28874,N_25622,N_25013);
or U28875 (N_28875,N_25505,N_27331);
nor U28876 (N_28876,N_25809,N_25400);
nor U28877 (N_28877,N_27149,N_25575);
nor U28878 (N_28878,N_27272,N_25601);
nor U28879 (N_28879,N_25174,N_27053);
and U28880 (N_28880,N_25437,N_26690);
and U28881 (N_28881,N_27000,N_25744);
xnor U28882 (N_28882,N_25263,N_26429);
nor U28883 (N_28883,N_27441,N_25951);
nor U28884 (N_28884,N_25914,N_25321);
xor U28885 (N_28885,N_25743,N_25264);
nor U28886 (N_28886,N_26920,N_25769);
xnor U28887 (N_28887,N_25623,N_27281);
and U28888 (N_28888,N_26700,N_26750);
nand U28889 (N_28889,N_26310,N_25066);
nand U28890 (N_28890,N_26479,N_26506);
xor U28891 (N_28891,N_25867,N_25551);
nand U28892 (N_28892,N_25983,N_26544);
nand U28893 (N_28893,N_25558,N_26118);
nand U28894 (N_28894,N_26899,N_25923);
or U28895 (N_28895,N_27358,N_25642);
nor U28896 (N_28896,N_26442,N_25593);
or U28897 (N_28897,N_27195,N_25983);
nand U28898 (N_28898,N_26752,N_26641);
or U28899 (N_28899,N_25102,N_26997);
or U28900 (N_28900,N_25580,N_27308);
and U28901 (N_28901,N_25055,N_25294);
xnor U28902 (N_28902,N_27078,N_25095);
or U28903 (N_28903,N_27111,N_25991);
xor U28904 (N_28904,N_25507,N_27226);
and U28905 (N_28905,N_25643,N_26302);
xnor U28906 (N_28906,N_27187,N_25787);
or U28907 (N_28907,N_27459,N_27198);
nand U28908 (N_28908,N_25992,N_25071);
and U28909 (N_28909,N_26995,N_26085);
or U28910 (N_28910,N_25250,N_26947);
xnor U28911 (N_28911,N_26296,N_25524);
and U28912 (N_28912,N_25519,N_25361);
and U28913 (N_28913,N_25897,N_26313);
or U28914 (N_28914,N_26164,N_25758);
nand U28915 (N_28915,N_25609,N_27000);
or U28916 (N_28916,N_27034,N_27474);
or U28917 (N_28917,N_26479,N_27260);
xor U28918 (N_28918,N_26582,N_25669);
and U28919 (N_28919,N_25998,N_25938);
or U28920 (N_28920,N_26135,N_26645);
xor U28921 (N_28921,N_26846,N_27054);
or U28922 (N_28922,N_27469,N_25790);
and U28923 (N_28923,N_26099,N_25242);
nor U28924 (N_28924,N_27148,N_26617);
nand U28925 (N_28925,N_27105,N_27059);
xnor U28926 (N_28926,N_27156,N_27423);
nor U28927 (N_28927,N_25734,N_26328);
and U28928 (N_28928,N_27394,N_25400);
nor U28929 (N_28929,N_27220,N_25597);
xnor U28930 (N_28930,N_25120,N_25926);
and U28931 (N_28931,N_27225,N_25296);
and U28932 (N_28932,N_25925,N_27111);
xnor U28933 (N_28933,N_25888,N_27213);
nand U28934 (N_28934,N_26276,N_25879);
xor U28935 (N_28935,N_25150,N_26333);
or U28936 (N_28936,N_27494,N_26335);
and U28937 (N_28937,N_25443,N_26167);
and U28938 (N_28938,N_26372,N_27066);
nor U28939 (N_28939,N_26001,N_26974);
xnor U28940 (N_28940,N_27080,N_26116);
nand U28941 (N_28941,N_26052,N_26106);
nand U28942 (N_28942,N_25910,N_26374);
nand U28943 (N_28943,N_25045,N_26796);
nor U28944 (N_28944,N_25350,N_25718);
xnor U28945 (N_28945,N_25519,N_27072);
nand U28946 (N_28946,N_25599,N_25946);
and U28947 (N_28947,N_26203,N_27019);
and U28948 (N_28948,N_26089,N_25315);
nand U28949 (N_28949,N_26052,N_25263);
nor U28950 (N_28950,N_26869,N_26097);
and U28951 (N_28951,N_25568,N_27243);
nand U28952 (N_28952,N_25537,N_25450);
nor U28953 (N_28953,N_27486,N_26961);
xnor U28954 (N_28954,N_26260,N_26485);
xor U28955 (N_28955,N_27200,N_26690);
xnor U28956 (N_28956,N_26961,N_26092);
or U28957 (N_28957,N_26083,N_26784);
nor U28958 (N_28958,N_26172,N_26674);
or U28959 (N_28959,N_27252,N_25717);
nor U28960 (N_28960,N_25034,N_25396);
nand U28961 (N_28961,N_26572,N_26692);
or U28962 (N_28962,N_26392,N_25028);
nand U28963 (N_28963,N_25165,N_25818);
nor U28964 (N_28964,N_26231,N_25970);
or U28965 (N_28965,N_25419,N_25291);
or U28966 (N_28966,N_25997,N_25077);
nor U28967 (N_28967,N_25060,N_26571);
and U28968 (N_28968,N_27161,N_25640);
and U28969 (N_28969,N_25650,N_26704);
xor U28970 (N_28970,N_25439,N_25451);
and U28971 (N_28971,N_26247,N_27402);
or U28972 (N_28972,N_27274,N_25463);
and U28973 (N_28973,N_25773,N_27411);
and U28974 (N_28974,N_27304,N_25807);
xnor U28975 (N_28975,N_27194,N_27308);
xor U28976 (N_28976,N_26314,N_26332);
or U28977 (N_28977,N_25226,N_25876);
nand U28978 (N_28978,N_27041,N_27175);
and U28979 (N_28979,N_25261,N_26959);
or U28980 (N_28980,N_25659,N_26856);
xor U28981 (N_28981,N_25035,N_26191);
and U28982 (N_28982,N_25455,N_26894);
or U28983 (N_28983,N_26546,N_25332);
nand U28984 (N_28984,N_26442,N_25470);
or U28985 (N_28985,N_25738,N_27166);
nand U28986 (N_28986,N_27085,N_25189);
or U28987 (N_28987,N_26317,N_26123);
and U28988 (N_28988,N_26232,N_26416);
xor U28989 (N_28989,N_25254,N_26799);
and U28990 (N_28990,N_26536,N_26006);
nand U28991 (N_28991,N_27317,N_26886);
or U28992 (N_28992,N_26609,N_27488);
nor U28993 (N_28993,N_26962,N_25412);
nor U28994 (N_28994,N_26036,N_27026);
and U28995 (N_28995,N_26323,N_26261);
nor U28996 (N_28996,N_26840,N_25237);
and U28997 (N_28997,N_26926,N_25341);
or U28998 (N_28998,N_25717,N_27016);
nand U28999 (N_28999,N_27424,N_26954);
nand U29000 (N_29000,N_25134,N_26140);
or U29001 (N_29001,N_25336,N_25370);
xnor U29002 (N_29002,N_25449,N_26237);
nand U29003 (N_29003,N_25558,N_27453);
xnor U29004 (N_29004,N_25719,N_27030);
xor U29005 (N_29005,N_25699,N_27244);
xnor U29006 (N_29006,N_25978,N_25285);
nor U29007 (N_29007,N_27363,N_26528);
or U29008 (N_29008,N_27140,N_25165);
xnor U29009 (N_29009,N_27238,N_25406);
nor U29010 (N_29010,N_27042,N_26217);
and U29011 (N_29011,N_25647,N_26093);
and U29012 (N_29012,N_25922,N_27346);
nand U29013 (N_29013,N_27029,N_26706);
or U29014 (N_29014,N_26774,N_25846);
or U29015 (N_29015,N_25852,N_25245);
nand U29016 (N_29016,N_26033,N_25331);
nand U29017 (N_29017,N_25672,N_25239);
xor U29018 (N_29018,N_25098,N_25611);
and U29019 (N_29019,N_26133,N_25247);
nand U29020 (N_29020,N_27067,N_26766);
or U29021 (N_29021,N_26026,N_27406);
nor U29022 (N_29022,N_25241,N_25814);
xor U29023 (N_29023,N_25811,N_25611);
or U29024 (N_29024,N_26954,N_25183);
or U29025 (N_29025,N_27456,N_26734);
or U29026 (N_29026,N_26231,N_25319);
nand U29027 (N_29027,N_26610,N_26618);
and U29028 (N_29028,N_26690,N_27260);
xor U29029 (N_29029,N_25926,N_25621);
and U29030 (N_29030,N_25244,N_25107);
xnor U29031 (N_29031,N_26892,N_25575);
xor U29032 (N_29032,N_25217,N_27281);
xnor U29033 (N_29033,N_26242,N_26749);
or U29034 (N_29034,N_26461,N_25520);
or U29035 (N_29035,N_26845,N_26328);
nand U29036 (N_29036,N_25797,N_26035);
or U29037 (N_29037,N_25226,N_26194);
nor U29038 (N_29038,N_26488,N_25099);
or U29039 (N_29039,N_26478,N_26985);
xnor U29040 (N_29040,N_25894,N_27083);
or U29041 (N_29041,N_26635,N_25944);
and U29042 (N_29042,N_26985,N_26605);
and U29043 (N_29043,N_26528,N_26861);
and U29044 (N_29044,N_27169,N_25027);
or U29045 (N_29045,N_26487,N_27473);
or U29046 (N_29046,N_27368,N_25194);
nor U29047 (N_29047,N_26387,N_25882);
and U29048 (N_29048,N_25734,N_27135);
xor U29049 (N_29049,N_26860,N_26420);
nand U29050 (N_29050,N_27039,N_25578);
xor U29051 (N_29051,N_25433,N_25440);
or U29052 (N_29052,N_25806,N_26604);
nand U29053 (N_29053,N_26305,N_25369);
nand U29054 (N_29054,N_26401,N_27137);
or U29055 (N_29055,N_26326,N_25559);
and U29056 (N_29056,N_25726,N_27199);
or U29057 (N_29057,N_27072,N_25688);
nor U29058 (N_29058,N_25635,N_26260);
nand U29059 (N_29059,N_26263,N_25081);
and U29060 (N_29060,N_26116,N_25534);
xor U29061 (N_29061,N_25413,N_25689);
and U29062 (N_29062,N_25991,N_27173);
nor U29063 (N_29063,N_26508,N_27484);
xnor U29064 (N_29064,N_25186,N_26117);
xor U29065 (N_29065,N_26037,N_25136);
xor U29066 (N_29066,N_25259,N_27055);
or U29067 (N_29067,N_25430,N_25876);
nand U29068 (N_29068,N_26975,N_26004);
nor U29069 (N_29069,N_26902,N_27099);
nand U29070 (N_29070,N_25427,N_26296);
xnor U29071 (N_29071,N_25591,N_25973);
nand U29072 (N_29072,N_26339,N_25392);
nor U29073 (N_29073,N_26712,N_26518);
or U29074 (N_29074,N_26248,N_25629);
nor U29075 (N_29075,N_25064,N_25603);
nand U29076 (N_29076,N_25737,N_25436);
nand U29077 (N_29077,N_27266,N_26387);
nand U29078 (N_29078,N_25805,N_25213);
xor U29079 (N_29079,N_26472,N_26468);
and U29080 (N_29080,N_27499,N_26791);
or U29081 (N_29081,N_25800,N_25331);
nor U29082 (N_29082,N_25863,N_26898);
or U29083 (N_29083,N_26260,N_25071);
xor U29084 (N_29084,N_26031,N_25103);
xor U29085 (N_29085,N_27156,N_27075);
nand U29086 (N_29086,N_26637,N_26603);
xnor U29087 (N_29087,N_25430,N_26756);
or U29088 (N_29088,N_27404,N_26517);
nor U29089 (N_29089,N_27432,N_27355);
nand U29090 (N_29090,N_27430,N_26236);
and U29091 (N_29091,N_26871,N_25619);
or U29092 (N_29092,N_25329,N_25478);
nand U29093 (N_29093,N_25990,N_25854);
nand U29094 (N_29094,N_25226,N_27088);
or U29095 (N_29095,N_25747,N_27225);
xor U29096 (N_29096,N_26822,N_26109);
or U29097 (N_29097,N_25044,N_26889);
or U29098 (N_29098,N_26057,N_27123);
or U29099 (N_29099,N_25278,N_27413);
nor U29100 (N_29100,N_27412,N_27459);
nor U29101 (N_29101,N_26177,N_25006);
xnor U29102 (N_29102,N_26623,N_26904);
and U29103 (N_29103,N_26429,N_25691);
and U29104 (N_29104,N_27044,N_26423);
nand U29105 (N_29105,N_26654,N_26129);
nor U29106 (N_29106,N_26538,N_26396);
or U29107 (N_29107,N_25759,N_27155);
xnor U29108 (N_29108,N_25342,N_25815);
and U29109 (N_29109,N_25695,N_25099);
nand U29110 (N_29110,N_25746,N_26257);
nand U29111 (N_29111,N_26736,N_26104);
or U29112 (N_29112,N_25390,N_25166);
nand U29113 (N_29113,N_26876,N_26461);
and U29114 (N_29114,N_25480,N_26423);
xnor U29115 (N_29115,N_25333,N_25912);
nand U29116 (N_29116,N_26899,N_26024);
nand U29117 (N_29117,N_25846,N_27165);
nand U29118 (N_29118,N_26998,N_27046);
and U29119 (N_29119,N_26705,N_25929);
and U29120 (N_29120,N_25936,N_25346);
or U29121 (N_29121,N_26529,N_27082);
or U29122 (N_29122,N_26247,N_26404);
and U29123 (N_29123,N_25124,N_26296);
and U29124 (N_29124,N_26087,N_25606);
or U29125 (N_29125,N_26326,N_27380);
and U29126 (N_29126,N_25861,N_26160);
nor U29127 (N_29127,N_25291,N_27221);
nor U29128 (N_29128,N_25610,N_25520);
xor U29129 (N_29129,N_25923,N_27292);
xnor U29130 (N_29130,N_27499,N_26965);
xnor U29131 (N_29131,N_26476,N_26672);
xnor U29132 (N_29132,N_26019,N_25760);
nand U29133 (N_29133,N_25285,N_26116);
nor U29134 (N_29134,N_26230,N_25386);
and U29135 (N_29135,N_27311,N_25284);
and U29136 (N_29136,N_26360,N_26840);
or U29137 (N_29137,N_26316,N_27033);
nand U29138 (N_29138,N_26569,N_25237);
or U29139 (N_29139,N_26014,N_26666);
xnor U29140 (N_29140,N_26180,N_26538);
xor U29141 (N_29141,N_26442,N_26348);
xor U29142 (N_29142,N_26398,N_25313);
xor U29143 (N_29143,N_27308,N_26087);
and U29144 (N_29144,N_25817,N_25837);
nand U29145 (N_29145,N_26743,N_26605);
or U29146 (N_29146,N_25016,N_25622);
nand U29147 (N_29147,N_26159,N_27269);
xor U29148 (N_29148,N_27198,N_25713);
xor U29149 (N_29149,N_25157,N_26349);
nor U29150 (N_29150,N_27216,N_26429);
or U29151 (N_29151,N_26953,N_25555);
nor U29152 (N_29152,N_25602,N_26798);
and U29153 (N_29153,N_25181,N_25963);
and U29154 (N_29154,N_25371,N_26020);
or U29155 (N_29155,N_25672,N_27104);
and U29156 (N_29156,N_25451,N_26216);
nor U29157 (N_29157,N_26650,N_26603);
and U29158 (N_29158,N_26438,N_26372);
nor U29159 (N_29159,N_26666,N_25154);
or U29160 (N_29160,N_25828,N_25619);
or U29161 (N_29161,N_26820,N_25205);
or U29162 (N_29162,N_26795,N_27381);
xnor U29163 (N_29163,N_27019,N_25566);
nand U29164 (N_29164,N_25185,N_27402);
or U29165 (N_29165,N_26969,N_26535);
xor U29166 (N_29166,N_26719,N_25485);
xnor U29167 (N_29167,N_26176,N_25492);
and U29168 (N_29168,N_25924,N_27209);
nor U29169 (N_29169,N_26314,N_25944);
and U29170 (N_29170,N_25921,N_25433);
nand U29171 (N_29171,N_27192,N_25959);
nand U29172 (N_29172,N_26277,N_25215);
xor U29173 (N_29173,N_27229,N_26464);
xnor U29174 (N_29174,N_26363,N_25964);
nor U29175 (N_29175,N_25885,N_25639);
nand U29176 (N_29176,N_25911,N_26676);
nand U29177 (N_29177,N_27165,N_25377);
or U29178 (N_29178,N_26337,N_26826);
and U29179 (N_29179,N_26789,N_27022);
nor U29180 (N_29180,N_25251,N_26088);
or U29181 (N_29181,N_27029,N_25908);
xnor U29182 (N_29182,N_26354,N_26536);
or U29183 (N_29183,N_25368,N_26036);
xnor U29184 (N_29184,N_25102,N_25565);
nor U29185 (N_29185,N_25346,N_26525);
and U29186 (N_29186,N_25073,N_25564);
or U29187 (N_29187,N_27059,N_26525);
nor U29188 (N_29188,N_26741,N_25910);
nand U29189 (N_29189,N_26376,N_26003);
or U29190 (N_29190,N_27285,N_25008);
nor U29191 (N_29191,N_26103,N_25736);
xor U29192 (N_29192,N_27360,N_26714);
nand U29193 (N_29193,N_25705,N_26885);
or U29194 (N_29194,N_27302,N_25321);
nor U29195 (N_29195,N_26729,N_25081);
or U29196 (N_29196,N_25911,N_25128);
xnor U29197 (N_29197,N_26820,N_26079);
or U29198 (N_29198,N_25007,N_27075);
nand U29199 (N_29199,N_25457,N_27225);
and U29200 (N_29200,N_25302,N_26918);
or U29201 (N_29201,N_26093,N_25713);
nor U29202 (N_29202,N_26478,N_26875);
nor U29203 (N_29203,N_25969,N_25010);
and U29204 (N_29204,N_25807,N_25938);
or U29205 (N_29205,N_26742,N_25053);
xor U29206 (N_29206,N_25129,N_26416);
xor U29207 (N_29207,N_26109,N_25356);
xnor U29208 (N_29208,N_25876,N_25930);
nand U29209 (N_29209,N_25914,N_27040);
nor U29210 (N_29210,N_27329,N_25448);
and U29211 (N_29211,N_27078,N_25140);
or U29212 (N_29212,N_25907,N_27165);
and U29213 (N_29213,N_27071,N_26462);
nand U29214 (N_29214,N_27089,N_26958);
nand U29215 (N_29215,N_26532,N_27402);
nand U29216 (N_29216,N_26532,N_25810);
nor U29217 (N_29217,N_27375,N_25168);
nor U29218 (N_29218,N_26260,N_26127);
or U29219 (N_29219,N_25500,N_26477);
nand U29220 (N_29220,N_27128,N_26234);
xor U29221 (N_29221,N_27357,N_27286);
and U29222 (N_29222,N_26656,N_27270);
nand U29223 (N_29223,N_25442,N_26124);
nand U29224 (N_29224,N_25036,N_25535);
nand U29225 (N_29225,N_25499,N_25367);
nand U29226 (N_29226,N_25807,N_26937);
nand U29227 (N_29227,N_27145,N_26247);
or U29228 (N_29228,N_25446,N_25686);
and U29229 (N_29229,N_25073,N_25865);
or U29230 (N_29230,N_25375,N_25595);
nor U29231 (N_29231,N_25411,N_26094);
xnor U29232 (N_29232,N_26231,N_25096);
and U29233 (N_29233,N_26335,N_27072);
or U29234 (N_29234,N_26333,N_25655);
or U29235 (N_29235,N_25103,N_26043);
nor U29236 (N_29236,N_25733,N_26899);
nor U29237 (N_29237,N_26150,N_26580);
nor U29238 (N_29238,N_27016,N_26649);
xnor U29239 (N_29239,N_26133,N_26257);
xnor U29240 (N_29240,N_27030,N_26361);
or U29241 (N_29241,N_27245,N_25061);
nor U29242 (N_29242,N_25728,N_26385);
xor U29243 (N_29243,N_25591,N_26637);
nor U29244 (N_29244,N_25844,N_26737);
nand U29245 (N_29245,N_25705,N_27373);
and U29246 (N_29246,N_26849,N_26019);
or U29247 (N_29247,N_27052,N_26615);
and U29248 (N_29248,N_26827,N_26272);
nor U29249 (N_29249,N_26919,N_27202);
xnor U29250 (N_29250,N_26497,N_26912);
and U29251 (N_29251,N_25712,N_27155);
xor U29252 (N_29252,N_25717,N_25414);
nor U29253 (N_29253,N_26746,N_26717);
nand U29254 (N_29254,N_27400,N_25002);
or U29255 (N_29255,N_27157,N_25686);
nor U29256 (N_29256,N_25155,N_25878);
nand U29257 (N_29257,N_25042,N_26432);
xnor U29258 (N_29258,N_25953,N_26911);
or U29259 (N_29259,N_25769,N_25099);
or U29260 (N_29260,N_27169,N_26761);
nor U29261 (N_29261,N_26780,N_26234);
nor U29262 (N_29262,N_26405,N_25122);
nor U29263 (N_29263,N_26896,N_26463);
and U29264 (N_29264,N_27377,N_26584);
xnor U29265 (N_29265,N_25681,N_26427);
and U29266 (N_29266,N_27079,N_26674);
nor U29267 (N_29267,N_27252,N_26420);
nor U29268 (N_29268,N_26711,N_25730);
xor U29269 (N_29269,N_25269,N_26198);
and U29270 (N_29270,N_25270,N_26046);
nand U29271 (N_29271,N_27449,N_25902);
nand U29272 (N_29272,N_25223,N_25886);
nand U29273 (N_29273,N_26107,N_26409);
or U29274 (N_29274,N_25605,N_26360);
nand U29275 (N_29275,N_26392,N_26322);
or U29276 (N_29276,N_26548,N_27174);
xnor U29277 (N_29277,N_27145,N_26746);
nand U29278 (N_29278,N_27034,N_27228);
or U29279 (N_29279,N_25681,N_27470);
nor U29280 (N_29280,N_26199,N_26348);
nor U29281 (N_29281,N_26065,N_26608);
and U29282 (N_29282,N_26616,N_26139);
nor U29283 (N_29283,N_25510,N_26206);
or U29284 (N_29284,N_25320,N_25733);
nand U29285 (N_29285,N_26949,N_26614);
or U29286 (N_29286,N_25264,N_26597);
nor U29287 (N_29287,N_25278,N_25466);
nor U29288 (N_29288,N_27055,N_26013);
nand U29289 (N_29289,N_26467,N_26188);
or U29290 (N_29290,N_26020,N_25715);
xnor U29291 (N_29291,N_25745,N_26267);
xor U29292 (N_29292,N_26600,N_25066);
nand U29293 (N_29293,N_26347,N_27365);
and U29294 (N_29294,N_26858,N_25176);
nand U29295 (N_29295,N_26055,N_25812);
or U29296 (N_29296,N_25473,N_25206);
and U29297 (N_29297,N_27460,N_26160);
nor U29298 (N_29298,N_25759,N_26132);
nand U29299 (N_29299,N_25626,N_25664);
or U29300 (N_29300,N_27455,N_25155);
or U29301 (N_29301,N_27228,N_25417);
or U29302 (N_29302,N_25159,N_25599);
and U29303 (N_29303,N_25595,N_27335);
and U29304 (N_29304,N_27388,N_25305);
nor U29305 (N_29305,N_25257,N_26614);
nand U29306 (N_29306,N_25881,N_26050);
xor U29307 (N_29307,N_25640,N_25481);
xor U29308 (N_29308,N_26187,N_27268);
nand U29309 (N_29309,N_26980,N_26559);
or U29310 (N_29310,N_25278,N_25040);
or U29311 (N_29311,N_26301,N_25320);
or U29312 (N_29312,N_27149,N_27174);
nor U29313 (N_29313,N_27492,N_26962);
and U29314 (N_29314,N_26056,N_25172);
or U29315 (N_29315,N_27012,N_25587);
and U29316 (N_29316,N_26976,N_26309);
xor U29317 (N_29317,N_26129,N_26134);
or U29318 (N_29318,N_25768,N_27474);
nor U29319 (N_29319,N_26702,N_26538);
or U29320 (N_29320,N_26643,N_26736);
nand U29321 (N_29321,N_25385,N_25975);
or U29322 (N_29322,N_26459,N_25384);
nand U29323 (N_29323,N_25067,N_25809);
or U29324 (N_29324,N_27177,N_26171);
nor U29325 (N_29325,N_27495,N_26526);
and U29326 (N_29326,N_25811,N_25405);
or U29327 (N_29327,N_26324,N_26819);
nor U29328 (N_29328,N_26347,N_25391);
or U29329 (N_29329,N_25164,N_26259);
or U29330 (N_29330,N_26080,N_25403);
or U29331 (N_29331,N_26238,N_25464);
or U29332 (N_29332,N_25925,N_26231);
and U29333 (N_29333,N_25684,N_25020);
nor U29334 (N_29334,N_27209,N_26066);
nor U29335 (N_29335,N_25614,N_27441);
xnor U29336 (N_29336,N_27379,N_25398);
or U29337 (N_29337,N_26797,N_25247);
nor U29338 (N_29338,N_26519,N_26681);
or U29339 (N_29339,N_26027,N_26550);
and U29340 (N_29340,N_26234,N_26058);
xor U29341 (N_29341,N_26108,N_26556);
nand U29342 (N_29342,N_26368,N_25999);
nand U29343 (N_29343,N_26419,N_25678);
nand U29344 (N_29344,N_26769,N_26185);
and U29345 (N_29345,N_26483,N_27050);
nand U29346 (N_29346,N_25787,N_25643);
nand U29347 (N_29347,N_27151,N_26261);
or U29348 (N_29348,N_26587,N_25977);
and U29349 (N_29349,N_27260,N_25086);
nand U29350 (N_29350,N_27185,N_27311);
and U29351 (N_29351,N_26447,N_26193);
or U29352 (N_29352,N_26577,N_26088);
nor U29353 (N_29353,N_25350,N_26142);
xnor U29354 (N_29354,N_25799,N_25817);
and U29355 (N_29355,N_25609,N_26347);
and U29356 (N_29356,N_26436,N_25295);
xnor U29357 (N_29357,N_25966,N_25237);
and U29358 (N_29358,N_27380,N_26174);
or U29359 (N_29359,N_26108,N_26828);
xor U29360 (N_29360,N_26107,N_25593);
xor U29361 (N_29361,N_26255,N_26311);
xor U29362 (N_29362,N_26442,N_25387);
nand U29363 (N_29363,N_25790,N_25014);
nor U29364 (N_29364,N_25779,N_27152);
nand U29365 (N_29365,N_25171,N_25335);
nor U29366 (N_29366,N_26846,N_26795);
nand U29367 (N_29367,N_25190,N_27249);
nand U29368 (N_29368,N_26895,N_26111);
nor U29369 (N_29369,N_25244,N_26656);
nand U29370 (N_29370,N_25989,N_26304);
nor U29371 (N_29371,N_25769,N_26695);
nand U29372 (N_29372,N_27178,N_25984);
or U29373 (N_29373,N_26262,N_27005);
nand U29374 (N_29374,N_27431,N_27472);
xor U29375 (N_29375,N_26690,N_26300);
nand U29376 (N_29376,N_27302,N_26920);
nor U29377 (N_29377,N_25549,N_27254);
xnor U29378 (N_29378,N_25263,N_26564);
nor U29379 (N_29379,N_26405,N_26080);
nand U29380 (N_29380,N_26726,N_27403);
or U29381 (N_29381,N_25655,N_26684);
or U29382 (N_29382,N_27023,N_25399);
and U29383 (N_29383,N_26655,N_25298);
xor U29384 (N_29384,N_26374,N_25719);
nand U29385 (N_29385,N_25407,N_27454);
and U29386 (N_29386,N_25081,N_25920);
or U29387 (N_29387,N_26843,N_25370);
and U29388 (N_29388,N_26194,N_25643);
or U29389 (N_29389,N_27364,N_27139);
xnor U29390 (N_29390,N_27329,N_25086);
and U29391 (N_29391,N_25858,N_25450);
or U29392 (N_29392,N_26665,N_26040);
xnor U29393 (N_29393,N_25828,N_26362);
or U29394 (N_29394,N_26902,N_25213);
nor U29395 (N_29395,N_25314,N_25340);
nor U29396 (N_29396,N_26612,N_25199);
or U29397 (N_29397,N_27460,N_25604);
nor U29398 (N_29398,N_26366,N_25858);
nor U29399 (N_29399,N_25853,N_27115);
and U29400 (N_29400,N_26034,N_25842);
or U29401 (N_29401,N_26358,N_25029);
and U29402 (N_29402,N_26639,N_26323);
nand U29403 (N_29403,N_26989,N_25306);
and U29404 (N_29404,N_25532,N_26905);
nand U29405 (N_29405,N_25265,N_26048);
xnor U29406 (N_29406,N_25155,N_26409);
nor U29407 (N_29407,N_25897,N_25912);
or U29408 (N_29408,N_26055,N_25946);
or U29409 (N_29409,N_26246,N_26891);
xor U29410 (N_29410,N_25499,N_25902);
and U29411 (N_29411,N_25874,N_25034);
xor U29412 (N_29412,N_26344,N_25615);
and U29413 (N_29413,N_27089,N_25709);
xnor U29414 (N_29414,N_26565,N_25248);
or U29415 (N_29415,N_25415,N_25462);
nand U29416 (N_29416,N_25302,N_25751);
nand U29417 (N_29417,N_27134,N_26614);
xor U29418 (N_29418,N_26481,N_27290);
xor U29419 (N_29419,N_27196,N_25476);
nand U29420 (N_29420,N_26269,N_25701);
nor U29421 (N_29421,N_26983,N_26814);
and U29422 (N_29422,N_25046,N_27359);
nand U29423 (N_29423,N_26936,N_27413);
xor U29424 (N_29424,N_26119,N_25202);
or U29425 (N_29425,N_26851,N_25843);
nor U29426 (N_29426,N_26514,N_25761);
nor U29427 (N_29427,N_26046,N_27119);
or U29428 (N_29428,N_25204,N_25141);
nor U29429 (N_29429,N_25037,N_26725);
xor U29430 (N_29430,N_26009,N_25963);
xor U29431 (N_29431,N_26731,N_26804);
nand U29432 (N_29432,N_25404,N_25656);
xnor U29433 (N_29433,N_27108,N_25428);
and U29434 (N_29434,N_27002,N_26813);
nor U29435 (N_29435,N_26780,N_26103);
or U29436 (N_29436,N_26256,N_26681);
xor U29437 (N_29437,N_27286,N_25306);
nor U29438 (N_29438,N_25822,N_27297);
nor U29439 (N_29439,N_25771,N_26087);
nor U29440 (N_29440,N_25584,N_27335);
or U29441 (N_29441,N_25838,N_27185);
nand U29442 (N_29442,N_26499,N_26260);
nor U29443 (N_29443,N_26971,N_25494);
nor U29444 (N_29444,N_27426,N_26474);
and U29445 (N_29445,N_26871,N_26231);
nor U29446 (N_29446,N_26729,N_27137);
nor U29447 (N_29447,N_27001,N_25520);
or U29448 (N_29448,N_25283,N_26043);
xor U29449 (N_29449,N_26192,N_25271);
nor U29450 (N_29450,N_25789,N_27167);
and U29451 (N_29451,N_26890,N_25822);
or U29452 (N_29452,N_26569,N_26858);
or U29453 (N_29453,N_26761,N_25467);
and U29454 (N_29454,N_25521,N_25612);
and U29455 (N_29455,N_26675,N_26127);
xor U29456 (N_29456,N_27140,N_26413);
xnor U29457 (N_29457,N_26607,N_26223);
nor U29458 (N_29458,N_25463,N_27174);
xor U29459 (N_29459,N_27465,N_26307);
or U29460 (N_29460,N_26054,N_27210);
and U29461 (N_29461,N_26404,N_25803);
xor U29462 (N_29462,N_26310,N_25382);
nand U29463 (N_29463,N_25886,N_27133);
or U29464 (N_29464,N_27256,N_26808);
or U29465 (N_29465,N_25844,N_26206);
and U29466 (N_29466,N_25857,N_26239);
or U29467 (N_29467,N_26039,N_25274);
xnor U29468 (N_29468,N_25120,N_27430);
xor U29469 (N_29469,N_25642,N_27438);
and U29470 (N_29470,N_25733,N_26774);
xnor U29471 (N_29471,N_27101,N_25535);
xnor U29472 (N_29472,N_25138,N_25671);
nand U29473 (N_29473,N_26829,N_26347);
and U29474 (N_29474,N_26010,N_25551);
xor U29475 (N_29475,N_25490,N_26315);
nor U29476 (N_29476,N_26300,N_25783);
nor U29477 (N_29477,N_25126,N_25724);
nor U29478 (N_29478,N_25433,N_26584);
xnor U29479 (N_29479,N_25535,N_25240);
and U29480 (N_29480,N_26704,N_27427);
and U29481 (N_29481,N_26203,N_25580);
or U29482 (N_29482,N_26874,N_27461);
xor U29483 (N_29483,N_26981,N_25295);
and U29484 (N_29484,N_25813,N_26616);
xnor U29485 (N_29485,N_25876,N_26628);
nand U29486 (N_29486,N_26865,N_26106);
nor U29487 (N_29487,N_27070,N_25704);
or U29488 (N_29488,N_26031,N_25143);
nor U29489 (N_29489,N_27392,N_26784);
xnor U29490 (N_29490,N_26918,N_27323);
or U29491 (N_29491,N_27234,N_26302);
and U29492 (N_29492,N_25424,N_26804);
or U29493 (N_29493,N_27297,N_26858);
nand U29494 (N_29494,N_26333,N_26615);
and U29495 (N_29495,N_25176,N_25557);
and U29496 (N_29496,N_25548,N_26674);
nand U29497 (N_29497,N_27214,N_26791);
xor U29498 (N_29498,N_26439,N_27395);
nor U29499 (N_29499,N_25817,N_25150);
nor U29500 (N_29500,N_25543,N_26904);
or U29501 (N_29501,N_25691,N_27443);
and U29502 (N_29502,N_26698,N_25225);
or U29503 (N_29503,N_25751,N_26851);
or U29504 (N_29504,N_25487,N_25873);
or U29505 (N_29505,N_26758,N_25893);
xor U29506 (N_29506,N_25429,N_26954);
nor U29507 (N_29507,N_27268,N_25211);
and U29508 (N_29508,N_26833,N_25117);
and U29509 (N_29509,N_26432,N_27047);
nor U29510 (N_29510,N_25240,N_25196);
nor U29511 (N_29511,N_25925,N_25873);
xnor U29512 (N_29512,N_26303,N_25611);
nand U29513 (N_29513,N_26887,N_25578);
nand U29514 (N_29514,N_26364,N_25984);
or U29515 (N_29515,N_25741,N_26162);
nand U29516 (N_29516,N_26373,N_25492);
nor U29517 (N_29517,N_25176,N_26866);
nand U29518 (N_29518,N_25533,N_25046);
nand U29519 (N_29519,N_25060,N_27155);
nand U29520 (N_29520,N_26367,N_27420);
nor U29521 (N_29521,N_26345,N_27374);
nand U29522 (N_29522,N_26588,N_26436);
or U29523 (N_29523,N_26296,N_26079);
nor U29524 (N_29524,N_25670,N_25833);
nor U29525 (N_29525,N_27410,N_25279);
or U29526 (N_29526,N_26175,N_25249);
nand U29527 (N_29527,N_26672,N_25611);
nor U29528 (N_29528,N_25802,N_25850);
nor U29529 (N_29529,N_25084,N_27021);
or U29530 (N_29530,N_27100,N_25766);
xor U29531 (N_29531,N_26675,N_25341);
and U29532 (N_29532,N_27217,N_26484);
xnor U29533 (N_29533,N_25708,N_26883);
nand U29534 (N_29534,N_27063,N_26102);
xor U29535 (N_29535,N_25828,N_25270);
nand U29536 (N_29536,N_27425,N_27371);
nand U29537 (N_29537,N_26402,N_26579);
xnor U29538 (N_29538,N_26958,N_25145);
nor U29539 (N_29539,N_27413,N_25712);
or U29540 (N_29540,N_26903,N_27147);
or U29541 (N_29541,N_26847,N_26355);
nor U29542 (N_29542,N_25763,N_26113);
nand U29543 (N_29543,N_25942,N_26759);
nor U29544 (N_29544,N_26080,N_25141);
or U29545 (N_29545,N_26384,N_25179);
and U29546 (N_29546,N_26413,N_25240);
nand U29547 (N_29547,N_25412,N_26830);
xor U29548 (N_29548,N_26756,N_25002);
and U29549 (N_29549,N_25708,N_25461);
nand U29550 (N_29550,N_26853,N_26783);
nand U29551 (N_29551,N_26192,N_26941);
xor U29552 (N_29552,N_25427,N_25895);
and U29553 (N_29553,N_25464,N_25100);
nand U29554 (N_29554,N_26807,N_26531);
xor U29555 (N_29555,N_26173,N_25387);
and U29556 (N_29556,N_26511,N_25158);
and U29557 (N_29557,N_26105,N_27149);
or U29558 (N_29558,N_27381,N_25619);
or U29559 (N_29559,N_27038,N_27433);
nor U29560 (N_29560,N_26694,N_26807);
and U29561 (N_29561,N_27150,N_26081);
xnor U29562 (N_29562,N_26605,N_25901);
xor U29563 (N_29563,N_27045,N_27279);
nor U29564 (N_29564,N_26154,N_25376);
or U29565 (N_29565,N_25587,N_27465);
nand U29566 (N_29566,N_25196,N_25712);
nor U29567 (N_29567,N_26707,N_27354);
or U29568 (N_29568,N_27151,N_26848);
nand U29569 (N_29569,N_25242,N_25938);
or U29570 (N_29570,N_26202,N_25608);
xnor U29571 (N_29571,N_27387,N_26975);
nand U29572 (N_29572,N_26468,N_25812);
nand U29573 (N_29573,N_25485,N_26830);
nand U29574 (N_29574,N_25217,N_27141);
xor U29575 (N_29575,N_26818,N_25642);
nand U29576 (N_29576,N_25470,N_26254);
nor U29577 (N_29577,N_25068,N_25213);
nor U29578 (N_29578,N_26042,N_26928);
xor U29579 (N_29579,N_25275,N_26480);
nand U29580 (N_29580,N_26022,N_26579);
or U29581 (N_29581,N_26580,N_26575);
nand U29582 (N_29582,N_25997,N_25042);
or U29583 (N_29583,N_26127,N_25709);
or U29584 (N_29584,N_26070,N_26204);
nand U29585 (N_29585,N_25552,N_25834);
nor U29586 (N_29586,N_25181,N_26227);
or U29587 (N_29587,N_26077,N_27406);
nor U29588 (N_29588,N_26746,N_25167);
and U29589 (N_29589,N_26556,N_25957);
nor U29590 (N_29590,N_26991,N_26990);
nor U29591 (N_29591,N_25165,N_27187);
nor U29592 (N_29592,N_25260,N_25819);
or U29593 (N_29593,N_26766,N_26424);
or U29594 (N_29594,N_27109,N_26931);
nor U29595 (N_29595,N_26062,N_26715);
xnor U29596 (N_29596,N_25653,N_25023);
xnor U29597 (N_29597,N_25536,N_26943);
nor U29598 (N_29598,N_27339,N_26856);
or U29599 (N_29599,N_26987,N_27292);
xor U29600 (N_29600,N_25655,N_26976);
and U29601 (N_29601,N_26860,N_27248);
nor U29602 (N_29602,N_25109,N_26729);
nand U29603 (N_29603,N_25681,N_26774);
and U29604 (N_29604,N_26180,N_27282);
and U29605 (N_29605,N_26078,N_26519);
nor U29606 (N_29606,N_26931,N_25166);
nor U29607 (N_29607,N_26917,N_27294);
nor U29608 (N_29608,N_25712,N_26459);
nand U29609 (N_29609,N_26663,N_26207);
nor U29610 (N_29610,N_25673,N_27409);
nor U29611 (N_29611,N_26508,N_26556);
nand U29612 (N_29612,N_26126,N_25461);
or U29613 (N_29613,N_25320,N_25359);
nand U29614 (N_29614,N_27095,N_26800);
nor U29615 (N_29615,N_26541,N_26335);
xor U29616 (N_29616,N_26502,N_25699);
and U29617 (N_29617,N_25078,N_26318);
nand U29618 (N_29618,N_27067,N_25429);
xnor U29619 (N_29619,N_26341,N_25465);
xor U29620 (N_29620,N_25227,N_27309);
or U29621 (N_29621,N_27189,N_26864);
or U29622 (N_29622,N_27049,N_25667);
nor U29623 (N_29623,N_26302,N_25255);
nand U29624 (N_29624,N_25629,N_26016);
or U29625 (N_29625,N_25665,N_26184);
or U29626 (N_29626,N_26199,N_26416);
xor U29627 (N_29627,N_26556,N_26433);
xnor U29628 (N_29628,N_27134,N_26169);
and U29629 (N_29629,N_27121,N_25102);
or U29630 (N_29630,N_26177,N_25092);
and U29631 (N_29631,N_25445,N_25239);
or U29632 (N_29632,N_26310,N_27394);
xor U29633 (N_29633,N_25851,N_26431);
and U29634 (N_29634,N_27413,N_26958);
nor U29635 (N_29635,N_25449,N_26288);
xor U29636 (N_29636,N_25131,N_27393);
nand U29637 (N_29637,N_27282,N_27032);
and U29638 (N_29638,N_25896,N_25794);
and U29639 (N_29639,N_25189,N_26621);
and U29640 (N_29640,N_25537,N_25386);
nor U29641 (N_29641,N_26887,N_27210);
xnor U29642 (N_29642,N_26432,N_26563);
nand U29643 (N_29643,N_26464,N_25673);
or U29644 (N_29644,N_25128,N_27186);
or U29645 (N_29645,N_27482,N_27250);
and U29646 (N_29646,N_27351,N_26298);
nor U29647 (N_29647,N_25523,N_27138);
and U29648 (N_29648,N_26887,N_26856);
nand U29649 (N_29649,N_25223,N_26639);
and U29650 (N_29650,N_25089,N_25653);
nor U29651 (N_29651,N_26823,N_26676);
xnor U29652 (N_29652,N_27302,N_25481);
nand U29653 (N_29653,N_25565,N_27078);
nor U29654 (N_29654,N_27357,N_26012);
nand U29655 (N_29655,N_25705,N_27041);
nor U29656 (N_29656,N_25147,N_25857);
nor U29657 (N_29657,N_25444,N_27210);
or U29658 (N_29658,N_26071,N_26797);
nand U29659 (N_29659,N_26628,N_27103);
nor U29660 (N_29660,N_25153,N_26799);
nand U29661 (N_29661,N_26546,N_25236);
xor U29662 (N_29662,N_25267,N_26993);
nand U29663 (N_29663,N_27151,N_27140);
nor U29664 (N_29664,N_26453,N_25120);
nor U29665 (N_29665,N_25744,N_27485);
and U29666 (N_29666,N_25140,N_25340);
nand U29667 (N_29667,N_26091,N_25017);
nand U29668 (N_29668,N_26768,N_27095);
xor U29669 (N_29669,N_25433,N_25457);
nand U29670 (N_29670,N_26889,N_26397);
xor U29671 (N_29671,N_26674,N_25774);
xnor U29672 (N_29672,N_26290,N_25314);
nand U29673 (N_29673,N_26906,N_25228);
nand U29674 (N_29674,N_27230,N_26928);
xor U29675 (N_29675,N_26915,N_25189);
or U29676 (N_29676,N_25557,N_27339);
or U29677 (N_29677,N_25610,N_25467);
and U29678 (N_29678,N_26813,N_25951);
xor U29679 (N_29679,N_27250,N_27417);
nand U29680 (N_29680,N_27198,N_25947);
and U29681 (N_29681,N_25758,N_26373);
and U29682 (N_29682,N_26918,N_25256);
nor U29683 (N_29683,N_26999,N_26649);
nand U29684 (N_29684,N_27048,N_25844);
xor U29685 (N_29685,N_26048,N_26006);
or U29686 (N_29686,N_25336,N_27187);
xor U29687 (N_29687,N_25982,N_26840);
nand U29688 (N_29688,N_26874,N_26546);
or U29689 (N_29689,N_25636,N_26613);
nand U29690 (N_29690,N_26222,N_26593);
and U29691 (N_29691,N_25645,N_26496);
nor U29692 (N_29692,N_27360,N_27461);
or U29693 (N_29693,N_26936,N_26911);
and U29694 (N_29694,N_26957,N_26220);
xnor U29695 (N_29695,N_26575,N_25251);
nand U29696 (N_29696,N_25776,N_25884);
xnor U29697 (N_29697,N_27239,N_26790);
xor U29698 (N_29698,N_25063,N_26434);
nand U29699 (N_29699,N_26057,N_26447);
or U29700 (N_29700,N_25379,N_25420);
nand U29701 (N_29701,N_25198,N_25675);
or U29702 (N_29702,N_27268,N_27378);
and U29703 (N_29703,N_26104,N_25949);
nand U29704 (N_29704,N_27115,N_26064);
nand U29705 (N_29705,N_27248,N_25721);
nor U29706 (N_29706,N_25576,N_26772);
xor U29707 (N_29707,N_27008,N_25329);
and U29708 (N_29708,N_26089,N_27481);
and U29709 (N_29709,N_26248,N_27279);
xor U29710 (N_29710,N_26910,N_26184);
nand U29711 (N_29711,N_25203,N_25658);
nor U29712 (N_29712,N_26577,N_27007);
nor U29713 (N_29713,N_25280,N_26769);
and U29714 (N_29714,N_25156,N_25583);
nand U29715 (N_29715,N_27393,N_27349);
and U29716 (N_29716,N_26929,N_25006);
and U29717 (N_29717,N_26171,N_27127);
xnor U29718 (N_29718,N_26912,N_25075);
nor U29719 (N_29719,N_26390,N_27478);
xnor U29720 (N_29720,N_26271,N_25650);
nor U29721 (N_29721,N_26795,N_27434);
or U29722 (N_29722,N_25777,N_27456);
or U29723 (N_29723,N_26591,N_27488);
xor U29724 (N_29724,N_27015,N_26201);
or U29725 (N_29725,N_25999,N_27290);
xnor U29726 (N_29726,N_26200,N_26225);
nand U29727 (N_29727,N_26461,N_25024);
nor U29728 (N_29728,N_27118,N_26172);
and U29729 (N_29729,N_25351,N_25508);
nor U29730 (N_29730,N_25483,N_25889);
or U29731 (N_29731,N_25518,N_27083);
nor U29732 (N_29732,N_26647,N_26773);
xor U29733 (N_29733,N_25771,N_25001);
nand U29734 (N_29734,N_26599,N_26281);
nand U29735 (N_29735,N_26399,N_25967);
nand U29736 (N_29736,N_25568,N_25591);
and U29737 (N_29737,N_25632,N_26998);
or U29738 (N_29738,N_25604,N_25792);
nor U29739 (N_29739,N_26306,N_27251);
nand U29740 (N_29740,N_27197,N_26216);
nand U29741 (N_29741,N_26011,N_26996);
and U29742 (N_29742,N_25645,N_25868);
xnor U29743 (N_29743,N_26289,N_27246);
or U29744 (N_29744,N_26517,N_25544);
nand U29745 (N_29745,N_25238,N_26264);
and U29746 (N_29746,N_25619,N_27474);
nand U29747 (N_29747,N_26172,N_26384);
nor U29748 (N_29748,N_25757,N_25436);
nand U29749 (N_29749,N_26667,N_26995);
nor U29750 (N_29750,N_25582,N_25388);
or U29751 (N_29751,N_26360,N_25273);
nor U29752 (N_29752,N_25528,N_25511);
xnor U29753 (N_29753,N_25567,N_25059);
xnor U29754 (N_29754,N_26659,N_26326);
and U29755 (N_29755,N_25217,N_25701);
or U29756 (N_29756,N_26148,N_27251);
nor U29757 (N_29757,N_25693,N_25002);
nor U29758 (N_29758,N_25516,N_25223);
nor U29759 (N_29759,N_25963,N_25821);
nand U29760 (N_29760,N_27227,N_26978);
and U29761 (N_29761,N_25516,N_25952);
nor U29762 (N_29762,N_26136,N_25688);
nor U29763 (N_29763,N_25743,N_25171);
or U29764 (N_29764,N_26672,N_25213);
nor U29765 (N_29765,N_25745,N_26179);
and U29766 (N_29766,N_26189,N_25118);
xor U29767 (N_29767,N_26145,N_26584);
and U29768 (N_29768,N_25284,N_25330);
nor U29769 (N_29769,N_25757,N_26550);
nand U29770 (N_29770,N_25193,N_25973);
nor U29771 (N_29771,N_25753,N_25386);
and U29772 (N_29772,N_25951,N_25479);
xor U29773 (N_29773,N_26312,N_26079);
nand U29774 (N_29774,N_27037,N_25747);
and U29775 (N_29775,N_25163,N_26414);
xnor U29776 (N_29776,N_26578,N_25786);
or U29777 (N_29777,N_26045,N_25595);
nand U29778 (N_29778,N_26227,N_26315);
or U29779 (N_29779,N_26970,N_26077);
nor U29780 (N_29780,N_25892,N_26819);
xor U29781 (N_29781,N_25244,N_27490);
nor U29782 (N_29782,N_25504,N_26257);
or U29783 (N_29783,N_27487,N_25899);
nand U29784 (N_29784,N_26451,N_26304);
or U29785 (N_29785,N_27402,N_26656);
nand U29786 (N_29786,N_26797,N_26316);
xor U29787 (N_29787,N_26304,N_25051);
or U29788 (N_29788,N_26264,N_25745);
nand U29789 (N_29789,N_25903,N_26054);
or U29790 (N_29790,N_27037,N_26941);
nor U29791 (N_29791,N_27021,N_26669);
xnor U29792 (N_29792,N_25612,N_26948);
nor U29793 (N_29793,N_26338,N_25222);
nor U29794 (N_29794,N_26670,N_25056);
xor U29795 (N_29795,N_26901,N_26446);
nor U29796 (N_29796,N_26662,N_25614);
xor U29797 (N_29797,N_25124,N_26429);
xor U29798 (N_29798,N_26326,N_25748);
nor U29799 (N_29799,N_25593,N_26293);
nand U29800 (N_29800,N_25600,N_26869);
nor U29801 (N_29801,N_26084,N_27378);
or U29802 (N_29802,N_26750,N_25290);
xnor U29803 (N_29803,N_25824,N_25131);
nand U29804 (N_29804,N_27005,N_26593);
or U29805 (N_29805,N_26625,N_27188);
nand U29806 (N_29806,N_26200,N_25672);
nand U29807 (N_29807,N_25257,N_25779);
and U29808 (N_29808,N_27305,N_25565);
nor U29809 (N_29809,N_26797,N_26743);
nor U29810 (N_29810,N_26257,N_26322);
nand U29811 (N_29811,N_25400,N_26001);
xnor U29812 (N_29812,N_27254,N_25343);
or U29813 (N_29813,N_26928,N_26271);
nand U29814 (N_29814,N_26793,N_25618);
and U29815 (N_29815,N_26687,N_27113);
nor U29816 (N_29816,N_25668,N_27117);
nor U29817 (N_29817,N_25249,N_25211);
nand U29818 (N_29818,N_27477,N_25326);
and U29819 (N_29819,N_26290,N_25672);
and U29820 (N_29820,N_26169,N_26830);
xnor U29821 (N_29821,N_27425,N_25610);
xnor U29822 (N_29822,N_26161,N_27111);
xor U29823 (N_29823,N_25925,N_27298);
and U29824 (N_29824,N_25834,N_26906);
and U29825 (N_29825,N_25766,N_26278);
nand U29826 (N_29826,N_26616,N_26907);
xor U29827 (N_29827,N_26412,N_27075);
and U29828 (N_29828,N_26212,N_27220);
nor U29829 (N_29829,N_26826,N_26636);
or U29830 (N_29830,N_27125,N_27223);
or U29831 (N_29831,N_25094,N_26493);
xnor U29832 (N_29832,N_26973,N_26541);
xnor U29833 (N_29833,N_26981,N_25694);
nand U29834 (N_29834,N_26202,N_25620);
or U29835 (N_29835,N_25039,N_25446);
or U29836 (N_29836,N_26828,N_26513);
nand U29837 (N_29837,N_25982,N_27064);
or U29838 (N_29838,N_25578,N_27130);
nor U29839 (N_29839,N_25481,N_27301);
xnor U29840 (N_29840,N_27175,N_25697);
nand U29841 (N_29841,N_26378,N_25471);
xor U29842 (N_29842,N_26366,N_27269);
nand U29843 (N_29843,N_26872,N_26952);
and U29844 (N_29844,N_25107,N_26837);
nand U29845 (N_29845,N_26990,N_25489);
or U29846 (N_29846,N_27388,N_25664);
nand U29847 (N_29847,N_26775,N_25801);
or U29848 (N_29848,N_27212,N_27459);
nand U29849 (N_29849,N_25733,N_25098);
and U29850 (N_29850,N_26360,N_26238);
and U29851 (N_29851,N_25180,N_25569);
nand U29852 (N_29852,N_26674,N_27466);
xor U29853 (N_29853,N_26806,N_26394);
nand U29854 (N_29854,N_26091,N_25566);
or U29855 (N_29855,N_26392,N_26247);
xnor U29856 (N_29856,N_25563,N_26703);
and U29857 (N_29857,N_26272,N_26611);
xor U29858 (N_29858,N_25811,N_26598);
nor U29859 (N_29859,N_25588,N_26175);
and U29860 (N_29860,N_25265,N_25330);
xor U29861 (N_29861,N_27476,N_27244);
and U29862 (N_29862,N_26424,N_26865);
or U29863 (N_29863,N_27147,N_26092);
xnor U29864 (N_29864,N_25164,N_27197);
and U29865 (N_29865,N_25944,N_27168);
nand U29866 (N_29866,N_26941,N_26057);
nor U29867 (N_29867,N_26700,N_27268);
nand U29868 (N_29868,N_25642,N_25277);
xnor U29869 (N_29869,N_25091,N_27220);
and U29870 (N_29870,N_26999,N_25732);
nor U29871 (N_29871,N_26787,N_26478);
xor U29872 (N_29872,N_25261,N_26026);
or U29873 (N_29873,N_25939,N_26357);
nand U29874 (N_29874,N_25861,N_26569);
nor U29875 (N_29875,N_26850,N_27331);
nor U29876 (N_29876,N_25355,N_25182);
nor U29877 (N_29877,N_26116,N_25318);
xnor U29878 (N_29878,N_25820,N_25290);
nor U29879 (N_29879,N_25238,N_26367);
nand U29880 (N_29880,N_27059,N_26642);
and U29881 (N_29881,N_27115,N_26777);
and U29882 (N_29882,N_26174,N_25978);
nor U29883 (N_29883,N_27224,N_25470);
or U29884 (N_29884,N_26354,N_27466);
or U29885 (N_29885,N_26512,N_26271);
and U29886 (N_29886,N_25143,N_27402);
or U29887 (N_29887,N_26006,N_25141);
or U29888 (N_29888,N_25976,N_26345);
or U29889 (N_29889,N_25108,N_27310);
nand U29890 (N_29890,N_27113,N_26992);
nor U29891 (N_29891,N_25043,N_25763);
xnor U29892 (N_29892,N_25201,N_27059);
and U29893 (N_29893,N_26258,N_26618);
or U29894 (N_29894,N_26575,N_27304);
or U29895 (N_29895,N_26871,N_25818);
nand U29896 (N_29896,N_25948,N_25614);
or U29897 (N_29897,N_27154,N_25284);
or U29898 (N_29898,N_26626,N_27036);
nand U29899 (N_29899,N_26539,N_25755);
xor U29900 (N_29900,N_26476,N_26841);
nor U29901 (N_29901,N_25676,N_26988);
nor U29902 (N_29902,N_25948,N_27114);
nor U29903 (N_29903,N_26695,N_26156);
nand U29904 (N_29904,N_27210,N_26696);
nor U29905 (N_29905,N_25187,N_26779);
nor U29906 (N_29906,N_26498,N_27107);
or U29907 (N_29907,N_27004,N_25468);
nor U29908 (N_29908,N_26479,N_25239);
or U29909 (N_29909,N_26322,N_25943);
nand U29910 (N_29910,N_25046,N_26606);
xor U29911 (N_29911,N_26329,N_25193);
xnor U29912 (N_29912,N_25624,N_27221);
nand U29913 (N_29913,N_25089,N_25790);
and U29914 (N_29914,N_26893,N_26972);
xnor U29915 (N_29915,N_27473,N_26171);
nor U29916 (N_29916,N_26891,N_25507);
xnor U29917 (N_29917,N_27199,N_25632);
nor U29918 (N_29918,N_25263,N_26286);
and U29919 (N_29919,N_26576,N_25162);
xnor U29920 (N_29920,N_27378,N_26885);
and U29921 (N_29921,N_25116,N_25015);
or U29922 (N_29922,N_25699,N_27270);
or U29923 (N_29923,N_25146,N_26301);
nor U29924 (N_29924,N_25927,N_25380);
or U29925 (N_29925,N_25923,N_26515);
and U29926 (N_29926,N_26654,N_26506);
nand U29927 (N_29927,N_26962,N_26388);
nor U29928 (N_29928,N_27304,N_25512);
xnor U29929 (N_29929,N_25961,N_26784);
or U29930 (N_29930,N_25349,N_25101);
and U29931 (N_29931,N_25425,N_25324);
nor U29932 (N_29932,N_25214,N_27473);
and U29933 (N_29933,N_25105,N_25532);
nand U29934 (N_29934,N_25087,N_26293);
nand U29935 (N_29935,N_26361,N_26085);
or U29936 (N_29936,N_27263,N_26452);
nor U29937 (N_29937,N_25252,N_27297);
nor U29938 (N_29938,N_25053,N_26388);
and U29939 (N_29939,N_25161,N_25880);
xnor U29940 (N_29940,N_26410,N_26247);
nor U29941 (N_29941,N_25189,N_26398);
nand U29942 (N_29942,N_26542,N_25839);
nand U29943 (N_29943,N_27013,N_26792);
nor U29944 (N_29944,N_25262,N_25892);
xnor U29945 (N_29945,N_25790,N_25869);
nand U29946 (N_29946,N_27350,N_26966);
nand U29947 (N_29947,N_25287,N_25464);
and U29948 (N_29948,N_27377,N_25729);
xor U29949 (N_29949,N_26217,N_25944);
nor U29950 (N_29950,N_25066,N_25616);
nor U29951 (N_29951,N_27252,N_25852);
or U29952 (N_29952,N_25790,N_27457);
xnor U29953 (N_29953,N_26201,N_26161);
or U29954 (N_29954,N_27001,N_25255);
and U29955 (N_29955,N_25860,N_27003);
xor U29956 (N_29956,N_25876,N_26231);
nand U29957 (N_29957,N_26648,N_25354);
xnor U29958 (N_29958,N_26703,N_25027);
or U29959 (N_29959,N_27443,N_26215);
xnor U29960 (N_29960,N_27267,N_27413);
nor U29961 (N_29961,N_26126,N_26330);
or U29962 (N_29962,N_25642,N_26447);
xnor U29963 (N_29963,N_25185,N_25508);
or U29964 (N_29964,N_26470,N_25989);
nor U29965 (N_29965,N_26500,N_25663);
xor U29966 (N_29966,N_27024,N_25431);
and U29967 (N_29967,N_26312,N_26599);
nand U29968 (N_29968,N_26284,N_25711);
xnor U29969 (N_29969,N_25407,N_25662);
and U29970 (N_29970,N_26884,N_26890);
and U29971 (N_29971,N_25268,N_26287);
xnor U29972 (N_29972,N_25207,N_26988);
or U29973 (N_29973,N_26005,N_27273);
xor U29974 (N_29974,N_25996,N_26901);
or U29975 (N_29975,N_25637,N_26354);
and U29976 (N_29976,N_25112,N_26815);
or U29977 (N_29977,N_25271,N_25873);
xnor U29978 (N_29978,N_25849,N_26638);
and U29979 (N_29979,N_27211,N_26214);
or U29980 (N_29980,N_27150,N_26955);
xor U29981 (N_29981,N_26438,N_26617);
and U29982 (N_29982,N_26558,N_26740);
or U29983 (N_29983,N_26857,N_25811);
nand U29984 (N_29984,N_26629,N_27027);
nand U29985 (N_29985,N_26721,N_25619);
and U29986 (N_29986,N_26995,N_26519);
and U29987 (N_29987,N_26409,N_27287);
nand U29988 (N_29988,N_25584,N_25630);
nand U29989 (N_29989,N_26224,N_25025);
xor U29990 (N_29990,N_25318,N_26002);
xor U29991 (N_29991,N_27372,N_27461);
and U29992 (N_29992,N_26355,N_26225);
and U29993 (N_29993,N_26461,N_27166);
xnor U29994 (N_29994,N_25639,N_27114);
and U29995 (N_29995,N_26617,N_26567);
nor U29996 (N_29996,N_26124,N_27245);
or U29997 (N_29997,N_26128,N_25847);
or U29998 (N_29998,N_25967,N_27033);
nor U29999 (N_29999,N_25705,N_25766);
or U30000 (N_30000,N_29900,N_29599);
or U30001 (N_30001,N_29158,N_28769);
and U30002 (N_30002,N_28132,N_27679);
xnor U30003 (N_30003,N_29032,N_28122);
xnor U30004 (N_30004,N_27617,N_28442);
or U30005 (N_30005,N_27911,N_28817);
xnor U30006 (N_30006,N_28449,N_28073);
xor U30007 (N_30007,N_27820,N_28406);
xnor U30008 (N_30008,N_28945,N_28051);
xor U30009 (N_30009,N_27762,N_29263);
xor U30010 (N_30010,N_29901,N_28460);
nand U30011 (N_30011,N_27959,N_28111);
or U30012 (N_30012,N_28522,N_28480);
and U30013 (N_30013,N_28933,N_29115);
xnor U30014 (N_30014,N_28917,N_28355);
or U30015 (N_30015,N_28053,N_28342);
and U30016 (N_30016,N_28528,N_27924);
xor U30017 (N_30017,N_28395,N_28687);
and U30018 (N_30018,N_27974,N_28661);
nor U30019 (N_30019,N_29097,N_27545);
nand U30020 (N_30020,N_29002,N_29378);
and U30021 (N_30021,N_27616,N_29689);
or U30022 (N_30022,N_29077,N_29027);
nand U30023 (N_30023,N_29707,N_28981);
and U30024 (N_30024,N_27783,N_28199);
nand U30025 (N_30025,N_28949,N_29774);
or U30026 (N_30026,N_28784,N_27878);
xnor U30027 (N_30027,N_29369,N_27703);
nand U30028 (N_30028,N_27773,N_29005);
nand U30029 (N_30029,N_28363,N_28403);
xnor U30030 (N_30030,N_28693,N_27810);
nor U30031 (N_30031,N_29946,N_27771);
or U30032 (N_30032,N_27704,N_29699);
or U30033 (N_30033,N_27894,N_29355);
and U30034 (N_30034,N_29483,N_29376);
nand U30035 (N_30035,N_28035,N_29358);
or U30036 (N_30036,N_28594,N_29804);
xor U30037 (N_30037,N_28867,N_28181);
xnor U30038 (N_30038,N_28531,N_27666);
xnor U30039 (N_30039,N_29773,N_28851);
and U30040 (N_30040,N_29653,N_29989);
nor U30041 (N_30041,N_29180,N_28649);
nor U30042 (N_30042,N_28941,N_28162);
or U30043 (N_30043,N_29570,N_27850);
or U30044 (N_30044,N_27578,N_28151);
nand U30045 (N_30045,N_28525,N_29433);
nand U30046 (N_30046,N_27505,N_27780);
and U30047 (N_30047,N_28086,N_29863);
and U30048 (N_30048,N_28796,N_27744);
xnor U30049 (N_30049,N_29450,N_28643);
nor U30050 (N_30050,N_27613,N_28716);
xnor U30051 (N_30051,N_27579,N_29073);
nor U30052 (N_30052,N_29882,N_29210);
or U30053 (N_30053,N_28588,N_28198);
and U30054 (N_30054,N_28623,N_28744);
or U30055 (N_30055,N_28112,N_29347);
or U30056 (N_30056,N_28014,N_29669);
or U30057 (N_30057,N_29566,N_28314);
nand U30058 (N_30058,N_28562,N_29472);
xor U30059 (N_30059,N_27951,N_28517);
and U30060 (N_30060,N_27740,N_28156);
nor U30061 (N_30061,N_29822,N_28402);
xnor U30062 (N_30062,N_27693,N_28082);
or U30063 (N_30063,N_27657,N_28367);
nand U30064 (N_30064,N_29585,N_29892);
xnor U30065 (N_30065,N_28019,N_28072);
or U30066 (N_30066,N_29473,N_27520);
or U30067 (N_30067,N_29515,N_29326);
nand U30068 (N_30068,N_28630,N_28325);
nor U30069 (N_30069,N_28662,N_29996);
and U30070 (N_30070,N_29943,N_29240);
nand U30071 (N_30071,N_29364,N_29510);
or U30072 (N_30072,N_27995,N_27735);
and U30073 (N_30073,N_29716,N_29408);
or U30074 (N_30074,N_28147,N_27635);
or U30075 (N_30075,N_28879,N_29475);
nor U30076 (N_30076,N_29666,N_29143);
xnor U30077 (N_30077,N_28564,N_29982);
nor U30078 (N_30078,N_27663,N_27950);
xor U30079 (N_30079,N_27640,N_28380);
nor U30080 (N_30080,N_27947,N_28202);
nor U30081 (N_30081,N_28795,N_28002);
and U30082 (N_30082,N_29542,N_29020);
and U30083 (N_30083,N_28898,N_28253);
or U30084 (N_30084,N_27993,N_28389);
xor U30085 (N_30085,N_28241,N_27538);
nand U30086 (N_30086,N_29603,N_28088);
nand U30087 (N_30087,N_29929,N_28100);
xor U30088 (N_30088,N_29001,N_28209);
and U30089 (N_30089,N_29646,N_28144);
nor U30090 (N_30090,N_29883,N_29648);
nor U30091 (N_30091,N_27596,N_28766);
nor U30092 (N_30092,N_29903,N_28811);
nor U30093 (N_30093,N_29543,N_29644);
and U30094 (N_30094,N_29250,N_29761);
nand U30095 (N_30095,N_29282,N_29563);
nor U30096 (N_30096,N_29322,N_29815);
and U30097 (N_30097,N_29502,N_28560);
or U30098 (N_30098,N_28794,N_27586);
and U30099 (N_30099,N_29306,N_27511);
nor U30100 (N_30100,N_29051,N_29036);
nand U30101 (N_30101,N_28464,N_29862);
or U30102 (N_30102,N_27753,N_28606);
or U30103 (N_30103,N_28552,N_27732);
nand U30104 (N_30104,N_29851,N_28024);
and U30105 (N_30105,N_29148,N_27712);
nor U30106 (N_30106,N_27925,N_28930);
and U30107 (N_30107,N_28809,N_28860);
xnor U30108 (N_30108,N_28826,N_28033);
xnor U30109 (N_30109,N_29942,N_28948);
nor U30110 (N_30110,N_28428,N_28154);
nor U30111 (N_30111,N_27814,N_28921);
and U30112 (N_30112,N_28686,N_28277);
nand U30113 (N_30113,N_29086,N_28283);
and U30114 (N_30114,N_29301,N_29278);
or U30115 (N_30115,N_28074,N_27769);
or U30116 (N_30116,N_28328,N_29744);
nor U30117 (N_30117,N_28773,N_29791);
and U30118 (N_30118,N_27557,N_27670);
and U30119 (N_30119,N_28441,N_29736);
and U30120 (N_30120,N_28967,N_28959);
or U30121 (N_30121,N_29676,N_28400);
xor U30122 (N_30122,N_29275,N_29190);
and U30123 (N_30123,N_28837,N_27842);
nor U30124 (N_30124,N_29065,N_28998);
nor U30125 (N_30125,N_27652,N_29714);
nor U30126 (N_30126,N_27790,N_28108);
or U30127 (N_30127,N_27718,N_28504);
nand U30128 (N_30128,N_28756,N_28094);
xnor U30129 (N_30129,N_29192,N_28276);
xor U30130 (N_30130,N_29448,N_28495);
or U30131 (N_30131,N_29198,N_27881);
or U30132 (N_30132,N_29695,N_29601);
nand U30133 (N_30133,N_27595,N_27509);
xor U30134 (N_30134,N_29541,N_29269);
xor U30135 (N_30135,N_28045,N_29485);
and U30136 (N_30136,N_28532,N_29911);
xnor U30137 (N_30137,N_27563,N_28566);
nor U30138 (N_30138,N_27831,N_29488);
nor U30139 (N_30139,N_28671,N_29303);
nor U30140 (N_30140,N_27943,N_27873);
nor U30141 (N_30141,N_29067,N_29308);
or U30142 (N_30142,N_27559,N_29746);
nand U30143 (N_30143,N_29954,N_29909);
and U30144 (N_30144,N_29368,N_28393);
nand U30145 (N_30145,N_28565,N_28150);
and U30146 (N_30146,N_27904,N_29110);
nand U30147 (N_30147,N_28250,N_27521);
nand U30148 (N_30148,N_28260,N_28281);
nor U30149 (N_30149,N_28884,N_28106);
or U30150 (N_30150,N_28071,N_27837);
nand U30151 (N_30151,N_28349,N_29517);
or U30152 (N_30152,N_27706,N_28865);
xnor U30153 (N_30153,N_27932,N_29516);
or U30154 (N_30154,N_29796,N_27705);
or U30155 (N_30155,N_27589,N_28059);
or U30156 (N_30156,N_28081,N_29486);
xor U30157 (N_30157,N_29589,N_28780);
nand U30158 (N_30158,N_29697,N_27664);
or U30159 (N_30159,N_29393,N_29343);
xor U30160 (N_30160,N_29017,N_29482);
nor U30161 (N_30161,N_28821,N_27689);
nor U30162 (N_30162,N_27877,N_29068);
and U30163 (N_30163,N_29614,N_29010);
nor U30164 (N_30164,N_28539,N_29569);
and U30165 (N_30165,N_29479,N_27685);
and U30166 (N_30166,N_28515,N_29135);
nor U30167 (N_30167,N_28842,N_27884);
xor U30168 (N_30168,N_28483,N_29767);
xnor U30169 (N_30169,N_27567,N_28477);
nand U30170 (N_30170,N_29604,N_29897);
nor U30171 (N_30171,N_27708,N_28688);
or U30172 (N_30172,N_29388,N_28484);
and U30173 (N_30173,N_28507,N_28702);
nor U30174 (N_30174,N_27998,N_28749);
nand U30175 (N_30175,N_29576,N_28203);
and U30176 (N_30176,N_28284,N_28412);
nor U30177 (N_30177,N_28740,N_28233);
nor U30178 (N_30178,N_28078,N_28801);
xnor U30179 (N_30179,N_29035,N_28447);
and U30180 (N_30180,N_27772,N_29532);
xor U30181 (N_30181,N_28899,N_28294);
nand U30182 (N_30182,N_27824,N_28908);
xor U30183 (N_30183,N_27898,N_27751);
and U30184 (N_30184,N_27677,N_29584);
xnor U30185 (N_30185,N_27817,N_29986);
nand U30186 (N_30186,N_29823,N_29772);
or U30187 (N_30187,N_28007,N_29285);
and U30188 (N_30188,N_27978,N_29613);
nor U30189 (N_30189,N_28500,N_28157);
nand U30190 (N_30190,N_29420,N_29317);
nand U30191 (N_30191,N_29212,N_29324);
nand U30192 (N_30192,N_27930,N_29867);
xnor U30193 (N_30193,N_28387,N_27870);
or U30194 (N_30194,N_29933,N_29089);
and U30195 (N_30195,N_28943,N_28624);
and U30196 (N_30196,N_29152,N_29012);
nor U30197 (N_30197,N_29905,N_29553);
and U30198 (N_30198,N_29164,N_29630);
nor U30199 (N_30199,N_29581,N_29749);
nand U30200 (N_30200,N_28476,N_29501);
xnor U30201 (N_30201,N_28365,N_28607);
nand U30202 (N_30202,N_28220,N_27671);
nor U30203 (N_30203,N_28788,N_28992);
xor U30204 (N_30204,N_28222,N_28267);
xnor U30205 (N_30205,N_29910,N_29594);
nor U30206 (N_30206,N_27886,N_27786);
xor U30207 (N_30207,N_29592,N_28559);
or U30208 (N_30208,N_28571,N_29498);
and U30209 (N_30209,N_29265,N_28734);
and U30210 (N_30210,N_28183,N_27902);
nand U30211 (N_30211,N_28543,N_27523);
nor U30212 (N_30212,N_29504,N_29264);
nor U30213 (N_30213,N_29559,N_27795);
xnor U30214 (N_30214,N_28574,N_27601);
nor U30215 (N_30215,N_28721,N_29527);
xor U30216 (N_30216,N_29865,N_28922);
xor U30217 (N_30217,N_27788,N_28771);
nor U30218 (N_30218,N_29023,N_27987);
nand U30219 (N_30219,N_27913,N_28416);
nand U30220 (N_30220,N_28603,N_28700);
xor U30221 (N_30221,N_29964,N_28980);
and U30222 (N_30222,N_28548,N_28118);
and U30223 (N_30223,N_28783,N_28168);
nand U30224 (N_30224,N_27848,N_28208);
and U30225 (N_30225,N_28085,N_29939);
nor U30226 (N_30226,N_27841,N_28158);
nand U30227 (N_30227,N_28768,N_29505);
nand U30228 (N_30228,N_28870,N_29006);
and U30229 (N_30229,N_29224,N_27941);
xor U30230 (N_30230,N_29509,N_28335);
nor U30231 (N_30231,N_29290,N_29400);
or U30232 (N_30232,N_28025,N_28117);
xor U30233 (N_30233,N_29366,N_27517);
nand U30234 (N_30234,N_28720,N_29932);
nand U30235 (N_30235,N_29987,N_28143);
and U30236 (N_30236,N_28333,N_29380);
or U30237 (N_30237,N_29332,N_28715);
nor U30238 (N_30238,N_29593,N_27871);
or U30239 (N_30239,N_28804,N_27979);
and U30240 (N_30240,N_28591,N_29354);
nand U30241 (N_30241,N_29350,N_29337);
xnor U30242 (N_30242,N_28474,N_28070);
and U30243 (N_30243,N_29430,N_29323);
nand U30244 (N_30244,N_29060,N_29832);
and U30245 (N_30245,N_29824,N_28261);
xor U30246 (N_30246,N_29629,N_29363);
nor U30247 (N_30247,N_28391,N_28535);
xor U30248 (N_30248,N_27525,N_28360);
or U30249 (N_30249,N_27912,N_28555);
and U30250 (N_30250,N_28758,N_28755);
nand U30251 (N_30251,N_29703,N_29793);
nor U30252 (N_30252,N_28966,N_29467);
or U30253 (N_30253,N_29805,N_29175);
nor U30254 (N_30254,N_29904,N_28269);
and U30255 (N_30255,N_29191,N_28883);
or U30256 (N_30256,N_28844,N_27518);
nor U30257 (N_30257,N_29064,N_27603);
or U30258 (N_30258,N_29225,N_29199);
xnor U30259 (N_30259,N_27593,N_29452);
nor U30260 (N_30260,N_29321,N_28841);
xor U30261 (N_30261,N_28174,N_28938);
nor U30262 (N_30262,N_28689,N_29621);
or U30263 (N_30263,N_29095,N_29030);
xor U30264 (N_30264,N_29745,N_29154);
and U30265 (N_30265,N_29829,N_27969);
nand U30266 (N_30266,N_27936,N_29950);
or U30267 (N_30267,N_29840,N_29312);
xnor U30268 (N_30268,N_28358,N_28832);
or U30269 (N_30269,N_28770,N_29319);
and U30270 (N_30270,N_28617,N_28888);
xnor U30271 (N_30271,N_29870,N_27605);
and U30272 (N_30272,N_29427,N_29550);
nor U30273 (N_30273,N_29846,N_29812);
nand U30274 (N_30274,N_29887,N_28582);
or U30275 (N_30275,N_29742,N_29918);
nor U30276 (N_30276,N_29525,N_27801);
nand U30277 (N_30277,N_29920,N_29560);
and U30278 (N_30278,N_28690,N_28502);
xor U30279 (N_30279,N_29179,N_29620);
xnor U30280 (N_30280,N_28102,N_27650);
nand U30281 (N_30281,N_29116,N_27628);
or U30282 (N_30282,N_29397,N_27840);
nor U30283 (N_30283,N_29398,N_28709);
xnor U30284 (N_30284,N_29137,N_28414);
nor U30285 (N_30285,N_27785,N_28526);
nor U30286 (N_30286,N_28779,N_28332);
nor U30287 (N_30287,N_28723,N_27917);
or U30288 (N_30288,N_28494,N_28904);
nand U30289 (N_30289,N_28044,N_29000);
xor U30290 (N_30290,N_28285,N_29552);
xnor U30291 (N_30291,N_28800,N_27519);
xor U30292 (N_30292,N_28853,N_29948);
and U30293 (N_30293,N_28429,N_28475);
nand U30294 (N_30294,N_27734,N_29792);
nor U30295 (N_30295,N_28994,N_28458);
or U30296 (N_30296,N_27639,N_29808);
and U30297 (N_30297,N_28608,N_28030);
or U30298 (N_30298,N_27526,N_29385);
xnor U30299 (N_30299,N_28834,N_29777);
nand U30300 (N_30300,N_28602,N_27606);
nand U30301 (N_30301,N_29723,N_29019);
nor U30302 (N_30302,N_27581,N_29710);
xor U30303 (N_30303,N_29582,N_29048);
nor U30304 (N_30304,N_28774,N_29281);
or U30305 (N_30305,N_28718,N_29302);
and U30306 (N_30306,N_28468,N_27592);
nand U30307 (N_30307,N_29133,N_28816);
xor U30308 (N_30308,N_29539,N_29186);
nand U30309 (N_30309,N_27763,N_29465);
and U30310 (N_30310,N_29720,N_29715);
and U30311 (N_30311,N_28644,N_29436);
or U30312 (N_30312,N_28159,N_29187);
xnor U30313 (N_30313,N_29880,N_29927);
and U30314 (N_30314,N_27674,N_27872);
and U30315 (N_30315,N_28371,N_29854);
or U30316 (N_30316,N_28558,N_27696);
nand U30317 (N_30317,N_29146,N_29026);
nor U30318 (N_30318,N_29174,N_28488);
nand U30319 (N_30319,N_28292,N_29480);
or U30320 (N_30320,N_29348,N_29349);
or U30321 (N_30321,N_29843,N_29114);
nor U30322 (N_30322,N_29518,N_29218);
xor U30323 (N_30323,N_29329,N_28009);
xor U30324 (N_30324,N_28553,N_27636);
and U30325 (N_30325,N_28300,N_28064);
xor U30326 (N_30326,N_28595,N_29864);
and U30327 (N_30327,N_27940,N_29841);
xor U30328 (N_30328,N_28954,N_29375);
xor U30329 (N_30329,N_28136,N_29298);
and U30330 (N_30330,N_29588,N_29468);
nand U30331 (N_30331,N_27667,N_29083);
nor U30332 (N_30332,N_29181,N_27745);
nor U30333 (N_30333,N_29776,N_28991);
xnor U30334 (N_30334,N_29770,N_29737);
nor U30335 (N_30335,N_29837,N_28704);
and U30336 (N_30336,N_29984,N_29222);
and U30337 (N_30337,N_28893,N_29506);
or U30338 (N_30338,N_29916,N_28972);
nor U30339 (N_30339,N_28829,N_29784);
nand U30340 (N_30340,N_28096,N_28694);
and U30341 (N_30341,N_29974,N_29196);
nor U30342 (N_30342,N_29658,N_28635);
xnor U30343 (N_30343,N_29995,N_28459);
or U30344 (N_30344,N_28211,N_28592);
and U30345 (N_30345,N_28481,N_29280);
nor U30346 (N_30346,N_28388,N_29262);
xor U30347 (N_30347,N_28666,N_28729);
xor U30348 (N_30348,N_28452,N_27514);
and U30349 (N_30349,N_27544,N_29670);
and U30350 (N_30350,N_29526,N_28383);
or U30351 (N_30351,N_28713,N_27991);
and U30352 (N_30352,N_27937,N_28145);
xnor U30353 (N_30353,N_29702,N_27737);
or U30354 (N_30354,N_28858,N_28316);
nand U30355 (N_30355,N_29674,N_29229);
or U30356 (N_30356,N_28301,N_28538);
xnor U30357 (N_30357,N_28152,N_28066);
or U30358 (N_30358,N_28748,N_28239);
nor U30359 (N_30359,N_29523,N_28750);
nor U30360 (N_30360,N_27632,N_28659);
xor U30361 (N_30361,N_27561,N_29411);
xor U30362 (N_30362,N_29320,N_27627);
or U30363 (N_30363,N_29660,N_29627);
nor U30364 (N_30364,N_29356,N_28008);
xnor U30365 (N_30365,N_29546,N_29463);
nor U30366 (N_30366,N_28172,N_27988);
nand U30367 (N_30367,N_28217,N_29561);
and U30368 (N_30368,N_28974,N_28519);
nand U30369 (N_30369,N_29980,N_29299);
xnor U30370 (N_30370,N_29925,N_27515);
and U30371 (N_30371,N_28485,N_28710);
nand U30372 (N_30372,N_29241,N_27507);
xor U30373 (N_30373,N_27854,N_29610);
and U30374 (N_30374,N_29979,N_27875);
and U30375 (N_30375,N_29432,N_29643);
or U30376 (N_30376,N_28196,N_29803);
nand U30377 (N_30377,N_28970,N_29171);
xor U30378 (N_30378,N_27680,N_27608);
nor U30379 (N_30379,N_28681,N_29100);
or U30380 (N_30380,N_29884,N_28576);
nor U30381 (N_30381,N_28663,N_29652);
nor U30382 (N_30382,N_28288,N_29247);
and U30383 (N_30383,N_29425,N_28337);
nand U30384 (N_30384,N_29845,N_27789);
or U30385 (N_30385,N_28141,N_28952);
nor U30386 (N_30386,N_27822,N_27760);
and U30387 (N_30387,N_28498,N_27836);
nor U30388 (N_30388,N_28180,N_27568);
nand U30389 (N_30389,N_29046,N_28736);
nand U30390 (N_30390,N_28937,N_27599);
nor U30391 (N_30391,N_29147,N_27710);
and U30392 (N_30392,N_29930,N_28712);
and U30393 (N_30393,N_27535,N_29300);
nand U30394 (N_30394,N_27956,N_29997);
nand U30395 (N_30395,N_28775,N_27825);
nor U30396 (N_30396,N_29415,N_28069);
or U30397 (N_30397,N_29284,N_29419);
nand U30398 (N_30398,N_28089,N_28385);
nor U30399 (N_30399,N_28242,N_28296);
nor U30400 (N_30400,N_29850,N_28423);
xnor U30401 (N_30401,N_27747,N_27591);
nor U30402 (N_30402,N_28909,N_28572);
xor U30403 (N_30403,N_28493,N_27803);
or U30404 (N_30404,N_29188,N_28808);
nand U30405 (N_30405,N_28651,N_29969);
xnor U30406 (N_30406,N_29434,N_29311);
nor U30407 (N_30407,N_28175,N_27725);
or U30408 (N_30408,N_28953,N_29216);
nor U30409 (N_30409,N_29693,N_29586);
nor U30410 (N_30410,N_29081,N_29912);
nor U30411 (N_30411,N_29287,N_28319);
and U30412 (N_30412,N_29888,N_29176);
nor U30413 (N_30413,N_27716,N_29377);
nor U30414 (N_30414,N_29968,N_28639);
xor U30415 (N_30415,N_29305,N_29600);
nand U30416 (N_30416,N_28581,N_28989);
nor U30417 (N_30417,N_29371,N_28955);
nor U30418 (N_30418,N_28999,N_29082);
nand U30419 (N_30419,N_28286,N_29106);
xor U30420 (N_30420,N_29608,N_27903);
or U30421 (N_30421,N_28184,N_27853);
nor U30422 (N_30422,N_29103,N_29474);
and U30423 (N_30423,N_27553,N_28121);
or U30424 (N_30424,N_28609,N_27975);
or U30425 (N_30425,N_29712,N_28633);
xor U30426 (N_30426,N_27990,N_28231);
and U30427 (N_30427,N_29072,N_28021);
and U30428 (N_30428,N_27529,N_29958);
nor U30429 (N_30429,N_29294,N_28062);
xnor U30430 (N_30430,N_29053,N_29978);
xnor U30431 (N_30431,N_29022,N_27598);
or U30432 (N_30432,N_27659,N_28219);
or U30433 (N_30433,N_29238,N_29437);
and U30434 (N_30434,N_28854,N_28445);
nand U30435 (N_30435,N_29858,N_28962);
xnor U30436 (N_30436,N_29748,N_29252);
nand U30437 (N_30437,N_28247,N_29220);
xor U30438 (N_30438,N_28900,N_28505);
nand U30439 (N_30439,N_28372,N_28944);
xor U30440 (N_30440,N_27742,N_29966);
nor U30441 (N_30441,N_29507,N_29551);
nand U30442 (N_30442,N_28964,N_29827);
and U30443 (N_30443,N_28031,N_28620);
xor U30444 (N_30444,N_28246,N_28448);
xor U30445 (N_30445,N_27893,N_29571);
and U30446 (N_30446,N_29835,N_27921);
xor U30447 (N_30447,N_27565,N_29047);
xor U30448 (N_30448,N_29424,N_29991);
or U30449 (N_30449,N_29395,N_29325);
nand U30450 (N_30450,N_29833,N_29664);
nor U30451 (N_30451,N_28965,N_27963);
and U30452 (N_30452,N_29780,N_29806);
nor U30453 (N_30453,N_29129,N_28824);
and U30454 (N_30454,N_27746,N_28119);
and U30455 (N_30455,N_28146,N_29149);
nor U30456 (N_30456,N_28266,N_28023);
xor U30457 (N_30457,N_27508,N_28664);
nand U30458 (N_30458,N_27889,N_28629);
nor U30459 (N_30459,N_28204,N_29800);
nor U30460 (N_30460,N_29766,N_29204);
or U30461 (N_30461,N_29487,N_28278);
nor U30462 (N_30462,N_28334,N_27855);
or U30463 (N_30463,N_29183,N_28856);
nor U30464 (N_30464,N_29994,N_27999);
xnor U30465 (N_30465,N_27590,N_29998);
nand U30466 (N_30466,N_29442,N_27954);
and U30467 (N_30467,N_28323,N_29362);
nand U30468 (N_30468,N_29173,N_28579);
nand U30469 (N_30469,N_29202,N_27835);
nor U30470 (N_30470,N_28929,N_27923);
nand U30471 (N_30471,N_28374,N_28491);
xor U30472 (N_30472,N_29700,N_27966);
and U30473 (N_30473,N_28392,N_28792);
and U30474 (N_30474,N_29423,N_27512);
xor U30475 (N_30475,N_27768,N_29524);
xnor U30476 (N_30476,N_29726,N_28384);
and U30477 (N_30477,N_29331,N_27739);
nor U30478 (N_30478,N_29813,N_27804);
xnor U30479 (N_30479,N_28855,N_28593);
or U30480 (N_30480,N_28487,N_28626);
and U30481 (N_30481,N_28546,N_29208);
xor U30482 (N_30482,N_29228,N_27976);
xnor U30483 (N_30483,N_27629,N_28058);
nor U30484 (N_30484,N_29144,N_29798);
nor U30485 (N_30485,N_29690,N_28272);
nor U30486 (N_30486,N_29727,N_29685);
nor U30487 (N_30487,N_28224,N_27765);
or U30488 (N_30488,N_28996,N_28373);
xor U30489 (N_30489,N_27675,N_28580);
or U30490 (N_30490,N_27630,N_28336);
nor U30491 (N_30491,N_28091,N_29595);
and U30492 (N_30492,N_28960,N_28830);
nand U30493 (N_30493,N_28616,N_28732);
or U30494 (N_30494,N_28754,N_28343);
or U30495 (N_30495,N_28437,N_29628);
nand U30496 (N_30496,N_27556,N_28223);
and U30497 (N_30497,N_27575,N_29557);
xnor U30498 (N_30498,N_28850,N_27624);
or U30499 (N_30499,N_29315,N_27953);
nand U30500 (N_30500,N_28719,N_28655);
xnor U30501 (N_30501,N_27916,N_29031);
nand U30502 (N_30502,N_27811,N_29227);
xor U30503 (N_30503,N_28864,N_29261);
nor U30504 (N_30504,N_29295,N_28273);
and U30505 (N_30505,N_27713,N_27736);
and U30506 (N_30506,N_29359,N_29492);
nor U30507 (N_30507,N_27543,N_29283);
xor U30508 (N_30508,N_29456,N_29038);
nand U30509 (N_30509,N_28497,N_29447);
or U30510 (N_30510,N_29965,N_29915);
nand U30511 (N_30511,N_29960,N_29536);
or U30512 (N_30512,N_27600,N_28728);
or U30513 (N_30513,N_29816,N_28596);
xor U30514 (N_30514,N_28701,N_29890);
xnor U30515 (N_30515,N_29616,N_29639);
xnor U30516 (N_30516,N_28262,N_29079);
and U30517 (N_30517,N_27516,N_28020);
xnor U30518 (N_30518,N_27815,N_28315);
and U30519 (N_30519,N_29008,N_28523);
nor U30520 (N_30520,N_29579,N_28310);
or U30521 (N_30521,N_29574,N_28248);
nor U30522 (N_30522,N_28382,N_28550);
nor U30523 (N_30523,N_28191,N_27660);
nand U30524 (N_30524,N_27564,N_28648);
nor U30525 (N_30525,N_27784,N_29878);
or U30526 (N_30526,N_28461,N_29041);
and U30527 (N_30527,N_28669,N_29399);
nand U30528 (N_30528,N_29678,N_28573);
nor U30529 (N_30529,N_29417,N_29454);
xnor U30530 (N_30530,N_29014,N_29522);
or U30531 (N_30531,N_28887,N_28645);
or U30532 (N_30532,N_29540,N_27702);
nor U30533 (N_30533,N_27727,N_29821);
nor U30534 (N_30534,N_27972,N_29394);
and U30535 (N_30535,N_27864,N_29092);
nand U30536 (N_30536,N_28492,N_29372);
and U30537 (N_30537,N_28149,N_27682);
nor U30538 (N_30538,N_28351,N_28984);
nand U30539 (N_30539,N_28129,N_29548);
nor U30540 (N_30540,N_27661,N_29093);
or U30541 (N_30541,N_28977,N_28785);
nand U30542 (N_30542,N_28257,N_27722);
or U30543 (N_30543,N_28983,N_27621);
and U30544 (N_30544,N_27571,N_29421);
nor U30545 (N_30545,N_28006,N_29839);
nand U30546 (N_30546,N_29743,N_28619);
nand U30547 (N_30547,N_29528,N_29963);
xnor U30548 (N_30548,N_29874,N_29131);
nand U30549 (N_30549,N_28894,N_27749);
or U30550 (N_30550,N_29206,N_27709);
nor U30551 (N_30551,N_29671,N_29453);
and U30552 (N_30552,N_29245,N_27918);
nor U30553 (N_30553,N_27692,N_28287);
xor U30554 (N_30554,N_29945,N_29127);
xor U30555 (N_30555,N_28611,N_28444);
xnor U30556 (N_30556,N_29799,N_27908);
and U30557 (N_30557,N_29769,N_29731);
or U30558 (N_30558,N_28182,N_29531);
nor U30559 (N_30559,N_27827,N_27909);
nor U30560 (N_30560,N_29957,N_27588);
or U30561 (N_30561,N_29713,N_28653);
and U30562 (N_30562,N_28760,N_28055);
and U30563 (N_30563,N_28741,N_27843);
xor U30564 (N_30564,N_29217,N_27607);
or U30565 (N_30565,N_27922,N_29439);
nand U30566 (N_30566,N_28311,N_28462);
nor U30567 (N_30567,N_28765,N_29213);
xor U30568 (N_30568,N_27996,N_28212);
nor U30569 (N_30569,N_28115,N_28435);
nand U30570 (N_30570,N_28379,N_27550);
nand U30571 (N_30571,N_28915,N_29209);
nand U30572 (N_30572,N_27750,N_28997);
nand U30573 (N_30573,N_29367,N_28583);
nor U30574 (N_30574,N_28434,N_28802);
and U30575 (N_30575,N_27847,N_28271);
nor U30576 (N_30576,N_28813,N_27539);
nand U30577 (N_30577,N_28703,N_28650);
or U30578 (N_30578,N_27962,N_27759);
nor U30579 (N_30579,N_28987,N_28003);
nor U30580 (N_30580,N_28040,N_29402);
or U30581 (N_30581,N_27558,N_29379);
or U30582 (N_30582,N_27860,N_29967);
xor U30583 (N_30583,N_29640,N_28421);
or U30584 (N_30584,N_29651,N_28105);
nor U30585 (N_30585,N_29215,N_29691);
nand U30586 (N_30586,N_28339,N_28407);
xor U30587 (N_30587,N_29338,N_28698);
nand U30588 (N_30588,N_27584,N_29617);
or U30589 (N_30589,N_28369,N_29902);
nand U30590 (N_30590,N_28932,N_28465);
and U30591 (N_30591,N_27994,N_29675);
nand U30592 (N_30592,N_28501,N_29908);
and U30593 (N_30593,N_29169,N_28309);
nand U30594 (N_30594,N_28782,N_28872);
and U30595 (N_30595,N_28846,N_28046);
and U30596 (N_30596,N_27668,N_29641);
and U30597 (N_30597,N_27501,N_28726);
or U30598 (N_30598,N_29830,N_28886);
nor U30599 (N_30599,N_29844,N_28737);
nand U30600 (N_30600,N_28575,N_29871);
or U30601 (N_30601,N_29386,N_27694);
nor U30602 (N_30602,N_29735,N_28496);
or U30603 (N_30603,N_27569,N_28187);
or U30604 (N_30604,N_28614,N_28752);
and U30605 (N_30605,N_28919,N_28889);
xor U30606 (N_30606,N_27541,N_28052);
and U30607 (N_30607,N_29751,N_28280);
nor U30608 (N_30608,N_29831,N_29396);
xor U30609 (N_30609,N_28724,N_28654);
xnor U30610 (N_30610,N_28450,N_29919);
nand U30611 (N_30611,N_29470,N_27819);
xnor U30612 (N_30612,N_29314,N_29373);
nand U30613 (N_30613,N_28628,N_29159);
or U30614 (N_30614,N_28544,N_28364);
nand U30615 (N_30615,N_29622,N_28098);
or U30616 (N_30616,N_28227,N_28797);
nand U30617 (N_30617,N_28652,N_27641);
and U30618 (N_30618,N_28398,N_29941);
nand U30619 (N_30619,N_29276,N_27821);
nand U30620 (N_30620,N_28759,N_27604);
and U30621 (N_30621,N_28988,N_28000);
xor U30622 (N_30622,N_29624,N_27698);
or U30623 (N_30623,N_29657,N_27961);
and U30624 (N_30624,N_28295,N_28969);
or U30625 (N_30625,N_28022,N_27882);
or U30626 (N_30626,N_29701,N_27555);
nand U30627 (N_30627,N_27551,N_29462);
nor U30628 (N_30628,N_29555,N_28104);
and U30629 (N_30629,N_28307,N_28142);
or U30630 (N_30630,N_29949,N_29330);
xnor U30631 (N_30631,N_27942,N_28345);
or U30632 (N_30632,N_29961,N_27948);
xor U30633 (N_30633,N_27676,N_27752);
nor U30634 (N_30634,N_29292,N_28430);
nor U30635 (N_30635,N_28397,N_28049);
nor U30636 (N_30636,N_28165,N_27546);
or U30637 (N_30637,N_29271,N_29661);
nand U30638 (N_30638,N_29221,N_29665);
nand U30639 (N_30639,N_29255,N_27834);
nor U30640 (N_30640,N_28290,N_28971);
nor U30641 (N_30641,N_29403,N_28054);
or U30642 (N_30642,N_29410,N_28926);
nand U30643 (N_30643,N_27929,N_29015);
nor U30644 (N_30644,N_29374,N_29272);
nand U30645 (N_30645,N_29977,N_27794);
and U30646 (N_30646,N_28679,N_27580);
nor U30647 (N_30647,N_29928,N_28197);
xor U30648 (N_30648,N_28895,N_29836);
and U30649 (N_30649,N_29931,N_27513);
nor U30650 (N_30650,N_29849,N_29534);
xor U30651 (N_30651,N_27920,N_28600);
and U30652 (N_30652,N_28490,N_27612);
nand U30653 (N_30653,N_28353,N_29170);
xnor U30654 (N_30654,N_28668,N_27868);
nand U30655 (N_30655,N_29580,N_28205);
nor U30656 (N_30656,N_28682,N_28015);
or U30657 (N_30657,N_29045,N_27900);
xnor U30658 (N_30658,N_29503,N_29404);
and U30659 (N_30659,N_27787,N_28786);
or U30660 (N_30660,N_29361,N_28951);
and U30661 (N_30661,N_29981,N_27833);
and U30662 (N_30662,N_29021,N_28957);
or U30663 (N_30663,N_29645,N_29441);
or U30664 (N_30664,N_29814,N_28123);
xnor U30665 (N_30665,N_28252,N_29786);
or U30666 (N_30666,N_27576,N_27828);
or U30667 (N_30667,N_29156,N_29316);
nand U30668 (N_30668,N_29681,N_29938);
nor U30669 (N_30669,N_29344,N_29304);
or U30670 (N_30670,N_28348,N_29426);
nand U30671 (N_30671,N_28245,N_28124);
and U30672 (N_30672,N_28413,N_27684);
or U30673 (N_30673,N_28320,N_28511);
or U30674 (N_30674,N_27823,N_29752);
and U30675 (N_30675,N_28376,N_29838);
xnor U30676 (N_30676,N_28299,N_28420);
nand U30677 (N_30677,N_28903,N_29054);
nand U30678 (N_30678,N_29230,N_28849);
nor U30679 (N_30679,N_28696,N_27754);
or U30680 (N_30680,N_28456,N_29070);
and U30681 (N_30681,N_29341,N_28210);
nor U30682 (N_30682,N_29273,N_27945);
nor U30683 (N_30683,N_28264,N_29891);
and U30684 (N_30684,N_28390,N_28767);
nor U30685 (N_30685,N_29917,N_27813);
nor U30686 (N_30686,N_29659,N_28885);
nor U30687 (N_30687,N_27662,N_28536);
and U30688 (N_30688,N_28961,N_28417);
and U30689 (N_30689,N_29688,N_28344);
or U30690 (N_30690,N_28327,N_27619);
nor U30691 (N_30691,N_27967,N_28790);
nor U30692 (N_30692,N_27719,N_28254);
nor U30693 (N_30693,N_28297,N_28293);
nand U30694 (N_30694,N_29893,N_29074);
nand U30695 (N_30695,N_29232,N_27934);
nand U30696 (N_30696,N_28394,N_28833);
and U30697 (N_30697,N_28090,N_29983);
nand U30698 (N_30698,N_29828,N_28274);
nor U30699 (N_30699,N_28179,N_27585);
and U30700 (N_30700,N_29759,N_27548);
and U30701 (N_30701,N_28258,N_29214);
or U30702 (N_30702,N_28330,N_27615);
nor U30703 (N_30703,N_27678,N_28680);
nand U30704 (N_30704,N_28137,N_29112);
nor U30705 (N_30705,N_29567,N_29168);
nand U30706 (N_30706,N_28561,N_28839);
xnor U30707 (N_30707,N_29868,N_29165);
or U30708 (N_30708,N_29236,N_27755);
or U30709 (N_30709,N_29512,N_28905);
xor U30710 (N_30710,N_28503,N_29059);
and U30711 (N_30711,N_27919,N_28079);
nand U30712 (N_30712,N_29732,N_27770);
and U30713 (N_30713,N_27861,N_27715);
xnor U30714 (N_30714,N_28975,N_27968);
nor U30715 (N_30715,N_28818,N_28130);
xor U30716 (N_30716,N_27970,N_29662);
nor U30717 (N_30717,N_29725,N_28516);
nand U30718 (N_30718,N_29099,N_29673);
nand U30719 (N_30719,N_28026,N_28057);
nor U30720 (N_30720,N_28510,N_29683);
nand U30721 (N_30721,N_28113,N_29826);
nand U30722 (N_30722,N_28167,N_27533);
nor U30723 (N_30723,N_28454,N_28861);
nor U30724 (N_30724,N_29952,N_29811);
nand U30725 (N_30725,N_28524,N_29605);
or U30726 (N_30726,N_29817,N_28578);
nand U30727 (N_30727,N_28587,N_27547);
nor U30728 (N_30728,N_29136,N_28169);
nor U30729 (N_30729,N_29872,N_28869);
nor U30730 (N_30730,N_27965,N_29360);
or U30731 (N_30731,N_29876,N_28831);
or U30732 (N_30732,N_28139,N_29856);
nor U30733 (N_30733,N_27989,N_29161);
xnor U30734 (N_30734,N_28289,N_28218);
xnor U30735 (N_30735,N_29547,N_29705);
nand U30736 (N_30736,N_27534,N_27985);
or U30737 (N_30737,N_29496,N_28268);
xnor U30738 (N_30738,N_28902,N_28585);
or U30739 (N_30739,N_28692,N_28746);
xor U30740 (N_30740,N_28727,N_28466);
nand U30741 (N_30741,N_28331,N_27933);
or U30742 (N_30742,N_28352,N_29063);
xnor U30743 (N_30743,N_28056,N_28995);
nor U30744 (N_30744,N_28225,N_29286);
nand U30745 (N_30745,N_27748,N_28541);
or U30746 (N_30746,N_28375,N_29788);
nand U30747 (N_30747,N_28092,N_29637);
or U30748 (N_30748,N_29018,N_28270);
xor U30749 (N_30749,N_27572,N_28791);
nand U30750 (N_30750,N_29677,N_27949);
nor U30751 (N_30751,N_28037,N_27764);
xnor U30752 (N_30752,N_28920,N_28979);
or U30753 (N_30753,N_28486,N_27594);
or U30754 (N_30754,N_29392,N_28647);
nor U30755 (N_30755,N_28127,N_28097);
or U30756 (N_30756,N_28799,N_29556);
xnor U30757 (N_30757,N_27807,N_29043);
nor U30758 (N_30758,N_27609,N_29591);
or U30759 (N_30759,N_28415,N_28632);
nand U30760 (N_30760,N_29999,N_27743);
or U30761 (N_30761,N_29632,N_28263);
nand U30762 (N_30762,N_29460,N_28793);
or U30763 (N_30763,N_29866,N_28660);
nand U30764 (N_30764,N_28916,N_27980);
nand U30765 (N_30765,N_27767,N_29383);
or U30766 (N_30766,N_29564,N_29993);
xnor U30767 (N_30767,N_29040,N_29268);
xor U30768 (N_30768,N_29758,N_28646);
and U30769 (N_30769,N_27914,N_28047);
nor U30770 (N_30770,N_28193,N_29500);
or U30771 (N_30771,N_28615,N_27844);
or U30772 (N_30772,N_28326,N_28370);
nor U30773 (N_30773,N_27901,N_27981);
and U30774 (N_30774,N_29078,N_29013);
and U30775 (N_30775,N_27611,N_29123);
and U30776 (N_30776,N_27733,N_27885);
or U30777 (N_30777,N_28016,N_29130);
or U30778 (N_30778,N_28757,N_28446);
nor U30779 (N_30779,N_28479,N_29606);
nand U30780 (N_30780,N_29708,N_28563);
nand U30781 (N_30781,N_29642,N_28171);
nand U30782 (N_30782,N_28230,N_27633);
and U30783 (N_30783,N_27537,N_28318);
nand U30784 (N_30784,N_29416,N_27646);
nor U30785 (N_30785,N_27879,N_27766);
or U30786 (N_30786,N_27738,N_29195);
nand U30787 (N_30787,N_29254,N_28739);
nand U30788 (N_30788,N_29738,N_29193);
nor U30789 (N_30789,N_28521,N_27758);
xor U30790 (N_30790,N_28673,N_29406);
or U30791 (N_30791,N_28812,N_29121);
nor U30792 (N_30792,N_29692,N_29687);
xor U30793 (N_30793,N_29297,N_29719);
xnor U30794 (N_30794,N_27683,N_28438);
nor U30795 (N_30795,N_29924,N_29698);
nand U30796 (N_30796,N_28063,N_27506);
or U30797 (N_30797,N_29973,N_28625);
and U30798 (N_30798,N_28968,N_28418);
nor U30799 (N_30799,N_29755,N_28569);
and U30800 (N_30800,N_28329,N_29775);
nor U30801 (N_30801,N_27960,N_28527);
xor U30802 (N_30802,N_27977,N_28243);
or U30803 (N_30803,N_29565,N_29233);
nand U30804 (N_30804,N_28599,N_29418);
or U30805 (N_30805,N_28419,N_28422);
and U30806 (N_30806,N_27731,N_27686);
or U30807 (N_30807,N_29650,N_29003);
xor U30808 (N_30808,N_28312,N_27729);
nor U30809 (N_30809,N_27644,N_29992);
nor U30810 (N_30810,N_28843,N_27863);
xor U30811 (N_30811,N_28549,N_29508);
xnor U30812 (N_30812,N_28717,N_27892);
nand U30813 (N_30813,N_28451,N_27928);
xnor U30814 (N_30814,N_27587,N_27812);
and U30815 (N_30815,N_29122,N_28163);
and U30816 (N_30816,N_28936,N_29655);
or U30817 (N_30817,N_28234,N_28471);
nor U30818 (N_30818,N_27876,N_29656);
nor U30819 (N_30819,N_29109,N_29970);
nand U30820 (N_30820,N_29401,N_28554);
nand U30821 (N_30821,N_28401,N_28776);
nand U30822 (N_30822,N_27573,N_29537);
nand U30823 (N_30823,N_29234,N_29061);
nand U30824 (N_30824,N_28236,N_28356);
nor U30825 (N_30825,N_29050,N_28282);
nand U30826 (N_30826,N_28923,N_27992);
and U30827 (N_30827,N_28381,N_27648);
nand U30828 (N_30828,N_29785,N_28973);
nand U30829 (N_30829,N_28805,N_28148);
nor U30830 (N_30830,N_29270,N_28279);
xor U30831 (N_30831,N_28001,N_28866);
nor U30832 (N_30832,N_28584,N_28806);
nand U30833 (N_30833,N_28133,N_29085);
and U30834 (N_30834,N_28906,N_29484);
and U30835 (N_30835,N_28787,N_29717);
and U30836 (N_30836,N_28506,N_29105);
or U30837 (N_30837,N_29107,N_29150);
xnor U30838 (N_30838,N_28568,N_27510);
nor U30839 (N_30839,N_28781,N_27890);
nand U30840 (N_30840,N_28076,N_29153);
or U30841 (N_30841,N_28017,N_27638);
and U30842 (N_30842,N_28508,N_28947);
xnor U30843 (N_30843,N_28912,N_28513);
and U30844 (N_30844,N_28963,N_29037);
nand U30845 (N_30845,N_28733,N_29921);
xor U30846 (N_30846,N_27910,N_29944);
nor U30847 (N_30847,N_29704,N_28924);
xnor U30848 (N_30848,N_28237,N_28306);
and U30849 (N_30849,N_27717,N_28347);
nand U30850 (N_30850,N_28814,N_28674);
and U30851 (N_30851,N_28892,N_29935);
nor U30852 (N_30852,N_29049,N_29291);
xor U30853 (N_30853,N_29985,N_28041);
xnor U30854 (N_30854,N_29583,N_28453);
or U30855 (N_30855,N_28170,N_28706);
nor U30856 (N_30856,N_28321,N_27699);
and U30857 (N_30857,N_29789,N_29899);
xor U30858 (N_30858,N_29869,N_29481);
xor U30859 (N_30859,N_28101,N_28638);
xnor U30860 (N_30860,N_28598,N_28520);
and U30861 (N_30861,N_27697,N_29988);
nor U30862 (N_30862,N_27955,N_28847);
nor U30863 (N_30863,N_28738,N_28178);
and U30864 (N_30864,N_29200,N_28730);
nand U30865 (N_30865,N_28881,N_29223);
xnor U30866 (N_30866,N_27846,N_27973);
nor U30867 (N_30867,N_27741,N_28067);
nand U30868 (N_30868,N_27634,N_28424);
nor U30869 (N_30869,N_27528,N_27527);
and U30870 (N_30870,N_28880,N_27711);
nor U30871 (N_30871,N_29219,N_28910);
xor U30872 (N_30872,N_28838,N_27701);
or U30873 (N_30873,N_28399,N_28114);
and U30874 (N_30874,N_27761,N_29444);
xor U30875 (N_30875,N_29724,N_28291);
or U30876 (N_30876,N_29926,N_29797);
nor U30877 (N_30877,N_29151,N_27938);
or U30878 (N_30878,N_27805,N_27797);
and U30879 (N_30879,N_28061,N_28827);
nand U30880 (N_30880,N_29087,N_29029);
xnor U30881 (N_30881,N_29184,N_29577);
or U30882 (N_30882,N_27798,N_28173);
and U30883 (N_30883,N_29457,N_29672);
or U30884 (N_30884,N_27658,N_29544);
nor U30885 (N_30885,N_29101,N_28534);
nand U30886 (N_30886,N_29801,N_28436);
nand U30887 (N_30887,N_27983,N_29310);
xor U30888 (N_30888,N_28093,N_28226);
nor U30889 (N_30889,N_27649,N_28443);
or U30890 (N_30890,N_28190,N_29499);
nor U30891 (N_30891,N_28126,N_28823);
or U30892 (N_30892,N_28641,N_27905);
nand U30893 (N_30893,N_27642,N_29145);
or U30894 (N_30894,N_29327,N_29455);
nand U30895 (N_30895,N_28762,N_27582);
or U30896 (N_30896,N_29721,N_28747);
and U30897 (N_30897,N_29446,N_27574);
nor U30898 (N_30898,N_29842,N_29134);
nor U30899 (N_30899,N_27887,N_28313);
xnor U30900 (N_30900,N_29011,N_28431);
nor U30901 (N_30901,N_29203,N_29848);
xor U30902 (N_30902,N_28134,N_28135);
or U30903 (N_30903,N_29108,N_28868);
nand U30904 (N_30904,N_29201,N_28533);
and U30905 (N_30905,N_29353,N_29119);
xor U30906 (N_30906,N_28707,N_29113);
xnor U30907 (N_30907,N_29042,N_29771);
xor U30908 (N_30908,N_28457,N_29923);
xor U30909 (N_30909,N_29818,N_29489);
nand U30910 (N_30910,N_29680,N_27554);
nand U30911 (N_30911,N_28695,N_29293);
xnor U30912 (N_30912,N_29913,N_28828);
or U30913 (N_30913,N_29118,N_29494);
xor U30914 (N_30914,N_28405,N_27927);
and U30915 (N_30915,N_27982,N_27793);
xor U30916 (N_30916,N_27852,N_28032);
nor U30917 (N_30917,N_29258,N_27653);
xnor U30918 (N_30918,N_28862,N_28404);
nand U30919 (N_30919,N_28499,N_29753);
nor U30920 (N_30920,N_27536,N_29609);
and U30921 (N_30921,N_29529,N_29231);
nand U30922 (N_30922,N_29873,N_28857);
nand U30923 (N_30923,N_29084,N_29384);
xor U30924 (N_30924,N_29936,N_28874);
or U30925 (N_30925,N_28873,N_28897);
and U30926 (N_30926,N_28545,N_28302);
nor U30927 (N_30927,N_28194,N_27891);
nand U30928 (N_30928,N_29340,N_29971);
or U30929 (N_30929,N_28518,N_27637);
or U30930 (N_30930,N_27957,N_28478);
nor U30931 (N_30931,N_29513,N_29471);
or U30932 (N_30932,N_27756,N_28004);
nand U30933 (N_30933,N_27799,N_29852);
or U30934 (N_30934,N_28354,N_29429);
xor U30935 (N_30935,N_27867,N_29934);
nor U30936 (N_30936,N_29497,N_27622);
nor U30937 (N_30937,N_28540,N_28612);
nand U30938 (N_30938,N_27687,N_28228);
nor U30939 (N_30939,N_29094,N_27874);
xnor U30940 (N_30940,N_29313,N_29351);
nand U30941 (N_30941,N_28845,N_28763);
nand U30942 (N_30942,N_28745,N_27845);
xor U30943 (N_30943,N_29590,N_28396);
or U30944 (N_30944,N_29469,N_27654);
nand U30945 (N_30945,N_29266,N_28820);
xor U30946 (N_30946,N_28107,N_29449);
and U30947 (N_30947,N_27560,N_28631);
nand U30948 (N_30948,N_29625,N_28697);
or U30949 (N_30949,N_29391,N_29157);
xor U30950 (N_30950,N_27935,N_28470);
xnor U30951 (N_30951,N_27583,N_29861);
nand U30952 (N_30952,N_29431,N_28034);
nor U30953 (N_30953,N_27880,N_27944);
or U30954 (N_30954,N_29328,N_29679);
and U30955 (N_30955,N_27723,N_28128);
or U30956 (N_30956,N_27778,N_28080);
xor U30957 (N_30957,N_27500,N_29167);
nand U30958 (N_30958,N_27645,N_29464);
and U30959 (N_30959,N_27899,N_27707);
xnor U30960 (N_30960,N_29795,N_28621);
or U30961 (N_30961,N_29886,N_29477);
nand U30962 (N_30962,N_28176,N_28927);
xnor U30963 (N_30963,N_28425,N_29091);
xor U30964 (N_30964,N_27832,N_29572);
nand U30965 (N_30965,N_28742,N_29575);
xor U30966 (N_30966,N_29649,N_27774);
or U30967 (N_30967,N_29959,N_29251);
nor U30968 (N_30968,N_29493,N_29155);
nor U30969 (N_30969,N_28099,N_27669);
nor U30970 (N_30970,N_29573,N_27964);
and U30971 (N_30971,N_29765,N_29768);
xor U30972 (N_30972,N_29289,N_29194);
xor U30973 (N_30973,N_29104,N_29602);
nor U30974 (N_30974,N_29879,N_27896);
nor U30975 (N_30975,N_27728,N_28083);
nand U30976 (N_30976,N_27623,N_28878);
nand U30977 (N_30977,N_28232,N_27779);
xnor U30978 (N_30978,N_28368,N_27796);
nand U30979 (N_30979,N_29847,N_29117);
nor U30980 (N_30980,N_29407,N_29618);
nor U30981 (N_30981,N_28950,N_28985);
and U30982 (N_30982,N_29098,N_28012);
xor U30983 (N_30983,N_27926,N_29519);
and U30984 (N_30984,N_27504,N_29318);
and U30985 (N_30985,N_28840,N_29102);
nor U30986 (N_30986,N_28803,N_28201);
or U30987 (N_30987,N_28155,N_27802);
nand U30988 (N_30988,N_28675,N_29587);
nor U30989 (N_30989,N_28634,N_27838);
xnor U30990 (N_30990,N_29956,N_28472);
nor U30991 (N_30991,N_29382,N_28308);
nor U30992 (N_30992,N_28618,N_29111);
nor U30993 (N_30993,N_29596,N_27522);
nor U30994 (N_30994,N_28275,N_28986);
nor U30995 (N_30995,N_28557,N_28362);
nand U30996 (N_30996,N_28542,N_27700);
or U30997 (N_30997,N_28725,N_29667);
nand U30998 (N_30998,N_29336,N_29730);
nand U30999 (N_30999,N_29189,N_28409);
nand U31000 (N_31000,N_28529,N_27907);
or U31001 (N_31001,N_28577,N_28590);
and U31002 (N_31002,N_29623,N_28439);
nand U31003 (N_31003,N_29389,N_28377);
or U31004 (N_31004,N_29459,N_27866);
nand U31005 (N_31005,N_27830,N_29825);
nand U31006 (N_31006,N_27958,N_29249);
or U31007 (N_31007,N_28216,N_29807);
xnor U31008 (N_31008,N_29779,N_29342);
and U31009 (N_31009,N_28939,N_29062);
nor U31010 (N_31010,N_29694,N_28240);
and U31011 (N_31011,N_27883,N_29728);
and U31012 (N_31012,N_28891,N_29257);
xnor U31013 (N_31013,N_29440,N_29538);
and U31014 (N_31014,N_29686,N_29663);
nor U31015 (N_31015,N_28341,N_28029);
and U31016 (N_31016,N_28551,N_29451);
or U31017 (N_31017,N_28340,N_28677);
or U31018 (N_31018,N_29860,N_29747);
and U31019 (N_31019,N_29741,N_28361);
or U31020 (N_31020,N_28901,N_27829);
nor U31021 (N_31021,N_28772,N_27816);
and U31022 (N_31022,N_28613,N_27726);
or U31023 (N_31023,N_28160,N_28039);
xor U31024 (N_31024,N_28065,N_27906);
or U31025 (N_31025,N_27695,N_27577);
nand U31026 (N_31026,N_28601,N_29740);
nand U31027 (N_31027,N_29533,N_29562);
nand U31028 (N_31028,N_28931,N_29057);
nand U31029 (N_31029,N_28670,N_27997);
nand U31030 (N_31030,N_29090,N_28683);
xnor U31031 (N_31031,N_29024,N_28303);
and U31032 (N_31032,N_29668,N_27651);
nand U31033 (N_31033,N_28798,N_29877);
and U31034 (N_31034,N_29160,N_28586);
or U31035 (N_31035,N_29096,N_28547);
nand U31036 (N_31036,N_27856,N_27809);
xor U31037 (N_31037,N_28684,N_28200);
nor U31038 (N_31038,N_28125,N_28489);
and U31039 (N_31039,N_29185,N_29857);
nand U31040 (N_31040,N_28836,N_28567);
xor U31041 (N_31041,N_28863,N_29080);
or U31042 (N_31042,N_29834,N_28982);
and U31043 (N_31043,N_29052,N_28244);
and U31044 (N_31044,N_28469,N_29783);
or U31045 (N_31045,N_29413,N_28077);
nor U31046 (N_31046,N_28907,N_29763);
and U31047 (N_31047,N_29940,N_29511);
or U31048 (N_31048,N_29554,N_28043);
and U31049 (N_31049,N_29033,N_28789);
nand U31050 (N_31050,N_27570,N_28038);
xor U31051 (N_31051,N_28530,N_28978);
and U31052 (N_31052,N_27730,N_29296);
nand U31053 (N_31053,N_28189,N_29009);
xor U31054 (N_31054,N_28935,N_28778);
and U31055 (N_31055,N_28570,N_29242);
xor U31056 (N_31056,N_28676,N_29055);
xor U31057 (N_31057,N_28743,N_28048);
xnor U31058 (N_31058,N_28512,N_27800);
nor U31059 (N_31059,N_27806,N_29764);
or U31060 (N_31060,N_27714,N_28140);
and U31061 (N_31061,N_29976,N_28622);
or U31062 (N_31062,N_28640,N_28060);
nand U31063 (N_31063,N_28807,N_28657);
nor U31064 (N_31064,N_28514,N_27681);
nor U31065 (N_31065,N_27691,N_29140);
and U31066 (N_31066,N_28463,N_27839);
and U31067 (N_31067,N_28256,N_28359);
xnor U31068 (N_31068,N_29458,N_28976);
and U31069 (N_31069,N_28213,N_27897);
or U31070 (N_31070,N_29345,N_28028);
or U31071 (N_31071,N_29476,N_28050);
or U31072 (N_31072,N_29235,N_28467);
nor U31073 (N_31073,N_28940,N_27782);
xnor U31074 (N_31074,N_27724,N_29568);
nand U31075 (N_31075,N_29207,N_28610);
xor U31076 (N_31076,N_27939,N_27859);
and U31077 (N_31077,N_29962,N_28642);
xnor U31078 (N_31078,N_29778,N_28131);
nand U31079 (N_31079,N_29922,N_28761);
and U31080 (N_31080,N_27971,N_29025);
xnor U31081 (N_31081,N_29520,N_28084);
xor U31082 (N_31082,N_29756,N_29288);
nand U31083 (N_31083,N_29889,N_28848);
nand U31084 (N_31084,N_28656,N_28011);
xor U31085 (N_31085,N_27566,N_29636);
xor U31086 (N_31086,N_27524,N_29438);
xnor U31087 (N_31087,N_27620,N_27540);
xnor U31088 (N_31088,N_29346,N_29445);
nand U31089 (N_31089,N_29390,N_28433);
or U31090 (N_31090,N_29937,N_27656);
nand U31091 (N_31091,N_29875,N_29237);
xor U31092 (N_31092,N_29066,N_29514);
xnor U31093 (N_31093,N_29243,N_28192);
xnor U31094 (N_31094,N_29253,N_27818);
nand U31095 (N_31095,N_28426,N_28699);
or U31096 (N_31096,N_27915,N_29125);
xor U31097 (N_31097,N_28877,N_28317);
or U31098 (N_31098,N_29684,N_29781);
nand U31099 (N_31099,N_27986,N_29859);
nor U31100 (N_31100,N_28928,N_27826);
and U31101 (N_31101,N_27672,N_27647);
or U31102 (N_31102,N_28195,N_28005);
or U31103 (N_31103,N_29635,N_27757);
or U31104 (N_31104,N_28138,N_28338);
and U31105 (N_31105,N_29260,N_28672);
xor U31106 (N_31106,N_28215,N_27857);
and U31107 (N_31107,N_27888,N_28186);
or U31108 (N_31108,N_29896,N_29357);
nand U31109 (N_31109,N_28161,N_29182);
or U31110 (N_31110,N_29016,N_28537);
nand U31111 (N_31111,N_29535,N_28010);
or U31112 (N_31112,N_29088,N_29244);
or U31113 (N_31113,N_28822,N_28605);
xor U31114 (N_31114,N_29787,N_29142);
nand U31115 (N_31115,N_29696,N_28597);
xor U31116 (N_31116,N_29139,N_29558);
nand U31117 (N_31117,N_27618,N_29132);
or U31118 (N_31118,N_28229,N_28238);
xnor U31119 (N_31119,N_27808,N_29124);
xnor U31120 (N_31120,N_29975,N_28322);
and U31121 (N_31121,N_29370,N_29007);
xnor U31122 (N_31122,N_27502,N_29898);
xnor U31123 (N_31123,N_28731,N_29709);
nor U31124 (N_31124,N_29820,N_28753);
nand U31125 (N_31125,N_28116,N_28604);
or U31126 (N_31126,N_29028,N_28153);
nor U31127 (N_31127,N_28075,N_28636);
xor U31128 (N_31128,N_28589,N_29762);
xor U31129 (N_31129,N_28859,N_27614);
or U31130 (N_31130,N_27720,N_29138);
nor U31131 (N_31131,N_29058,N_28925);
xnor U31132 (N_31132,N_27655,N_27643);
and U31133 (N_31133,N_28378,N_29647);
nand U31134 (N_31134,N_28890,N_28188);
and U31135 (N_31135,N_29075,N_29166);
and U31136 (N_31136,N_28914,N_27775);
nand U31137 (N_31137,N_28087,N_27777);
nor U31138 (N_31138,N_29172,N_28708);
and U31139 (N_31139,N_28473,N_29120);
and U31140 (N_31140,N_29711,N_29853);
xnor U31141 (N_31141,N_27610,N_29972);
nand U31142 (N_31142,N_28255,N_28411);
xnor U31143 (N_31143,N_29428,N_29521);
xnor U31144 (N_31144,N_29335,N_29729);
nor U31145 (N_31145,N_28298,N_27631);
xor U31146 (N_31146,N_28027,N_29478);
nand U31147 (N_31147,N_28455,N_27625);
xnor U31148 (N_31148,N_28120,N_29461);
and U31149 (N_31149,N_27984,N_29443);
or U31150 (N_31150,N_29633,N_28815);
and U31151 (N_31151,N_29333,N_29733);
or U31152 (N_31152,N_28324,N_29990);
nor U31153 (N_31153,N_27858,N_28185);
or U31154 (N_31154,N_28835,N_28304);
nor U31155 (N_31155,N_29895,N_29638);
xor U31156 (N_31156,N_29405,N_29381);
nand U31157 (N_31157,N_29466,N_27530);
and U31158 (N_31158,N_28685,N_28265);
nor U31159 (N_31159,N_29307,N_28691);
and U31160 (N_31160,N_28207,N_27851);
nor U31161 (N_31161,N_29631,N_29619);
nor U31162 (N_31162,N_29734,N_29760);
and U31163 (N_31163,N_28882,N_29069);
or U31164 (N_31164,N_29239,N_27532);
xnor U31165 (N_31165,N_29750,N_28259);
nand U31166 (N_31166,N_29722,N_28627);
nor U31167 (N_31167,N_29352,N_28913);
or U31168 (N_31168,N_29126,N_29248);
nor U31169 (N_31169,N_29615,N_29626);
nand U31170 (N_31170,N_29211,N_28357);
xnor U31171 (N_31171,N_29490,N_29739);
and U31172 (N_31172,N_27665,N_28103);
or U31173 (N_31173,N_29809,N_28705);
or U31174 (N_31174,N_28667,N_28956);
nand U31175 (N_31175,N_29682,N_28735);
and U31176 (N_31176,N_28875,N_28432);
xnor U31177 (N_31177,N_27946,N_29819);
nor U31178 (N_31178,N_29414,N_29162);
or U31179 (N_31179,N_29197,N_28386);
or U31180 (N_31180,N_29279,N_29309);
xor U31181 (N_31181,N_29906,N_29409);
or U31182 (N_31182,N_29277,N_28825);
nor U31183 (N_31183,N_27849,N_28440);
or U31184 (N_31184,N_28946,N_29530);
and U31185 (N_31185,N_28658,N_27626);
nand U31186 (N_31186,N_29706,N_28018);
nand U31187 (N_31187,N_29578,N_29004);
or U31188 (N_31188,N_29071,N_29612);
nor U31189 (N_31189,N_29654,N_28346);
nand U31190 (N_31190,N_28993,N_27792);
nand U31191 (N_31191,N_27531,N_28164);
nor U31192 (N_31192,N_29246,N_29267);
nor U31193 (N_31193,N_27688,N_29545);
nor U31194 (N_31194,N_28764,N_28042);
or U31195 (N_31195,N_27931,N_28166);
xor U31196 (N_31196,N_28556,N_28871);
nand U31197 (N_31197,N_29141,N_29894);
or U31198 (N_31198,N_28852,N_29491);
or U31199 (N_31199,N_29056,N_27503);
xnor U31200 (N_31200,N_28249,N_29274);
nand U31201 (N_31201,N_29914,N_29802);
xor U31202 (N_31202,N_28366,N_28896);
and U31203 (N_31203,N_29951,N_29855);
nor U31204 (N_31204,N_28714,N_28110);
or U31205 (N_31205,N_28427,N_28482);
nand U31206 (N_31206,N_28214,N_28221);
and U31207 (N_31207,N_29947,N_29634);
and U31208 (N_31208,N_29422,N_27673);
xnor U31209 (N_31209,N_28918,N_29718);
or U31210 (N_31210,N_28711,N_27562);
and U31211 (N_31211,N_29598,N_29256);
xor U31212 (N_31212,N_27869,N_28408);
nand U31213 (N_31213,N_28942,N_27952);
nor U31214 (N_31214,N_29365,N_28665);
and U31215 (N_31215,N_29607,N_29034);
nor U31216 (N_31216,N_29177,N_27690);
xor U31217 (N_31217,N_28722,N_27602);
xor U31218 (N_31218,N_29881,N_28911);
and U31219 (N_31219,N_28810,N_27776);
or U31220 (N_31220,N_29754,N_29794);
nor U31221 (N_31221,N_28305,N_29339);
nand U31222 (N_31222,N_29782,N_29597);
xnor U31223 (N_31223,N_28095,N_28751);
or U31224 (N_31224,N_29955,N_28177);
and U31225 (N_31225,N_29790,N_29259);
or U31226 (N_31226,N_28235,N_27549);
nor U31227 (N_31227,N_28777,N_29205);
nand U31228 (N_31228,N_28637,N_27895);
or U31229 (N_31229,N_29885,N_29128);
xnor U31230 (N_31230,N_27791,N_27597);
xor U31231 (N_31231,N_28509,N_27865);
nand U31232 (N_31232,N_27862,N_28109);
or U31233 (N_31233,N_29953,N_29334);
and U31234 (N_31234,N_29757,N_29387);
or U31235 (N_31235,N_27781,N_28206);
nand U31236 (N_31236,N_29178,N_27552);
and U31237 (N_31237,N_29044,N_28934);
and U31238 (N_31238,N_29810,N_29495);
xnor U31239 (N_31239,N_28036,N_27542);
and U31240 (N_31240,N_28013,N_29435);
or U31241 (N_31241,N_27721,N_28876);
and U31242 (N_31242,N_28350,N_28410);
xor U31243 (N_31243,N_29163,N_28678);
xnor U31244 (N_31244,N_28251,N_29611);
xor U31245 (N_31245,N_29907,N_28068);
and U31246 (N_31246,N_29412,N_29549);
xor U31247 (N_31247,N_29076,N_28958);
and U31248 (N_31248,N_29226,N_28990);
nand U31249 (N_31249,N_29039,N_28819);
or U31250 (N_31250,N_28241,N_29345);
and U31251 (N_31251,N_27562,N_28406);
or U31252 (N_31252,N_29049,N_27866);
and U31253 (N_31253,N_28762,N_28353);
or U31254 (N_31254,N_29874,N_28129);
or U31255 (N_31255,N_29811,N_28992);
nor U31256 (N_31256,N_29560,N_28418);
or U31257 (N_31257,N_27834,N_28114);
and U31258 (N_31258,N_27983,N_28978);
nor U31259 (N_31259,N_29292,N_28160);
and U31260 (N_31260,N_28338,N_27789);
xor U31261 (N_31261,N_29154,N_27510);
nor U31262 (N_31262,N_28849,N_29440);
or U31263 (N_31263,N_27517,N_28662);
and U31264 (N_31264,N_27946,N_27947);
or U31265 (N_31265,N_29479,N_29738);
xor U31266 (N_31266,N_27666,N_29602);
xnor U31267 (N_31267,N_27802,N_28720);
and U31268 (N_31268,N_27860,N_29796);
nand U31269 (N_31269,N_28143,N_29629);
or U31270 (N_31270,N_28867,N_29197);
nor U31271 (N_31271,N_29831,N_28139);
and U31272 (N_31272,N_28839,N_27648);
and U31273 (N_31273,N_29788,N_29282);
nor U31274 (N_31274,N_29562,N_28131);
or U31275 (N_31275,N_28588,N_29858);
xnor U31276 (N_31276,N_29259,N_29753);
xor U31277 (N_31277,N_29515,N_28054);
nand U31278 (N_31278,N_29192,N_28764);
xor U31279 (N_31279,N_29983,N_28936);
nand U31280 (N_31280,N_29362,N_27578);
xnor U31281 (N_31281,N_28050,N_28621);
and U31282 (N_31282,N_29438,N_27890);
and U31283 (N_31283,N_28783,N_29963);
xor U31284 (N_31284,N_27604,N_29705);
or U31285 (N_31285,N_29260,N_28640);
xor U31286 (N_31286,N_29352,N_29817);
nand U31287 (N_31287,N_28884,N_29667);
nand U31288 (N_31288,N_27577,N_28927);
nand U31289 (N_31289,N_29273,N_29795);
or U31290 (N_31290,N_27839,N_29837);
or U31291 (N_31291,N_29327,N_29927);
and U31292 (N_31292,N_29165,N_28904);
nor U31293 (N_31293,N_28918,N_29001);
nand U31294 (N_31294,N_29037,N_29878);
nand U31295 (N_31295,N_29427,N_29739);
and U31296 (N_31296,N_28645,N_27759);
nand U31297 (N_31297,N_27626,N_29826);
nor U31298 (N_31298,N_28773,N_28536);
nand U31299 (N_31299,N_29241,N_29791);
or U31300 (N_31300,N_28744,N_28567);
nor U31301 (N_31301,N_28503,N_27550);
nor U31302 (N_31302,N_29195,N_29200);
and U31303 (N_31303,N_27635,N_29804);
nand U31304 (N_31304,N_28604,N_28545);
nand U31305 (N_31305,N_29445,N_29410);
and U31306 (N_31306,N_29202,N_27597);
and U31307 (N_31307,N_27639,N_28413);
xnor U31308 (N_31308,N_27951,N_28209);
xnor U31309 (N_31309,N_28262,N_28017);
xor U31310 (N_31310,N_27817,N_29849);
nand U31311 (N_31311,N_27838,N_27983);
and U31312 (N_31312,N_28629,N_29954);
or U31313 (N_31313,N_28571,N_27936);
xnor U31314 (N_31314,N_27625,N_29614);
or U31315 (N_31315,N_28416,N_28134);
or U31316 (N_31316,N_29693,N_28657);
and U31317 (N_31317,N_28365,N_29862);
nor U31318 (N_31318,N_28739,N_29892);
xor U31319 (N_31319,N_28670,N_29526);
nand U31320 (N_31320,N_27928,N_27891);
or U31321 (N_31321,N_29567,N_28930);
nand U31322 (N_31322,N_28110,N_28598);
nor U31323 (N_31323,N_29445,N_28006);
nand U31324 (N_31324,N_28820,N_29231);
and U31325 (N_31325,N_27525,N_28443);
or U31326 (N_31326,N_29117,N_27935);
or U31327 (N_31327,N_28080,N_27752);
nor U31328 (N_31328,N_28993,N_29642);
and U31329 (N_31329,N_28711,N_29855);
and U31330 (N_31330,N_29416,N_27867);
xor U31331 (N_31331,N_29352,N_28413);
or U31332 (N_31332,N_27913,N_28887);
and U31333 (N_31333,N_28380,N_28199);
nor U31334 (N_31334,N_27921,N_28718);
nor U31335 (N_31335,N_29899,N_29587);
xor U31336 (N_31336,N_28957,N_29792);
nand U31337 (N_31337,N_28105,N_29007);
nand U31338 (N_31338,N_29987,N_28312);
nand U31339 (N_31339,N_27924,N_28521);
nor U31340 (N_31340,N_29477,N_28652);
xnor U31341 (N_31341,N_29041,N_29318);
xnor U31342 (N_31342,N_27793,N_27666);
xnor U31343 (N_31343,N_28905,N_29934);
nand U31344 (N_31344,N_29837,N_27814);
xnor U31345 (N_31345,N_27968,N_28765);
and U31346 (N_31346,N_28461,N_27882);
nor U31347 (N_31347,N_29517,N_27557);
xnor U31348 (N_31348,N_29284,N_29575);
xor U31349 (N_31349,N_29285,N_28244);
nor U31350 (N_31350,N_29001,N_28265);
xor U31351 (N_31351,N_28598,N_28951);
and U31352 (N_31352,N_27687,N_29335);
or U31353 (N_31353,N_28960,N_28543);
xnor U31354 (N_31354,N_29596,N_29392);
xnor U31355 (N_31355,N_29386,N_29951);
xnor U31356 (N_31356,N_28855,N_29170);
and U31357 (N_31357,N_29000,N_29573);
nor U31358 (N_31358,N_27517,N_28669);
and U31359 (N_31359,N_28352,N_28577);
and U31360 (N_31360,N_27961,N_29060);
or U31361 (N_31361,N_29696,N_27851);
or U31362 (N_31362,N_29648,N_29087);
nand U31363 (N_31363,N_28708,N_28606);
nand U31364 (N_31364,N_28909,N_28570);
or U31365 (N_31365,N_28688,N_28800);
and U31366 (N_31366,N_27996,N_28543);
and U31367 (N_31367,N_29431,N_28327);
or U31368 (N_31368,N_29558,N_27559);
nor U31369 (N_31369,N_28128,N_28669);
xnor U31370 (N_31370,N_29912,N_29720);
and U31371 (N_31371,N_29268,N_28784);
xnor U31372 (N_31372,N_28617,N_29734);
xor U31373 (N_31373,N_28742,N_28189);
and U31374 (N_31374,N_29887,N_29866);
or U31375 (N_31375,N_29151,N_28343);
and U31376 (N_31376,N_28376,N_28039);
nor U31377 (N_31377,N_29365,N_29620);
nand U31378 (N_31378,N_27991,N_28889);
xnor U31379 (N_31379,N_27755,N_29888);
xnor U31380 (N_31380,N_28478,N_29625);
nor U31381 (N_31381,N_29870,N_27709);
or U31382 (N_31382,N_28441,N_28503);
or U31383 (N_31383,N_27830,N_28732);
or U31384 (N_31384,N_27910,N_28866);
nand U31385 (N_31385,N_29092,N_28055);
xnor U31386 (N_31386,N_27929,N_28314);
xnor U31387 (N_31387,N_29584,N_29128);
nor U31388 (N_31388,N_29136,N_29773);
nor U31389 (N_31389,N_27868,N_27538);
and U31390 (N_31390,N_28025,N_28705);
nor U31391 (N_31391,N_28865,N_29735);
or U31392 (N_31392,N_28109,N_28684);
or U31393 (N_31393,N_28529,N_27518);
and U31394 (N_31394,N_29202,N_29564);
nand U31395 (N_31395,N_29209,N_28377);
nor U31396 (N_31396,N_27726,N_27563);
or U31397 (N_31397,N_27671,N_28333);
or U31398 (N_31398,N_28201,N_28062);
nand U31399 (N_31399,N_28508,N_29892);
nor U31400 (N_31400,N_29967,N_27507);
or U31401 (N_31401,N_27675,N_28031);
nand U31402 (N_31402,N_28284,N_29056);
and U31403 (N_31403,N_28455,N_29531);
and U31404 (N_31404,N_28458,N_28998);
or U31405 (N_31405,N_28346,N_28528);
and U31406 (N_31406,N_28871,N_29023);
xor U31407 (N_31407,N_28640,N_28083);
nand U31408 (N_31408,N_27856,N_27925);
or U31409 (N_31409,N_27823,N_27794);
and U31410 (N_31410,N_28658,N_29691);
and U31411 (N_31411,N_27733,N_28971);
or U31412 (N_31412,N_28011,N_29695);
nor U31413 (N_31413,N_29159,N_28210);
nand U31414 (N_31414,N_28311,N_28190);
or U31415 (N_31415,N_29947,N_29891);
or U31416 (N_31416,N_28841,N_27984);
and U31417 (N_31417,N_29255,N_28813);
and U31418 (N_31418,N_28277,N_29858);
nand U31419 (N_31419,N_29385,N_29564);
nand U31420 (N_31420,N_27995,N_29169);
nor U31421 (N_31421,N_29198,N_29861);
or U31422 (N_31422,N_27946,N_29274);
nor U31423 (N_31423,N_27702,N_28734);
or U31424 (N_31424,N_29444,N_29965);
and U31425 (N_31425,N_29991,N_29931);
nor U31426 (N_31426,N_28629,N_28739);
and U31427 (N_31427,N_28224,N_29067);
nand U31428 (N_31428,N_29903,N_27683);
or U31429 (N_31429,N_29950,N_29423);
nor U31430 (N_31430,N_29559,N_28748);
or U31431 (N_31431,N_27596,N_27502);
nor U31432 (N_31432,N_29620,N_29635);
and U31433 (N_31433,N_28570,N_28015);
nand U31434 (N_31434,N_28591,N_27559);
xnor U31435 (N_31435,N_27532,N_29873);
and U31436 (N_31436,N_29290,N_27728);
or U31437 (N_31437,N_27554,N_29213);
nor U31438 (N_31438,N_27542,N_28987);
xor U31439 (N_31439,N_27891,N_29407);
or U31440 (N_31440,N_27750,N_27500);
nor U31441 (N_31441,N_29455,N_29638);
and U31442 (N_31442,N_27844,N_29920);
xnor U31443 (N_31443,N_28289,N_29687);
xnor U31444 (N_31444,N_28114,N_28434);
and U31445 (N_31445,N_28255,N_28808);
and U31446 (N_31446,N_28271,N_27618);
and U31447 (N_31447,N_29928,N_28151);
or U31448 (N_31448,N_28588,N_29005);
nor U31449 (N_31449,N_29927,N_27608);
xor U31450 (N_31450,N_28241,N_29785);
or U31451 (N_31451,N_28551,N_28511);
nor U31452 (N_31452,N_27840,N_27580);
nor U31453 (N_31453,N_29602,N_27541);
or U31454 (N_31454,N_29044,N_27788);
nor U31455 (N_31455,N_29115,N_29867);
nand U31456 (N_31456,N_28662,N_29208);
nor U31457 (N_31457,N_28816,N_27763);
or U31458 (N_31458,N_29239,N_29790);
or U31459 (N_31459,N_29233,N_29936);
nand U31460 (N_31460,N_28979,N_29421);
xnor U31461 (N_31461,N_28123,N_27748);
and U31462 (N_31462,N_29798,N_29878);
xor U31463 (N_31463,N_29344,N_27955);
nand U31464 (N_31464,N_28710,N_28069);
xnor U31465 (N_31465,N_28703,N_29323);
and U31466 (N_31466,N_28778,N_29005);
nand U31467 (N_31467,N_29260,N_29421);
or U31468 (N_31468,N_28238,N_28676);
or U31469 (N_31469,N_29856,N_29384);
nor U31470 (N_31470,N_29871,N_29715);
nand U31471 (N_31471,N_29384,N_28702);
xor U31472 (N_31472,N_28002,N_28234);
xor U31473 (N_31473,N_29453,N_29963);
and U31474 (N_31474,N_28525,N_28890);
xor U31475 (N_31475,N_27983,N_27792);
and U31476 (N_31476,N_29528,N_28124);
or U31477 (N_31477,N_28385,N_29815);
nor U31478 (N_31478,N_29588,N_27816);
nor U31479 (N_31479,N_29339,N_27803);
nand U31480 (N_31480,N_29723,N_29299);
nand U31481 (N_31481,N_27570,N_29020);
xnor U31482 (N_31482,N_28879,N_29167);
nor U31483 (N_31483,N_28906,N_29447);
or U31484 (N_31484,N_29044,N_29936);
and U31485 (N_31485,N_29116,N_29481);
and U31486 (N_31486,N_29854,N_27880);
or U31487 (N_31487,N_28557,N_28017);
nand U31488 (N_31488,N_28125,N_29315);
xnor U31489 (N_31489,N_28535,N_29013);
xor U31490 (N_31490,N_29357,N_29364);
or U31491 (N_31491,N_28500,N_28576);
or U31492 (N_31492,N_28143,N_28199);
or U31493 (N_31493,N_29975,N_28525);
nand U31494 (N_31494,N_28159,N_28541);
and U31495 (N_31495,N_28465,N_28013);
nand U31496 (N_31496,N_27619,N_28174);
and U31497 (N_31497,N_29729,N_29384);
or U31498 (N_31498,N_28861,N_29526);
xor U31499 (N_31499,N_28696,N_29069);
and U31500 (N_31500,N_28867,N_29082);
nand U31501 (N_31501,N_29558,N_28254);
nand U31502 (N_31502,N_27937,N_28758);
or U31503 (N_31503,N_29025,N_27610);
or U31504 (N_31504,N_27612,N_29416);
xnor U31505 (N_31505,N_29601,N_29094);
xor U31506 (N_31506,N_29018,N_29161);
or U31507 (N_31507,N_29522,N_28448);
nor U31508 (N_31508,N_28874,N_28097);
nand U31509 (N_31509,N_27758,N_29456);
nand U31510 (N_31510,N_28898,N_27972);
nand U31511 (N_31511,N_27613,N_29225);
and U31512 (N_31512,N_29829,N_28028);
nor U31513 (N_31513,N_29216,N_27900);
and U31514 (N_31514,N_28185,N_27939);
or U31515 (N_31515,N_27548,N_28389);
or U31516 (N_31516,N_27670,N_28321);
or U31517 (N_31517,N_29738,N_27703);
nor U31518 (N_31518,N_27980,N_27894);
nor U31519 (N_31519,N_29580,N_29619);
nor U31520 (N_31520,N_29702,N_28799);
nand U31521 (N_31521,N_29826,N_27945);
nor U31522 (N_31522,N_28708,N_27598);
and U31523 (N_31523,N_27641,N_29205);
xor U31524 (N_31524,N_27998,N_27503);
and U31525 (N_31525,N_27719,N_29977);
or U31526 (N_31526,N_27781,N_29902);
nand U31527 (N_31527,N_28352,N_29555);
xor U31528 (N_31528,N_27669,N_28000);
nand U31529 (N_31529,N_27821,N_29875);
nor U31530 (N_31530,N_28021,N_29306);
xor U31531 (N_31531,N_29338,N_28839);
nand U31532 (N_31532,N_28382,N_29393);
nand U31533 (N_31533,N_27649,N_28598);
or U31534 (N_31534,N_28307,N_28804);
xor U31535 (N_31535,N_27887,N_29379);
nand U31536 (N_31536,N_29024,N_28168);
or U31537 (N_31537,N_29611,N_29767);
and U31538 (N_31538,N_27905,N_28494);
or U31539 (N_31539,N_27625,N_29049);
nor U31540 (N_31540,N_28074,N_29882);
xnor U31541 (N_31541,N_27571,N_29949);
nor U31542 (N_31542,N_28081,N_29361);
nor U31543 (N_31543,N_27588,N_28595);
xor U31544 (N_31544,N_28649,N_28973);
nor U31545 (N_31545,N_29268,N_27997);
or U31546 (N_31546,N_29136,N_28323);
or U31547 (N_31547,N_28141,N_28868);
nand U31548 (N_31548,N_28449,N_27808);
or U31549 (N_31549,N_27865,N_27651);
or U31550 (N_31550,N_28950,N_28071);
and U31551 (N_31551,N_28527,N_28876);
nand U31552 (N_31552,N_29578,N_29511);
and U31553 (N_31553,N_29404,N_28319);
or U31554 (N_31554,N_28711,N_29923);
nor U31555 (N_31555,N_27521,N_27637);
nand U31556 (N_31556,N_28595,N_29193);
and U31557 (N_31557,N_28726,N_28880);
xor U31558 (N_31558,N_28539,N_29798);
or U31559 (N_31559,N_29442,N_29142);
or U31560 (N_31560,N_27866,N_28842);
and U31561 (N_31561,N_28630,N_27720);
or U31562 (N_31562,N_29634,N_29879);
xnor U31563 (N_31563,N_27770,N_28928);
xor U31564 (N_31564,N_28943,N_27888);
nor U31565 (N_31565,N_27648,N_27805);
xnor U31566 (N_31566,N_29576,N_28156);
nand U31567 (N_31567,N_29780,N_28016);
nor U31568 (N_31568,N_29278,N_27931);
xnor U31569 (N_31569,N_29412,N_27826);
xor U31570 (N_31570,N_28886,N_28475);
nand U31571 (N_31571,N_27784,N_29824);
nor U31572 (N_31572,N_28954,N_27878);
nand U31573 (N_31573,N_28939,N_29600);
and U31574 (N_31574,N_28691,N_29555);
and U31575 (N_31575,N_27896,N_29894);
or U31576 (N_31576,N_29583,N_28373);
and U31577 (N_31577,N_28793,N_28689);
xnor U31578 (N_31578,N_28076,N_28651);
nand U31579 (N_31579,N_29907,N_29052);
or U31580 (N_31580,N_27609,N_28701);
nor U31581 (N_31581,N_29153,N_29126);
or U31582 (N_31582,N_28645,N_28220);
and U31583 (N_31583,N_28495,N_28861);
nor U31584 (N_31584,N_27915,N_29265);
nor U31585 (N_31585,N_28605,N_29531);
nor U31586 (N_31586,N_27958,N_28904);
or U31587 (N_31587,N_28939,N_28269);
or U31588 (N_31588,N_27520,N_29516);
and U31589 (N_31589,N_28454,N_28674);
nand U31590 (N_31590,N_29954,N_29826);
nand U31591 (N_31591,N_28191,N_29508);
and U31592 (N_31592,N_29134,N_27965);
or U31593 (N_31593,N_29307,N_28097);
nor U31594 (N_31594,N_28338,N_28430);
nand U31595 (N_31595,N_28695,N_28846);
nand U31596 (N_31596,N_29078,N_28656);
and U31597 (N_31597,N_28769,N_28836);
nand U31598 (N_31598,N_29261,N_29567);
nand U31599 (N_31599,N_28915,N_29037);
nand U31600 (N_31600,N_29477,N_29128);
nor U31601 (N_31601,N_27673,N_29106);
nand U31602 (N_31602,N_27715,N_28607);
xor U31603 (N_31603,N_28519,N_28002);
xnor U31604 (N_31604,N_29984,N_27762);
or U31605 (N_31605,N_27709,N_28473);
nand U31606 (N_31606,N_28485,N_28714);
and U31607 (N_31607,N_27699,N_28380);
nand U31608 (N_31608,N_28356,N_28074);
nand U31609 (N_31609,N_29423,N_27629);
nor U31610 (N_31610,N_28555,N_27994);
nor U31611 (N_31611,N_29086,N_29981);
xnor U31612 (N_31612,N_28444,N_28329);
and U31613 (N_31613,N_28194,N_29342);
nand U31614 (N_31614,N_29196,N_28946);
nor U31615 (N_31615,N_28732,N_27502);
or U31616 (N_31616,N_29471,N_29865);
nand U31617 (N_31617,N_29642,N_28678);
nor U31618 (N_31618,N_28911,N_29347);
and U31619 (N_31619,N_29695,N_28141);
nand U31620 (N_31620,N_29522,N_28479);
or U31621 (N_31621,N_28834,N_29580);
nor U31622 (N_31622,N_29625,N_27802);
and U31623 (N_31623,N_28500,N_29698);
or U31624 (N_31624,N_28767,N_27984);
nor U31625 (N_31625,N_27865,N_27790);
and U31626 (N_31626,N_29166,N_27821);
or U31627 (N_31627,N_28255,N_29241);
or U31628 (N_31628,N_28464,N_27867);
xor U31629 (N_31629,N_28811,N_28429);
nor U31630 (N_31630,N_29885,N_28508);
or U31631 (N_31631,N_27968,N_29981);
nand U31632 (N_31632,N_29640,N_28226);
nand U31633 (N_31633,N_28938,N_28889);
or U31634 (N_31634,N_28878,N_28443);
and U31635 (N_31635,N_28263,N_28605);
nor U31636 (N_31636,N_29113,N_28539);
or U31637 (N_31637,N_29963,N_27912);
and U31638 (N_31638,N_29603,N_28668);
nand U31639 (N_31639,N_29133,N_27843);
xor U31640 (N_31640,N_29811,N_29495);
xor U31641 (N_31641,N_28986,N_27822);
nor U31642 (N_31642,N_28695,N_28321);
and U31643 (N_31643,N_28400,N_28932);
nand U31644 (N_31644,N_28210,N_27702);
nor U31645 (N_31645,N_29395,N_29178);
or U31646 (N_31646,N_29606,N_27757);
or U31647 (N_31647,N_28783,N_29498);
nor U31648 (N_31648,N_28709,N_29650);
nand U31649 (N_31649,N_28682,N_28327);
or U31650 (N_31650,N_28028,N_29180);
nor U31651 (N_31651,N_28684,N_29626);
nor U31652 (N_31652,N_28197,N_28207);
and U31653 (N_31653,N_27592,N_29419);
nand U31654 (N_31654,N_27814,N_28299);
or U31655 (N_31655,N_28016,N_28397);
xnor U31656 (N_31656,N_29183,N_29710);
or U31657 (N_31657,N_28878,N_28475);
xor U31658 (N_31658,N_27991,N_28515);
nor U31659 (N_31659,N_28372,N_28277);
or U31660 (N_31660,N_29186,N_29808);
nor U31661 (N_31661,N_29076,N_28663);
nand U31662 (N_31662,N_28526,N_28658);
nor U31663 (N_31663,N_27715,N_27506);
and U31664 (N_31664,N_27723,N_29101);
nand U31665 (N_31665,N_28741,N_27818);
nor U31666 (N_31666,N_27866,N_28180);
nor U31667 (N_31667,N_29770,N_28485);
xor U31668 (N_31668,N_29935,N_28893);
and U31669 (N_31669,N_28432,N_27516);
nand U31670 (N_31670,N_27931,N_28505);
xnor U31671 (N_31671,N_28663,N_29205);
xnor U31672 (N_31672,N_29165,N_29172);
nand U31673 (N_31673,N_29721,N_28870);
or U31674 (N_31674,N_27672,N_27660);
xnor U31675 (N_31675,N_27703,N_27803);
nand U31676 (N_31676,N_29776,N_27782);
xnor U31677 (N_31677,N_28271,N_28053);
or U31678 (N_31678,N_29181,N_27614);
nand U31679 (N_31679,N_29240,N_28076);
or U31680 (N_31680,N_29621,N_27508);
and U31681 (N_31681,N_28274,N_29905);
nand U31682 (N_31682,N_29827,N_28459);
or U31683 (N_31683,N_28189,N_29683);
and U31684 (N_31684,N_29001,N_28053);
or U31685 (N_31685,N_27875,N_29601);
nand U31686 (N_31686,N_28011,N_28471);
nor U31687 (N_31687,N_29272,N_28472);
nor U31688 (N_31688,N_29099,N_27985);
nand U31689 (N_31689,N_29620,N_29589);
and U31690 (N_31690,N_29380,N_27933);
or U31691 (N_31691,N_28694,N_28334);
xnor U31692 (N_31692,N_28606,N_27899);
nor U31693 (N_31693,N_29515,N_29154);
xnor U31694 (N_31694,N_29440,N_27862);
nor U31695 (N_31695,N_27713,N_29549);
or U31696 (N_31696,N_29907,N_27687);
nor U31697 (N_31697,N_29789,N_28218);
and U31698 (N_31698,N_29537,N_28800);
nor U31699 (N_31699,N_28590,N_28980);
and U31700 (N_31700,N_29857,N_28956);
and U31701 (N_31701,N_28995,N_28269);
and U31702 (N_31702,N_29845,N_28461);
nor U31703 (N_31703,N_28009,N_28889);
nand U31704 (N_31704,N_28474,N_28055);
or U31705 (N_31705,N_28544,N_28582);
and U31706 (N_31706,N_27796,N_29646);
and U31707 (N_31707,N_28303,N_27506);
and U31708 (N_31708,N_28716,N_29420);
nand U31709 (N_31709,N_28767,N_28634);
nand U31710 (N_31710,N_29104,N_27972);
xor U31711 (N_31711,N_28047,N_27847);
and U31712 (N_31712,N_28968,N_29365);
or U31713 (N_31713,N_29119,N_28509);
or U31714 (N_31714,N_29148,N_29334);
and U31715 (N_31715,N_29270,N_29773);
and U31716 (N_31716,N_28678,N_29455);
or U31717 (N_31717,N_29087,N_29506);
xnor U31718 (N_31718,N_28731,N_27692);
or U31719 (N_31719,N_29389,N_27849);
nor U31720 (N_31720,N_27684,N_27549);
and U31721 (N_31721,N_29309,N_29533);
nand U31722 (N_31722,N_27735,N_29535);
nand U31723 (N_31723,N_27978,N_29576);
nor U31724 (N_31724,N_29226,N_28356);
nor U31725 (N_31725,N_28041,N_27886);
nor U31726 (N_31726,N_28031,N_27705);
nor U31727 (N_31727,N_29182,N_29608);
nor U31728 (N_31728,N_28038,N_28197);
nand U31729 (N_31729,N_29804,N_27884);
nor U31730 (N_31730,N_29949,N_28697);
xor U31731 (N_31731,N_29724,N_28842);
xnor U31732 (N_31732,N_29209,N_29455);
and U31733 (N_31733,N_27874,N_28363);
and U31734 (N_31734,N_27911,N_27759);
xnor U31735 (N_31735,N_28852,N_28428);
nor U31736 (N_31736,N_28886,N_27863);
nand U31737 (N_31737,N_28629,N_28860);
xor U31738 (N_31738,N_27581,N_28068);
nand U31739 (N_31739,N_28896,N_28889);
and U31740 (N_31740,N_27748,N_29783);
or U31741 (N_31741,N_28208,N_29477);
and U31742 (N_31742,N_28722,N_28103);
nand U31743 (N_31743,N_28758,N_27536);
nor U31744 (N_31744,N_29671,N_28722);
or U31745 (N_31745,N_28328,N_29606);
or U31746 (N_31746,N_29049,N_28150);
and U31747 (N_31747,N_28695,N_29457);
nor U31748 (N_31748,N_28914,N_29093);
and U31749 (N_31749,N_27667,N_29637);
or U31750 (N_31750,N_29483,N_28740);
nor U31751 (N_31751,N_28849,N_28746);
nor U31752 (N_31752,N_28398,N_27987);
or U31753 (N_31753,N_27959,N_29860);
xor U31754 (N_31754,N_29924,N_28871);
xnor U31755 (N_31755,N_29535,N_29051);
xor U31756 (N_31756,N_29906,N_28514);
or U31757 (N_31757,N_29363,N_27820);
xnor U31758 (N_31758,N_27838,N_28135);
nand U31759 (N_31759,N_29747,N_28165);
xor U31760 (N_31760,N_29102,N_29825);
or U31761 (N_31761,N_28246,N_28754);
xnor U31762 (N_31762,N_28191,N_28848);
or U31763 (N_31763,N_29628,N_29546);
xor U31764 (N_31764,N_27963,N_28142);
nor U31765 (N_31765,N_28366,N_27603);
xor U31766 (N_31766,N_29384,N_28196);
or U31767 (N_31767,N_28046,N_27923);
nand U31768 (N_31768,N_28651,N_29653);
nor U31769 (N_31769,N_29342,N_28814);
or U31770 (N_31770,N_28548,N_29761);
xnor U31771 (N_31771,N_28748,N_28126);
nor U31772 (N_31772,N_28323,N_28402);
or U31773 (N_31773,N_28605,N_28244);
nor U31774 (N_31774,N_29937,N_29159);
xor U31775 (N_31775,N_29733,N_28741);
or U31776 (N_31776,N_29858,N_27915);
xnor U31777 (N_31777,N_28855,N_29799);
xor U31778 (N_31778,N_28539,N_28892);
xnor U31779 (N_31779,N_29597,N_28882);
xor U31780 (N_31780,N_29626,N_28177);
and U31781 (N_31781,N_29368,N_28043);
and U31782 (N_31782,N_29491,N_29694);
xnor U31783 (N_31783,N_28305,N_28203);
and U31784 (N_31784,N_29499,N_29893);
and U31785 (N_31785,N_28140,N_28838);
xnor U31786 (N_31786,N_29267,N_28623);
or U31787 (N_31787,N_29427,N_28142);
nand U31788 (N_31788,N_28502,N_29765);
xor U31789 (N_31789,N_27950,N_28326);
xnor U31790 (N_31790,N_28865,N_27557);
nor U31791 (N_31791,N_29629,N_27938);
and U31792 (N_31792,N_28222,N_29939);
nor U31793 (N_31793,N_29036,N_28071);
nand U31794 (N_31794,N_29653,N_28076);
xnor U31795 (N_31795,N_27563,N_29779);
nand U31796 (N_31796,N_28290,N_28013);
or U31797 (N_31797,N_29198,N_28821);
nor U31798 (N_31798,N_29395,N_28106);
nor U31799 (N_31799,N_28574,N_28614);
xor U31800 (N_31800,N_27802,N_28829);
or U31801 (N_31801,N_28226,N_27761);
xnor U31802 (N_31802,N_29767,N_28062);
xor U31803 (N_31803,N_28248,N_29932);
xor U31804 (N_31804,N_29963,N_29695);
and U31805 (N_31805,N_27947,N_28138);
xor U31806 (N_31806,N_29904,N_29068);
nand U31807 (N_31807,N_27918,N_29848);
or U31808 (N_31808,N_29125,N_28135);
and U31809 (N_31809,N_28965,N_28400);
nor U31810 (N_31810,N_29778,N_29458);
xnor U31811 (N_31811,N_27550,N_29261);
nand U31812 (N_31812,N_29343,N_29611);
xor U31813 (N_31813,N_27956,N_29727);
nand U31814 (N_31814,N_29873,N_27791);
nand U31815 (N_31815,N_27852,N_27507);
xor U31816 (N_31816,N_27997,N_28054);
xor U31817 (N_31817,N_28640,N_28619);
nand U31818 (N_31818,N_28705,N_28841);
and U31819 (N_31819,N_28461,N_29249);
xor U31820 (N_31820,N_27885,N_28511);
xor U31821 (N_31821,N_28629,N_27560);
or U31822 (N_31822,N_29945,N_29902);
nor U31823 (N_31823,N_28571,N_28435);
xor U31824 (N_31824,N_27770,N_28810);
xnor U31825 (N_31825,N_28835,N_27660);
nand U31826 (N_31826,N_29070,N_29111);
or U31827 (N_31827,N_29342,N_27582);
xnor U31828 (N_31828,N_29585,N_29101);
xnor U31829 (N_31829,N_29723,N_29266);
and U31830 (N_31830,N_29198,N_28167);
and U31831 (N_31831,N_27682,N_28303);
nor U31832 (N_31832,N_28186,N_29293);
xnor U31833 (N_31833,N_29059,N_29235);
and U31834 (N_31834,N_29811,N_27945);
or U31835 (N_31835,N_27859,N_29682);
xor U31836 (N_31836,N_29354,N_29274);
nor U31837 (N_31837,N_27602,N_27839);
nand U31838 (N_31838,N_29402,N_28439);
or U31839 (N_31839,N_29675,N_29300);
nor U31840 (N_31840,N_28558,N_29008);
xnor U31841 (N_31841,N_28803,N_28005);
and U31842 (N_31842,N_27986,N_29422);
and U31843 (N_31843,N_28575,N_28756);
nor U31844 (N_31844,N_28977,N_27602);
or U31845 (N_31845,N_27856,N_28102);
nand U31846 (N_31846,N_28170,N_27936);
nor U31847 (N_31847,N_29880,N_28459);
nand U31848 (N_31848,N_29245,N_27859);
nor U31849 (N_31849,N_28898,N_27968);
xor U31850 (N_31850,N_28133,N_28879);
xnor U31851 (N_31851,N_28112,N_29125);
xnor U31852 (N_31852,N_28559,N_29497);
xor U31853 (N_31853,N_27979,N_29152);
nand U31854 (N_31854,N_28513,N_29751);
and U31855 (N_31855,N_29619,N_29430);
or U31856 (N_31856,N_28655,N_28682);
xnor U31857 (N_31857,N_29941,N_28252);
xor U31858 (N_31858,N_29274,N_29392);
and U31859 (N_31859,N_28263,N_27511);
xnor U31860 (N_31860,N_28939,N_28938);
or U31861 (N_31861,N_28621,N_29618);
xnor U31862 (N_31862,N_27979,N_28611);
nand U31863 (N_31863,N_29501,N_28031);
xor U31864 (N_31864,N_29655,N_27509);
nor U31865 (N_31865,N_27601,N_28158);
or U31866 (N_31866,N_28259,N_28112);
xnor U31867 (N_31867,N_29349,N_28804);
nand U31868 (N_31868,N_27984,N_27524);
xor U31869 (N_31869,N_28321,N_28478);
or U31870 (N_31870,N_27820,N_29944);
nand U31871 (N_31871,N_27981,N_29350);
xnor U31872 (N_31872,N_29977,N_28307);
and U31873 (N_31873,N_28687,N_29512);
nand U31874 (N_31874,N_29390,N_29479);
and U31875 (N_31875,N_28134,N_29433);
nand U31876 (N_31876,N_27565,N_27869);
nand U31877 (N_31877,N_29853,N_27901);
and U31878 (N_31878,N_27539,N_29181);
xnor U31879 (N_31879,N_27820,N_27923);
nand U31880 (N_31880,N_28092,N_27929);
xor U31881 (N_31881,N_28605,N_28137);
or U31882 (N_31882,N_27521,N_29422);
nor U31883 (N_31883,N_29950,N_28115);
and U31884 (N_31884,N_27802,N_29774);
or U31885 (N_31885,N_28492,N_28978);
nand U31886 (N_31886,N_27758,N_29400);
nand U31887 (N_31887,N_29963,N_29355);
and U31888 (N_31888,N_29689,N_29645);
or U31889 (N_31889,N_29287,N_27530);
or U31890 (N_31890,N_29287,N_28020);
nand U31891 (N_31891,N_29817,N_28080);
xor U31892 (N_31892,N_28242,N_28992);
nor U31893 (N_31893,N_29450,N_28732);
nand U31894 (N_31894,N_29793,N_29728);
xor U31895 (N_31895,N_28476,N_29620);
nor U31896 (N_31896,N_27722,N_28861);
or U31897 (N_31897,N_28579,N_27676);
nor U31898 (N_31898,N_29270,N_29940);
nand U31899 (N_31899,N_27646,N_29949);
nand U31900 (N_31900,N_28842,N_29773);
or U31901 (N_31901,N_28130,N_29676);
nand U31902 (N_31902,N_28634,N_29413);
and U31903 (N_31903,N_28364,N_28764);
and U31904 (N_31904,N_28153,N_28023);
or U31905 (N_31905,N_29702,N_28152);
or U31906 (N_31906,N_27864,N_28858);
nor U31907 (N_31907,N_28958,N_29595);
nor U31908 (N_31908,N_29741,N_27875);
or U31909 (N_31909,N_28973,N_27847);
and U31910 (N_31910,N_28024,N_28708);
nand U31911 (N_31911,N_28564,N_29932);
or U31912 (N_31912,N_27545,N_28509);
xnor U31913 (N_31913,N_28444,N_27968);
nand U31914 (N_31914,N_29109,N_29779);
and U31915 (N_31915,N_27586,N_29782);
xnor U31916 (N_31916,N_29281,N_29631);
nor U31917 (N_31917,N_27640,N_27585);
nand U31918 (N_31918,N_29483,N_27745);
or U31919 (N_31919,N_28500,N_29378);
xnor U31920 (N_31920,N_28206,N_28438);
nor U31921 (N_31921,N_29120,N_29974);
or U31922 (N_31922,N_29155,N_28118);
or U31923 (N_31923,N_28544,N_28304);
and U31924 (N_31924,N_28794,N_27778);
xor U31925 (N_31925,N_28099,N_28248);
nand U31926 (N_31926,N_29658,N_29553);
nor U31927 (N_31927,N_28812,N_28107);
and U31928 (N_31928,N_27965,N_27692);
and U31929 (N_31929,N_29405,N_29176);
nor U31930 (N_31930,N_29311,N_28706);
nand U31931 (N_31931,N_28674,N_27501);
and U31932 (N_31932,N_29154,N_28893);
or U31933 (N_31933,N_29351,N_29111);
or U31934 (N_31934,N_27958,N_28139);
and U31935 (N_31935,N_28351,N_29876);
nor U31936 (N_31936,N_29673,N_27842);
and U31937 (N_31937,N_28825,N_27784);
nand U31938 (N_31938,N_28285,N_27538);
or U31939 (N_31939,N_28662,N_29730);
xnor U31940 (N_31940,N_27850,N_28212);
nand U31941 (N_31941,N_28737,N_29172);
xor U31942 (N_31942,N_28245,N_28924);
xor U31943 (N_31943,N_28496,N_28822);
xnor U31944 (N_31944,N_27741,N_29406);
xor U31945 (N_31945,N_28079,N_27564);
nor U31946 (N_31946,N_27579,N_29487);
xor U31947 (N_31947,N_29064,N_28984);
and U31948 (N_31948,N_29997,N_28272);
nand U31949 (N_31949,N_29475,N_28889);
and U31950 (N_31950,N_28076,N_28748);
or U31951 (N_31951,N_28445,N_28620);
nand U31952 (N_31952,N_28543,N_27906);
nand U31953 (N_31953,N_29935,N_28770);
nand U31954 (N_31954,N_27962,N_27528);
nor U31955 (N_31955,N_29003,N_28540);
nor U31956 (N_31956,N_29042,N_29536);
nor U31957 (N_31957,N_28976,N_29873);
nand U31958 (N_31958,N_29527,N_28738);
xnor U31959 (N_31959,N_29039,N_28028);
and U31960 (N_31960,N_28426,N_29670);
xnor U31961 (N_31961,N_27847,N_28126);
or U31962 (N_31962,N_29855,N_28105);
and U31963 (N_31963,N_29367,N_28644);
or U31964 (N_31964,N_27786,N_28238);
or U31965 (N_31965,N_28553,N_28781);
or U31966 (N_31966,N_29328,N_28709);
nor U31967 (N_31967,N_28767,N_28855);
and U31968 (N_31968,N_29076,N_29742);
nor U31969 (N_31969,N_28309,N_28962);
and U31970 (N_31970,N_29480,N_28428);
xnor U31971 (N_31971,N_29848,N_27682);
and U31972 (N_31972,N_29293,N_27572);
xor U31973 (N_31973,N_27840,N_29971);
xor U31974 (N_31974,N_27852,N_27812);
nor U31975 (N_31975,N_29352,N_28517);
nor U31976 (N_31976,N_28172,N_28437);
and U31977 (N_31977,N_28844,N_29964);
xnor U31978 (N_31978,N_27537,N_29828);
or U31979 (N_31979,N_27650,N_28118);
xnor U31980 (N_31980,N_29381,N_28189);
and U31981 (N_31981,N_28154,N_28181);
xor U31982 (N_31982,N_28283,N_29990);
nand U31983 (N_31983,N_28685,N_28889);
or U31984 (N_31984,N_28683,N_29081);
xnor U31985 (N_31985,N_27651,N_28772);
nand U31986 (N_31986,N_27720,N_28549);
xor U31987 (N_31987,N_27896,N_28285);
or U31988 (N_31988,N_29769,N_29761);
and U31989 (N_31989,N_29188,N_28970);
nand U31990 (N_31990,N_28580,N_27765);
nand U31991 (N_31991,N_27901,N_29115);
nand U31992 (N_31992,N_29259,N_27886);
nor U31993 (N_31993,N_28527,N_28149);
nor U31994 (N_31994,N_29826,N_27886);
nand U31995 (N_31995,N_29060,N_29275);
and U31996 (N_31996,N_29188,N_29676);
nand U31997 (N_31997,N_27793,N_29433);
nand U31998 (N_31998,N_29421,N_29098);
nor U31999 (N_31999,N_27561,N_28057);
and U32000 (N_32000,N_27849,N_28638);
xnor U32001 (N_32001,N_27913,N_28335);
nand U32002 (N_32002,N_28250,N_29365);
nand U32003 (N_32003,N_28833,N_27546);
nand U32004 (N_32004,N_29353,N_28652);
and U32005 (N_32005,N_29435,N_27591);
and U32006 (N_32006,N_29434,N_29092);
and U32007 (N_32007,N_29767,N_29716);
or U32008 (N_32008,N_28157,N_28992);
xnor U32009 (N_32009,N_29559,N_29635);
and U32010 (N_32010,N_28327,N_28395);
and U32011 (N_32011,N_29849,N_28948);
or U32012 (N_32012,N_28864,N_28942);
nand U32013 (N_32013,N_27820,N_27880);
or U32014 (N_32014,N_29081,N_28016);
xnor U32015 (N_32015,N_29618,N_28574);
nand U32016 (N_32016,N_27701,N_28705);
nor U32017 (N_32017,N_28900,N_28800);
xor U32018 (N_32018,N_28566,N_27630);
xor U32019 (N_32019,N_28364,N_29951);
xnor U32020 (N_32020,N_29209,N_29940);
xnor U32021 (N_32021,N_28946,N_27896);
nand U32022 (N_32022,N_27790,N_29479);
nor U32023 (N_32023,N_29397,N_27662);
nor U32024 (N_32024,N_29190,N_28436);
or U32025 (N_32025,N_27568,N_28480);
nand U32026 (N_32026,N_29110,N_28990);
and U32027 (N_32027,N_27799,N_28646);
xnor U32028 (N_32028,N_27771,N_27781);
nand U32029 (N_32029,N_29596,N_29969);
or U32030 (N_32030,N_28675,N_28780);
nor U32031 (N_32031,N_28815,N_28776);
nor U32032 (N_32032,N_29252,N_27567);
nor U32033 (N_32033,N_29873,N_28496);
nor U32034 (N_32034,N_29222,N_28470);
xnor U32035 (N_32035,N_27983,N_28881);
or U32036 (N_32036,N_28494,N_27567);
and U32037 (N_32037,N_29568,N_29561);
and U32038 (N_32038,N_27914,N_28325);
nand U32039 (N_32039,N_29393,N_29706);
nand U32040 (N_32040,N_28429,N_29188);
and U32041 (N_32041,N_29870,N_27677);
nor U32042 (N_32042,N_29715,N_28710);
and U32043 (N_32043,N_28521,N_28199);
and U32044 (N_32044,N_28611,N_28517);
or U32045 (N_32045,N_27550,N_27528);
and U32046 (N_32046,N_27638,N_29204);
or U32047 (N_32047,N_28116,N_28918);
or U32048 (N_32048,N_29378,N_29861);
nor U32049 (N_32049,N_29182,N_28602);
xor U32050 (N_32050,N_27718,N_29177);
xnor U32051 (N_32051,N_28010,N_28742);
and U32052 (N_32052,N_28215,N_27723);
xnor U32053 (N_32053,N_28656,N_28052);
nand U32054 (N_32054,N_29323,N_29683);
xnor U32055 (N_32055,N_29080,N_28809);
nand U32056 (N_32056,N_29272,N_27605);
and U32057 (N_32057,N_27726,N_29706);
or U32058 (N_32058,N_29645,N_28899);
xnor U32059 (N_32059,N_29175,N_27960);
xnor U32060 (N_32060,N_27988,N_29362);
nor U32061 (N_32061,N_29791,N_27807);
or U32062 (N_32062,N_29686,N_28659);
xor U32063 (N_32063,N_29632,N_29044);
xnor U32064 (N_32064,N_29149,N_28785);
and U32065 (N_32065,N_29210,N_29994);
nand U32066 (N_32066,N_28726,N_28534);
nor U32067 (N_32067,N_27897,N_29609);
and U32068 (N_32068,N_27773,N_29889);
or U32069 (N_32069,N_27741,N_28602);
nor U32070 (N_32070,N_29991,N_28908);
and U32071 (N_32071,N_28214,N_28293);
nor U32072 (N_32072,N_27683,N_28811);
nor U32073 (N_32073,N_28052,N_27822);
nor U32074 (N_32074,N_29482,N_27978);
or U32075 (N_32075,N_28606,N_29792);
or U32076 (N_32076,N_29305,N_29744);
or U32077 (N_32077,N_28324,N_27997);
nand U32078 (N_32078,N_29501,N_29180);
or U32079 (N_32079,N_28519,N_29560);
and U32080 (N_32080,N_29859,N_28866);
nor U32081 (N_32081,N_28849,N_28341);
or U32082 (N_32082,N_27770,N_28537);
nor U32083 (N_32083,N_27857,N_28831);
and U32084 (N_32084,N_29083,N_29088);
and U32085 (N_32085,N_29841,N_29648);
and U32086 (N_32086,N_29439,N_27957);
xnor U32087 (N_32087,N_29111,N_28581);
or U32088 (N_32088,N_27926,N_28667);
nor U32089 (N_32089,N_28464,N_28101);
or U32090 (N_32090,N_28079,N_28926);
nand U32091 (N_32091,N_29378,N_29364);
nor U32092 (N_32092,N_28038,N_28851);
xnor U32093 (N_32093,N_28896,N_28880);
xor U32094 (N_32094,N_28632,N_27835);
or U32095 (N_32095,N_27773,N_29188);
xnor U32096 (N_32096,N_29499,N_29671);
xnor U32097 (N_32097,N_28307,N_28459);
nor U32098 (N_32098,N_28549,N_29257);
nor U32099 (N_32099,N_28612,N_29075);
and U32100 (N_32100,N_28965,N_28589);
nor U32101 (N_32101,N_28190,N_29260);
nor U32102 (N_32102,N_29386,N_28501);
and U32103 (N_32103,N_27581,N_27804);
or U32104 (N_32104,N_28313,N_29678);
nand U32105 (N_32105,N_29667,N_28367);
nand U32106 (N_32106,N_28812,N_29255);
nor U32107 (N_32107,N_28965,N_28849);
nand U32108 (N_32108,N_29491,N_29325);
or U32109 (N_32109,N_29580,N_29902);
xor U32110 (N_32110,N_28564,N_29504);
nor U32111 (N_32111,N_28967,N_29261);
nor U32112 (N_32112,N_28933,N_29704);
xor U32113 (N_32113,N_27760,N_29768);
nor U32114 (N_32114,N_29525,N_29740);
or U32115 (N_32115,N_29574,N_29591);
nand U32116 (N_32116,N_29635,N_27902);
xor U32117 (N_32117,N_29473,N_28378);
xnor U32118 (N_32118,N_29913,N_28292);
nand U32119 (N_32119,N_29391,N_29138);
xnor U32120 (N_32120,N_29837,N_28773);
nor U32121 (N_32121,N_27804,N_27692);
xor U32122 (N_32122,N_29331,N_28438);
nor U32123 (N_32123,N_28116,N_28305);
nor U32124 (N_32124,N_28093,N_28889);
and U32125 (N_32125,N_29592,N_29966);
nand U32126 (N_32126,N_28749,N_28759);
or U32127 (N_32127,N_29987,N_28388);
xnor U32128 (N_32128,N_29367,N_27619);
xnor U32129 (N_32129,N_27844,N_27904);
and U32130 (N_32130,N_29090,N_28557);
nand U32131 (N_32131,N_27875,N_28638);
nand U32132 (N_32132,N_28913,N_28564);
nor U32133 (N_32133,N_28458,N_29974);
nor U32134 (N_32134,N_28965,N_28765);
or U32135 (N_32135,N_29930,N_28850);
nand U32136 (N_32136,N_27879,N_29866);
nand U32137 (N_32137,N_28734,N_28574);
and U32138 (N_32138,N_29991,N_28109);
xor U32139 (N_32139,N_27791,N_28407);
or U32140 (N_32140,N_27674,N_28501);
nor U32141 (N_32141,N_28459,N_28425);
nor U32142 (N_32142,N_27692,N_29267);
and U32143 (N_32143,N_28612,N_29659);
nand U32144 (N_32144,N_29101,N_29398);
xnor U32145 (N_32145,N_28188,N_29409);
or U32146 (N_32146,N_28742,N_29093);
and U32147 (N_32147,N_29445,N_28214);
and U32148 (N_32148,N_29835,N_27945);
and U32149 (N_32149,N_27647,N_28769);
nand U32150 (N_32150,N_29199,N_28144);
and U32151 (N_32151,N_29231,N_29188);
or U32152 (N_32152,N_27735,N_28502);
nand U32153 (N_32153,N_27714,N_29997);
nor U32154 (N_32154,N_28653,N_27769);
xor U32155 (N_32155,N_28061,N_29820);
xnor U32156 (N_32156,N_27768,N_28173);
and U32157 (N_32157,N_29240,N_28579);
or U32158 (N_32158,N_27595,N_28949);
xnor U32159 (N_32159,N_28102,N_29773);
xnor U32160 (N_32160,N_29626,N_28362);
xor U32161 (N_32161,N_28392,N_28859);
nor U32162 (N_32162,N_27657,N_27841);
nand U32163 (N_32163,N_29051,N_28761);
or U32164 (N_32164,N_28098,N_28479);
nand U32165 (N_32165,N_28603,N_29787);
nand U32166 (N_32166,N_28023,N_28006);
nand U32167 (N_32167,N_29852,N_28413);
nand U32168 (N_32168,N_28039,N_29996);
or U32169 (N_32169,N_29463,N_29843);
and U32170 (N_32170,N_29597,N_27815);
nor U32171 (N_32171,N_27534,N_28336);
or U32172 (N_32172,N_28980,N_27808);
and U32173 (N_32173,N_29015,N_28415);
nand U32174 (N_32174,N_29694,N_29689);
or U32175 (N_32175,N_28591,N_29446);
xnor U32176 (N_32176,N_28689,N_29273);
xor U32177 (N_32177,N_28983,N_28873);
and U32178 (N_32178,N_27784,N_28859);
nor U32179 (N_32179,N_28340,N_28164);
nand U32180 (N_32180,N_27526,N_28409);
or U32181 (N_32181,N_29085,N_28027);
or U32182 (N_32182,N_28338,N_28065);
nor U32183 (N_32183,N_28786,N_29958);
nor U32184 (N_32184,N_28750,N_28048);
and U32185 (N_32185,N_28075,N_28105);
xnor U32186 (N_32186,N_27559,N_29909);
or U32187 (N_32187,N_29053,N_28882);
and U32188 (N_32188,N_27521,N_29652);
nor U32189 (N_32189,N_28685,N_28785);
or U32190 (N_32190,N_28848,N_29341);
and U32191 (N_32191,N_27684,N_28022);
or U32192 (N_32192,N_29165,N_29146);
and U32193 (N_32193,N_28726,N_29592);
xor U32194 (N_32194,N_28214,N_29028);
nor U32195 (N_32195,N_28444,N_29553);
or U32196 (N_32196,N_28714,N_27848);
or U32197 (N_32197,N_29761,N_29349);
and U32198 (N_32198,N_27836,N_28301);
nand U32199 (N_32199,N_29057,N_28251);
xor U32200 (N_32200,N_28280,N_28538);
nor U32201 (N_32201,N_28742,N_28845);
and U32202 (N_32202,N_29779,N_29947);
nand U32203 (N_32203,N_28603,N_27553);
nor U32204 (N_32204,N_29249,N_27869);
xor U32205 (N_32205,N_27513,N_28303);
nand U32206 (N_32206,N_29642,N_27938);
nand U32207 (N_32207,N_28981,N_28283);
nor U32208 (N_32208,N_28097,N_28409);
nor U32209 (N_32209,N_27559,N_27983);
or U32210 (N_32210,N_27732,N_28522);
nor U32211 (N_32211,N_27989,N_29935);
xor U32212 (N_32212,N_28752,N_28753);
and U32213 (N_32213,N_27714,N_28681);
xor U32214 (N_32214,N_28280,N_29412);
xnor U32215 (N_32215,N_29141,N_28914);
and U32216 (N_32216,N_27688,N_29882);
nor U32217 (N_32217,N_29582,N_29558);
nor U32218 (N_32218,N_29336,N_28807);
nor U32219 (N_32219,N_28049,N_27527);
xnor U32220 (N_32220,N_29936,N_28406);
nand U32221 (N_32221,N_29603,N_27872);
or U32222 (N_32222,N_28860,N_29207);
and U32223 (N_32223,N_27557,N_29602);
nand U32224 (N_32224,N_28116,N_28012);
or U32225 (N_32225,N_27883,N_29277);
and U32226 (N_32226,N_28230,N_29695);
xor U32227 (N_32227,N_28203,N_29851);
nor U32228 (N_32228,N_28057,N_29880);
and U32229 (N_32229,N_29943,N_29064);
xor U32230 (N_32230,N_28773,N_28221);
nor U32231 (N_32231,N_29218,N_28901);
nor U32232 (N_32232,N_27627,N_28468);
or U32233 (N_32233,N_29030,N_28936);
or U32234 (N_32234,N_29300,N_28951);
or U32235 (N_32235,N_27702,N_29939);
nor U32236 (N_32236,N_28751,N_29289);
or U32237 (N_32237,N_28107,N_29692);
and U32238 (N_32238,N_29694,N_28808);
nand U32239 (N_32239,N_29698,N_29160);
xnor U32240 (N_32240,N_29076,N_29302);
and U32241 (N_32241,N_29376,N_27885);
or U32242 (N_32242,N_28488,N_29296);
or U32243 (N_32243,N_28614,N_29442);
and U32244 (N_32244,N_29937,N_27838);
nand U32245 (N_32245,N_28122,N_28528);
nor U32246 (N_32246,N_28193,N_28759);
nand U32247 (N_32247,N_27840,N_27624);
or U32248 (N_32248,N_29907,N_29855);
xnor U32249 (N_32249,N_27557,N_29354);
nor U32250 (N_32250,N_28842,N_28333);
and U32251 (N_32251,N_27699,N_28352);
or U32252 (N_32252,N_29155,N_29257);
nand U32253 (N_32253,N_27717,N_28888);
and U32254 (N_32254,N_29649,N_29816);
or U32255 (N_32255,N_27708,N_29635);
xor U32256 (N_32256,N_27578,N_27620);
nand U32257 (N_32257,N_28011,N_27608);
and U32258 (N_32258,N_28043,N_28959);
xnor U32259 (N_32259,N_27796,N_28761);
xnor U32260 (N_32260,N_29316,N_27684);
nor U32261 (N_32261,N_28101,N_28376);
or U32262 (N_32262,N_29618,N_29320);
and U32263 (N_32263,N_27510,N_28043);
nor U32264 (N_32264,N_27527,N_27975);
nor U32265 (N_32265,N_28372,N_28946);
xor U32266 (N_32266,N_28277,N_29305);
or U32267 (N_32267,N_28988,N_28065);
xor U32268 (N_32268,N_27871,N_27630);
nand U32269 (N_32269,N_29001,N_28570);
nand U32270 (N_32270,N_29778,N_27517);
xnor U32271 (N_32271,N_28743,N_28600);
or U32272 (N_32272,N_27708,N_28806);
or U32273 (N_32273,N_28033,N_28371);
or U32274 (N_32274,N_28591,N_27891);
or U32275 (N_32275,N_27747,N_27684);
nor U32276 (N_32276,N_29705,N_28693);
nor U32277 (N_32277,N_28658,N_28692);
or U32278 (N_32278,N_27702,N_29116);
or U32279 (N_32279,N_27848,N_27979);
xor U32280 (N_32280,N_28047,N_29821);
or U32281 (N_32281,N_27936,N_29144);
or U32282 (N_32282,N_27961,N_28607);
nand U32283 (N_32283,N_29674,N_28554);
and U32284 (N_32284,N_29202,N_27624);
and U32285 (N_32285,N_29226,N_29218);
or U32286 (N_32286,N_27936,N_27901);
and U32287 (N_32287,N_29830,N_29871);
and U32288 (N_32288,N_28158,N_29849);
or U32289 (N_32289,N_27624,N_27525);
nand U32290 (N_32290,N_27615,N_28411);
xor U32291 (N_32291,N_29780,N_28745);
nor U32292 (N_32292,N_27793,N_29693);
nor U32293 (N_32293,N_27898,N_29091);
or U32294 (N_32294,N_29729,N_28449);
nor U32295 (N_32295,N_28753,N_29241);
xor U32296 (N_32296,N_29271,N_27565);
xor U32297 (N_32297,N_28234,N_29019);
xor U32298 (N_32298,N_29766,N_28183);
nor U32299 (N_32299,N_28801,N_29539);
nor U32300 (N_32300,N_29450,N_29144);
nand U32301 (N_32301,N_28897,N_29075);
nor U32302 (N_32302,N_28532,N_28692);
xnor U32303 (N_32303,N_27989,N_28477);
xnor U32304 (N_32304,N_28574,N_28025);
nand U32305 (N_32305,N_28765,N_29353);
or U32306 (N_32306,N_28458,N_28449);
xor U32307 (N_32307,N_29363,N_28767);
xnor U32308 (N_32308,N_27876,N_29034);
or U32309 (N_32309,N_29539,N_29769);
or U32310 (N_32310,N_29233,N_28899);
and U32311 (N_32311,N_28869,N_27990);
nor U32312 (N_32312,N_28778,N_29888);
nand U32313 (N_32313,N_27868,N_27523);
nor U32314 (N_32314,N_29339,N_27700);
xnor U32315 (N_32315,N_29313,N_27766);
nor U32316 (N_32316,N_28016,N_29008);
nand U32317 (N_32317,N_28819,N_28230);
or U32318 (N_32318,N_29494,N_27799);
nor U32319 (N_32319,N_28383,N_29788);
and U32320 (N_32320,N_29607,N_28165);
nand U32321 (N_32321,N_29117,N_27988);
xnor U32322 (N_32322,N_28339,N_27980);
or U32323 (N_32323,N_27970,N_28064);
and U32324 (N_32324,N_28672,N_29428);
or U32325 (N_32325,N_28218,N_27880);
xnor U32326 (N_32326,N_29031,N_28224);
xor U32327 (N_32327,N_29760,N_28344);
or U32328 (N_32328,N_27662,N_28350);
nand U32329 (N_32329,N_27725,N_29821);
or U32330 (N_32330,N_29967,N_28756);
nand U32331 (N_32331,N_28148,N_29607);
nor U32332 (N_32332,N_28744,N_29236);
nor U32333 (N_32333,N_28601,N_27879);
and U32334 (N_32334,N_28251,N_29322);
or U32335 (N_32335,N_28400,N_29009);
and U32336 (N_32336,N_28732,N_28254);
nor U32337 (N_32337,N_28555,N_27884);
xnor U32338 (N_32338,N_27660,N_28749);
nor U32339 (N_32339,N_29242,N_28291);
xor U32340 (N_32340,N_28558,N_28486);
and U32341 (N_32341,N_28908,N_28531);
or U32342 (N_32342,N_29212,N_28793);
nor U32343 (N_32343,N_28150,N_29727);
nor U32344 (N_32344,N_29325,N_29481);
or U32345 (N_32345,N_28022,N_29926);
nor U32346 (N_32346,N_29033,N_28132);
xnor U32347 (N_32347,N_29051,N_27662);
or U32348 (N_32348,N_29642,N_28395);
and U32349 (N_32349,N_29427,N_29887);
and U32350 (N_32350,N_29248,N_28929);
xor U32351 (N_32351,N_27536,N_28424);
and U32352 (N_32352,N_28644,N_29175);
nand U32353 (N_32353,N_28060,N_27620);
or U32354 (N_32354,N_28932,N_29389);
nand U32355 (N_32355,N_27605,N_28440);
xnor U32356 (N_32356,N_28437,N_29694);
or U32357 (N_32357,N_27691,N_29070);
xor U32358 (N_32358,N_28521,N_28182);
nand U32359 (N_32359,N_28260,N_27730);
and U32360 (N_32360,N_28402,N_28880);
nor U32361 (N_32361,N_29771,N_28454);
nor U32362 (N_32362,N_29990,N_27748);
and U32363 (N_32363,N_29800,N_28965);
xnor U32364 (N_32364,N_28835,N_29566);
nor U32365 (N_32365,N_28851,N_29741);
nand U32366 (N_32366,N_29198,N_27813);
nand U32367 (N_32367,N_28271,N_29682);
nand U32368 (N_32368,N_29927,N_28815);
xor U32369 (N_32369,N_29511,N_29434);
or U32370 (N_32370,N_29673,N_27699);
nand U32371 (N_32371,N_29318,N_29126);
or U32372 (N_32372,N_28710,N_28006);
and U32373 (N_32373,N_28545,N_27993);
nor U32374 (N_32374,N_28724,N_29927);
nor U32375 (N_32375,N_28752,N_29083);
and U32376 (N_32376,N_29093,N_28060);
xnor U32377 (N_32377,N_28097,N_28400);
nand U32378 (N_32378,N_27998,N_27864);
or U32379 (N_32379,N_28488,N_28585);
and U32380 (N_32380,N_29915,N_27913);
nand U32381 (N_32381,N_29649,N_28866);
and U32382 (N_32382,N_29760,N_27536);
or U32383 (N_32383,N_29830,N_29187);
and U32384 (N_32384,N_28169,N_29308);
nor U32385 (N_32385,N_28565,N_29282);
or U32386 (N_32386,N_28638,N_29275);
nand U32387 (N_32387,N_29678,N_29536);
xnor U32388 (N_32388,N_27864,N_29788);
nor U32389 (N_32389,N_29686,N_28733);
and U32390 (N_32390,N_28781,N_28494);
xor U32391 (N_32391,N_29511,N_27681);
and U32392 (N_32392,N_28582,N_28490);
nor U32393 (N_32393,N_27839,N_29518);
nand U32394 (N_32394,N_28720,N_27585);
nor U32395 (N_32395,N_27832,N_28386);
xor U32396 (N_32396,N_28890,N_29412);
xnor U32397 (N_32397,N_28302,N_27548);
nand U32398 (N_32398,N_28021,N_27681);
and U32399 (N_32399,N_29629,N_29011);
or U32400 (N_32400,N_29038,N_29779);
nor U32401 (N_32401,N_27908,N_29433);
xor U32402 (N_32402,N_28722,N_28165);
and U32403 (N_32403,N_29395,N_29207);
or U32404 (N_32404,N_29717,N_28364);
or U32405 (N_32405,N_28251,N_28151);
or U32406 (N_32406,N_29939,N_28996);
xnor U32407 (N_32407,N_29535,N_29732);
xor U32408 (N_32408,N_28426,N_28937);
xnor U32409 (N_32409,N_28831,N_28020);
or U32410 (N_32410,N_29742,N_28919);
xnor U32411 (N_32411,N_29121,N_28669);
or U32412 (N_32412,N_28373,N_29355);
or U32413 (N_32413,N_28836,N_29085);
and U32414 (N_32414,N_29062,N_28854);
and U32415 (N_32415,N_28330,N_28534);
and U32416 (N_32416,N_29758,N_28777);
and U32417 (N_32417,N_29495,N_29120);
xor U32418 (N_32418,N_27568,N_29091);
nor U32419 (N_32419,N_27841,N_28833);
or U32420 (N_32420,N_29478,N_28892);
xor U32421 (N_32421,N_28706,N_28415);
and U32422 (N_32422,N_28320,N_27574);
nand U32423 (N_32423,N_29432,N_28208);
nor U32424 (N_32424,N_28275,N_29129);
nand U32425 (N_32425,N_29307,N_28447);
and U32426 (N_32426,N_27753,N_28563);
or U32427 (N_32427,N_28313,N_29677);
nand U32428 (N_32428,N_29764,N_27534);
and U32429 (N_32429,N_27655,N_28153);
or U32430 (N_32430,N_28770,N_28447);
or U32431 (N_32431,N_28862,N_27914);
xnor U32432 (N_32432,N_29737,N_27998);
nand U32433 (N_32433,N_29508,N_29947);
or U32434 (N_32434,N_28442,N_29208);
nand U32435 (N_32435,N_29734,N_29248);
xor U32436 (N_32436,N_28218,N_28669);
xor U32437 (N_32437,N_27844,N_28751);
nor U32438 (N_32438,N_29921,N_28418);
or U32439 (N_32439,N_27842,N_29555);
or U32440 (N_32440,N_29916,N_28111);
or U32441 (N_32441,N_29777,N_29593);
nor U32442 (N_32442,N_28842,N_28996);
xor U32443 (N_32443,N_29618,N_28805);
or U32444 (N_32444,N_28345,N_29329);
or U32445 (N_32445,N_28795,N_29537);
nand U32446 (N_32446,N_29344,N_27876);
and U32447 (N_32447,N_28004,N_28366);
or U32448 (N_32448,N_29323,N_27611);
or U32449 (N_32449,N_28217,N_27984);
xor U32450 (N_32450,N_28144,N_28384);
nor U32451 (N_32451,N_28893,N_28627);
xor U32452 (N_32452,N_28397,N_27977);
xor U32453 (N_32453,N_28437,N_29978);
xor U32454 (N_32454,N_27996,N_29856);
nor U32455 (N_32455,N_29044,N_28585);
or U32456 (N_32456,N_29519,N_27636);
nor U32457 (N_32457,N_28757,N_28943);
xnor U32458 (N_32458,N_28860,N_28976);
nand U32459 (N_32459,N_28781,N_28770);
nor U32460 (N_32460,N_28237,N_29097);
xnor U32461 (N_32461,N_28309,N_28269);
or U32462 (N_32462,N_29823,N_28179);
or U32463 (N_32463,N_28717,N_28890);
or U32464 (N_32464,N_27601,N_28154);
or U32465 (N_32465,N_28701,N_27717);
and U32466 (N_32466,N_28886,N_29064);
or U32467 (N_32467,N_28840,N_29395);
nand U32468 (N_32468,N_28394,N_29165);
nand U32469 (N_32469,N_29760,N_27895);
nor U32470 (N_32470,N_29882,N_29942);
or U32471 (N_32471,N_29096,N_29154);
xnor U32472 (N_32472,N_29382,N_28538);
and U32473 (N_32473,N_28482,N_29434);
or U32474 (N_32474,N_29127,N_28439);
xor U32475 (N_32475,N_29912,N_29934);
or U32476 (N_32476,N_28419,N_29826);
xor U32477 (N_32477,N_28027,N_27805);
nor U32478 (N_32478,N_28279,N_27683);
nand U32479 (N_32479,N_28404,N_27564);
or U32480 (N_32480,N_29251,N_29370);
or U32481 (N_32481,N_28347,N_28204);
nand U32482 (N_32482,N_29790,N_27705);
nand U32483 (N_32483,N_29153,N_28744);
nand U32484 (N_32484,N_27849,N_29236);
nor U32485 (N_32485,N_29764,N_28386);
and U32486 (N_32486,N_28662,N_29036);
or U32487 (N_32487,N_28015,N_28777);
nand U32488 (N_32488,N_29875,N_28625);
and U32489 (N_32489,N_28022,N_28598);
or U32490 (N_32490,N_28583,N_28025);
and U32491 (N_32491,N_28236,N_29931);
nand U32492 (N_32492,N_28068,N_28547);
xnor U32493 (N_32493,N_28510,N_27865);
or U32494 (N_32494,N_27780,N_29299);
or U32495 (N_32495,N_28460,N_28834);
xnor U32496 (N_32496,N_29584,N_27703);
nand U32497 (N_32497,N_27839,N_29205);
xnor U32498 (N_32498,N_27867,N_29725);
nor U32499 (N_32499,N_29010,N_29705);
or U32500 (N_32500,N_30918,N_31193);
and U32501 (N_32501,N_31990,N_32210);
or U32502 (N_32502,N_30877,N_32032);
and U32503 (N_32503,N_31330,N_30171);
or U32504 (N_32504,N_30035,N_32288);
or U32505 (N_32505,N_32265,N_31737);
nand U32506 (N_32506,N_30036,N_30747);
or U32507 (N_32507,N_31404,N_32191);
or U32508 (N_32508,N_32342,N_30486);
xnor U32509 (N_32509,N_31270,N_32377);
or U32510 (N_32510,N_31118,N_31750);
xnor U32511 (N_32511,N_31918,N_30619);
xor U32512 (N_32512,N_30915,N_30765);
xnor U32513 (N_32513,N_32408,N_31805);
and U32514 (N_32514,N_30124,N_31933);
xor U32515 (N_32515,N_31054,N_32156);
and U32516 (N_32516,N_31275,N_30611);
xnor U32517 (N_32517,N_31907,N_30851);
or U32518 (N_32518,N_32130,N_31149);
nand U32519 (N_32519,N_30345,N_31224);
and U32520 (N_32520,N_32178,N_31728);
xnor U32521 (N_32521,N_32325,N_32347);
and U32522 (N_32522,N_31354,N_31426);
nor U32523 (N_32523,N_30504,N_32078);
xnor U32524 (N_32524,N_30593,N_32431);
nand U32525 (N_32525,N_32261,N_31154);
nand U32526 (N_32526,N_32491,N_30587);
xnor U32527 (N_32527,N_30043,N_32297);
nand U32528 (N_32528,N_31243,N_30474);
nor U32529 (N_32529,N_32275,N_30317);
nand U32530 (N_32530,N_31019,N_32081);
and U32531 (N_32531,N_30320,N_32382);
or U32532 (N_32532,N_32292,N_31669);
nor U32533 (N_32533,N_31761,N_31518);
xnor U32534 (N_32534,N_30255,N_31186);
and U32535 (N_32535,N_30245,N_31626);
nor U32536 (N_32536,N_32317,N_30689);
and U32537 (N_32537,N_31047,N_32184);
nand U32538 (N_32538,N_31147,N_31748);
nor U32539 (N_32539,N_31241,N_31771);
nor U32540 (N_32540,N_32225,N_30104);
nand U32541 (N_32541,N_30189,N_30408);
or U32542 (N_32542,N_30353,N_32103);
nand U32543 (N_32543,N_31423,N_32387);
xnor U32544 (N_32544,N_31809,N_30943);
and U32545 (N_32545,N_31797,N_30973);
or U32546 (N_32546,N_30053,N_32234);
xnor U32547 (N_32547,N_31712,N_31845);
or U32548 (N_32548,N_30605,N_30076);
nand U32549 (N_32549,N_31714,N_30759);
nor U32550 (N_32550,N_30884,N_30718);
xor U32551 (N_32551,N_31636,N_31026);
nand U32552 (N_32552,N_31995,N_30283);
nand U32553 (N_32553,N_31848,N_30061);
xnor U32554 (N_32554,N_30694,N_30733);
or U32555 (N_32555,N_30792,N_30110);
or U32556 (N_32556,N_31098,N_30978);
and U32557 (N_32557,N_31260,N_31914);
xor U32558 (N_32558,N_31938,N_32131);
and U32559 (N_32559,N_30829,N_32009);
nor U32560 (N_32560,N_31841,N_31081);
or U32561 (N_32561,N_30824,N_31606);
nand U32562 (N_32562,N_30433,N_31656);
or U32563 (N_32563,N_32162,N_30365);
nor U32564 (N_32564,N_30821,N_31050);
and U32565 (N_32565,N_32366,N_31581);
or U32566 (N_32566,N_32049,N_30585);
nand U32567 (N_32567,N_32036,N_30022);
xnor U32568 (N_32568,N_30805,N_32085);
xnor U32569 (N_32569,N_30284,N_31795);
nand U32570 (N_32570,N_32395,N_31344);
xnor U32571 (N_32571,N_31202,N_30517);
nand U32572 (N_32572,N_30996,N_30967);
nand U32573 (N_32573,N_32152,N_31568);
nand U32574 (N_32574,N_31265,N_31483);
or U32575 (N_32575,N_31480,N_30767);
xnor U32576 (N_32576,N_31802,N_31171);
nor U32577 (N_32577,N_31791,N_30193);
nor U32578 (N_32578,N_32199,N_31025);
and U32579 (N_32579,N_30367,N_31548);
xor U32580 (N_32580,N_31706,N_31557);
and U32581 (N_32581,N_31371,N_32330);
nor U32582 (N_32582,N_31271,N_32179);
or U32583 (N_32583,N_31119,N_31095);
xor U32584 (N_32584,N_30502,N_30001);
nor U32585 (N_32585,N_30722,N_30222);
and U32586 (N_32586,N_32138,N_31390);
nor U32587 (N_32587,N_31309,N_32010);
nand U32588 (N_32588,N_31200,N_30966);
or U32589 (N_32589,N_32003,N_31168);
nand U32590 (N_32590,N_30914,N_30087);
nor U32591 (N_32591,N_30233,N_31691);
or U32592 (N_32592,N_32177,N_30908);
nor U32593 (N_32593,N_31259,N_31897);
nor U32594 (N_32594,N_32285,N_30420);
and U32595 (N_32595,N_32096,N_30258);
xnor U32596 (N_32596,N_30019,N_32211);
nand U32597 (N_32597,N_31664,N_32422);
nor U32598 (N_32598,N_30912,N_32467);
xnor U32599 (N_32599,N_31041,N_31704);
or U32600 (N_32600,N_30993,N_31400);
nor U32601 (N_32601,N_32104,N_30359);
xnor U32602 (N_32602,N_30146,N_31744);
and U32603 (N_32603,N_30923,N_31043);
or U32604 (N_32604,N_30772,N_31741);
and U32605 (N_32605,N_30190,N_32237);
and U32606 (N_32606,N_30134,N_31492);
nand U32607 (N_32607,N_30095,N_30447);
or U32608 (N_32608,N_32042,N_31916);
or U32609 (N_32609,N_30793,N_31343);
or U32610 (N_32610,N_31657,N_31756);
or U32611 (N_32611,N_32429,N_30819);
nor U32612 (N_32612,N_31208,N_31128);
nand U32613 (N_32613,N_30436,N_32338);
and U32614 (N_32614,N_30114,N_31954);
nor U32615 (N_32615,N_31236,N_30266);
nand U32616 (N_32616,N_31864,N_32067);
or U32617 (N_32617,N_31263,N_31974);
and U32618 (N_32618,N_32164,N_32361);
nand U32619 (N_32619,N_30898,N_32132);
nand U32620 (N_32620,N_30665,N_30054);
nor U32621 (N_32621,N_31770,N_31121);
nand U32622 (N_32622,N_30147,N_32017);
nand U32623 (N_32623,N_32129,N_30542);
or U32624 (N_32624,N_31865,N_31768);
and U32625 (N_32625,N_31803,N_31520);
and U32626 (N_32626,N_31951,N_32443);
or U32627 (N_32627,N_30835,N_30469);
or U32628 (N_32628,N_30964,N_31655);
nor U32629 (N_32629,N_32093,N_30904);
nand U32630 (N_32630,N_30512,N_32231);
nand U32631 (N_32631,N_31227,N_30487);
nand U32632 (N_32632,N_30895,N_31646);
nor U32633 (N_32633,N_31509,N_31488);
and U32634 (N_32634,N_31088,N_31724);
nor U32635 (N_32635,N_31798,N_32306);
nor U32636 (N_32636,N_32163,N_32428);
xor U32637 (N_32637,N_31485,N_32416);
or U32638 (N_32638,N_31563,N_30600);
or U32639 (N_32639,N_31240,N_32002);
nand U32640 (N_32640,N_30327,N_30228);
nor U32641 (N_32641,N_30157,N_31535);
nand U32642 (N_32642,N_32380,N_31014);
nand U32643 (N_32643,N_31576,N_30968);
or U32644 (N_32644,N_31837,N_31647);
or U32645 (N_32645,N_31829,N_30290);
nor U32646 (N_32646,N_30787,N_30720);
nand U32647 (N_32647,N_30012,N_31002);
xor U32648 (N_32648,N_30021,N_30702);
and U32649 (N_32649,N_31217,N_32397);
xor U32650 (N_32650,N_30782,N_30874);
nand U32651 (N_32651,N_32449,N_30913);
and U32652 (N_32652,N_31583,N_32180);
nand U32653 (N_32653,N_31876,N_30807);
and U32654 (N_32654,N_31759,N_30618);
nand U32655 (N_32655,N_30267,N_30868);
nor U32656 (N_32656,N_30601,N_31367);
xor U32657 (N_32657,N_32300,N_30238);
or U32658 (N_32658,N_32436,N_30778);
nand U32659 (N_32659,N_30341,N_30195);
nand U32660 (N_32660,N_31462,N_30540);
and U32661 (N_32661,N_30232,N_30595);
nand U32662 (N_32662,N_32186,N_30306);
xor U32663 (N_32663,N_31676,N_31327);
and U32664 (N_32664,N_31928,N_31064);
and U32665 (N_32665,N_30674,N_32358);
or U32666 (N_32666,N_31130,N_31823);
or U32667 (N_32667,N_31613,N_32020);
and U32668 (N_32668,N_30647,N_32398);
nor U32669 (N_32669,N_31955,N_30869);
or U32670 (N_32670,N_30501,N_32057);
nand U32671 (N_32671,N_32469,N_30634);
and U32672 (N_32672,N_32173,N_31325);
and U32673 (N_32673,N_31783,N_30450);
nand U32674 (N_32674,N_31678,N_30745);
nand U32675 (N_32675,N_31286,N_31383);
nand U32676 (N_32676,N_31328,N_32215);
xor U32677 (N_32677,N_31507,N_30208);
or U32678 (N_32678,N_32025,N_30183);
nand U32679 (N_32679,N_30957,N_30773);
or U32680 (N_32680,N_32301,N_30123);
xor U32681 (N_32681,N_31686,N_31475);
and U32682 (N_32682,N_31040,N_30607);
and U32683 (N_32683,N_31612,N_30198);
or U32684 (N_32684,N_32483,N_31818);
nor U32685 (N_32685,N_30264,N_32492);
xor U32686 (N_32686,N_31570,N_30920);
xor U32687 (N_32687,N_30201,N_32364);
nor U32688 (N_32688,N_30276,N_32474);
nand U32689 (N_32689,N_30513,N_32456);
nor U32690 (N_32690,N_30555,N_31450);
nor U32691 (N_32691,N_30399,N_30421);
nor U32692 (N_32692,N_30567,N_32294);
nor U32693 (N_32693,N_31196,N_31902);
xor U32694 (N_32694,N_31245,N_32247);
xnor U32695 (N_32695,N_30280,N_32465);
xnor U32696 (N_32696,N_31824,N_30308);
xor U32697 (N_32697,N_31873,N_30786);
nand U32698 (N_32698,N_31554,N_30620);
xor U32699 (N_32699,N_30314,N_31778);
nor U32700 (N_32700,N_32050,N_30435);
or U32701 (N_32701,N_31695,N_31861);
xnor U32702 (N_32702,N_31934,N_30931);
and U32703 (N_32703,N_31151,N_31156);
or U32704 (N_32704,N_31888,N_31197);
or U32705 (N_32705,N_31464,N_31775);
or U32706 (N_32706,N_31977,N_32043);
xor U32707 (N_32707,N_30818,N_32426);
or U32708 (N_32708,N_31209,N_30960);
xor U32709 (N_32709,N_30710,N_31603);
xor U32710 (N_32710,N_30571,N_31044);
xor U32711 (N_32711,N_32222,N_30641);
xor U32712 (N_32712,N_32457,N_30573);
nand U32713 (N_32713,N_30128,N_31523);
nand U32714 (N_32714,N_30418,N_31587);
nor U32715 (N_32715,N_32367,N_31436);
or U32716 (N_32716,N_32249,N_32430);
or U32717 (N_32717,N_30795,N_30669);
and U32718 (N_32718,N_32205,N_30566);
and U32719 (N_32719,N_30033,N_31295);
and U32720 (N_32720,N_31401,N_31037);
and U32721 (N_32721,N_30465,N_32484);
and U32722 (N_32722,N_30929,N_32077);
nor U32723 (N_32723,N_30074,N_32202);
or U32724 (N_32724,N_31495,N_31255);
and U32725 (N_32725,N_31429,N_30172);
or U32726 (N_32726,N_31484,N_31421);
or U32727 (N_32727,N_31572,N_30063);
nand U32728 (N_32728,N_31500,N_30385);
nor U32729 (N_32729,N_31297,N_32329);
nand U32730 (N_32730,N_30937,N_31164);
xor U32731 (N_32731,N_31068,N_32233);
or U32732 (N_32732,N_31828,N_30612);
or U32733 (N_32733,N_31308,N_31161);
nand U32734 (N_32734,N_31766,N_31472);
or U32735 (N_32735,N_31248,N_31703);
xnor U32736 (N_32736,N_30986,N_30906);
xor U32737 (N_32737,N_30160,N_31287);
nand U32738 (N_32738,N_31486,N_30386);
nand U32739 (N_32739,N_31122,N_31177);
or U32740 (N_32740,N_31264,N_32214);
nand U32741 (N_32741,N_31937,N_31380);
xor U32742 (N_32742,N_31942,N_30743);
nor U32743 (N_32743,N_30196,N_32011);
or U32744 (N_32744,N_30974,N_30192);
and U32745 (N_32745,N_32128,N_30143);
nand U32746 (N_32746,N_31639,N_30844);
nand U32747 (N_32747,N_30548,N_30006);
xor U32748 (N_32748,N_31979,N_30666);
or U32749 (N_32749,N_30606,N_31697);
xnor U32750 (N_32750,N_31854,N_31447);
nand U32751 (N_32751,N_31333,N_30551);
nand U32752 (N_32752,N_30148,N_30830);
and U32753 (N_32753,N_31641,N_30460);
and U32754 (N_32754,N_31490,N_31601);
xnor U32755 (N_32755,N_30464,N_31534);
and U32756 (N_32756,N_32256,N_30349);
nor U32757 (N_32757,N_31096,N_30203);
nand U32758 (N_32758,N_32280,N_31216);
nand U32759 (N_32759,N_31352,N_31762);
xnor U32760 (N_32760,N_31452,N_32113);
nor U32761 (N_32761,N_31533,N_30380);
or U32762 (N_32762,N_30439,N_30298);
nor U32763 (N_32763,N_30197,N_30018);
xnor U32764 (N_32764,N_31677,N_30791);
nand U32765 (N_32765,N_30191,N_32027);
nand U32766 (N_32766,N_30339,N_31135);
or U32767 (N_32767,N_30888,N_30882);
or U32768 (N_32768,N_31427,N_31921);
nor U32769 (N_32769,N_30543,N_30131);
xor U32770 (N_32770,N_31032,N_31710);
and U32771 (N_32771,N_32198,N_32331);
and U32772 (N_32772,N_31808,N_31785);
or U32773 (N_32773,N_30375,N_30936);
or U32774 (N_32774,N_30971,N_32235);
xnor U32775 (N_32775,N_30261,N_31769);
nand U32776 (N_32776,N_31957,N_32393);
or U32777 (N_32777,N_30933,N_31203);
and U32778 (N_32778,N_30262,N_32434);
and U32779 (N_32779,N_30972,N_32493);
nor U32780 (N_32780,N_30442,N_31060);
nor U32781 (N_32781,N_30944,N_32065);
and U32782 (N_32782,N_30758,N_31110);
or U32783 (N_32783,N_31443,N_31755);
nand U32784 (N_32784,N_30631,N_31299);
nand U32785 (N_32785,N_31395,N_31784);
and U32786 (N_32786,N_30369,N_30648);
nand U32787 (N_32787,N_32054,N_31635);
and U32788 (N_32788,N_31917,N_32480);
nand U32789 (N_32789,N_30212,N_30085);
nor U32790 (N_32790,N_30958,N_31467);
or U32791 (N_32791,N_31739,N_31623);
or U32792 (N_32792,N_31693,N_32033);
and U32793 (N_32793,N_30695,N_32120);
nor U32794 (N_32794,N_30862,N_32060);
nor U32795 (N_32795,N_30628,N_31307);
or U32796 (N_32796,N_30126,N_30377);
xor U32797 (N_32797,N_30458,N_31830);
and U32798 (N_32798,N_30871,N_31922);
nor U32799 (N_32799,N_30194,N_30922);
nand U32800 (N_32800,N_31011,N_30663);
xnor U32801 (N_32801,N_30397,N_31561);
nand U32802 (N_32802,N_32499,N_31145);
nor U32803 (N_32803,N_32182,N_31680);
and U32804 (N_32804,N_32105,N_30679);
or U32805 (N_32805,N_31849,N_30692);
nor U32806 (N_32806,N_31302,N_31494);
nor U32807 (N_32807,N_31718,N_31558);
or U32808 (N_32808,N_32304,N_31136);
nor U32809 (N_32809,N_32295,N_31034);
and U32810 (N_32810,N_31978,N_32135);
and U32811 (N_32811,N_31709,N_31970);
and U32812 (N_32812,N_32146,N_32296);
nand U32813 (N_32813,N_31511,N_32013);
nand U32814 (N_32814,N_30951,N_30569);
or U32815 (N_32815,N_30315,N_30272);
nand U32816 (N_32816,N_31036,N_31860);
nor U32817 (N_32817,N_31630,N_32477);
xor U32818 (N_32818,N_31621,N_30462);
and U32819 (N_32819,N_30581,N_32341);
xnor U32820 (N_32820,N_30640,N_32374);
or U32821 (N_32821,N_30133,N_32496);
xor U32822 (N_32822,N_30271,N_30603);
or U32823 (N_32823,N_31273,N_30338);
nor U32824 (N_32824,N_30831,N_30428);
nor U32825 (N_32825,N_32401,N_32171);
xor U32826 (N_32826,N_31000,N_30039);
or U32827 (N_32827,N_30062,N_31257);
or U32828 (N_32828,N_30816,N_30637);
nor U32829 (N_32829,N_32411,N_32343);
or U32830 (N_32830,N_32230,N_31430);
and U32831 (N_32831,N_32251,N_31679);
xnor U32832 (N_32832,N_30840,N_30776);
or U32833 (N_32833,N_30510,N_31094);
or U32834 (N_32834,N_30219,N_31411);
or U32835 (N_32835,N_30471,N_32352);
and U32836 (N_32836,N_30432,N_30246);
or U32837 (N_32837,N_32039,N_30107);
and U32838 (N_32838,N_30899,N_31109);
nand U32839 (N_32839,N_31223,N_31569);
and U32840 (N_32840,N_31634,N_30394);
xor U32841 (N_32841,N_30313,N_30749);
xor U32842 (N_32842,N_31713,N_31359);
or U32843 (N_32843,N_32250,N_31020);
nor U32844 (N_32844,N_32044,N_32437);
xnor U32845 (N_32845,N_32383,N_31996);
or U32846 (N_32846,N_31843,N_30524);
nand U32847 (N_32847,N_30166,N_31751);
nor U32848 (N_32848,N_30354,N_30708);
xnor U32849 (N_32849,N_31560,N_30356);
xnor U32850 (N_32850,N_32119,N_31522);
nor U32851 (N_32851,N_30590,N_31986);
xor U32852 (N_32852,N_31765,N_32409);
and U32853 (N_32853,N_31363,N_32095);
nand U32854 (N_32854,N_31434,N_30994);
and U32855 (N_32855,N_31878,N_30886);
and U32856 (N_32856,N_30655,N_30864);
xor U32857 (N_32857,N_32116,N_30690);
or U32858 (N_32858,N_31962,N_31442);
nand U32859 (N_32859,N_32174,N_31687);
xnor U32860 (N_32860,N_31456,N_32125);
xor U32861 (N_32861,N_30538,N_31372);
nor U32862 (N_32862,N_31850,N_31219);
and U32863 (N_32863,N_31251,N_31336);
nor U32864 (N_32864,N_30764,N_31321);
and U32865 (N_32865,N_31331,N_30627);
nor U32866 (N_32866,N_31407,N_30323);
and U32867 (N_32867,N_32240,N_31776);
or U32868 (N_32868,N_30503,N_30051);
and U32869 (N_32869,N_31496,N_30784);
and U32870 (N_32870,N_31651,N_31546);
xnor U32871 (N_32871,N_31760,N_32446);
xnor U32872 (N_32872,N_31015,N_31585);
nor U32873 (N_32873,N_31465,N_32227);
xor U32874 (N_32874,N_31182,N_31685);
and U32875 (N_32875,N_32269,N_30744);
nand U32876 (N_32876,N_31935,N_31174);
and U32877 (N_32877,N_32270,N_31090);
nor U32878 (N_32878,N_30179,N_31106);
xor U32879 (N_32879,N_30105,N_31432);
or U32880 (N_32880,N_30024,N_30533);
nor U32881 (N_32881,N_31529,N_31089);
xnor U32882 (N_32882,N_31422,N_32472);
nor U32883 (N_32883,N_31348,N_31945);
nand U32884 (N_32884,N_31622,N_31449);
nand U32885 (N_32885,N_31468,N_30358);
or U32886 (N_32886,N_31702,N_30329);
or U32887 (N_32887,N_31414,N_32056);
or U32888 (N_32888,N_30724,N_31593);
nand U32889 (N_32889,N_32318,N_30027);
and U32890 (N_32890,N_31129,N_30461);
xor U32891 (N_32891,N_30546,N_31301);
or U32892 (N_32892,N_32126,N_31833);
nand U32893 (N_32893,N_30325,N_31204);
nand U32894 (N_32894,N_31445,N_32026);
and U32895 (N_32895,N_30583,N_32302);
nor U32896 (N_32896,N_32045,N_31883);
nor U32897 (N_32897,N_30809,N_30878);
or U32898 (N_32898,N_30897,N_31479);
or U32899 (N_32899,N_30867,N_30981);
and U32900 (N_32900,N_32047,N_30234);
or U32901 (N_32901,N_30717,N_32345);
nand U32902 (N_32902,N_31502,N_30505);
nand U32903 (N_32903,N_30324,N_30484);
or U32904 (N_32904,N_30398,N_30950);
or U32905 (N_32905,N_31039,N_32217);
nor U32906 (N_32906,N_32333,N_31517);
nand U32907 (N_32907,N_32195,N_30662);
nor U32908 (N_32908,N_32169,N_31076);
and U32909 (N_32909,N_31001,N_32309);
and U32910 (N_32910,N_32485,N_30168);
xnor U32911 (N_32911,N_32281,N_30668);
nor U32912 (N_32912,N_32379,N_30336);
nor U32913 (N_32913,N_30064,N_31525);
nand U32914 (N_32914,N_31066,N_31056);
and U32915 (N_32915,N_31637,N_31879);
nand U32916 (N_32916,N_30736,N_31221);
and U32917 (N_32917,N_32299,N_30011);
or U32918 (N_32918,N_31872,N_30401);
xnor U32919 (N_32919,N_30090,N_32417);
nand U32920 (N_32920,N_31940,N_32092);
nand U32921 (N_32921,N_32445,N_31139);
and U32922 (N_32922,N_31253,N_31596);
nand U32923 (N_32923,N_32448,N_30523);
or U32924 (N_32924,N_30059,N_31545);
or U32925 (N_32925,N_31789,N_30941);
xor U32926 (N_32926,N_32037,N_31905);
xnor U32927 (N_32927,N_31586,N_31890);
and U32928 (N_32928,N_30350,N_31285);
or U32929 (N_32929,N_30297,N_30456);
and U32930 (N_32930,N_31786,N_32451);
nor U32931 (N_32931,N_30357,N_30970);
xor U32932 (N_32932,N_31377,N_32098);
nand U32933 (N_32933,N_30682,N_31364);
and U32934 (N_32934,N_30108,N_30376);
nor U32935 (N_32935,N_31117,N_30726);
and U32936 (N_32936,N_31987,N_31782);
and U32937 (N_32937,N_30843,N_30673);
or U32938 (N_32938,N_31575,N_30236);
nand U32939 (N_32939,N_31868,N_32123);
nor U32940 (N_32940,N_30697,N_31262);
or U32941 (N_32941,N_32087,N_30479);
nand U32942 (N_32942,N_30514,N_30156);
nand U32943 (N_32943,N_31323,N_32133);
nor U32944 (N_32944,N_30594,N_32052);
xor U32945 (N_32945,N_31510,N_32425);
or U32946 (N_32946,N_32442,N_30928);
and U32947 (N_32947,N_30506,N_30653);
nor U32948 (N_32948,N_32298,N_31440);
and U32949 (N_32949,N_31645,N_32089);
or U32950 (N_32950,N_30274,N_30400);
nand U32951 (N_32951,N_30558,N_31416);
and U32952 (N_32952,N_31875,N_30111);
and U32953 (N_32953,N_32316,N_30621);
xnor U32954 (N_32954,N_32410,N_31629);
xnor U32955 (N_32955,N_30268,N_30187);
xor U32956 (N_32956,N_31012,N_32310);
nor U32957 (N_32957,N_31294,N_30130);
nand U32958 (N_32958,N_31515,N_31296);
nand U32959 (N_32959,N_31555,N_31880);
and U32960 (N_32960,N_30169,N_30070);
xnor U32961 (N_32961,N_31070,N_31408);
nor U32962 (N_32962,N_31238,N_30909);
and U32963 (N_32963,N_30854,N_30221);
xnor U32964 (N_32964,N_30017,N_31201);
and U32965 (N_32965,N_31017,N_31289);
or U32966 (N_32966,N_31453,N_31108);
xnor U32967 (N_32967,N_31389,N_30925);
nor U32968 (N_32968,N_31425,N_32216);
xnor U32969 (N_32969,N_31250,N_32019);
nor U32970 (N_32970,N_31179,N_31249);
xor U32971 (N_32971,N_32391,N_32141);
or U32972 (N_32972,N_31983,N_32389);
nand U32973 (N_32973,N_30982,N_31016);
or U32974 (N_32974,N_30424,N_32319);
or U32975 (N_32975,N_30005,N_31029);
or U32976 (N_32976,N_30141,N_32069);
nor U32977 (N_32977,N_31514,N_31589);
xnor U32978 (N_32978,N_31619,N_30086);
xnor U32979 (N_32979,N_30303,N_32357);
nor U32980 (N_32980,N_32213,N_30522);
nand U32981 (N_32981,N_32167,N_32185);
nand U32982 (N_32982,N_32136,N_32454);
nand U32983 (N_32983,N_31796,N_31206);
xor U32984 (N_32984,N_30333,N_30241);
xnor U32985 (N_32985,N_30582,N_30256);
xnor U32986 (N_32986,N_31565,N_31045);
nand U32987 (N_32987,N_31144,N_30216);
nand U32988 (N_32988,N_30935,N_31582);
or U32989 (N_32989,N_30429,N_31303);
xnor U32990 (N_32990,N_32497,N_32143);
nor U32991 (N_32991,N_30707,N_32030);
or U32992 (N_32992,N_30188,N_30492);
or U32993 (N_32993,N_30737,N_32396);
xnor U32994 (N_32994,N_30837,N_31375);
or U32995 (N_32995,N_30846,N_32372);
or U32996 (N_32996,N_32353,N_31385);
and U32997 (N_32997,N_30122,N_30296);
nand U32998 (N_32998,N_32473,N_30446);
xor U32999 (N_32999,N_31906,N_31246);
or U33000 (N_33000,N_30227,N_31543);
xor U33001 (N_33001,N_31454,N_31895);
and U33002 (N_33002,N_30472,N_31007);
nor U33003 (N_33003,N_31335,N_30281);
xnor U33004 (N_33004,N_31670,N_32218);
nand U33005 (N_33005,N_30286,N_31022);
xor U33006 (N_33006,N_31715,N_30622);
and U33007 (N_33007,N_32490,N_31085);
and U33008 (N_33008,N_31721,N_32447);
or U33009 (N_33009,N_30073,N_30257);
nand U33010 (N_33010,N_31192,N_30518);
nor U33011 (N_33011,N_31887,N_32440);
xor U33012 (N_33012,N_32453,N_32328);
or U33013 (N_33013,N_31607,N_30406);
nand U33014 (N_33014,N_30557,N_32090);
nand U33015 (N_33015,N_30034,N_31757);
nand U33016 (N_33016,N_30534,N_31936);
or U33017 (N_33017,N_31617,N_32015);
or U33018 (N_33018,N_31931,N_30209);
nand U33019 (N_33019,N_30161,N_30879);
nor U33020 (N_33020,N_30466,N_30010);
xnor U33021 (N_33021,N_31567,N_31132);
xor U33022 (N_33022,N_31351,N_30788);
or U33023 (N_33023,N_30714,N_31313);
nand U33024 (N_33024,N_30919,N_31282);
nor U33025 (N_33025,N_31893,N_30393);
or U33026 (N_33026,N_31611,N_32405);
xor U33027 (N_33027,N_30288,N_31506);
xor U33028 (N_33028,N_30934,N_31175);
and U33029 (N_33029,N_31745,N_31459);
nand U33030 (N_33030,N_30529,N_30331);
xor U33031 (N_33031,N_31355,N_31382);
nand U33032 (N_33032,N_32076,N_31155);
nor U33033 (N_33033,N_31463,N_31315);
nand U33034 (N_33034,N_30162,N_30224);
xnor U33035 (N_33035,N_30734,N_31903);
or U33036 (N_33036,N_31925,N_31584);
nor U33037 (N_33037,N_30576,N_30638);
nor U33038 (N_33038,N_31790,N_31688);
xnor U33039 (N_33039,N_30541,N_30977);
and U33040 (N_33040,N_30178,N_31214);
or U33041 (N_33041,N_32158,N_30652);
or U33042 (N_33042,N_30954,N_31280);
xnor U33043 (N_33043,N_30760,N_31579);
nor U33044 (N_33044,N_30905,N_32356);
nor U33045 (N_33045,N_32204,N_30881);
nand U33046 (N_33046,N_31810,N_31074);
or U33047 (N_33047,N_32248,N_30117);
nor U33048 (N_33048,N_31350,N_31662);
or U33049 (N_33049,N_31242,N_30939);
or U33050 (N_33050,N_30302,N_30615);
nor U33051 (N_33051,N_31183,N_30030);
or U33052 (N_33052,N_30777,N_30211);
and U33053 (N_33053,N_30544,N_30371);
or U33054 (N_33054,N_31373,N_31091);
xor U33055 (N_33055,N_31732,N_32189);
xnor U33056 (N_33056,N_31773,N_31625);
and U33057 (N_33057,N_31058,N_30507);
or U33058 (N_33058,N_32363,N_32262);
or U33059 (N_33059,N_31727,N_31958);
xnor U33060 (N_33060,N_32305,N_30811);
xor U33061 (N_33061,N_31994,N_31820);
xor U33062 (N_33062,N_31141,N_32264);
xor U33063 (N_33063,N_30207,N_30938);
and U33064 (N_33064,N_30820,N_31923);
nand U33065 (N_33065,N_30999,N_32282);
xor U33066 (N_33066,N_32082,N_30137);
or U33067 (N_33067,N_32461,N_31403);
xnor U33068 (N_33068,N_31349,N_32165);
nand U33069 (N_33069,N_30766,N_30413);
xor U33070 (N_33070,N_30705,N_32421);
and U33071 (N_33071,N_30127,N_31077);
or U33072 (N_33072,N_30206,N_31065);
nand U33073 (N_33073,N_30630,N_32142);
and U33074 (N_33074,N_30330,N_30083);
nor U33075 (N_33075,N_31912,N_32390);
and U33076 (N_33076,N_31112,N_31230);
nand U33077 (N_33077,N_31832,N_30159);
nor U33078 (N_33078,N_32351,N_30992);
xnor U33079 (N_33079,N_30709,N_31381);
and U33080 (N_33080,N_31892,N_32086);
and U33081 (N_33081,N_30455,N_31746);
or U33082 (N_33082,N_32088,N_31512);
or U33083 (N_33083,N_30956,N_30152);
and U33084 (N_33084,N_30781,N_30532);
nand U33085 (N_33085,N_30476,N_31188);
or U33086 (N_33086,N_32267,N_32194);
or U33087 (N_33087,N_30949,N_30686);
and U33088 (N_33088,N_32097,N_31332);
xnor U33089 (N_33089,N_30057,N_32149);
and U33090 (N_33090,N_30101,N_30020);
nor U33091 (N_33091,N_30364,N_30140);
and U33092 (N_33092,N_31547,N_30817);
and U33093 (N_33093,N_30656,N_30050);
and U33094 (N_33094,N_30613,N_31314);
nand U33095 (N_33095,N_31886,N_30754);
nor U33096 (N_33096,N_32346,N_31527);
and U33097 (N_33097,N_31101,N_31731);
xor U33098 (N_33098,N_30346,N_32283);
and U33099 (N_33099,N_30556,N_32168);
nor U33100 (N_33100,N_31341,N_32460);
or U33101 (N_33101,N_32150,N_31811);
nor U33102 (N_33102,N_31717,N_32139);
nand U33103 (N_33103,N_30672,N_30080);
nand U33104 (N_33104,N_30516,N_31274);
nor U33105 (N_33105,N_32258,N_30307);
or U33106 (N_33106,N_30310,N_31650);
xnor U33107 (N_33107,N_31482,N_31105);
or U33108 (N_33108,N_31478,N_31102);
and U33109 (N_33109,N_30755,N_31959);
and U33110 (N_33110,N_31602,N_31080);
xnor U33111 (N_33111,N_30921,N_31781);
and U33112 (N_33112,N_31816,N_31807);
nand U33113 (N_33113,N_31965,N_30794);
or U33114 (N_33114,N_30803,N_30040);
and U33115 (N_33115,N_30000,N_30237);
nor U33116 (N_33116,N_31052,N_31093);
and U33117 (N_33117,N_31758,N_31476);
xor U33118 (N_33118,N_32284,N_32272);
or U33119 (N_33119,N_30158,N_31666);
nand U33120 (N_33120,N_30205,N_32108);
or U33121 (N_33121,N_30713,N_30890);
or U33122 (N_33122,N_32014,N_31291);
nand U33123 (N_33123,N_32290,N_30808);
nor U33124 (N_33124,N_31708,N_32432);
nand U33125 (N_33125,N_31346,N_30617);
xor U33126 (N_33126,N_30642,N_30804);
xnor U33127 (N_33127,N_30822,N_30438);
and U33128 (N_33128,N_32244,N_30826);
xor U33129 (N_33129,N_30322,N_31682);
or U33130 (N_33130,N_31675,N_30388);
and U33131 (N_33131,N_30866,N_31787);
or U33132 (N_33132,N_31774,N_31817);
xor U33133 (N_33133,N_31021,N_32161);
and U33134 (N_33134,N_32433,N_31852);
nor U33135 (N_33135,N_31859,N_31498);
or U33136 (N_33136,N_30563,N_30945);
and U33137 (N_33137,N_30165,N_30693);
xor U33138 (N_33138,N_31312,N_31471);
or U33139 (N_33139,N_32157,N_31552);
or U33140 (N_33140,N_31904,N_30748);
nor U33141 (N_33141,N_32424,N_32079);
and U33142 (N_33142,N_30102,N_30082);
and U33143 (N_33143,N_30423,N_32007);
nor U33144 (N_33144,N_31981,N_31146);
nand U33145 (N_33145,N_30235,N_30129);
nor U33146 (N_33146,N_30289,N_31305);
and U33147 (N_33147,N_31521,N_30865);
nor U33148 (N_33148,N_31329,N_31067);
and U33149 (N_33149,N_31877,N_32183);
nand U33150 (N_33150,N_30242,N_32495);
or U33151 (N_33151,N_31894,N_31437);
nand U33152 (N_33152,N_32326,N_30965);
nand U33153 (N_33153,N_30891,N_30381);
nor U33154 (N_33154,N_30883,N_31993);
xnor U33155 (N_33155,N_31181,N_30047);
nor U33156 (N_33156,N_31711,N_31627);
xor U33157 (N_33157,N_32115,N_30468);
nor U33158 (N_33158,N_30703,N_30810);
nor U33159 (N_33159,N_31424,N_30768);
or U33160 (N_33160,N_30252,N_32486);
nor U33161 (N_33161,N_32176,N_30677);
nor U33162 (N_33162,N_30355,N_31180);
xor U33163 (N_33163,N_30815,N_30535);
or U33164 (N_33164,N_30664,N_30598);
nor U33165 (N_33165,N_30383,N_32112);
nand U33166 (N_33166,N_32160,N_32106);
nand U33167 (N_33167,N_30742,N_32271);
or U33168 (N_33168,N_31092,N_32339);
nor U33169 (N_33169,N_32000,N_30559);
or U33170 (N_33170,N_30660,N_31701);
nand U33171 (N_33171,N_30136,N_32023);
or U33172 (N_33172,N_31665,N_31387);
nor U33173 (N_33173,N_30752,N_30292);
nor U33174 (N_33174,N_30550,N_31300);
nor U33175 (N_33175,N_30202,N_30214);
or U33176 (N_33176,N_30985,N_30348);
xnor U33177 (N_33177,N_30067,N_30218);
and U33178 (N_33178,N_30319,N_32220);
or U33179 (N_33179,N_30948,N_31428);
nor U33180 (N_33180,N_31663,N_30975);
nor U33181 (N_33181,N_32273,N_30564);
xor U33182 (N_33182,N_30723,N_30200);
and U33183 (N_33183,N_31767,N_30649);
nor U33184 (N_33184,N_31213,N_30407);
and U33185 (N_33185,N_30853,N_31920);
nand U33186 (N_33186,N_30841,N_31616);
and U33187 (N_33187,N_30250,N_31292);
nand U33188 (N_33188,N_31013,N_30263);
nor U33189 (N_33189,N_32091,N_30500);
xor U33190 (N_33190,N_30374,N_30071);
or U33191 (N_33191,N_30217,N_32208);
nand U33192 (N_33192,N_32212,N_30735);
and U33193 (N_33193,N_31163,N_32055);
or U33194 (N_33194,N_31600,N_31215);
and U33195 (N_33195,N_31358,N_30459);
nor U33196 (N_33196,N_32223,N_30636);
nor U33197 (N_33197,N_30545,N_31152);
or U33198 (N_33198,N_30387,N_30334);
and U33199 (N_33199,N_30552,N_30596);
and U33200 (N_33200,N_32291,N_30060);
xor U33201 (N_33201,N_30610,N_30991);
nand U33202 (N_33202,N_30260,N_30096);
nand U33203 (N_33203,N_32080,N_31266);
xnor U33204 (N_33204,N_32479,N_31801);
xor U33205 (N_33205,N_30037,N_32117);
nor U33206 (N_33206,N_31998,N_31244);
xnor U33207 (N_33207,N_30643,N_30889);
or U33208 (N_33208,N_31574,N_31620);
or U33209 (N_33209,N_30220,N_31749);
nand U33210 (N_33210,N_30395,N_31412);
and U33211 (N_33211,N_30659,N_32209);
nor U33212 (N_33212,N_30917,N_30983);
or U33213 (N_33213,N_30812,N_31322);
xor U33214 (N_33214,N_32148,N_30265);
nand U33215 (N_33215,N_30685,N_31005);
or U33216 (N_33216,N_32118,N_32170);
nor U33217 (N_33217,N_31858,N_32024);
nand U33218 (N_33218,N_31049,N_31288);
or U33219 (N_33219,N_31319,N_30930);
and U33220 (N_33220,N_32404,N_32450);
xor U33221 (N_33221,N_30463,N_31599);
nand U33222 (N_33222,N_30715,N_31062);
or U33223 (N_33223,N_31540,N_32413);
and U33224 (N_33224,N_31086,N_31410);
nand U33225 (N_33225,N_31393,N_31079);
and U33226 (N_33226,N_30493,N_31982);
xor U33227 (N_33227,N_30100,N_32083);
nor U33228 (N_33228,N_31698,N_32481);
and U33229 (N_33229,N_30175,N_31590);
and U33230 (N_33230,N_30570,N_30870);
nand U33231 (N_33231,N_30984,N_30646);
xnor U33232 (N_33232,N_30624,N_31386);
nor U33233 (N_33233,N_32084,N_31268);
or U33234 (N_33234,N_30761,N_31318);
and U33235 (N_33235,N_30711,N_31562);
nor U33236 (N_33236,N_30379,N_30412);
xnor U33237 (N_33237,N_30997,N_31239);
and U33238 (N_33238,N_31487,N_30041);
and U33239 (N_33239,N_30568,N_32075);
or U33240 (N_33240,N_30800,N_31405);
or U33241 (N_33241,N_30802,N_31794);
and U33242 (N_33242,N_31460,N_30031);
and U33243 (N_33243,N_31851,N_32279);
nor U33244 (N_33244,N_32277,N_32243);
nand U33245 (N_33245,N_31189,N_31822);
nand U33246 (N_33246,N_30528,N_30382);
and U33247 (N_33247,N_32475,N_31231);
or U33248 (N_33248,N_31800,N_30762);
nor U33249 (N_33249,N_31573,N_31597);
xor U33250 (N_33250,N_32094,N_32147);
nor U33251 (N_33251,N_31610,N_30243);
and U33252 (N_33252,N_30602,N_31176);
and U33253 (N_33253,N_31027,N_30592);
or U33254 (N_33254,N_30452,N_30589);
nand U33255 (N_33255,N_30625,N_30892);
nor U33256 (N_33256,N_31956,N_30769);
nand U33257 (N_33257,N_31267,N_30154);
nand U33258 (N_33258,N_31111,N_31360);
and U33259 (N_33259,N_31120,N_31448);
and U33260 (N_33260,N_30426,N_30496);
and U33261 (N_33261,N_30119,N_30499);
nand U33262 (N_33262,N_30396,N_30893);
nand U33263 (N_33263,N_32197,N_30417);
and U33264 (N_33264,N_31388,N_30093);
nor U33265 (N_33265,N_31293,N_30924);
and U33266 (N_33266,N_30309,N_30738);
or U33267 (N_33267,N_31126,N_32278);
or U33268 (N_33268,N_30470,N_30186);
and U33269 (N_33269,N_32489,N_32051);
or U33270 (N_33270,N_31024,N_32053);
nand U33271 (N_33271,N_32399,N_32312);
xnor U33272 (N_33272,N_31591,N_31730);
xnor U33273 (N_33273,N_32068,N_31819);
xor U33274 (N_33274,N_30293,N_30351);
xor U33275 (N_33275,N_31504,N_30609);
and U33276 (N_33276,N_32254,N_32028);
xnor U33277 (N_33277,N_31659,N_30990);
nand U33278 (N_33278,N_30454,N_31681);
and U33279 (N_33279,N_31559,N_30953);
nand U33280 (N_33280,N_30444,N_30683);
xnor U33281 (N_33281,N_32276,N_30304);
nand U33282 (N_33282,N_30940,N_31707);
or U33283 (N_33283,N_30482,N_30150);
xnor U33284 (N_33284,N_32187,N_31162);
and U33285 (N_33285,N_31138,N_31694);
nand U33286 (N_33286,N_32371,N_31549);
nor U33287 (N_33287,N_32239,N_31225);
nand U33288 (N_33288,N_30635,N_32360);
and U33289 (N_33289,N_30806,N_31944);
nand U33290 (N_33290,N_31237,N_32074);
and U33291 (N_33291,N_31753,N_30414);
xnor U33292 (N_33292,N_31072,N_31004);
nand U33293 (N_33293,N_30730,N_30857);
nand U33294 (N_33294,N_31191,N_30177);
xor U33295 (N_33295,N_31261,N_31324);
xnor U33296 (N_33296,N_31898,N_32321);
and U33297 (N_33297,N_31536,N_30498);
nor U33298 (N_33298,N_32462,N_31207);
or U33299 (N_33299,N_31588,N_31473);
nand U33300 (N_33300,N_30015,N_32349);
nor U33301 (N_33301,N_31455,N_30185);
xor U33302 (N_33302,N_30902,N_31985);
xnor U33303 (N_33303,N_31187,N_30632);
or U33304 (N_33304,N_30511,N_31550);
and U33305 (N_33305,N_31963,N_30342);
nor U33306 (N_33306,N_31172,N_31233);
or U33307 (N_33307,N_31391,N_30199);
and U33308 (N_33308,N_32252,N_31009);
xor U33309 (N_33309,N_31489,N_31624);
nand U33310 (N_33310,N_30299,N_31446);
or U33311 (N_33311,N_31648,N_32487);
and U33312 (N_33312,N_30494,N_30416);
nand U33313 (N_33313,N_32494,N_31142);
nor U33314 (N_33314,N_31413,N_30410);
nor U33315 (N_33315,N_30961,N_30825);
nand U33316 (N_33316,N_31777,N_32476);
nand U33317 (N_33317,N_31185,N_30473);
or U33318 (N_33318,N_30588,N_31279);
xor U33319 (N_33319,N_31073,N_30163);
or U33320 (N_33320,N_31719,N_30989);
nor U33321 (N_33321,N_31969,N_30626);
nor U33322 (N_33322,N_30419,N_30932);
and U33323 (N_33323,N_31673,N_30828);
and U33324 (N_33324,N_31915,N_30858);
nor U33325 (N_33325,N_31046,N_31409);
nand U33326 (N_33326,N_31884,N_31909);
nand U33327 (N_33327,N_32415,N_31184);
and U33328 (N_33328,N_30547,N_32470);
xnor U33329 (N_33329,N_30763,N_31866);
nor U33330 (N_33330,N_30706,N_30055);
and U33331 (N_33331,N_32012,N_31740);
or U33332 (N_33332,N_30149,N_30092);
and U33333 (N_33333,N_32412,N_32061);
xnor U33334 (N_33334,N_31087,N_30488);
and U33335 (N_33335,N_32072,N_30947);
or U33336 (N_33336,N_31551,N_32444);
nand U33337 (N_33337,N_30180,N_31960);
nand U33338 (N_33338,N_30827,N_31530);
nor U33339 (N_33339,N_31952,N_32155);
xor U33340 (N_33340,N_31672,N_31975);
and U33341 (N_33341,N_30430,N_30337);
nand U33342 (N_33342,N_31913,N_32018);
nor U33343 (N_33343,N_30856,N_30305);
or U33344 (N_33344,N_30483,N_31578);
nand U33345 (N_33345,N_30580,N_32439);
xor U33346 (N_33346,N_30519,N_30091);
nor U33347 (N_33347,N_31643,N_32246);
or U33348 (N_33348,N_30537,N_30979);
nor U33349 (N_33349,N_30575,N_32059);
and U33350 (N_33350,N_30845,N_31317);
nor U33351 (N_33351,N_32376,N_31752);
xnor U33352 (N_33352,N_30667,N_30294);
and U33353 (N_33353,N_30623,N_31930);
xnor U33354 (N_33354,N_31628,N_31160);
or U33355 (N_33355,N_30248,N_31167);
and U33356 (N_33356,N_31772,N_31742);
xnor U33357 (N_33357,N_30876,N_32022);
and U33358 (N_33358,N_31269,N_31173);
xor U33359 (N_33359,N_32464,N_30244);
nor U33360 (N_33360,N_32287,N_32420);
or U33361 (N_33361,N_30495,N_30437);
nand U33362 (N_33362,N_30056,N_30363);
and U33363 (N_33363,N_31997,N_30525);
and U33364 (N_33364,N_31469,N_30118);
nor U33365 (N_33365,N_30614,N_30392);
nor U33366 (N_33366,N_31481,N_30069);
and U33367 (N_33367,N_30894,N_32458);
nand U33368 (N_33368,N_31030,N_31896);
or U33369 (N_33369,N_31276,N_31491);
and U33370 (N_33370,N_32313,N_31284);
nand U33371 (N_33371,N_30721,N_30536);
nand U33372 (N_33372,N_31104,N_31170);
xor U33373 (N_33373,N_32441,N_30247);
xor U33374 (N_33374,N_31736,N_31311);
nand U33375 (N_33375,N_30783,N_30561);
or U33376 (N_33376,N_31061,N_32121);
xor U33377 (N_33377,N_31082,N_32314);
xnor U33378 (N_33378,N_30955,N_31148);
nand U33379 (N_33379,N_31519,N_30756);
or U33380 (N_33380,N_30004,N_30254);
or U33381 (N_33381,N_32181,N_32373);
and U33382 (N_33382,N_31618,N_32452);
and U33383 (N_33383,N_30089,N_30103);
or U33384 (N_33384,N_32021,N_31831);
and U33385 (N_33385,N_30741,N_32073);
or U33386 (N_33386,N_31838,N_32400);
nand U33387 (N_33387,N_32488,N_30680);
nor U33388 (N_33388,N_31825,N_30003);
and U33389 (N_33389,N_31059,N_30729);
nand U33390 (N_33390,N_30368,N_32407);
nand U33391 (N_33391,N_31631,N_30676);
xnor U33392 (N_33392,N_31376,N_30270);
nand U33393 (N_33393,N_30475,N_32001);
xor U33394 (N_33394,N_31042,N_30654);
and U33395 (N_33395,N_31228,N_31220);
nor U33396 (N_33396,N_31595,N_30174);
nor U33397 (N_33397,N_31435,N_30847);
nand U33398 (N_33398,N_30952,N_31474);
or U33399 (N_33399,N_30115,N_31316);
and U33400 (N_33400,N_30048,N_31814);
xor U33401 (N_33401,N_31870,N_30072);
xnor U33402 (N_33402,N_32140,N_30132);
nand U33403 (N_33403,N_30182,N_30732);
nand U33404 (N_33404,N_31143,N_31735);
nor U33405 (N_33405,N_31827,N_32008);
or U33406 (N_33406,N_32308,N_30880);
nor U33407 (N_33407,N_30120,N_31948);
or U33408 (N_33408,N_31638,N_30099);
xor U33409 (N_33409,N_31690,N_30790);
or U33410 (N_33410,N_31134,N_31891);
nor U33411 (N_33411,N_31415,N_32307);
or U33412 (N_33412,N_32402,N_30520);
nand U33413 (N_33413,N_31256,N_31114);
or U33414 (N_33414,N_30813,N_30253);
nor U33415 (N_33415,N_31342,N_30875);
nor U33416 (N_33416,N_30789,N_31006);
nand U33417 (N_33417,N_30775,N_32255);
xor U33418 (N_33418,N_32336,N_31406);
or U33419 (N_33419,N_30425,N_31212);
nand U33420 (N_33420,N_31949,N_31157);
nor U33421 (N_33421,N_31855,N_31980);
and U33422 (N_33422,N_32423,N_31964);
or U33423 (N_33423,N_30223,N_30927);
and U33424 (N_33424,N_32102,N_30135);
xor U33425 (N_33425,N_31115,N_31821);
nor U33426 (N_33426,N_30411,N_31889);
nor U33427 (N_33427,N_31684,N_30328);
nor U33428 (N_33428,N_30832,N_32145);
xor U33429 (N_33429,N_30449,N_31083);
nand U33430 (N_33430,N_31374,N_30490);
nand U33431 (N_33431,N_31420,N_31258);
or U33432 (N_33432,N_30145,N_31899);
nand U33433 (N_33433,N_30427,N_31556);
and U33434 (N_33434,N_32303,N_30138);
or U33435 (N_33435,N_31723,N_30530);
and U33436 (N_33436,N_30842,N_31477);
and U33437 (N_33437,N_30731,N_31444);
and U33438 (N_33438,N_31218,N_30712);
xnor U33439 (N_33439,N_30699,N_30515);
and U33440 (N_33440,N_31399,N_31379);
nor U33441 (N_33441,N_32153,N_30591);
xor U33442 (N_33442,N_31553,N_32365);
or U33443 (N_33443,N_32031,N_30282);
nor U33444 (N_33444,N_30852,N_30671);
and U33445 (N_33445,N_32175,N_32332);
xnor U33446 (N_33446,N_30485,N_31874);
nor U33447 (N_33447,N_30467,N_31431);
or U33448 (N_33448,N_31924,N_31283);
xor U33449 (N_33449,N_31857,N_31347);
or U33450 (N_33450,N_32203,N_31340);
or U33451 (N_33451,N_32381,N_31051);
nor U33452 (N_33452,N_30164,N_32063);
xnor U33453 (N_33453,N_30531,N_30976);
xor U33454 (N_33454,N_31653,N_31747);
xor U33455 (N_33455,N_31362,N_30098);
nand U33456 (N_33456,N_32344,N_31973);
xor U33457 (N_33457,N_30025,N_31835);
or U33458 (N_33458,N_30549,N_32459);
and U33459 (N_33459,N_31989,N_31658);
nor U33460 (N_33460,N_30344,N_31526);
nor U33461 (N_33461,N_30850,N_30579);
or U33462 (N_33462,N_31153,N_30045);
xor U33463 (N_33463,N_31392,N_32236);
nand U33464 (N_33464,N_30042,N_31532);
or U33465 (N_33465,N_30980,N_30757);
xnor U33466 (N_33466,N_30963,N_30277);
or U33467 (N_33467,N_30477,N_30834);
nor U33468 (N_33468,N_32100,N_30404);
nor U33469 (N_33469,N_30691,N_30448);
xor U33470 (N_33470,N_32238,N_32193);
xnor U33471 (N_33471,N_32166,N_31542);
or U33472 (N_33472,N_31158,N_31661);
or U33473 (N_33473,N_31689,N_31806);
xnor U33474 (N_33474,N_32274,N_31211);
or U33475 (N_33475,N_30002,N_30295);
or U33476 (N_33476,N_31457,N_31919);
nor U33477 (N_33477,N_31943,N_31839);
xor U33478 (N_33478,N_30916,N_31577);
and U33479 (N_33479,N_31226,N_32335);
nor U33480 (N_33480,N_32392,N_30887);
nor U33481 (N_33481,N_30409,N_32226);
or U33482 (N_33482,N_31729,N_31813);
and U33483 (N_33483,N_31116,N_30269);
or U33484 (N_33484,N_31493,N_30833);
and U33485 (N_33485,N_31418,N_32048);
nand U33486 (N_33486,N_31696,N_32435);
nand U33487 (N_33487,N_30650,N_31932);
xor U33488 (N_33488,N_31290,N_30687);
nand U33489 (N_33489,N_30727,N_30855);
and U33490 (N_33490,N_30684,N_32455);
and U33491 (N_33491,N_30014,N_32369);
xnor U33492 (N_33492,N_31812,N_32190);
and U33493 (N_33493,N_30678,N_30312);
xor U33494 (N_33494,N_31417,N_31609);
nor U33495 (N_33495,N_31524,N_31779);
nor U33496 (N_33496,N_31247,N_31804);
nor U33497 (N_33497,N_30489,N_30728);
or U33498 (N_33498,N_31856,N_31863);
and U33499 (N_33499,N_31836,N_30079);
nor U33500 (N_33500,N_32206,N_30077);
and U33501 (N_33501,N_32201,N_30440);
xor U33502 (N_33502,N_32064,N_32219);
nand U33503 (N_33503,N_30213,N_31867);
nor U33504 (N_33504,N_30016,N_30153);
or U33505 (N_33505,N_30044,N_30390);
and U33506 (N_33506,N_31433,N_30081);
or U33507 (N_33507,N_30109,N_30597);
or U33508 (N_33508,N_30023,N_31632);
and U33509 (N_33509,N_31326,N_30481);
or U33510 (N_33510,N_30629,N_30453);
nor U33511 (N_33511,N_31178,N_30167);
and U33512 (N_33512,N_30946,N_30801);
nor U33513 (N_33513,N_30301,N_30094);
and U33514 (N_33514,N_31929,N_31537);
xnor U33515 (N_33515,N_32378,N_32062);
nor U33516 (N_33516,N_31123,N_31720);
or U33517 (N_33517,N_32006,N_32289);
nand U33518 (N_33518,N_31539,N_30701);
nand U33519 (N_33519,N_30969,N_31598);
or U33520 (N_33520,N_32385,N_30774);
nor U33521 (N_33521,N_31402,N_30509);
xnor U33522 (N_33522,N_31513,N_30903);
and U33523 (N_33523,N_31232,N_31649);
or U33524 (N_33524,N_32406,N_30422);
or U33525 (N_33525,N_30084,N_31834);
nand U33526 (N_33526,N_31205,N_32034);
xnor U33527 (N_33527,N_31234,N_30225);
and U33528 (N_33528,N_31439,N_31125);
or U33529 (N_33529,N_30480,N_30849);
xor U33530 (N_33530,N_31222,N_30670);
or U33531 (N_33531,N_30885,N_31604);
nor U33532 (N_33532,N_32107,N_31815);
and U33533 (N_33533,N_31743,N_30343);
or U33534 (N_33534,N_31853,N_32368);
or U33535 (N_33535,N_31366,N_31615);
and U33536 (N_33536,N_30861,N_30347);
or U33537 (N_33537,N_30962,N_32498);
nor U33538 (N_33538,N_30173,N_30009);
and U33539 (N_33539,N_30046,N_31683);
nand U33540 (N_33540,N_30698,N_30998);
and U33541 (N_33541,N_30251,N_31028);
nor U33542 (N_33542,N_30599,N_30240);
nand U33543 (N_33543,N_30725,N_32370);
or U33544 (N_33544,N_30075,N_31871);
nor U33545 (N_33545,N_31320,N_31564);
or U33546 (N_33546,N_32196,N_30644);
or U33547 (N_33547,N_31972,N_30391);
nand U33548 (N_33548,N_31594,N_31725);
nand U33549 (N_33549,N_31939,N_32005);
or U33550 (N_33550,N_31195,N_32286);
or U33551 (N_33551,N_31113,N_31338);
or U33552 (N_33552,N_31946,N_30508);
and U33553 (N_33553,N_30901,N_30739);
xor U33554 (N_33554,N_30326,N_31793);
nor U33555 (N_33555,N_31501,N_31075);
and U33556 (N_33556,N_30770,N_30318);
and U33557 (N_33557,N_31198,N_30926);
nor U33558 (N_33558,N_31356,N_31396);
and U33559 (N_33559,N_31281,N_30497);
xnor U33560 (N_33560,N_32046,N_32029);
nor U33561 (N_33561,N_32122,N_30574);
nand U33562 (N_33562,N_31976,N_31165);
nand U33563 (N_33563,N_31277,N_32293);
or U33564 (N_33564,N_31078,N_30527);
nand U33565 (N_33565,N_30112,N_30521);
and U33566 (N_33566,N_30780,N_32221);
nand U33567 (N_33567,N_30362,N_32224);
and U33568 (N_33568,N_32192,N_30370);
xor U33569 (N_33569,N_30750,N_31908);
and U33570 (N_33570,N_30366,N_32228);
nand U33571 (N_33571,N_31763,N_32110);
xor U33572 (N_33572,N_30389,N_30013);
nand U33573 (N_33573,N_32482,N_30907);
or U33574 (N_33574,N_32154,N_31497);
nor U33575 (N_33575,N_32362,N_31927);
nand U33576 (N_33576,N_31229,N_31541);
nand U33577 (N_33577,N_30372,N_30170);
and U33578 (N_33578,N_32355,N_31640);
nand U33579 (N_33579,N_32324,N_32257);
and U33580 (N_33580,N_30068,N_31953);
xor U33581 (N_33581,N_31700,N_31357);
or U33582 (N_33582,N_31642,N_31961);
xor U33583 (N_33583,N_31847,N_32315);
nor U33584 (N_33584,N_30696,N_31528);
or U33585 (N_33585,N_31166,N_30554);
or U33586 (N_33586,N_31699,N_30751);
and U33587 (N_33587,N_30443,N_32386);
and U33588 (N_33588,N_30796,N_31667);
or U33589 (N_33589,N_31137,N_32109);
and U33590 (N_33590,N_32463,N_30719);
or U33591 (N_33591,N_31900,N_31353);
and U33592 (N_33592,N_30577,N_30278);
and U33593 (N_33593,N_31398,N_32058);
or U33594 (N_33594,N_32418,N_30058);
nand U33595 (N_33595,N_30139,N_32016);
nor U33596 (N_33596,N_30553,N_30539);
or U33597 (N_33597,N_31660,N_31754);
or U33598 (N_33598,N_30360,N_31644);
or U33599 (N_33599,N_30942,N_32137);
and U33600 (N_33600,N_30291,N_31842);
nand U33601 (N_33601,N_32111,N_30779);
nand U33602 (N_33602,N_30184,N_31461);
xnor U33603 (N_33603,N_30097,N_31053);
and U33604 (N_33604,N_31911,N_30798);
xor U33605 (N_33605,N_30836,N_31531);
nor U33606 (N_33606,N_30661,N_30273);
or U33607 (N_33607,N_31881,N_31654);
nor U33608 (N_33608,N_30287,N_31988);
nor U33609 (N_33609,N_30402,N_31140);
or U33610 (N_33610,N_31369,N_31306);
nor U33611 (N_33611,N_30478,N_30088);
xnor U33612 (N_33612,N_30560,N_31069);
nand U33613 (N_33613,N_30911,N_32127);
or U33614 (N_33614,N_30645,N_31018);
xor U33615 (N_33615,N_31097,N_30361);
and U33616 (N_33616,N_32323,N_30526);
and U33617 (N_33617,N_30681,N_30771);
or U33618 (N_33618,N_32038,N_32327);
nor U33619 (N_33619,N_30675,N_31733);
xor U33620 (N_33620,N_31035,N_30340);
nand U33621 (N_33621,N_31984,N_31345);
xnor U33622 (N_33622,N_31592,N_32354);
nand U33623 (N_33623,N_31516,N_30052);
nand U33624 (N_33624,N_30658,N_31384);
xnor U33625 (N_33625,N_31099,N_31438);
nand U33626 (N_33626,N_31278,N_30181);
xor U33627 (N_33627,N_31947,N_31544);
or U33628 (N_33628,N_30896,N_30300);
and U33629 (N_33629,N_31966,N_31780);
xnor U33630 (N_33630,N_32066,N_32259);
xnor U33631 (N_33631,N_30065,N_31668);
nor U33632 (N_33632,N_31055,N_31470);
nor U33633 (N_33633,N_31566,N_30838);
or U33634 (N_33634,N_31008,N_31722);
xor U33635 (N_33635,N_32245,N_30704);
nor U33636 (N_33636,N_32266,N_32322);
or U33637 (N_33637,N_32151,N_30797);
nand U33638 (N_33638,N_32260,N_30823);
or U33639 (N_33639,N_30848,N_30078);
nand U33640 (N_33640,N_30431,N_32268);
xnor U33641 (N_33641,N_30335,N_31503);
or U33642 (N_33642,N_31716,N_32478);
xnor U33643 (N_33643,N_31023,N_31441);
nor U33644 (N_33644,N_32340,N_30113);
and U33645 (N_33645,N_30008,N_31370);
nand U33646 (N_33646,N_32384,N_30155);
xor U33647 (N_33647,N_32144,N_31190);
nor U33648 (N_33648,N_30403,N_30176);
nand U33649 (N_33649,N_32207,N_30125);
and U33650 (N_33650,N_31458,N_31084);
nand U33651 (N_33651,N_32188,N_30028);
xnor U33652 (N_33652,N_30657,N_30785);
or U33653 (N_33653,N_31466,N_30007);
and U33654 (N_33654,N_30872,N_30716);
and U33655 (N_33655,N_30910,N_30373);
xnor U33656 (N_33656,N_31764,N_31941);
or U33657 (N_33657,N_31840,N_31169);
and U33658 (N_33658,N_31991,N_30572);
or U33659 (N_33659,N_31633,N_30215);
xor U33660 (N_33660,N_31124,N_30988);
and U33661 (N_33661,N_30445,N_32159);
nor U33662 (N_33662,N_31298,N_31499);
nor U33663 (N_33663,N_31538,N_30639);
nor U33664 (N_33664,N_31846,N_30451);
or U33665 (N_33665,N_31010,N_31133);
or U33666 (N_33666,N_30753,N_32099);
xnor U33667 (N_33667,N_30032,N_30457);
nor U33668 (N_33668,N_32241,N_30210);
nor U33669 (N_33669,N_32375,N_32040);
and U33670 (N_33670,N_30586,N_31397);
xnor U33671 (N_33671,N_31159,N_31826);
xor U33672 (N_33672,N_32200,N_30230);
nor U33673 (N_33673,N_30231,N_32471);
nor U33674 (N_33674,N_31885,N_31950);
nand U33675 (N_33675,N_30415,N_32004);
xor U33676 (N_33676,N_32253,N_32388);
nor U33677 (N_33677,N_32134,N_30352);
or U33678 (N_33678,N_31580,N_32359);
nand U33679 (N_33679,N_31272,N_30275);
xor U33680 (N_33680,N_31671,N_31799);
and U33681 (N_33681,N_31788,N_30608);
nand U33682 (N_33682,N_32337,N_30959);
nand U33683 (N_33683,N_31235,N_30578);
nor U33684 (N_33684,N_31508,N_32035);
and U33685 (N_33685,N_31692,N_30279);
nor U33686 (N_33686,N_30860,N_30226);
and U33687 (N_33687,N_30405,N_30316);
xor U33688 (N_33688,N_30332,N_31131);
nor U33689 (N_33689,N_32350,N_31614);
and U33690 (N_33690,N_31968,N_30584);
and U33691 (N_33691,N_32242,N_31057);
nand U33692 (N_33692,N_31705,N_30839);
or U33693 (N_33693,N_31505,N_32311);
xor U33694 (N_33694,N_32320,N_32071);
and U33695 (N_33695,N_31199,N_30746);
and U33696 (N_33696,N_30378,N_31033);
or U33697 (N_33697,N_30863,N_32468);
and U33698 (N_33698,N_31926,N_30633);
and U33699 (N_33699,N_31862,N_32403);
xor U33700 (N_33700,N_30239,N_31210);
nand U33701 (N_33701,N_31726,N_30900);
and U33702 (N_33702,N_32101,N_30562);
xnor U33703 (N_33703,N_31901,N_31882);
xnor U33704 (N_33704,N_30285,N_31150);
nor U33705 (N_33705,N_32041,N_30026);
nand U33706 (N_33706,N_30049,N_31365);
nor U33707 (N_33707,N_32124,N_31967);
xor U33708 (N_33708,N_32229,N_32263);
and U33709 (N_33709,N_31734,N_31605);
nor U33710 (N_33710,N_31608,N_31127);
nand U33711 (N_33711,N_31337,N_31048);
or U33712 (N_33712,N_32466,N_31254);
xor U33713 (N_33713,N_31063,N_30229);
nand U33714 (N_33714,N_30066,N_30604);
nand U33715 (N_33715,N_31107,N_30688);
nor U33716 (N_33716,N_30311,N_31334);
nor U33717 (N_33717,N_30814,N_31910);
nor U33718 (N_33718,N_31103,N_31368);
and U33719 (N_33719,N_30204,N_30029);
or U33720 (N_33720,N_31003,N_30121);
or U33721 (N_33721,N_30142,N_32232);
and U33722 (N_33722,N_31971,N_31792);
nor U33723 (N_33723,N_31038,N_31394);
xor U33724 (N_33724,N_30799,N_31304);
or U33725 (N_33725,N_31999,N_30491);
nand U33726 (N_33726,N_31992,N_31844);
or U33727 (N_33727,N_32334,N_30106);
nor U33728 (N_33728,N_30651,N_31100);
nor U33729 (N_33729,N_31869,N_32348);
nand U33730 (N_33730,N_31378,N_30987);
xor U33731 (N_33731,N_32172,N_30441);
and U33732 (N_33732,N_30873,N_30116);
nand U33733 (N_33733,N_30249,N_31252);
or U33734 (N_33734,N_30259,N_30616);
nand U33735 (N_33735,N_32394,N_32114);
nor U33736 (N_33736,N_31674,N_30859);
nor U33737 (N_33737,N_32414,N_30740);
or U33738 (N_33738,N_31339,N_32419);
nand U33739 (N_33739,N_30038,N_30151);
and U33740 (N_33740,N_30144,N_30434);
xnor U33741 (N_33741,N_31031,N_31738);
or U33742 (N_33742,N_31451,N_30384);
and U33743 (N_33743,N_30321,N_31071);
or U33744 (N_33744,N_32070,N_30700);
xor U33745 (N_33745,N_32438,N_31310);
xor U33746 (N_33746,N_31652,N_31419);
nor U33747 (N_33747,N_30995,N_31361);
xor U33748 (N_33748,N_31194,N_30565);
nor U33749 (N_33749,N_31571,N_32427);
nand U33750 (N_33750,N_32378,N_30706);
and U33751 (N_33751,N_30336,N_31986);
xnor U33752 (N_33752,N_32273,N_31618);
and U33753 (N_33753,N_31843,N_30715);
and U33754 (N_33754,N_30829,N_31964);
or U33755 (N_33755,N_32216,N_31503);
and U33756 (N_33756,N_30863,N_30145);
xnor U33757 (N_33757,N_30713,N_31286);
nand U33758 (N_33758,N_31853,N_30482);
or U33759 (N_33759,N_30439,N_31932);
or U33760 (N_33760,N_31215,N_30867);
and U33761 (N_33761,N_31577,N_31229);
xor U33762 (N_33762,N_31669,N_32091);
or U33763 (N_33763,N_30591,N_31148);
nand U33764 (N_33764,N_30284,N_30505);
nor U33765 (N_33765,N_31238,N_32140);
and U33766 (N_33766,N_32118,N_32062);
xnor U33767 (N_33767,N_31363,N_31493);
or U33768 (N_33768,N_31519,N_30589);
nor U33769 (N_33769,N_31854,N_30175);
or U33770 (N_33770,N_30618,N_31993);
or U33771 (N_33771,N_31846,N_30728);
nor U33772 (N_33772,N_32306,N_30375);
and U33773 (N_33773,N_31781,N_30014);
or U33774 (N_33774,N_31131,N_30385);
and U33775 (N_33775,N_31961,N_31097);
nand U33776 (N_33776,N_31910,N_30151);
or U33777 (N_33777,N_31775,N_30336);
nand U33778 (N_33778,N_32467,N_31913);
nand U33779 (N_33779,N_31861,N_30831);
nor U33780 (N_33780,N_31343,N_31250);
and U33781 (N_33781,N_31304,N_31939);
and U33782 (N_33782,N_30382,N_31604);
xor U33783 (N_33783,N_32102,N_31388);
nor U33784 (N_33784,N_30189,N_31756);
nand U33785 (N_33785,N_32271,N_30431);
xor U33786 (N_33786,N_31339,N_31551);
or U33787 (N_33787,N_31333,N_30444);
nand U33788 (N_33788,N_31310,N_31540);
nor U33789 (N_33789,N_30076,N_31460);
nand U33790 (N_33790,N_30843,N_31716);
nor U33791 (N_33791,N_31364,N_30922);
nor U33792 (N_33792,N_32374,N_30784);
xnor U33793 (N_33793,N_31093,N_31278);
nor U33794 (N_33794,N_31411,N_31105);
nor U33795 (N_33795,N_32225,N_30906);
xor U33796 (N_33796,N_31893,N_31821);
xnor U33797 (N_33797,N_30068,N_31344);
and U33798 (N_33798,N_30700,N_31937);
and U33799 (N_33799,N_30905,N_32060);
and U33800 (N_33800,N_32208,N_30125);
xor U33801 (N_33801,N_32102,N_30123);
nor U33802 (N_33802,N_30558,N_30583);
and U33803 (N_33803,N_32077,N_30463);
nor U33804 (N_33804,N_31111,N_30499);
or U33805 (N_33805,N_30106,N_30724);
and U33806 (N_33806,N_31868,N_30176);
and U33807 (N_33807,N_30910,N_32265);
and U33808 (N_33808,N_32150,N_31942);
xor U33809 (N_33809,N_30255,N_30870);
xor U33810 (N_33810,N_30529,N_30919);
nor U33811 (N_33811,N_31118,N_31204);
xor U33812 (N_33812,N_30591,N_32269);
and U33813 (N_33813,N_31812,N_30318);
nand U33814 (N_33814,N_31053,N_31972);
xor U33815 (N_33815,N_32102,N_31092);
xnor U33816 (N_33816,N_30120,N_31120);
or U33817 (N_33817,N_32034,N_31315);
or U33818 (N_33818,N_31538,N_32148);
nand U33819 (N_33819,N_30507,N_30608);
or U33820 (N_33820,N_31684,N_31014);
nor U33821 (N_33821,N_32113,N_30398);
and U33822 (N_33822,N_31531,N_32179);
nand U33823 (N_33823,N_30829,N_31368);
nor U33824 (N_33824,N_31454,N_31451);
xor U33825 (N_33825,N_30781,N_31326);
xnor U33826 (N_33826,N_30534,N_32021);
nor U33827 (N_33827,N_31744,N_32371);
and U33828 (N_33828,N_30010,N_31002);
or U33829 (N_33829,N_31624,N_30663);
and U33830 (N_33830,N_31198,N_31140);
and U33831 (N_33831,N_31037,N_31330);
nand U33832 (N_33832,N_30568,N_32434);
or U33833 (N_33833,N_31174,N_30296);
and U33834 (N_33834,N_32257,N_32319);
and U33835 (N_33835,N_31696,N_30433);
nor U33836 (N_33836,N_30565,N_30166);
nand U33837 (N_33837,N_30981,N_30640);
nand U33838 (N_33838,N_31856,N_30286);
nand U33839 (N_33839,N_30935,N_32312);
or U33840 (N_33840,N_31801,N_31874);
and U33841 (N_33841,N_32338,N_30170);
or U33842 (N_33842,N_31879,N_32050);
nand U33843 (N_33843,N_31808,N_31862);
nand U33844 (N_33844,N_31887,N_30200);
nor U33845 (N_33845,N_30734,N_32396);
nand U33846 (N_33846,N_30954,N_31782);
nand U33847 (N_33847,N_31652,N_30128);
nor U33848 (N_33848,N_30363,N_31732);
and U33849 (N_33849,N_31483,N_30912);
nor U33850 (N_33850,N_32318,N_32177);
xor U33851 (N_33851,N_31552,N_31353);
and U33852 (N_33852,N_30983,N_31118);
nand U33853 (N_33853,N_30605,N_30193);
nor U33854 (N_33854,N_31055,N_31269);
xnor U33855 (N_33855,N_30702,N_31471);
or U33856 (N_33856,N_31808,N_32385);
or U33857 (N_33857,N_31732,N_30020);
nor U33858 (N_33858,N_32490,N_30177);
and U33859 (N_33859,N_30370,N_32355);
xnor U33860 (N_33860,N_30561,N_31925);
and U33861 (N_33861,N_31181,N_32270);
xnor U33862 (N_33862,N_30167,N_30460);
and U33863 (N_33863,N_31311,N_30665);
xnor U33864 (N_33864,N_32389,N_31500);
and U33865 (N_33865,N_31053,N_30721);
xnor U33866 (N_33866,N_30111,N_30193);
nand U33867 (N_33867,N_32163,N_30551);
or U33868 (N_33868,N_32343,N_31312);
xnor U33869 (N_33869,N_32057,N_31589);
xor U33870 (N_33870,N_30227,N_30147);
nor U33871 (N_33871,N_32057,N_31656);
xor U33872 (N_33872,N_30148,N_31962);
xnor U33873 (N_33873,N_30125,N_30599);
nor U33874 (N_33874,N_30280,N_31564);
nand U33875 (N_33875,N_31846,N_31464);
and U33876 (N_33876,N_30789,N_30755);
or U33877 (N_33877,N_30083,N_31343);
nand U33878 (N_33878,N_30121,N_30490);
xor U33879 (N_33879,N_30940,N_30029);
or U33880 (N_33880,N_32221,N_30988);
nand U33881 (N_33881,N_32036,N_31486);
or U33882 (N_33882,N_30700,N_30991);
nor U33883 (N_33883,N_31911,N_30080);
xnor U33884 (N_33884,N_32330,N_32295);
xnor U33885 (N_33885,N_30099,N_30913);
nor U33886 (N_33886,N_30029,N_30042);
or U33887 (N_33887,N_30510,N_31020);
xnor U33888 (N_33888,N_30611,N_32378);
nand U33889 (N_33889,N_31626,N_32438);
and U33890 (N_33890,N_30541,N_31073);
xor U33891 (N_33891,N_31206,N_32374);
nand U33892 (N_33892,N_30104,N_31806);
nand U33893 (N_33893,N_31945,N_30643);
xnor U33894 (N_33894,N_32366,N_32075);
nor U33895 (N_33895,N_30980,N_30633);
or U33896 (N_33896,N_30965,N_31000);
or U33897 (N_33897,N_30727,N_31110);
xor U33898 (N_33898,N_31850,N_31735);
nor U33899 (N_33899,N_32177,N_30118);
nand U33900 (N_33900,N_30164,N_31556);
xor U33901 (N_33901,N_30396,N_31182);
xnor U33902 (N_33902,N_31789,N_30029);
xor U33903 (N_33903,N_30532,N_30595);
nor U33904 (N_33904,N_31274,N_31020);
nor U33905 (N_33905,N_32109,N_31894);
and U33906 (N_33906,N_30323,N_31855);
or U33907 (N_33907,N_32001,N_32333);
nor U33908 (N_33908,N_32171,N_31611);
xor U33909 (N_33909,N_31210,N_30352);
and U33910 (N_33910,N_32135,N_31202);
and U33911 (N_33911,N_30716,N_31418);
or U33912 (N_33912,N_30185,N_31210);
and U33913 (N_33913,N_31611,N_32371);
xor U33914 (N_33914,N_30973,N_32123);
or U33915 (N_33915,N_32283,N_31492);
or U33916 (N_33916,N_31299,N_31973);
nor U33917 (N_33917,N_31258,N_30602);
or U33918 (N_33918,N_31915,N_30523);
and U33919 (N_33919,N_30004,N_30985);
nand U33920 (N_33920,N_30011,N_31024);
nand U33921 (N_33921,N_30847,N_30482);
nand U33922 (N_33922,N_30076,N_31563);
xor U33923 (N_33923,N_31657,N_30827);
nor U33924 (N_33924,N_30621,N_31038);
nor U33925 (N_33925,N_32258,N_31250);
and U33926 (N_33926,N_32095,N_31120);
nand U33927 (N_33927,N_30031,N_31243);
nand U33928 (N_33928,N_30498,N_30523);
or U33929 (N_33929,N_31587,N_31610);
and U33930 (N_33930,N_30851,N_30531);
xor U33931 (N_33931,N_30541,N_30759);
and U33932 (N_33932,N_30853,N_31065);
xnor U33933 (N_33933,N_30393,N_30728);
xnor U33934 (N_33934,N_30231,N_31690);
or U33935 (N_33935,N_31417,N_30261);
xnor U33936 (N_33936,N_31176,N_30227);
xnor U33937 (N_33937,N_32088,N_31041);
xor U33938 (N_33938,N_30879,N_31924);
and U33939 (N_33939,N_30465,N_31211);
and U33940 (N_33940,N_31682,N_30822);
xnor U33941 (N_33941,N_30901,N_31585);
nor U33942 (N_33942,N_31302,N_32308);
nor U33943 (N_33943,N_32269,N_31389);
xor U33944 (N_33944,N_31924,N_30255);
nand U33945 (N_33945,N_32471,N_30225);
xor U33946 (N_33946,N_31788,N_30354);
nand U33947 (N_33947,N_32369,N_31044);
xor U33948 (N_33948,N_30325,N_32471);
and U33949 (N_33949,N_30620,N_31368);
and U33950 (N_33950,N_31561,N_30426);
or U33951 (N_33951,N_30561,N_32264);
nor U33952 (N_33952,N_32484,N_30271);
or U33953 (N_33953,N_31581,N_30182);
nor U33954 (N_33954,N_30205,N_30280);
and U33955 (N_33955,N_31543,N_31702);
or U33956 (N_33956,N_31060,N_31976);
or U33957 (N_33957,N_31811,N_31499);
nor U33958 (N_33958,N_30152,N_30978);
and U33959 (N_33959,N_30853,N_31789);
and U33960 (N_33960,N_32032,N_32464);
and U33961 (N_33961,N_30556,N_31317);
and U33962 (N_33962,N_32457,N_32174);
xor U33963 (N_33963,N_32245,N_30910);
nor U33964 (N_33964,N_30598,N_31644);
xnor U33965 (N_33965,N_32443,N_30022);
nand U33966 (N_33966,N_31704,N_31676);
and U33967 (N_33967,N_31412,N_32314);
or U33968 (N_33968,N_31391,N_30699);
or U33969 (N_33969,N_32052,N_31392);
nor U33970 (N_33970,N_30418,N_31205);
nor U33971 (N_33971,N_31218,N_31888);
xor U33972 (N_33972,N_30105,N_32269);
and U33973 (N_33973,N_31147,N_32256);
and U33974 (N_33974,N_30244,N_30553);
nor U33975 (N_33975,N_32491,N_30840);
or U33976 (N_33976,N_32118,N_30561);
nor U33977 (N_33977,N_31007,N_30062);
or U33978 (N_33978,N_30522,N_31709);
nand U33979 (N_33979,N_30392,N_30517);
xor U33980 (N_33980,N_30798,N_30071);
nand U33981 (N_33981,N_32200,N_31195);
or U33982 (N_33982,N_31084,N_30581);
xor U33983 (N_33983,N_30872,N_30100);
or U33984 (N_33984,N_30119,N_30442);
nor U33985 (N_33985,N_30188,N_32341);
and U33986 (N_33986,N_30395,N_31351);
or U33987 (N_33987,N_31712,N_30474);
and U33988 (N_33988,N_30451,N_30802);
nor U33989 (N_33989,N_31840,N_30350);
xor U33990 (N_33990,N_32027,N_32460);
xnor U33991 (N_33991,N_30924,N_30671);
nand U33992 (N_33992,N_31475,N_31473);
or U33993 (N_33993,N_31385,N_30090);
xnor U33994 (N_33994,N_31543,N_30053);
nor U33995 (N_33995,N_30470,N_32141);
nor U33996 (N_33996,N_31431,N_31442);
nor U33997 (N_33997,N_31792,N_31475);
or U33998 (N_33998,N_30843,N_31358);
xor U33999 (N_33999,N_32264,N_30927);
nor U34000 (N_34000,N_32253,N_31905);
or U34001 (N_34001,N_31341,N_30584);
or U34002 (N_34002,N_30916,N_30343);
or U34003 (N_34003,N_30840,N_31401);
nand U34004 (N_34004,N_32390,N_30554);
or U34005 (N_34005,N_31443,N_30488);
or U34006 (N_34006,N_30536,N_32434);
nor U34007 (N_34007,N_31058,N_30544);
and U34008 (N_34008,N_31051,N_31164);
xnor U34009 (N_34009,N_30200,N_30085);
or U34010 (N_34010,N_30110,N_30220);
nor U34011 (N_34011,N_30470,N_30047);
nand U34012 (N_34012,N_31901,N_31318);
nor U34013 (N_34013,N_31208,N_31932);
and U34014 (N_34014,N_31121,N_31667);
or U34015 (N_34015,N_30560,N_30051);
nor U34016 (N_34016,N_31885,N_31694);
nor U34017 (N_34017,N_31799,N_32072);
or U34018 (N_34018,N_32093,N_31666);
and U34019 (N_34019,N_31454,N_30300);
nand U34020 (N_34020,N_32390,N_32089);
xnor U34021 (N_34021,N_30958,N_30171);
or U34022 (N_34022,N_31009,N_31764);
or U34023 (N_34023,N_31420,N_31098);
nand U34024 (N_34024,N_32334,N_31844);
and U34025 (N_34025,N_31679,N_30623);
or U34026 (N_34026,N_30398,N_31847);
or U34027 (N_34027,N_31189,N_30161);
and U34028 (N_34028,N_32018,N_32032);
xnor U34029 (N_34029,N_32375,N_31838);
nor U34030 (N_34030,N_30404,N_31139);
nand U34031 (N_34031,N_31878,N_30981);
nor U34032 (N_34032,N_30720,N_30898);
and U34033 (N_34033,N_32228,N_31329);
or U34034 (N_34034,N_30908,N_31914);
or U34035 (N_34035,N_32049,N_31867);
nand U34036 (N_34036,N_30763,N_31420);
nor U34037 (N_34037,N_31865,N_31736);
nor U34038 (N_34038,N_32206,N_31493);
xor U34039 (N_34039,N_31357,N_31687);
and U34040 (N_34040,N_30012,N_31776);
xnor U34041 (N_34041,N_31239,N_32300);
or U34042 (N_34042,N_30893,N_31611);
and U34043 (N_34043,N_30861,N_30404);
nand U34044 (N_34044,N_30747,N_31724);
xor U34045 (N_34045,N_30497,N_30799);
nor U34046 (N_34046,N_31334,N_31266);
or U34047 (N_34047,N_31575,N_32483);
nand U34048 (N_34048,N_31329,N_30992);
and U34049 (N_34049,N_31067,N_32244);
and U34050 (N_34050,N_31802,N_30224);
or U34051 (N_34051,N_30337,N_32106);
or U34052 (N_34052,N_31093,N_31999);
nand U34053 (N_34053,N_31255,N_30694);
or U34054 (N_34054,N_32172,N_30826);
and U34055 (N_34055,N_32469,N_30018);
or U34056 (N_34056,N_30137,N_30663);
xor U34057 (N_34057,N_31014,N_30181);
and U34058 (N_34058,N_31948,N_30376);
or U34059 (N_34059,N_32499,N_30093);
and U34060 (N_34060,N_32460,N_30152);
xor U34061 (N_34061,N_31193,N_32006);
xor U34062 (N_34062,N_30417,N_30881);
xor U34063 (N_34063,N_31759,N_32027);
and U34064 (N_34064,N_30486,N_31761);
or U34065 (N_34065,N_31464,N_30003);
nor U34066 (N_34066,N_30486,N_31176);
and U34067 (N_34067,N_31180,N_31244);
xnor U34068 (N_34068,N_30976,N_30549);
nand U34069 (N_34069,N_32022,N_30399);
xor U34070 (N_34070,N_31708,N_31125);
nor U34071 (N_34071,N_31468,N_30270);
and U34072 (N_34072,N_31072,N_30020);
or U34073 (N_34073,N_31687,N_31143);
nor U34074 (N_34074,N_32465,N_30363);
nand U34075 (N_34075,N_30602,N_31034);
nand U34076 (N_34076,N_32163,N_31973);
or U34077 (N_34077,N_31632,N_30701);
xnor U34078 (N_34078,N_31957,N_30547);
nand U34079 (N_34079,N_30992,N_30155);
or U34080 (N_34080,N_31544,N_31105);
or U34081 (N_34081,N_30745,N_31832);
nor U34082 (N_34082,N_31816,N_31765);
and U34083 (N_34083,N_30807,N_31594);
nand U34084 (N_34084,N_30327,N_31278);
and U34085 (N_34085,N_30553,N_31610);
xnor U34086 (N_34086,N_32350,N_31959);
nor U34087 (N_34087,N_30900,N_30785);
or U34088 (N_34088,N_31332,N_31264);
or U34089 (N_34089,N_31439,N_32378);
nor U34090 (N_34090,N_31914,N_30110);
or U34091 (N_34091,N_31877,N_30578);
or U34092 (N_34092,N_31903,N_31802);
nand U34093 (N_34093,N_30225,N_30624);
nand U34094 (N_34094,N_32309,N_32131);
nand U34095 (N_34095,N_30853,N_31393);
and U34096 (N_34096,N_32266,N_31933);
nor U34097 (N_34097,N_30229,N_30721);
nand U34098 (N_34098,N_31087,N_30397);
xor U34099 (N_34099,N_30711,N_30242);
xnor U34100 (N_34100,N_31915,N_32408);
or U34101 (N_34101,N_31984,N_30981);
xor U34102 (N_34102,N_30240,N_32350);
and U34103 (N_34103,N_30431,N_32284);
xnor U34104 (N_34104,N_30517,N_32328);
xnor U34105 (N_34105,N_31041,N_32086);
or U34106 (N_34106,N_30141,N_31689);
and U34107 (N_34107,N_31989,N_30955);
and U34108 (N_34108,N_30123,N_31441);
and U34109 (N_34109,N_30003,N_31566);
nor U34110 (N_34110,N_31131,N_31915);
nor U34111 (N_34111,N_30792,N_32435);
xor U34112 (N_34112,N_30555,N_32135);
nand U34113 (N_34113,N_30741,N_32136);
xor U34114 (N_34114,N_31570,N_30238);
xnor U34115 (N_34115,N_31749,N_32294);
or U34116 (N_34116,N_31923,N_30835);
nand U34117 (N_34117,N_30714,N_30124);
xnor U34118 (N_34118,N_30001,N_31747);
and U34119 (N_34119,N_30355,N_32227);
xnor U34120 (N_34120,N_30393,N_30356);
and U34121 (N_34121,N_31215,N_32278);
xnor U34122 (N_34122,N_32044,N_30605);
or U34123 (N_34123,N_30985,N_31866);
xor U34124 (N_34124,N_31852,N_31085);
nor U34125 (N_34125,N_31119,N_30936);
and U34126 (N_34126,N_30050,N_30358);
or U34127 (N_34127,N_31982,N_30211);
nand U34128 (N_34128,N_32089,N_32017);
and U34129 (N_34129,N_31330,N_30935);
nor U34130 (N_34130,N_30433,N_32096);
nor U34131 (N_34131,N_30150,N_31369);
xor U34132 (N_34132,N_30996,N_31574);
or U34133 (N_34133,N_31603,N_32439);
and U34134 (N_34134,N_31324,N_31600);
xnor U34135 (N_34135,N_32054,N_31644);
and U34136 (N_34136,N_31648,N_30615);
nand U34137 (N_34137,N_30130,N_30776);
or U34138 (N_34138,N_31675,N_32159);
xnor U34139 (N_34139,N_31635,N_31780);
or U34140 (N_34140,N_31185,N_30931);
and U34141 (N_34141,N_30347,N_31710);
and U34142 (N_34142,N_30305,N_32233);
nor U34143 (N_34143,N_30580,N_30680);
nand U34144 (N_34144,N_31790,N_32481);
xor U34145 (N_34145,N_31434,N_30231);
nand U34146 (N_34146,N_31377,N_31337);
or U34147 (N_34147,N_31367,N_32180);
nor U34148 (N_34148,N_31449,N_32344);
or U34149 (N_34149,N_31555,N_31962);
and U34150 (N_34150,N_31058,N_30032);
or U34151 (N_34151,N_31234,N_31325);
and U34152 (N_34152,N_31311,N_30626);
nand U34153 (N_34153,N_31744,N_30677);
xnor U34154 (N_34154,N_31574,N_30099);
or U34155 (N_34155,N_30888,N_30185);
nor U34156 (N_34156,N_32223,N_30483);
xnor U34157 (N_34157,N_31534,N_31207);
and U34158 (N_34158,N_30859,N_32058);
nor U34159 (N_34159,N_30347,N_31718);
and U34160 (N_34160,N_31624,N_31935);
nor U34161 (N_34161,N_30848,N_30905);
or U34162 (N_34162,N_32127,N_30748);
xnor U34163 (N_34163,N_30135,N_31835);
or U34164 (N_34164,N_30991,N_30251);
nand U34165 (N_34165,N_30850,N_32479);
xor U34166 (N_34166,N_31305,N_30830);
or U34167 (N_34167,N_31433,N_32331);
nand U34168 (N_34168,N_32228,N_31572);
xnor U34169 (N_34169,N_32263,N_30983);
nand U34170 (N_34170,N_31950,N_30809);
nor U34171 (N_34171,N_30014,N_30816);
or U34172 (N_34172,N_32191,N_31448);
and U34173 (N_34173,N_30467,N_32349);
xor U34174 (N_34174,N_31191,N_31327);
nand U34175 (N_34175,N_30669,N_31440);
xor U34176 (N_34176,N_30679,N_31335);
xnor U34177 (N_34177,N_32455,N_32425);
xor U34178 (N_34178,N_32219,N_31581);
nor U34179 (N_34179,N_30190,N_32356);
and U34180 (N_34180,N_32160,N_30862);
and U34181 (N_34181,N_30821,N_30924);
or U34182 (N_34182,N_31431,N_31937);
nand U34183 (N_34183,N_32386,N_30772);
and U34184 (N_34184,N_31768,N_31050);
or U34185 (N_34185,N_32363,N_30267);
nor U34186 (N_34186,N_30153,N_32262);
or U34187 (N_34187,N_32228,N_31911);
or U34188 (N_34188,N_30569,N_32110);
and U34189 (N_34189,N_31169,N_30417);
xnor U34190 (N_34190,N_30544,N_31847);
and U34191 (N_34191,N_31864,N_31838);
nor U34192 (N_34192,N_31388,N_31628);
xor U34193 (N_34193,N_30451,N_31962);
and U34194 (N_34194,N_31753,N_30771);
xnor U34195 (N_34195,N_32341,N_31343);
or U34196 (N_34196,N_30869,N_30331);
or U34197 (N_34197,N_30367,N_31241);
and U34198 (N_34198,N_32032,N_32220);
nand U34199 (N_34199,N_31238,N_32358);
or U34200 (N_34200,N_30593,N_31726);
nor U34201 (N_34201,N_31929,N_31506);
xor U34202 (N_34202,N_30894,N_30994);
and U34203 (N_34203,N_31660,N_32093);
xnor U34204 (N_34204,N_30692,N_31238);
and U34205 (N_34205,N_32373,N_30317);
nor U34206 (N_34206,N_32034,N_32305);
nor U34207 (N_34207,N_30948,N_31282);
and U34208 (N_34208,N_31205,N_30755);
and U34209 (N_34209,N_30709,N_30604);
nand U34210 (N_34210,N_31469,N_31346);
or U34211 (N_34211,N_32207,N_30466);
nand U34212 (N_34212,N_32317,N_30869);
nand U34213 (N_34213,N_30859,N_31736);
or U34214 (N_34214,N_30869,N_31898);
and U34215 (N_34215,N_30244,N_31794);
nand U34216 (N_34216,N_30988,N_31281);
xnor U34217 (N_34217,N_31856,N_31787);
or U34218 (N_34218,N_30129,N_30698);
or U34219 (N_34219,N_30038,N_30842);
xnor U34220 (N_34220,N_31099,N_30936);
xor U34221 (N_34221,N_30754,N_30880);
and U34222 (N_34222,N_32145,N_31650);
nor U34223 (N_34223,N_31208,N_30283);
and U34224 (N_34224,N_30775,N_32179);
nand U34225 (N_34225,N_32262,N_31205);
nand U34226 (N_34226,N_31853,N_32161);
nor U34227 (N_34227,N_30065,N_32455);
xor U34228 (N_34228,N_32087,N_30387);
nor U34229 (N_34229,N_30452,N_32346);
xnor U34230 (N_34230,N_30622,N_30707);
or U34231 (N_34231,N_31055,N_30491);
or U34232 (N_34232,N_30871,N_32086);
xor U34233 (N_34233,N_31852,N_32314);
or U34234 (N_34234,N_31856,N_30750);
and U34235 (N_34235,N_31993,N_30772);
nor U34236 (N_34236,N_30609,N_31894);
nor U34237 (N_34237,N_31532,N_32073);
or U34238 (N_34238,N_31990,N_30741);
nand U34239 (N_34239,N_30990,N_31809);
and U34240 (N_34240,N_30179,N_30747);
xnor U34241 (N_34241,N_32433,N_31209);
xnor U34242 (N_34242,N_30356,N_30276);
xor U34243 (N_34243,N_31248,N_30770);
or U34244 (N_34244,N_30700,N_30261);
or U34245 (N_34245,N_31285,N_31381);
xnor U34246 (N_34246,N_31812,N_30411);
xor U34247 (N_34247,N_30964,N_30380);
and U34248 (N_34248,N_30735,N_30773);
and U34249 (N_34249,N_30717,N_30441);
nand U34250 (N_34250,N_30081,N_30341);
xor U34251 (N_34251,N_30356,N_30646);
nand U34252 (N_34252,N_30107,N_30801);
nand U34253 (N_34253,N_32394,N_31966);
nor U34254 (N_34254,N_30814,N_30848);
and U34255 (N_34255,N_30848,N_31056);
and U34256 (N_34256,N_32301,N_32268);
nand U34257 (N_34257,N_31627,N_32384);
and U34258 (N_34258,N_31289,N_31338);
and U34259 (N_34259,N_31730,N_30927);
nor U34260 (N_34260,N_32417,N_31465);
or U34261 (N_34261,N_31730,N_31338);
or U34262 (N_34262,N_31459,N_30063);
xnor U34263 (N_34263,N_31254,N_30566);
nand U34264 (N_34264,N_32324,N_31547);
or U34265 (N_34265,N_30939,N_32371);
nand U34266 (N_34266,N_30671,N_32313);
xor U34267 (N_34267,N_30248,N_32146);
nor U34268 (N_34268,N_30652,N_31430);
xor U34269 (N_34269,N_31234,N_31263);
or U34270 (N_34270,N_31285,N_31265);
nor U34271 (N_34271,N_31637,N_31927);
or U34272 (N_34272,N_30605,N_32481);
or U34273 (N_34273,N_31567,N_31549);
or U34274 (N_34274,N_31482,N_30114);
xor U34275 (N_34275,N_31811,N_31321);
and U34276 (N_34276,N_30608,N_30128);
xnor U34277 (N_34277,N_30765,N_31778);
or U34278 (N_34278,N_31733,N_31785);
xnor U34279 (N_34279,N_32063,N_30801);
or U34280 (N_34280,N_31822,N_30386);
xnor U34281 (N_34281,N_30894,N_30380);
xnor U34282 (N_34282,N_30450,N_31680);
nand U34283 (N_34283,N_30606,N_31130);
and U34284 (N_34284,N_31213,N_30052);
xor U34285 (N_34285,N_31743,N_31302);
and U34286 (N_34286,N_31458,N_30117);
nor U34287 (N_34287,N_30669,N_30073);
or U34288 (N_34288,N_31870,N_30116);
or U34289 (N_34289,N_30015,N_30660);
or U34290 (N_34290,N_32266,N_31077);
nor U34291 (N_34291,N_30704,N_31418);
nand U34292 (N_34292,N_32074,N_32246);
nor U34293 (N_34293,N_31446,N_30247);
nand U34294 (N_34294,N_31972,N_30205);
and U34295 (N_34295,N_32231,N_30225);
xnor U34296 (N_34296,N_31634,N_30449);
nor U34297 (N_34297,N_30501,N_30023);
nor U34298 (N_34298,N_31091,N_31150);
nor U34299 (N_34299,N_31740,N_31925);
and U34300 (N_34300,N_31259,N_30999);
and U34301 (N_34301,N_30866,N_32103);
nand U34302 (N_34302,N_31373,N_30158);
nor U34303 (N_34303,N_32210,N_31958);
nor U34304 (N_34304,N_30611,N_32354);
or U34305 (N_34305,N_30993,N_30743);
nor U34306 (N_34306,N_31826,N_31912);
nor U34307 (N_34307,N_30417,N_32235);
nor U34308 (N_34308,N_31528,N_30334);
and U34309 (N_34309,N_32458,N_30280);
or U34310 (N_34310,N_31889,N_30947);
or U34311 (N_34311,N_30560,N_30299);
and U34312 (N_34312,N_30190,N_32142);
xor U34313 (N_34313,N_32401,N_30962);
or U34314 (N_34314,N_30544,N_30335);
nand U34315 (N_34315,N_30926,N_30849);
nand U34316 (N_34316,N_31572,N_31085);
nor U34317 (N_34317,N_30762,N_30125);
nor U34318 (N_34318,N_31064,N_30720);
or U34319 (N_34319,N_31853,N_31500);
nor U34320 (N_34320,N_32485,N_30749);
nor U34321 (N_34321,N_30724,N_31007);
xnor U34322 (N_34322,N_32234,N_32366);
xnor U34323 (N_34323,N_31981,N_32182);
xnor U34324 (N_34324,N_31781,N_32362);
nor U34325 (N_34325,N_30948,N_31963);
xnor U34326 (N_34326,N_30013,N_32431);
and U34327 (N_34327,N_32406,N_31574);
and U34328 (N_34328,N_31467,N_32334);
and U34329 (N_34329,N_31520,N_30161);
and U34330 (N_34330,N_31342,N_30869);
xor U34331 (N_34331,N_31907,N_30353);
nor U34332 (N_34332,N_30779,N_31663);
nor U34333 (N_34333,N_30932,N_31435);
and U34334 (N_34334,N_30729,N_30815);
or U34335 (N_34335,N_30669,N_31669);
xnor U34336 (N_34336,N_32194,N_31782);
xor U34337 (N_34337,N_30973,N_32300);
xor U34338 (N_34338,N_32374,N_32234);
nand U34339 (N_34339,N_32254,N_30676);
xor U34340 (N_34340,N_32056,N_31313);
or U34341 (N_34341,N_30773,N_32057);
nand U34342 (N_34342,N_32187,N_31332);
nand U34343 (N_34343,N_32259,N_31042);
and U34344 (N_34344,N_31709,N_32019);
or U34345 (N_34345,N_30601,N_31448);
nand U34346 (N_34346,N_30079,N_30199);
and U34347 (N_34347,N_30922,N_30625);
nor U34348 (N_34348,N_32339,N_31036);
nand U34349 (N_34349,N_30919,N_32087);
or U34350 (N_34350,N_30614,N_31816);
and U34351 (N_34351,N_31502,N_30156);
nor U34352 (N_34352,N_30455,N_32142);
xor U34353 (N_34353,N_30713,N_31281);
xor U34354 (N_34354,N_31682,N_31105);
nor U34355 (N_34355,N_31133,N_31481);
nor U34356 (N_34356,N_30380,N_30841);
and U34357 (N_34357,N_31413,N_30500);
and U34358 (N_34358,N_30062,N_30963);
xnor U34359 (N_34359,N_30679,N_30830);
nand U34360 (N_34360,N_31545,N_32196);
or U34361 (N_34361,N_30178,N_31499);
nor U34362 (N_34362,N_31994,N_32395);
xor U34363 (N_34363,N_31186,N_32386);
nand U34364 (N_34364,N_32401,N_31831);
nor U34365 (N_34365,N_30730,N_31305);
nand U34366 (N_34366,N_30074,N_31366);
nor U34367 (N_34367,N_30288,N_31529);
and U34368 (N_34368,N_30730,N_31323);
or U34369 (N_34369,N_31028,N_30361);
nand U34370 (N_34370,N_30298,N_30808);
or U34371 (N_34371,N_31077,N_31688);
or U34372 (N_34372,N_31884,N_32174);
nor U34373 (N_34373,N_30078,N_31960);
nor U34374 (N_34374,N_31931,N_30844);
nand U34375 (N_34375,N_31456,N_31718);
nand U34376 (N_34376,N_32310,N_31051);
xor U34377 (N_34377,N_30132,N_32245);
xor U34378 (N_34378,N_30773,N_31329);
xor U34379 (N_34379,N_30631,N_31381);
or U34380 (N_34380,N_31312,N_32100);
xnor U34381 (N_34381,N_30485,N_31574);
xor U34382 (N_34382,N_30797,N_31253);
xor U34383 (N_34383,N_32012,N_31170);
nand U34384 (N_34384,N_32163,N_31652);
nand U34385 (N_34385,N_30112,N_31233);
nand U34386 (N_34386,N_31987,N_31719);
nand U34387 (N_34387,N_30238,N_31613);
xnor U34388 (N_34388,N_31312,N_30026);
or U34389 (N_34389,N_31796,N_31907);
nor U34390 (N_34390,N_31881,N_32482);
nor U34391 (N_34391,N_30480,N_31063);
nor U34392 (N_34392,N_30695,N_31273);
nand U34393 (N_34393,N_30697,N_32082);
nor U34394 (N_34394,N_30396,N_31277);
xor U34395 (N_34395,N_31480,N_31130);
or U34396 (N_34396,N_30273,N_31407);
and U34397 (N_34397,N_30080,N_31499);
xnor U34398 (N_34398,N_31491,N_30349);
nor U34399 (N_34399,N_30914,N_32170);
nor U34400 (N_34400,N_30503,N_31040);
nand U34401 (N_34401,N_32180,N_31555);
or U34402 (N_34402,N_31243,N_31287);
xor U34403 (N_34403,N_32060,N_30387);
or U34404 (N_34404,N_30760,N_32352);
xor U34405 (N_34405,N_32416,N_30304);
xor U34406 (N_34406,N_31761,N_30548);
nor U34407 (N_34407,N_31534,N_31614);
nor U34408 (N_34408,N_30243,N_30316);
nor U34409 (N_34409,N_30593,N_31436);
nor U34410 (N_34410,N_32059,N_32258);
or U34411 (N_34411,N_30371,N_31520);
and U34412 (N_34412,N_31666,N_30341);
nor U34413 (N_34413,N_31209,N_30130);
nand U34414 (N_34414,N_30187,N_31192);
or U34415 (N_34415,N_32438,N_30501);
and U34416 (N_34416,N_30502,N_30631);
xor U34417 (N_34417,N_32014,N_31961);
xnor U34418 (N_34418,N_32464,N_31728);
and U34419 (N_34419,N_32240,N_30596);
xor U34420 (N_34420,N_31210,N_30435);
or U34421 (N_34421,N_32172,N_32353);
and U34422 (N_34422,N_31391,N_30222);
nand U34423 (N_34423,N_30531,N_31625);
nand U34424 (N_34424,N_31145,N_30478);
or U34425 (N_34425,N_31819,N_30473);
nand U34426 (N_34426,N_30364,N_31486);
or U34427 (N_34427,N_31972,N_30017);
nand U34428 (N_34428,N_30773,N_31943);
xor U34429 (N_34429,N_31846,N_30850);
or U34430 (N_34430,N_32337,N_30844);
and U34431 (N_34431,N_31683,N_31095);
or U34432 (N_34432,N_31558,N_32265);
or U34433 (N_34433,N_32383,N_31335);
nand U34434 (N_34434,N_30791,N_32099);
nor U34435 (N_34435,N_30478,N_30915);
nand U34436 (N_34436,N_32470,N_30382);
xor U34437 (N_34437,N_31553,N_31588);
xor U34438 (N_34438,N_30711,N_32066);
nand U34439 (N_34439,N_31733,N_30596);
nand U34440 (N_34440,N_31014,N_30304);
nand U34441 (N_34441,N_30962,N_30736);
nand U34442 (N_34442,N_30323,N_30729);
xnor U34443 (N_34443,N_32403,N_30164);
nand U34444 (N_34444,N_31119,N_30883);
xor U34445 (N_34445,N_31733,N_30156);
nor U34446 (N_34446,N_30479,N_30862);
and U34447 (N_34447,N_31375,N_31809);
nor U34448 (N_34448,N_30430,N_31562);
nor U34449 (N_34449,N_32242,N_31486);
or U34450 (N_34450,N_32266,N_31015);
nand U34451 (N_34451,N_32449,N_30543);
nand U34452 (N_34452,N_30715,N_30841);
xor U34453 (N_34453,N_31075,N_30699);
and U34454 (N_34454,N_31094,N_31835);
and U34455 (N_34455,N_30276,N_31179);
or U34456 (N_34456,N_30093,N_32258);
xnor U34457 (N_34457,N_30891,N_32247);
nand U34458 (N_34458,N_32272,N_31221);
nor U34459 (N_34459,N_32331,N_31574);
nor U34460 (N_34460,N_30048,N_31850);
and U34461 (N_34461,N_30585,N_31545);
nor U34462 (N_34462,N_31441,N_31160);
xor U34463 (N_34463,N_30824,N_31464);
and U34464 (N_34464,N_31059,N_31394);
or U34465 (N_34465,N_30805,N_30239);
nand U34466 (N_34466,N_31602,N_31339);
xor U34467 (N_34467,N_31901,N_30768);
nand U34468 (N_34468,N_31712,N_30635);
and U34469 (N_34469,N_30947,N_31321);
xor U34470 (N_34470,N_30194,N_31368);
xnor U34471 (N_34471,N_31511,N_32381);
or U34472 (N_34472,N_32288,N_30047);
xnor U34473 (N_34473,N_30573,N_32496);
and U34474 (N_34474,N_32082,N_30583);
xor U34475 (N_34475,N_30381,N_31378);
nor U34476 (N_34476,N_30369,N_30985);
xnor U34477 (N_34477,N_30766,N_32314);
xnor U34478 (N_34478,N_30325,N_31176);
nand U34479 (N_34479,N_32104,N_30409);
and U34480 (N_34480,N_31804,N_31979);
and U34481 (N_34481,N_32342,N_30132);
xor U34482 (N_34482,N_32196,N_30709);
xor U34483 (N_34483,N_32367,N_30696);
and U34484 (N_34484,N_32108,N_32389);
nand U34485 (N_34485,N_31963,N_31691);
nand U34486 (N_34486,N_30531,N_31759);
nor U34487 (N_34487,N_30524,N_32295);
or U34488 (N_34488,N_32039,N_31622);
and U34489 (N_34489,N_31376,N_30709);
and U34490 (N_34490,N_31801,N_30632);
nor U34491 (N_34491,N_31672,N_31173);
and U34492 (N_34492,N_30364,N_30733);
xor U34493 (N_34493,N_31874,N_31588);
or U34494 (N_34494,N_31934,N_32223);
nand U34495 (N_34495,N_31414,N_31001);
or U34496 (N_34496,N_31584,N_31294);
or U34497 (N_34497,N_31582,N_31610);
or U34498 (N_34498,N_30292,N_31484);
xor U34499 (N_34499,N_32185,N_30719);
nor U34500 (N_34500,N_31758,N_31520);
nand U34501 (N_34501,N_31371,N_31009);
nor U34502 (N_34502,N_30639,N_31629);
xnor U34503 (N_34503,N_30507,N_30497);
nor U34504 (N_34504,N_32354,N_32200);
xor U34505 (N_34505,N_32473,N_32362);
xnor U34506 (N_34506,N_30087,N_31606);
nand U34507 (N_34507,N_30822,N_30237);
xor U34508 (N_34508,N_31173,N_32064);
nor U34509 (N_34509,N_30618,N_31966);
and U34510 (N_34510,N_32238,N_30766);
xnor U34511 (N_34511,N_30032,N_31122);
xor U34512 (N_34512,N_31082,N_31697);
xnor U34513 (N_34513,N_32487,N_31447);
nor U34514 (N_34514,N_32464,N_31886);
or U34515 (N_34515,N_31277,N_32290);
xnor U34516 (N_34516,N_30438,N_30692);
xor U34517 (N_34517,N_31878,N_30916);
nor U34518 (N_34518,N_30412,N_31726);
xnor U34519 (N_34519,N_31239,N_31750);
nand U34520 (N_34520,N_30949,N_32126);
or U34521 (N_34521,N_30198,N_32477);
nand U34522 (N_34522,N_30846,N_32401);
or U34523 (N_34523,N_30252,N_31398);
and U34524 (N_34524,N_31852,N_31270);
or U34525 (N_34525,N_30617,N_31404);
xnor U34526 (N_34526,N_32243,N_31487);
or U34527 (N_34527,N_30945,N_31901);
or U34528 (N_34528,N_31597,N_32335);
nand U34529 (N_34529,N_31641,N_31995);
nand U34530 (N_34530,N_30861,N_30239);
nor U34531 (N_34531,N_30648,N_31811);
xor U34532 (N_34532,N_30210,N_30577);
and U34533 (N_34533,N_31456,N_32103);
xor U34534 (N_34534,N_30563,N_30929);
or U34535 (N_34535,N_32037,N_32368);
nor U34536 (N_34536,N_31344,N_30627);
xnor U34537 (N_34537,N_31464,N_30760);
xnor U34538 (N_34538,N_30068,N_32043);
or U34539 (N_34539,N_31078,N_30898);
xnor U34540 (N_34540,N_31155,N_31365);
nor U34541 (N_34541,N_31472,N_30057);
nor U34542 (N_34542,N_31787,N_30571);
nand U34543 (N_34543,N_30241,N_31971);
nand U34544 (N_34544,N_31630,N_30071);
nand U34545 (N_34545,N_31679,N_30951);
or U34546 (N_34546,N_31014,N_32153);
nor U34547 (N_34547,N_31625,N_31015);
or U34548 (N_34548,N_30246,N_32129);
and U34549 (N_34549,N_31367,N_32214);
nand U34550 (N_34550,N_31904,N_31328);
or U34551 (N_34551,N_30279,N_30165);
nor U34552 (N_34552,N_30120,N_30743);
xnor U34553 (N_34553,N_31392,N_32306);
or U34554 (N_34554,N_30158,N_31878);
or U34555 (N_34555,N_30506,N_30832);
nor U34556 (N_34556,N_31781,N_31200);
and U34557 (N_34557,N_31010,N_32353);
or U34558 (N_34558,N_31326,N_30298);
and U34559 (N_34559,N_30313,N_31171);
and U34560 (N_34560,N_31917,N_31707);
or U34561 (N_34561,N_30299,N_30342);
xor U34562 (N_34562,N_30178,N_32120);
and U34563 (N_34563,N_30102,N_31197);
nand U34564 (N_34564,N_31020,N_30716);
or U34565 (N_34565,N_31301,N_31661);
or U34566 (N_34566,N_31231,N_30359);
nand U34567 (N_34567,N_32113,N_32258);
nand U34568 (N_34568,N_31481,N_32109);
or U34569 (N_34569,N_30865,N_31062);
nor U34570 (N_34570,N_31038,N_30929);
nand U34571 (N_34571,N_30211,N_30371);
nand U34572 (N_34572,N_32394,N_31414);
or U34573 (N_34573,N_32294,N_32452);
nand U34574 (N_34574,N_30321,N_31453);
xor U34575 (N_34575,N_30372,N_31887);
nand U34576 (N_34576,N_32298,N_31046);
xor U34577 (N_34577,N_31733,N_32358);
and U34578 (N_34578,N_31685,N_30266);
nor U34579 (N_34579,N_30202,N_30862);
xor U34580 (N_34580,N_32020,N_30778);
nor U34581 (N_34581,N_31136,N_30925);
nand U34582 (N_34582,N_31854,N_32378);
nand U34583 (N_34583,N_30259,N_30009);
nor U34584 (N_34584,N_30026,N_30380);
xor U34585 (N_34585,N_31920,N_30269);
xor U34586 (N_34586,N_30294,N_30551);
or U34587 (N_34587,N_31482,N_30203);
and U34588 (N_34588,N_30485,N_31895);
or U34589 (N_34589,N_30752,N_32327);
xor U34590 (N_34590,N_32065,N_30614);
xor U34591 (N_34591,N_32478,N_30902);
nand U34592 (N_34592,N_32004,N_30047);
and U34593 (N_34593,N_31280,N_32133);
and U34594 (N_34594,N_31818,N_32076);
nor U34595 (N_34595,N_31142,N_30210);
nor U34596 (N_34596,N_31019,N_31011);
xor U34597 (N_34597,N_30013,N_30339);
nand U34598 (N_34598,N_31548,N_31804);
xnor U34599 (N_34599,N_30823,N_30439);
nor U34600 (N_34600,N_30887,N_30953);
nor U34601 (N_34601,N_30710,N_31575);
nor U34602 (N_34602,N_30485,N_30495);
xnor U34603 (N_34603,N_31649,N_31369);
nor U34604 (N_34604,N_31626,N_30856);
or U34605 (N_34605,N_32367,N_31074);
and U34606 (N_34606,N_30362,N_30690);
nor U34607 (N_34607,N_31663,N_30527);
or U34608 (N_34608,N_32430,N_30068);
or U34609 (N_34609,N_30923,N_30701);
nor U34610 (N_34610,N_32074,N_32148);
nor U34611 (N_34611,N_32231,N_30085);
and U34612 (N_34612,N_31907,N_30445);
nand U34613 (N_34613,N_30885,N_30225);
or U34614 (N_34614,N_31845,N_31753);
or U34615 (N_34615,N_30034,N_30851);
xnor U34616 (N_34616,N_30518,N_31529);
xnor U34617 (N_34617,N_32270,N_31334);
nand U34618 (N_34618,N_31847,N_30838);
nand U34619 (N_34619,N_31022,N_31297);
nor U34620 (N_34620,N_31411,N_31669);
nand U34621 (N_34621,N_30239,N_30388);
xnor U34622 (N_34622,N_32473,N_30349);
nand U34623 (N_34623,N_30842,N_31318);
or U34624 (N_34624,N_31877,N_32384);
nand U34625 (N_34625,N_31625,N_30609);
xnor U34626 (N_34626,N_30454,N_31769);
xor U34627 (N_34627,N_30794,N_32335);
or U34628 (N_34628,N_31756,N_31387);
or U34629 (N_34629,N_32434,N_30793);
nor U34630 (N_34630,N_32207,N_30309);
xnor U34631 (N_34631,N_31896,N_32292);
nand U34632 (N_34632,N_30642,N_32149);
nor U34633 (N_34633,N_31492,N_31437);
and U34634 (N_34634,N_31303,N_31968);
nor U34635 (N_34635,N_31972,N_30223);
and U34636 (N_34636,N_30299,N_30851);
or U34637 (N_34637,N_30261,N_31260);
and U34638 (N_34638,N_31887,N_31094);
nor U34639 (N_34639,N_32065,N_30513);
or U34640 (N_34640,N_30603,N_31126);
xor U34641 (N_34641,N_30434,N_30219);
or U34642 (N_34642,N_31458,N_31709);
xnor U34643 (N_34643,N_32481,N_30250);
xnor U34644 (N_34644,N_30036,N_32231);
xnor U34645 (N_34645,N_31775,N_32232);
nand U34646 (N_34646,N_32013,N_30065);
nor U34647 (N_34647,N_31896,N_31849);
and U34648 (N_34648,N_31583,N_32457);
nor U34649 (N_34649,N_31584,N_32470);
nand U34650 (N_34650,N_31875,N_30732);
or U34651 (N_34651,N_30092,N_30624);
nor U34652 (N_34652,N_30078,N_30446);
nand U34653 (N_34653,N_31660,N_30103);
xnor U34654 (N_34654,N_32150,N_30002);
xor U34655 (N_34655,N_30789,N_31994);
nor U34656 (N_34656,N_30658,N_31712);
nand U34657 (N_34657,N_30738,N_31716);
nand U34658 (N_34658,N_32115,N_32043);
xnor U34659 (N_34659,N_30943,N_30376);
or U34660 (N_34660,N_31217,N_30908);
nand U34661 (N_34661,N_31446,N_30499);
nor U34662 (N_34662,N_32291,N_31166);
and U34663 (N_34663,N_30216,N_31005);
nand U34664 (N_34664,N_30635,N_32259);
nand U34665 (N_34665,N_31282,N_31583);
nor U34666 (N_34666,N_30513,N_30361);
and U34667 (N_34667,N_30004,N_30186);
or U34668 (N_34668,N_30238,N_30497);
and U34669 (N_34669,N_31350,N_31193);
xor U34670 (N_34670,N_31314,N_32378);
xnor U34671 (N_34671,N_32202,N_30408);
nand U34672 (N_34672,N_30399,N_30456);
and U34673 (N_34673,N_32195,N_31555);
or U34674 (N_34674,N_32139,N_30484);
and U34675 (N_34675,N_30964,N_31381);
or U34676 (N_34676,N_30709,N_30251);
xnor U34677 (N_34677,N_30187,N_32447);
xor U34678 (N_34678,N_30829,N_30355);
nor U34679 (N_34679,N_32162,N_30988);
nor U34680 (N_34680,N_30425,N_30807);
or U34681 (N_34681,N_30761,N_30337);
and U34682 (N_34682,N_31513,N_30919);
xor U34683 (N_34683,N_32160,N_31633);
and U34684 (N_34684,N_31331,N_32077);
and U34685 (N_34685,N_30621,N_31404);
and U34686 (N_34686,N_31016,N_32472);
or U34687 (N_34687,N_30358,N_31526);
and U34688 (N_34688,N_31264,N_31086);
or U34689 (N_34689,N_31026,N_32338);
nand U34690 (N_34690,N_32250,N_31721);
and U34691 (N_34691,N_32225,N_30477);
nand U34692 (N_34692,N_30703,N_30816);
and U34693 (N_34693,N_31339,N_32046);
and U34694 (N_34694,N_31652,N_31812);
nand U34695 (N_34695,N_30751,N_30112);
or U34696 (N_34696,N_31594,N_31285);
nor U34697 (N_34697,N_30989,N_32440);
xor U34698 (N_34698,N_30194,N_30264);
nand U34699 (N_34699,N_31300,N_32168);
xor U34700 (N_34700,N_31908,N_31560);
and U34701 (N_34701,N_30042,N_30497);
or U34702 (N_34702,N_30283,N_32046);
xor U34703 (N_34703,N_31368,N_32280);
and U34704 (N_34704,N_31710,N_31133);
xnor U34705 (N_34705,N_30365,N_30430);
nor U34706 (N_34706,N_32239,N_32376);
and U34707 (N_34707,N_30247,N_30804);
nand U34708 (N_34708,N_30034,N_30626);
nor U34709 (N_34709,N_30860,N_31636);
xnor U34710 (N_34710,N_31556,N_30322);
and U34711 (N_34711,N_31065,N_31555);
or U34712 (N_34712,N_30856,N_30011);
and U34713 (N_34713,N_31796,N_30042);
xor U34714 (N_34714,N_30396,N_30302);
nand U34715 (N_34715,N_32363,N_30749);
and U34716 (N_34716,N_30061,N_30513);
nand U34717 (N_34717,N_30751,N_31024);
or U34718 (N_34718,N_32375,N_30103);
or U34719 (N_34719,N_30683,N_30394);
xor U34720 (N_34720,N_32367,N_32427);
or U34721 (N_34721,N_30834,N_31562);
xor U34722 (N_34722,N_30071,N_31908);
nand U34723 (N_34723,N_31978,N_30445);
nor U34724 (N_34724,N_32270,N_31616);
or U34725 (N_34725,N_31601,N_32207);
and U34726 (N_34726,N_31229,N_31138);
nor U34727 (N_34727,N_31583,N_31754);
xor U34728 (N_34728,N_31601,N_32025);
nor U34729 (N_34729,N_30627,N_30068);
xnor U34730 (N_34730,N_31545,N_30336);
xnor U34731 (N_34731,N_30511,N_31909);
nor U34732 (N_34732,N_32210,N_30783);
or U34733 (N_34733,N_30062,N_31203);
and U34734 (N_34734,N_30246,N_31828);
nor U34735 (N_34735,N_31926,N_30038);
and U34736 (N_34736,N_31740,N_31200);
nor U34737 (N_34737,N_31770,N_30845);
xor U34738 (N_34738,N_31479,N_30262);
or U34739 (N_34739,N_32137,N_30433);
nor U34740 (N_34740,N_30226,N_31882);
xor U34741 (N_34741,N_31249,N_30661);
or U34742 (N_34742,N_30671,N_30131);
nor U34743 (N_34743,N_30277,N_30348);
nand U34744 (N_34744,N_31384,N_30135);
nand U34745 (N_34745,N_32023,N_31246);
nand U34746 (N_34746,N_30189,N_32139);
and U34747 (N_34747,N_31561,N_32001);
and U34748 (N_34748,N_32099,N_31205);
nor U34749 (N_34749,N_30387,N_31480);
xnor U34750 (N_34750,N_30723,N_32136);
nand U34751 (N_34751,N_31665,N_32463);
nor U34752 (N_34752,N_31778,N_30802);
nand U34753 (N_34753,N_32204,N_31928);
nor U34754 (N_34754,N_32291,N_31462);
nand U34755 (N_34755,N_30112,N_32423);
and U34756 (N_34756,N_30881,N_31458);
or U34757 (N_34757,N_30103,N_31735);
nand U34758 (N_34758,N_30731,N_32008);
xnor U34759 (N_34759,N_32466,N_30174);
xor U34760 (N_34760,N_31922,N_30532);
or U34761 (N_34761,N_32143,N_30974);
nor U34762 (N_34762,N_30898,N_30064);
nand U34763 (N_34763,N_31083,N_30217);
and U34764 (N_34764,N_31031,N_32426);
nand U34765 (N_34765,N_32290,N_30433);
xnor U34766 (N_34766,N_31437,N_31926);
nand U34767 (N_34767,N_31245,N_31201);
or U34768 (N_34768,N_31451,N_31719);
nand U34769 (N_34769,N_30819,N_30621);
and U34770 (N_34770,N_30451,N_30869);
nand U34771 (N_34771,N_31363,N_31771);
xor U34772 (N_34772,N_31732,N_32268);
and U34773 (N_34773,N_31225,N_30367);
xor U34774 (N_34774,N_30803,N_31769);
nor U34775 (N_34775,N_31644,N_31041);
nor U34776 (N_34776,N_30953,N_32470);
nor U34777 (N_34777,N_31251,N_31567);
nand U34778 (N_34778,N_30991,N_31549);
nand U34779 (N_34779,N_30619,N_32201);
nand U34780 (N_34780,N_31131,N_30086);
nand U34781 (N_34781,N_32317,N_31887);
or U34782 (N_34782,N_31282,N_31488);
nor U34783 (N_34783,N_31127,N_31588);
and U34784 (N_34784,N_30098,N_31784);
or U34785 (N_34785,N_30786,N_30915);
nand U34786 (N_34786,N_32184,N_32277);
nor U34787 (N_34787,N_31425,N_31288);
nand U34788 (N_34788,N_32113,N_30722);
nor U34789 (N_34789,N_30221,N_30373);
or U34790 (N_34790,N_30112,N_30286);
nand U34791 (N_34791,N_30467,N_31991);
nand U34792 (N_34792,N_31089,N_32144);
nand U34793 (N_34793,N_30370,N_31947);
or U34794 (N_34794,N_31247,N_31126);
and U34795 (N_34795,N_32073,N_32046);
nor U34796 (N_34796,N_30375,N_31654);
xnor U34797 (N_34797,N_31329,N_30850);
xor U34798 (N_34798,N_30531,N_31624);
nor U34799 (N_34799,N_31581,N_30951);
nor U34800 (N_34800,N_30616,N_30982);
or U34801 (N_34801,N_30281,N_30558);
and U34802 (N_34802,N_30168,N_32148);
xor U34803 (N_34803,N_30833,N_31763);
or U34804 (N_34804,N_31268,N_31506);
or U34805 (N_34805,N_30622,N_31175);
nand U34806 (N_34806,N_31907,N_30822);
xor U34807 (N_34807,N_30287,N_31184);
nor U34808 (N_34808,N_31276,N_32281);
and U34809 (N_34809,N_30199,N_32459);
or U34810 (N_34810,N_30288,N_31137);
or U34811 (N_34811,N_31098,N_31043);
nand U34812 (N_34812,N_31552,N_32275);
nand U34813 (N_34813,N_31669,N_31156);
xnor U34814 (N_34814,N_31956,N_31265);
nand U34815 (N_34815,N_30957,N_31467);
nor U34816 (N_34816,N_31046,N_30188);
or U34817 (N_34817,N_31841,N_32126);
xor U34818 (N_34818,N_30741,N_31184);
nor U34819 (N_34819,N_31738,N_31411);
nor U34820 (N_34820,N_31354,N_32137);
nor U34821 (N_34821,N_31679,N_30235);
nand U34822 (N_34822,N_31845,N_30880);
xnor U34823 (N_34823,N_31037,N_32233);
nand U34824 (N_34824,N_30057,N_30952);
and U34825 (N_34825,N_31064,N_31004);
nor U34826 (N_34826,N_30491,N_30774);
nand U34827 (N_34827,N_30278,N_30798);
and U34828 (N_34828,N_30996,N_31666);
xor U34829 (N_34829,N_31571,N_31623);
and U34830 (N_34830,N_30853,N_31644);
or U34831 (N_34831,N_31753,N_30330);
or U34832 (N_34832,N_31890,N_31306);
nand U34833 (N_34833,N_30951,N_31311);
xnor U34834 (N_34834,N_30611,N_30707);
and U34835 (N_34835,N_31268,N_30023);
or U34836 (N_34836,N_30365,N_30141);
nand U34837 (N_34837,N_32465,N_30076);
nor U34838 (N_34838,N_31085,N_31631);
nor U34839 (N_34839,N_32000,N_32057);
nor U34840 (N_34840,N_30021,N_30886);
nand U34841 (N_34841,N_31898,N_31703);
xor U34842 (N_34842,N_30246,N_32200);
xnor U34843 (N_34843,N_32416,N_31787);
and U34844 (N_34844,N_32216,N_31563);
nor U34845 (N_34845,N_31721,N_31778);
and U34846 (N_34846,N_30871,N_30081);
xnor U34847 (N_34847,N_30548,N_30174);
or U34848 (N_34848,N_31077,N_32168);
nand U34849 (N_34849,N_30815,N_31346);
or U34850 (N_34850,N_32481,N_30732);
xor U34851 (N_34851,N_31343,N_30107);
and U34852 (N_34852,N_30095,N_31721);
and U34853 (N_34853,N_30416,N_31933);
nand U34854 (N_34854,N_31284,N_31092);
nor U34855 (N_34855,N_30508,N_30457);
and U34856 (N_34856,N_32320,N_30528);
nor U34857 (N_34857,N_31376,N_31485);
and U34858 (N_34858,N_31637,N_30899);
or U34859 (N_34859,N_32087,N_30688);
nand U34860 (N_34860,N_31669,N_31202);
nand U34861 (N_34861,N_31847,N_30435);
and U34862 (N_34862,N_30236,N_31895);
nor U34863 (N_34863,N_31786,N_30649);
and U34864 (N_34864,N_30738,N_31041);
xor U34865 (N_34865,N_32114,N_30811);
nor U34866 (N_34866,N_32171,N_32009);
or U34867 (N_34867,N_32219,N_30584);
or U34868 (N_34868,N_31108,N_31654);
xor U34869 (N_34869,N_30753,N_31738);
and U34870 (N_34870,N_32380,N_30145);
nor U34871 (N_34871,N_30211,N_30190);
and U34872 (N_34872,N_30659,N_30697);
nor U34873 (N_34873,N_31059,N_30851);
nor U34874 (N_34874,N_30500,N_30615);
and U34875 (N_34875,N_30454,N_30556);
nand U34876 (N_34876,N_31542,N_32423);
nand U34877 (N_34877,N_30581,N_31395);
xnor U34878 (N_34878,N_30864,N_30508);
xnor U34879 (N_34879,N_30796,N_30794);
and U34880 (N_34880,N_30267,N_32297);
nor U34881 (N_34881,N_32477,N_31383);
nand U34882 (N_34882,N_31221,N_32273);
nand U34883 (N_34883,N_32105,N_30396);
or U34884 (N_34884,N_32393,N_30215);
xnor U34885 (N_34885,N_31479,N_31589);
and U34886 (N_34886,N_31111,N_30534);
xor U34887 (N_34887,N_30077,N_32200);
nor U34888 (N_34888,N_31595,N_32428);
nand U34889 (N_34889,N_32216,N_32066);
nand U34890 (N_34890,N_30248,N_31750);
nand U34891 (N_34891,N_30391,N_31031);
and U34892 (N_34892,N_32233,N_30615);
xor U34893 (N_34893,N_31247,N_31284);
and U34894 (N_34894,N_32217,N_31086);
nor U34895 (N_34895,N_30501,N_30745);
or U34896 (N_34896,N_30548,N_31288);
nor U34897 (N_34897,N_31987,N_31663);
or U34898 (N_34898,N_32082,N_31594);
xor U34899 (N_34899,N_31065,N_31409);
nor U34900 (N_34900,N_30189,N_31781);
nor U34901 (N_34901,N_31360,N_30519);
nor U34902 (N_34902,N_32150,N_30746);
xor U34903 (N_34903,N_31639,N_30942);
or U34904 (N_34904,N_31904,N_30864);
nor U34905 (N_34905,N_30124,N_30071);
or U34906 (N_34906,N_31553,N_30240);
and U34907 (N_34907,N_30127,N_30143);
nand U34908 (N_34908,N_32345,N_30474);
and U34909 (N_34909,N_32279,N_30622);
or U34910 (N_34910,N_30716,N_31281);
xnor U34911 (N_34911,N_30092,N_31237);
xnor U34912 (N_34912,N_30725,N_30478);
nand U34913 (N_34913,N_31484,N_32257);
or U34914 (N_34914,N_32339,N_31689);
or U34915 (N_34915,N_30125,N_30108);
or U34916 (N_34916,N_31406,N_31609);
nand U34917 (N_34917,N_30745,N_32183);
or U34918 (N_34918,N_30882,N_31273);
nor U34919 (N_34919,N_30291,N_30102);
xor U34920 (N_34920,N_30492,N_31956);
xnor U34921 (N_34921,N_32230,N_31941);
nand U34922 (N_34922,N_31480,N_31525);
nor U34923 (N_34923,N_32306,N_30800);
xor U34924 (N_34924,N_30127,N_31753);
and U34925 (N_34925,N_32265,N_31200);
nor U34926 (N_34926,N_32076,N_31059);
xor U34927 (N_34927,N_31967,N_30291);
and U34928 (N_34928,N_30255,N_31810);
nor U34929 (N_34929,N_31336,N_32145);
xnor U34930 (N_34930,N_30807,N_31544);
xnor U34931 (N_34931,N_32452,N_31697);
nor U34932 (N_34932,N_30422,N_30943);
nor U34933 (N_34933,N_32287,N_31301);
nor U34934 (N_34934,N_32488,N_30183);
or U34935 (N_34935,N_32370,N_31815);
or U34936 (N_34936,N_31248,N_32046);
or U34937 (N_34937,N_31352,N_30260);
or U34938 (N_34938,N_30207,N_30570);
nor U34939 (N_34939,N_31474,N_31991);
and U34940 (N_34940,N_31540,N_30810);
nand U34941 (N_34941,N_32332,N_31404);
and U34942 (N_34942,N_30747,N_31327);
xnor U34943 (N_34943,N_31020,N_31752);
and U34944 (N_34944,N_31322,N_30977);
or U34945 (N_34945,N_32145,N_31097);
nor U34946 (N_34946,N_30138,N_30350);
and U34947 (N_34947,N_32099,N_31174);
nor U34948 (N_34948,N_31201,N_31052);
nor U34949 (N_34949,N_30030,N_31577);
xnor U34950 (N_34950,N_31988,N_31920);
or U34951 (N_34951,N_30413,N_30449);
xor U34952 (N_34952,N_32021,N_31431);
and U34953 (N_34953,N_30409,N_32358);
nor U34954 (N_34954,N_30522,N_31299);
or U34955 (N_34955,N_31163,N_32217);
nand U34956 (N_34956,N_30408,N_30763);
nand U34957 (N_34957,N_32051,N_32076);
or U34958 (N_34958,N_32103,N_31504);
nor U34959 (N_34959,N_32028,N_30425);
xnor U34960 (N_34960,N_30062,N_32078);
nor U34961 (N_34961,N_30184,N_32447);
xnor U34962 (N_34962,N_32393,N_32125);
nand U34963 (N_34963,N_30200,N_30408);
and U34964 (N_34964,N_30309,N_31055);
xor U34965 (N_34965,N_31169,N_30871);
xnor U34966 (N_34966,N_30494,N_30005);
and U34967 (N_34967,N_30400,N_30335);
or U34968 (N_34968,N_30353,N_30520);
and U34969 (N_34969,N_31986,N_30948);
nand U34970 (N_34970,N_31642,N_31172);
nor U34971 (N_34971,N_31342,N_32357);
and U34972 (N_34972,N_31392,N_31807);
xnor U34973 (N_34973,N_30975,N_31432);
and U34974 (N_34974,N_31509,N_31213);
xor U34975 (N_34975,N_32061,N_31234);
nand U34976 (N_34976,N_31813,N_32054);
nand U34977 (N_34977,N_32473,N_30331);
nor U34978 (N_34978,N_32244,N_30341);
xnor U34979 (N_34979,N_31179,N_30413);
nand U34980 (N_34980,N_30500,N_31939);
nand U34981 (N_34981,N_30925,N_32249);
nand U34982 (N_34982,N_31090,N_31456);
xnor U34983 (N_34983,N_30004,N_31106);
nand U34984 (N_34984,N_31381,N_30326);
nand U34985 (N_34985,N_32015,N_31327);
nand U34986 (N_34986,N_32300,N_31462);
or U34987 (N_34987,N_30961,N_30111);
xnor U34988 (N_34988,N_31763,N_31516);
nor U34989 (N_34989,N_31515,N_30114);
nor U34990 (N_34990,N_32338,N_32031);
nand U34991 (N_34991,N_32111,N_30162);
nor U34992 (N_34992,N_32128,N_31795);
and U34993 (N_34993,N_31114,N_31128);
nor U34994 (N_34994,N_30196,N_30639);
and U34995 (N_34995,N_30831,N_30669);
nor U34996 (N_34996,N_31042,N_31410);
and U34997 (N_34997,N_31666,N_30578);
xnor U34998 (N_34998,N_31274,N_32439);
nand U34999 (N_34999,N_30195,N_32013);
and U35000 (N_35000,N_34226,N_33111);
or U35001 (N_35001,N_32520,N_33188);
nor U35002 (N_35002,N_33904,N_32690);
xnor U35003 (N_35003,N_34302,N_33594);
nand U35004 (N_35004,N_34559,N_32847);
nor U35005 (N_35005,N_34317,N_32915);
or U35006 (N_35006,N_32609,N_33093);
and U35007 (N_35007,N_32934,N_33176);
nand U35008 (N_35008,N_34982,N_34715);
nand U35009 (N_35009,N_34497,N_33551);
nand U35010 (N_35010,N_34456,N_32704);
and U35011 (N_35011,N_33925,N_32948);
and U35012 (N_35012,N_34015,N_32578);
nor U35013 (N_35013,N_34315,N_33761);
and U35014 (N_35014,N_34657,N_33617);
nor U35015 (N_35015,N_33201,N_32619);
nor U35016 (N_35016,N_34759,N_32631);
xor U35017 (N_35017,N_33395,N_34427);
or U35018 (N_35018,N_33776,N_32831);
nor U35019 (N_35019,N_34784,N_34314);
xnor U35020 (N_35020,N_33820,N_34174);
or U35021 (N_35021,N_32627,N_33935);
xnor U35022 (N_35022,N_33012,N_32679);
and U35023 (N_35023,N_32504,N_32559);
xnor U35024 (N_35024,N_33623,N_33908);
xnor U35025 (N_35025,N_34186,N_34989);
nand U35026 (N_35026,N_33689,N_32860);
xor U35027 (N_35027,N_34956,N_33031);
xnor U35028 (N_35028,N_33785,N_33157);
xor U35029 (N_35029,N_33678,N_33947);
nor U35030 (N_35030,N_33651,N_33252);
and U35031 (N_35031,N_33948,N_33044);
and U35032 (N_35032,N_32621,N_32606);
xnor U35033 (N_35033,N_33493,N_33106);
xor U35034 (N_35034,N_33185,N_34493);
nor U35035 (N_35035,N_34350,N_33489);
xor U35036 (N_35036,N_34138,N_34475);
and U35037 (N_35037,N_34899,N_33177);
nor U35038 (N_35038,N_33887,N_32507);
xor U35039 (N_35039,N_34184,N_33049);
nand U35040 (N_35040,N_32931,N_32634);
nor U35041 (N_35041,N_33876,N_32872);
and U35042 (N_35042,N_34041,N_34096);
nor U35043 (N_35043,N_34908,N_34901);
or U35044 (N_35044,N_33241,N_33076);
or U35045 (N_35045,N_33530,N_33636);
nor U35046 (N_35046,N_32577,N_34631);
xor U35047 (N_35047,N_33903,N_34697);
nor U35048 (N_35048,N_34794,N_33764);
xnor U35049 (N_35049,N_33618,N_34380);
or U35050 (N_35050,N_34419,N_34867);
nor U35051 (N_35051,N_34799,N_34240);
and U35052 (N_35052,N_33810,N_34248);
nor U35053 (N_35053,N_33500,N_32898);
xnor U35054 (N_35054,N_33403,N_32607);
nand U35055 (N_35055,N_33867,N_33021);
or U35056 (N_35056,N_33824,N_34798);
nand U35057 (N_35057,N_34047,N_34010);
and U35058 (N_35058,N_34454,N_32971);
xor U35059 (N_35059,N_33152,N_33909);
or U35060 (N_35060,N_33945,N_32626);
or U35061 (N_35061,N_34824,N_33601);
or U35062 (N_35062,N_34034,N_32549);
and U35063 (N_35063,N_34820,N_34059);
nor U35064 (N_35064,N_32593,N_32664);
xnor U35065 (N_35065,N_33606,N_33751);
nand U35066 (N_35066,N_33516,N_33470);
nand U35067 (N_35067,N_33787,N_33672);
or U35068 (N_35068,N_34868,N_32982);
or U35069 (N_35069,N_33183,N_34938);
nor U35070 (N_35070,N_34676,N_34936);
xnor U35071 (N_35071,N_33992,N_33557);
xor U35072 (N_35072,N_33913,N_32822);
and U35073 (N_35073,N_34461,N_34738);
xnor U35074 (N_35074,N_34575,N_33314);
or U35075 (N_35075,N_34374,N_32984);
xor U35076 (N_35076,N_34133,N_32942);
or U35077 (N_35077,N_34352,N_32735);
or U35078 (N_35078,N_33225,N_34349);
and U35079 (N_35079,N_34109,N_34050);
nor U35080 (N_35080,N_33303,N_33575);
and U35081 (N_35081,N_33409,N_33608);
xnor U35082 (N_35082,N_33206,N_34455);
and U35083 (N_35083,N_33224,N_33015);
xor U35084 (N_35084,N_34073,N_33569);
nor U35085 (N_35085,N_33479,N_34628);
xnor U35086 (N_35086,N_33704,N_32674);
and U35087 (N_35087,N_34627,N_33864);
and U35088 (N_35088,N_32892,N_33496);
nand U35089 (N_35089,N_33717,N_34215);
nor U35090 (N_35090,N_34655,N_34487);
or U35091 (N_35091,N_34690,N_33022);
or U35092 (N_35092,N_33006,N_32616);
or U35093 (N_35093,N_33349,N_34859);
or U35094 (N_35094,N_33644,N_32895);
and U35095 (N_35095,N_34217,N_33167);
nor U35096 (N_35096,N_34346,N_34939);
nand U35097 (N_35097,N_34760,N_32715);
nor U35098 (N_35098,N_33546,N_33124);
or U35099 (N_35099,N_33577,N_32779);
xor U35100 (N_35100,N_32623,N_33961);
nand U35101 (N_35101,N_33590,N_34209);
nor U35102 (N_35102,N_34363,N_34603);
and U35103 (N_35103,N_33816,N_34616);
nand U35104 (N_35104,N_32827,N_34845);
nor U35105 (N_35105,N_34301,N_33494);
or U35106 (N_35106,N_33216,N_33930);
nor U35107 (N_35107,N_34661,N_34071);
or U35108 (N_35108,N_32981,N_33918);
xnor U35109 (N_35109,N_34529,N_32820);
and U35110 (N_35110,N_32807,N_34612);
nand U35111 (N_35111,N_34724,N_33626);
nor U35112 (N_35112,N_33178,N_34749);
and U35113 (N_35113,N_34926,N_32937);
xor U35114 (N_35114,N_33629,N_33650);
and U35115 (N_35115,N_33294,N_33736);
or U35116 (N_35116,N_33217,N_33249);
nor U35117 (N_35117,N_34923,N_32502);
and U35118 (N_35118,N_34143,N_34643);
nor U35119 (N_35119,N_32696,N_33426);
xor U35120 (N_35120,N_33251,N_33633);
nand U35121 (N_35121,N_32750,N_34785);
or U35122 (N_35122,N_33790,N_33611);
nor U35123 (N_35123,N_32579,N_33030);
and U35124 (N_35124,N_34806,N_33112);
nor U35125 (N_35125,N_34505,N_33166);
and U35126 (N_35126,N_33207,N_32646);
and U35127 (N_35127,N_34020,N_32712);
xnor U35128 (N_35128,N_32673,N_33316);
xnor U35129 (N_35129,N_32535,N_34390);
or U35130 (N_35130,N_33813,N_34391);
nand U35131 (N_35131,N_34563,N_34500);
nor U35132 (N_35132,N_34453,N_34921);
or U35133 (N_35133,N_34610,N_33513);
xnor U35134 (N_35134,N_32657,N_32655);
nor U35135 (N_35135,N_34517,N_33994);
xnor U35136 (N_35136,N_32918,N_33372);
or U35137 (N_35137,N_33986,N_34665);
or U35138 (N_35138,N_32736,N_34422);
nand U35139 (N_35139,N_32661,N_33467);
nor U35140 (N_35140,N_33615,N_34489);
nor U35141 (N_35141,N_33807,N_34864);
xnor U35142 (N_35142,N_33688,N_33812);
nand U35143 (N_35143,N_34694,N_32710);
and U35144 (N_35144,N_32772,N_34823);
nor U35145 (N_35145,N_34407,N_33881);
and U35146 (N_35146,N_34995,N_33118);
or U35147 (N_35147,N_34025,N_33270);
or U35148 (N_35148,N_33090,N_33682);
nor U35149 (N_35149,N_33694,N_33845);
and U35150 (N_35150,N_33995,N_32826);
or U35151 (N_35151,N_32632,N_33000);
and U35152 (N_35152,N_34394,N_33019);
xnor U35153 (N_35153,N_34687,N_33315);
or U35154 (N_35154,N_33671,N_32806);
nand U35155 (N_35155,N_34365,N_33326);
and U35156 (N_35156,N_34637,N_32614);
or U35157 (N_35157,N_34731,N_34581);
or U35158 (N_35158,N_34112,N_33410);
or U35159 (N_35159,N_33684,N_34998);
or U35160 (N_35160,N_33237,N_32729);
and U35161 (N_35161,N_32746,N_34980);
and U35162 (N_35162,N_33210,N_34742);
xor U35163 (N_35163,N_32840,N_33724);
and U35164 (N_35164,N_34647,N_34764);
or U35165 (N_35165,N_32768,N_34651);
nor U35166 (N_35166,N_34592,N_33013);
or U35167 (N_35167,N_33480,N_33744);
nor U35168 (N_35168,N_34105,N_33839);
or U35169 (N_35169,N_34035,N_32983);
xnor U35170 (N_35170,N_32534,N_34291);
nor U35171 (N_35171,N_34658,N_34644);
or U35172 (N_35172,N_32944,N_33998);
nand U35173 (N_35173,N_34728,N_34323);
or U35174 (N_35174,N_33777,N_32687);
or U35175 (N_35175,N_34558,N_34984);
or U35176 (N_35176,N_32846,N_33701);
or U35177 (N_35177,N_34905,N_34622);
nor U35178 (N_35178,N_34305,N_34477);
nor U35179 (N_35179,N_33970,N_33681);
and U35180 (N_35180,N_34538,N_34070);
or U35181 (N_35181,N_33665,N_34316);
nand U35182 (N_35182,N_33953,N_33318);
xnor U35183 (N_35183,N_33975,N_33784);
nor U35184 (N_35184,N_34464,N_33028);
nand U35185 (N_35185,N_34987,N_34668);
and U35186 (N_35186,N_34682,N_34796);
nand U35187 (N_35187,N_34652,N_34153);
or U35188 (N_35188,N_33313,N_32727);
xor U35189 (N_35189,N_33794,N_34404);
nand U35190 (N_35190,N_33946,N_32836);
or U35191 (N_35191,N_33804,N_34932);
nand U35192 (N_35192,N_33127,N_33833);
or U35193 (N_35193,N_33831,N_34044);
nor U35194 (N_35194,N_33691,N_34045);
xor U35195 (N_35195,N_33852,N_34773);
or U35196 (N_35196,N_33203,N_34460);
nand U35197 (N_35197,N_34950,N_32992);
and U35198 (N_35198,N_33085,N_34698);
xnor U35199 (N_35199,N_33039,N_34421);
xnor U35200 (N_35200,N_33635,N_33956);
and U35201 (N_35201,N_32849,N_33829);
nand U35202 (N_35202,N_34278,N_34091);
nor U35203 (N_35203,N_33340,N_34147);
nor U35204 (N_35204,N_33630,N_33668);
nand U35205 (N_35205,N_34832,N_34928);
or U35206 (N_35206,N_33967,N_33305);
and U35207 (N_35207,N_33233,N_34108);
xor U35208 (N_35208,N_34418,N_32555);
and U35209 (N_35209,N_34854,N_32835);
and U35210 (N_35210,N_33711,N_32901);
nand U35211 (N_35211,N_33614,N_34384);
xor U35212 (N_35212,N_33540,N_32967);
nor U35213 (N_35213,N_34192,N_33838);
nand U35214 (N_35214,N_34338,N_33074);
nor U35215 (N_35215,N_33158,N_33828);
nor U35216 (N_35216,N_34378,N_33430);
or U35217 (N_35217,N_32999,N_32963);
or U35218 (N_35218,N_34113,N_34907);
or U35219 (N_35219,N_32728,N_33705);
xor U35220 (N_35220,N_34256,N_34746);
nor U35221 (N_35221,N_33043,N_32794);
nor U35222 (N_35222,N_32802,N_33104);
nand U35223 (N_35223,N_32582,N_33125);
nand U35224 (N_35224,N_34874,N_32688);
and U35225 (N_35225,N_32595,N_34855);
and U35226 (N_35226,N_34260,N_32740);
nor U35227 (N_35227,N_34355,N_33685);
nor U35228 (N_35228,N_33311,N_33610);
and U35229 (N_35229,N_34792,N_32838);
and U35230 (N_35230,N_33285,N_34289);
and U35231 (N_35231,N_33827,N_33466);
xor U35232 (N_35232,N_32884,N_33433);
or U35233 (N_35233,N_32526,N_33057);
nor U35234 (N_35234,N_33299,N_33860);
nand U35235 (N_35235,N_33740,N_34426);
or U35236 (N_35236,N_32516,N_33054);
xnor U35237 (N_35237,N_34183,N_32528);
nor U35238 (N_35238,N_33096,N_33312);
and U35239 (N_35239,N_33002,N_33379);
xor U35240 (N_35240,N_34595,N_32945);
nand U35241 (N_35241,N_34333,N_32813);
nand U35242 (N_35242,N_34442,N_32900);
and U35243 (N_35243,N_34815,N_34827);
and U35244 (N_35244,N_33747,N_33389);
nor U35245 (N_35245,N_33843,N_34400);
nand U35246 (N_35246,N_34159,N_33756);
and U35247 (N_35247,N_34021,N_33745);
nor U35248 (N_35248,N_33418,N_33718);
xor U35249 (N_35249,N_33084,N_32979);
or U35250 (N_35250,N_34437,N_34339);
nand U35251 (N_35251,N_33604,N_32897);
nor U35252 (N_35252,N_34398,N_34534);
nor U35253 (N_35253,N_34848,N_33102);
nand U35254 (N_35254,N_33593,N_32683);
or U35255 (N_35255,N_34739,N_33655);
or U35256 (N_35256,N_33055,N_32854);
or U35257 (N_35257,N_34079,N_32801);
nor U35258 (N_35258,N_34379,N_34249);
nand U35259 (N_35259,N_34648,N_33679);
or U35260 (N_35260,N_34841,N_34282);
or U35261 (N_35261,N_32702,N_34269);
xnor U35262 (N_35262,N_34863,N_34170);
nor U35263 (N_35263,N_32745,N_33170);
and U35264 (N_35264,N_33435,N_34683);
nand U35265 (N_35265,N_33149,N_33431);
nor U35266 (N_35266,N_33733,N_33154);
xnor U35267 (N_35267,N_33246,N_33713);
and U35268 (N_35268,N_34948,N_33268);
xor U35269 (N_35269,N_33215,N_32953);
nand U35270 (N_35270,N_32537,N_34341);
xor U35271 (N_35271,N_32642,N_33164);
nor U35272 (N_35272,N_32777,N_32685);
or U35273 (N_35273,N_34725,N_33261);
and U35274 (N_35274,N_34231,N_33750);
xor U35275 (N_35275,N_34941,N_33844);
nor U35276 (N_35276,N_34205,N_34325);
nand U35277 (N_35277,N_32681,N_34320);
nand U35278 (N_35278,N_34872,N_34416);
and U35279 (N_35279,N_34039,N_34801);
xor U35280 (N_35280,N_34252,N_34840);
xnor U35281 (N_35281,N_33400,N_34934);
or U35282 (N_35282,N_33487,N_32625);
nand U35283 (N_35283,N_33708,N_33979);
xnor U35284 (N_35284,N_34803,N_32701);
xnor U35285 (N_35285,N_34036,N_32828);
nor U35286 (N_35286,N_32639,N_33854);
nor U35287 (N_35287,N_32996,N_34604);
or U35288 (N_35288,N_32969,N_32771);
or U35289 (N_35289,N_33539,N_34897);
and U35290 (N_35290,N_32864,N_34942);
nand U35291 (N_35291,N_33365,N_34970);
nor U35292 (N_35292,N_32960,N_33003);
and U35293 (N_35293,N_34880,N_34735);
xnor U35294 (N_35294,N_33906,N_32697);
nand U35295 (N_35295,N_34608,N_33515);
or U35296 (N_35296,N_33646,N_34467);
or U35297 (N_35297,N_32525,N_34031);
nor U35298 (N_35298,N_34213,N_33574);
nand U35299 (N_35299,N_33440,N_34227);
nor U35300 (N_35300,N_34817,N_32719);
nor U35301 (N_35301,N_33597,N_33136);
nand U35302 (N_35302,N_34568,N_34247);
nor U35303 (N_35303,N_33137,N_34001);
nor U35304 (N_35304,N_32584,N_34369);
and U35305 (N_35305,N_33809,N_32695);
nand U35306 (N_35306,N_34413,N_33638);
nor U35307 (N_35307,N_33073,N_33017);
xnor U35308 (N_35308,N_33707,N_33563);
xnor U35309 (N_35309,N_33455,N_34555);
and U35310 (N_35310,N_32599,N_33194);
or U35311 (N_35311,N_33197,N_33079);
and U35312 (N_35312,N_34206,N_34714);
nand U35313 (N_35313,N_32908,N_34614);
nor U35314 (N_35314,N_33570,N_34005);
xnor U35315 (N_35315,N_34829,N_34567);
xor U35316 (N_35316,N_33011,N_34944);
nor U35317 (N_35317,N_34717,N_33212);
and U35318 (N_35318,N_33083,N_34465);
xnor U35319 (N_35319,N_33266,N_34546);
or U35320 (N_35320,N_32709,N_32924);
nor U35321 (N_35321,N_33748,N_34721);
nor U35322 (N_35322,N_32612,N_33041);
xor U35323 (N_35323,N_33107,N_34107);
or U35324 (N_35324,N_34046,N_34027);
nand U35325 (N_35325,N_32783,N_34755);
nor U35326 (N_35326,N_34789,N_34571);
or U35327 (N_35327,N_33439,N_34667);
and U35328 (N_35328,N_33066,N_34123);
nand U35329 (N_35329,N_34167,N_33499);
xor U35330 (N_35330,N_34808,N_33663);
and U35331 (N_35331,N_34539,N_33898);
nand U35332 (N_35332,N_34300,N_33902);
xnor U35333 (N_35333,N_32909,N_33156);
nor U35334 (N_35334,N_33976,N_33622);
or U35335 (N_35335,N_34635,N_34412);
or U35336 (N_35336,N_34891,N_34620);
nand U35337 (N_35337,N_33588,N_33327);
nand U35338 (N_35338,N_32926,N_33703);
and U35339 (N_35339,N_34064,N_33339);
nand U35340 (N_35340,N_34521,N_33388);
nor U35341 (N_35341,N_34584,N_32692);
nand U35342 (N_35342,N_33958,N_33460);
xnor U35343 (N_35343,N_33005,N_33583);
or U35344 (N_35344,N_33847,N_32568);
and U35345 (N_35345,N_33652,N_34494);
xnor U35346 (N_35346,N_34666,N_33585);
nor U35347 (N_35347,N_33959,N_33631);
or U35348 (N_35348,N_34003,N_33556);
and U35349 (N_35349,N_34011,N_33320);
nor U35350 (N_35350,N_32869,N_33376);
nand U35351 (N_35351,N_34586,N_33180);
nor U35352 (N_35352,N_34244,N_33738);
xor U35353 (N_35353,N_33397,N_32622);
and U35354 (N_35354,N_32651,N_33126);
and U35355 (N_35355,N_33086,N_33234);
xor U35356 (N_35356,N_34937,N_34187);
and U35357 (N_35357,N_34570,N_33269);
nor U35358 (N_35358,N_33147,N_33105);
and U35359 (N_35359,N_34328,N_33328);
and U35360 (N_35360,N_34700,N_32891);
or U35361 (N_35361,N_34364,N_34862);
xor U35362 (N_35362,N_34142,N_33230);
nor U35363 (N_35363,N_33661,N_34788);
or U35364 (N_35364,N_34996,N_33800);
nand U35365 (N_35365,N_33714,N_33542);
nand U35366 (N_35366,N_34572,N_33335);
and U35367 (N_35367,N_32851,N_34719);
and U35368 (N_35368,N_33566,N_33934);
and U35369 (N_35369,N_32879,N_34214);
xor U35370 (N_35370,N_33609,N_34639);
and U35371 (N_35371,N_33595,N_33442);
nand U35372 (N_35372,N_33307,N_34599);
xor U35373 (N_35373,N_33464,N_34104);
and U35374 (N_35374,N_34411,N_33357);
and U35375 (N_35375,N_34747,N_34791);
nand U35376 (N_35376,N_34161,N_32993);
nand U35377 (N_35377,N_33619,N_34125);
xor U35378 (N_35378,N_32604,N_33402);
or U35379 (N_35379,N_32788,N_34561);
nor U35380 (N_35380,N_33468,N_32640);
xnor U35381 (N_35381,N_34472,N_34136);
xnor U35382 (N_35382,N_34446,N_32961);
nor U35383 (N_35383,N_34495,N_34288);
or U35384 (N_35384,N_33443,N_32596);
and U35385 (N_35385,N_32876,N_34367);
nor U35386 (N_35386,N_34624,N_33508);
xnor U35387 (N_35387,N_32571,N_33666);
and U35388 (N_35388,N_33071,N_33599);
nand U35389 (N_35389,N_33232,N_32672);
and U35390 (N_35390,N_34957,N_34381);
xor U35391 (N_35391,N_34018,N_34902);
nand U35392 (N_35392,N_34383,N_34322);
nor U35393 (N_35393,N_34512,N_32956);
or U35394 (N_35394,N_33331,N_33475);
or U35395 (N_35395,N_34710,N_34765);
xor U35396 (N_35396,N_33477,N_34182);
xnor U35397 (N_35397,N_32671,N_34116);
and U35398 (N_35398,N_33427,N_33915);
or U35399 (N_35399,N_33890,N_33978);
and U35400 (N_35400,N_32691,N_34157);
xor U35401 (N_35401,N_32628,N_34836);
nor U35402 (N_35402,N_34433,N_34882);
xnor U35403 (N_35403,N_33901,N_33667);
nand U35404 (N_35404,N_32545,N_33150);
nand U35405 (N_35405,N_32991,N_33457);
nand U35406 (N_35406,N_33250,N_34155);
and U35407 (N_35407,N_34137,N_33371);
xor U35408 (N_35408,N_33363,N_34342);
or U35409 (N_35409,N_32837,N_33135);
and U35410 (N_35410,N_32734,N_34985);
xnor U35411 (N_35411,N_33647,N_33720);
or U35412 (N_35412,N_34933,N_33192);
or U35413 (N_35413,N_32567,N_33352);
xor U35414 (N_35414,N_32682,N_34826);
nor U35415 (N_35415,N_33760,N_34033);
or U35416 (N_35416,N_32732,N_34525);
nand U35417 (N_35417,N_34988,N_33990);
and U35418 (N_35418,N_34869,N_34330);
nor U35419 (N_35419,N_33380,N_34955);
nor U35420 (N_35420,N_34327,N_33360);
and U35421 (N_35421,N_32780,N_34115);
nor U35422 (N_35422,N_32659,N_34618);
and U35423 (N_35423,N_34431,N_34276);
and U35424 (N_35424,N_34629,N_34134);
nor U35425 (N_35425,N_33461,N_32601);
nand U35426 (N_35426,N_32814,N_32543);
and U35427 (N_35427,N_34201,N_34967);
and U35428 (N_35428,N_34522,N_34062);
or U35429 (N_35429,N_34946,N_33868);
or U35430 (N_35430,N_33119,N_34833);
or U35431 (N_35431,N_32747,N_34259);
nand U35432 (N_35432,N_34782,N_33336);
nor U35433 (N_35433,N_33301,N_34898);
and U35434 (N_35434,N_33875,N_33016);
and U35435 (N_35435,N_33300,N_32749);
xnor U35436 (N_35436,N_32731,N_34615);
and U35437 (N_35437,N_33554,N_34818);
or U35438 (N_35438,N_34524,N_33428);
nand U35439 (N_35439,N_34254,N_34310);
and U35440 (N_35440,N_33725,N_33545);
nor U35441 (N_35441,N_33193,N_32573);
xor U35442 (N_35442,N_33347,N_33757);
and U35443 (N_35443,N_32561,N_34781);
nand U35444 (N_35444,N_33398,N_34444);
nand U35445 (N_35445,N_34219,N_34922);
xor U35446 (N_35446,N_34130,N_34417);
xnor U35447 (N_35447,N_34663,N_33732);
nand U35448 (N_35448,N_33884,N_33628);
or U35449 (N_35449,N_33123,N_32603);
or U35450 (N_35450,N_33907,N_33368);
nor U35451 (N_35451,N_34630,N_33100);
or U35452 (N_35452,N_33983,N_32974);
or U35453 (N_35453,N_33385,N_33417);
or U35454 (N_35454,N_34602,N_33337);
and U35455 (N_35455,N_33871,N_33739);
nand U35456 (N_35456,N_33406,N_33755);
xnor U35457 (N_35457,N_34345,N_33295);
nand U35458 (N_35458,N_32656,N_33855);
nor U35459 (N_35459,N_34387,N_32751);
and U35460 (N_35460,N_33896,N_34993);
or U35461 (N_35461,N_33429,N_34587);
nor U35462 (N_35462,N_33065,N_32600);
xor U35463 (N_35463,N_32778,N_32726);
and U35464 (N_35464,N_33026,N_34106);
or U35465 (N_35465,N_32620,N_34963);
and U35466 (N_35466,N_32796,N_32586);
xor U35467 (N_35467,N_34152,N_34466);
nand U35468 (N_35468,N_33792,N_32737);
or U35469 (N_35469,N_34774,N_34619);
xnor U35470 (N_35470,N_34311,N_34262);
and U35471 (N_35471,N_33448,N_33228);
nand U35472 (N_35472,N_33345,N_34347);
nand U35473 (N_35473,N_32698,N_34429);
nor U35474 (N_35474,N_33142,N_33659);
and U35475 (N_35475,N_34294,N_34973);
xnor U35476 (N_35476,N_34479,N_34360);
or U35477 (N_35477,N_33605,N_32793);
and U35478 (N_35478,N_33236,N_33805);
nand U35479 (N_35479,N_34366,N_32800);
and U35480 (N_35480,N_34204,N_33742);
xor U35481 (N_35481,N_34793,N_33706);
or U35482 (N_35482,N_34689,N_33949);
nand U35483 (N_35483,N_33632,N_34230);
nand U35484 (N_35484,N_32654,N_33826);
xor U35485 (N_35485,N_33173,N_32686);
or U35486 (N_35486,N_34769,N_32738);
and U35487 (N_35487,N_33553,N_34709);
and U35488 (N_35488,N_34168,N_33941);
or U35489 (N_35489,N_33374,N_33227);
xor U35490 (N_35490,N_33064,N_32693);
or U35491 (N_35491,N_32583,N_34674);
nand U35492 (N_35492,N_33288,N_32741);
or U35493 (N_35493,N_34156,N_34893);
nand U35494 (N_35494,N_34049,N_34900);
or U35495 (N_35495,N_32760,N_33245);
or U35496 (N_35496,N_34532,N_33254);
and U35497 (N_35497,N_32865,N_33895);
nor U35498 (N_35498,N_34669,N_34752);
or U35499 (N_35499,N_34382,N_34207);
and U35500 (N_35500,N_33933,N_33561);
nor U35501 (N_35501,N_33710,N_34858);
nor U35502 (N_35502,N_34488,N_32513);
xor U35503 (N_35503,N_34179,N_34238);
xnor U35504 (N_35504,N_32830,N_34280);
nand U35505 (N_35505,N_34353,N_33133);
or U35506 (N_35506,N_32575,N_33483);
and U35507 (N_35507,N_33795,N_33437);
and U35508 (N_35508,N_34800,N_32964);
nor U35509 (N_35509,N_32832,N_34006);
or U35510 (N_35510,N_32587,N_34385);
xnor U35511 (N_35511,N_33798,N_32733);
or U35512 (N_35512,N_33159,N_34609);
or U35513 (N_35513,N_32580,N_34068);
xor U35514 (N_35514,N_34758,N_33103);
nand U35515 (N_35515,N_33968,N_34055);
nand U35516 (N_35516,N_33541,N_34450);
nor U35517 (N_35517,N_32650,N_33473);
nor U35518 (N_35518,N_32989,N_32532);
and U35519 (N_35519,N_34290,N_34850);
xor U35520 (N_35520,N_33399,N_34951);
nand U35521 (N_35521,N_32770,N_33050);
nor U35522 (N_35522,N_33278,N_32711);
xor U35523 (N_35523,N_34098,N_32803);
or U35524 (N_35524,N_34560,N_34975);
xnor U35525 (N_35525,N_33524,N_34030);
or U35526 (N_35526,N_33488,N_34090);
nor U35527 (N_35527,N_34711,N_33921);
xnor U35528 (N_35528,N_32913,N_34362);
nand U35529 (N_35529,N_33229,N_32684);
and U35530 (N_35530,N_34660,N_32660);
xnor U35531 (N_35531,N_33558,N_33730);
or U35532 (N_35532,N_34593,N_34918);
and U35533 (N_35533,N_34139,N_33560);
nor U35534 (N_35534,N_33520,N_34335);
or U35535 (N_35535,N_33687,N_32668);
or U35536 (N_35536,N_32533,N_32853);
xor U35537 (N_35537,N_34258,N_32677);
nor U35538 (N_35538,N_34780,N_34958);
nand U35539 (N_35539,N_34312,N_34763);
nor U35540 (N_35540,N_32790,N_33624);
or U35541 (N_35541,N_34514,N_33413);
and U35542 (N_35542,N_34216,N_34686);
or U35543 (N_35543,N_34208,N_33926);
nand U35544 (N_35544,N_33920,N_33143);
or U35545 (N_35545,N_33068,N_33023);
nand U35546 (N_35546,N_33674,N_33658);
xnor U35547 (N_35547,N_34253,N_34974);
or U35548 (N_35548,N_33793,N_33894);
or U35549 (N_35549,N_34935,N_34239);
and U35550 (N_35550,N_34641,N_33879);
nand U35551 (N_35551,N_32680,N_33582);
nand U35552 (N_35552,N_34636,N_33160);
nor U35553 (N_35553,N_33344,N_33195);
nor U35554 (N_35554,N_32724,N_32868);
xnor U35555 (N_35555,N_34410,N_34476);
and U35556 (N_35556,N_32888,N_33432);
and U35557 (N_35557,N_34978,N_33223);
nand U35558 (N_35558,N_34720,N_34439);
and U35559 (N_35559,N_33559,N_32844);
and U35560 (N_35560,N_33010,N_32859);
nor U35561 (N_35561,N_33145,N_33988);
xor U35562 (N_35562,N_33053,N_33492);
nand U35563 (N_35563,N_34701,N_33247);
or U35564 (N_35564,N_34722,N_32919);
or U35565 (N_35565,N_33491,N_34979);
nor U35566 (N_35566,N_34086,N_34723);
nand U35567 (N_35567,N_34991,N_34757);
or U35568 (N_35568,N_34813,N_32666);
and U35569 (N_35569,N_34358,N_34075);
nor U35570 (N_35570,N_33361,N_32718);
and U35571 (N_35571,N_32590,N_33444);
or U35572 (N_35572,N_34255,N_33572);
xnor U35573 (N_35573,N_33944,N_32597);
xnor U35574 (N_35574,N_33260,N_33098);
nor U35575 (N_35575,N_33529,N_33434);
or U35576 (N_35576,N_34878,N_33505);
nand U35577 (N_35577,N_32523,N_33356);
nand U35578 (N_35578,N_34678,N_32529);
nor U35579 (N_35579,N_33752,N_34195);
nor U35580 (N_35580,N_34693,N_34541);
nor U35581 (N_35581,N_32972,N_33743);
nor U35582 (N_35582,N_34332,N_33931);
or U35583 (N_35583,N_32817,N_34816);
and U35584 (N_35584,N_33174,N_33997);
xor U35585 (N_35585,N_33726,N_34607);
or U35586 (N_35586,N_33686,N_34331);
nor U35587 (N_35587,N_32557,N_33394);
xor U35588 (N_35588,N_34585,N_34528);
or U35589 (N_35589,N_32758,N_34072);
or U35590 (N_35590,N_33034,N_34992);
xor U35591 (N_35591,N_32550,N_34547);
or U35592 (N_35592,N_32739,N_32910);
and U35593 (N_35593,N_33391,N_32899);
nand U35594 (N_35594,N_34054,N_34582);
or U35595 (N_35595,N_32885,N_32706);
nor U35596 (N_35596,N_34009,N_34076);
and U35597 (N_35597,N_32857,N_33129);
xor U35598 (N_35598,N_33382,N_34122);
or U35599 (N_35599,N_34553,N_33256);
nor U35600 (N_35600,N_34014,N_33421);
nand U35601 (N_35601,N_33091,N_34653);
nand U35602 (N_35602,N_33351,N_32598);
nor U35603 (N_35603,N_33669,N_33128);
and U35604 (N_35604,N_33702,N_32954);
nand U35605 (N_35605,N_33221,N_34052);
nand U35606 (N_35606,N_32815,N_33565);
nor U35607 (N_35607,N_34606,N_33842);
nor U35608 (N_35608,N_32896,N_34396);
nand U35609 (N_35609,N_32789,N_33734);
nor U35610 (N_35610,N_33536,N_33329);
xor U35611 (N_35611,N_33202,N_34861);
or U35612 (N_35612,N_33244,N_34810);
nand U35613 (N_35613,N_34199,N_33310);
and U35614 (N_35614,N_33490,N_34692);
and U35615 (N_35615,N_33097,N_34078);
nand U35616 (N_35616,N_33965,N_33171);
xor U35617 (N_35617,N_33184,N_33991);
or U35618 (N_35618,N_32722,N_34480);
nand U35619 (N_35619,N_34095,N_32667);
or U35620 (N_35620,N_34890,N_33070);
or U35621 (N_35621,N_34819,N_34129);
nor U35622 (N_35622,N_32645,N_33700);
nand U35623 (N_35623,N_33051,N_33841);
xor U35624 (N_35624,N_34994,N_34856);
nor U35625 (N_35625,N_32703,N_34457);
or U35626 (N_35626,N_33045,N_33779);
or U35627 (N_35627,N_32527,N_34783);
and U35628 (N_35628,N_32515,N_32530);
nor U35629 (N_35629,N_34304,N_34297);
nand U35630 (N_35630,N_33454,N_33075);
nand U35631 (N_35631,N_34947,N_32965);
nand U35632 (N_35632,N_33690,N_34016);
and U35633 (N_35633,N_33450,N_33873);
or U35634 (N_35634,N_33304,N_34679);
xnor U35635 (N_35635,N_33486,N_33257);
or U35636 (N_35636,N_33891,N_34750);
and U35637 (N_35637,N_33298,N_33059);
and U35638 (N_35638,N_34340,N_34275);
and U35639 (N_35639,N_34811,N_33272);
nand U35640 (N_35640,N_33281,N_32503);
nand U35641 (N_35641,N_34236,N_32975);
or U35642 (N_35642,N_33797,N_34931);
or U35643 (N_35643,N_34440,N_34000);
or U35644 (N_35644,N_32766,N_34083);
or U35645 (N_35645,N_32861,N_32608);
nand U35646 (N_35646,N_33025,N_34057);
nand U35647 (N_35647,N_33819,N_33484);
nor U35648 (N_35648,N_32767,N_34029);
and U35649 (N_35649,N_34449,N_32611);
xnor U35650 (N_35650,N_33547,N_33035);
nor U35651 (N_35651,N_32883,N_33168);
xor U35652 (N_35652,N_33200,N_34074);
and U35653 (N_35653,N_34509,N_33419);
nor U35654 (N_35654,N_34084,N_34502);
or U35655 (N_35655,N_34251,N_34484);
and U35656 (N_35656,N_33323,N_32878);
nor U35657 (N_35657,N_34754,N_33029);
nand U35658 (N_35658,N_32786,N_34914);
nand U35659 (N_35659,N_33048,N_34726);
and U35660 (N_35660,N_33122,N_34596);
or U35661 (N_35661,N_32591,N_34751);
xnor U35662 (N_35662,N_33153,N_33627);
or U35663 (N_35663,N_34943,N_34839);
or U35664 (N_35664,N_33791,N_33568);
or U35665 (N_35665,N_33535,N_33982);
or U35666 (N_35666,N_34492,N_33849);
or U35667 (N_35667,N_34229,N_33007);
and U35668 (N_35668,N_33578,N_33077);
nand U35669 (N_35669,N_34220,N_34212);
nand U35670 (N_35670,N_34225,N_34837);
xor U35671 (N_35671,N_32863,N_34625);
nand U35672 (N_35672,N_34144,N_32843);
and U35673 (N_35673,N_32904,N_32570);
and U35674 (N_35674,N_34857,N_34913);
nand U35675 (N_35675,N_34172,N_34344);
or U35676 (N_35676,N_32588,N_34223);
nor U35677 (N_35677,N_32638,N_34284);
nand U35678 (N_35678,N_32792,N_33660);
or U35679 (N_35679,N_32730,N_34243);
nand U35680 (N_35680,N_34888,N_33392);
nor U35681 (N_35681,N_32753,N_33469);
and U35682 (N_35682,N_34272,N_34688);
xnor U35683 (N_35683,N_33753,N_34318);
and U35684 (N_35684,N_33456,N_33047);
xor U35685 (N_35685,N_34038,N_34736);
xor U35686 (N_35686,N_34740,N_32893);
nor U35687 (N_35687,N_34151,N_34348);
and U35688 (N_35688,N_32713,N_33420);
and U35689 (N_35689,N_32958,N_34911);
and U35690 (N_35690,N_34732,N_33858);
nand U35691 (N_35691,N_34202,N_33424);
nor U35692 (N_35692,N_33676,N_32922);
and U35693 (N_35693,N_32705,N_33972);
xnor U35694 (N_35694,N_33275,N_32505);
nand U35695 (N_35695,N_33869,N_34189);
and U35696 (N_35696,N_32565,N_32548);
xnor U35697 (N_35697,N_32784,N_32976);
nor U35698 (N_35698,N_34954,N_32987);
nand U35699 (N_35699,N_34040,N_34042);
nor U35700 (N_35700,N_33693,N_33099);
and U35701 (N_35701,N_33977,N_34504);
nor U35702 (N_35702,N_34100,N_33411);
nand U35703 (N_35703,N_34704,N_32652);
xnor U35704 (N_35704,N_34797,N_33656);
and U35705 (N_35705,N_33497,N_34562);
and U35706 (N_35706,N_33498,N_34126);
or U35707 (N_35707,N_33865,N_32643);
or U35708 (N_35708,N_34600,N_33573);
nor U35709 (N_35709,N_34458,N_34023);
nand U35710 (N_35710,N_34513,N_33032);
or U35711 (N_35711,N_33186,N_34149);
nand U35712 (N_35712,N_34420,N_32717);
or U35713 (N_35713,N_34481,N_34279);
and U35714 (N_35714,N_32716,N_34415);
and U35715 (N_35715,N_34671,N_34131);
or U35716 (N_35716,N_34530,N_32930);
xor U35717 (N_35717,N_33503,N_32506);
nor U35718 (N_35718,N_34730,N_34778);
xnor U35719 (N_35719,N_33625,N_32812);
nand U35720 (N_35720,N_34702,N_33731);
and U35721 (N_35721,N_34632,N_33696);
nand U35722 (N_35722,N_33087,N_34397);
nor U35723 (N_35723,N_34904,N_34319);
and U35724 (N_35724,N_34471,N_34424);
nor U35725 (N_35725,N_32658,N_32995);
xor U35726 (N_35726,N_34640,N_34879);
nand U35727 (N_35727,N_34633,N_33811);
and U35728 (N_35728,N_32866,N_33544);
and U35729 (N_35729,N_34447,N_33781);
xor U35730 (N_35730,N_33770,N_32524);
and U35731 (N_35731,N_33375,N_34443);
nor U35732 (N_35732,N_32572,N_34463);
xor U35733 (N_35733,N_32602,N_33286);
xnor U35734 (N_35734,N_34673,N_34462);
nand U35735 (N_35735,N_34966,N_34695);
xor U35736 (N_35736,N_33191,N_34672);
xnor U35737 (N_35737,N_33822,N_33446);
nand U35738 (N_35738,N_33148,N_34886);
and U35739 (N_35739,N_33808,N_33451);
nand U35740 (N_35740,N_32743,N_33893);
nand U35741 (N_35741,N_34087,N_33187);
nand U35742 (N_35742,N_34866,N_34295);
nor U35743 (N_35743,N_34028,N_34598);
or U35744 (N_35744,N_34556,N_34729);
nand U35745 (N_35745,N_33161,N_32787);
nor U35746 (N_35746,N_33683,N_33366);
or U35747 (N_35747,N_33835,N_34916);
or U35748 (N_35748,N_32804,N_32742);
or U35749 (N_35749,N_34777,N_34067);
nand U35750 (N_35750,N_34656,N_32955);
or U35751 (N_35751,N_33175,N_32882);
and U35752 (N_35752,N_34677,N_33653);
xor U35753 (N_35753,N_33141,N_34924);
nand U35754 (N_35754,N_34077,N_32769);
and U35755 (N_35755,N_34441,N_33637);
and U35756 (N_35756,N_34779,N_33531);
nand U35757 (N_35757,N_33042,N_34140);
and U35758 (N_35758,N_32636,N_34313);
xor U35759 (N_35759,N_33052,N_32852);
and U35760 (N_35760,N_33350,N_33603);
nor U35761 (N_35761,N_32764,N_33190);
xor U35762 (N_35762,N_33196,N_34434);
nor U35763 (N_35763,N_34919,N_33384);
and U35764 (N_35764,N_33208,N_32950);
nor U35765 (N_35765,N_33297,N_33078);
xor U35766 (N_35766,N_33680,N_32774);
or U35767 (N_35767,N_34889,N_33642);
and U35768 (N_35768,N_34579,N_33877);
nor U35769 (N_35769,N_32675,N_32917);
nand U35770 (N_35770,N_33289,N_32850);
nand U35771 (N_35771,N_33600,N_32594);
nor U35772 (N_35772,N_34825,N_33981);
nor U35773 (N_35773,N_33806,N_33131);
xnor U35774 (N_35774,N_33001,N_32635);
nand U35775 (N_35775,N_32902,N_34964);
xor U35776 (N_35776,N_34713,N_34523);
and U35777 (N_35777,N_34681,N_34588);
nor U35778 (N_35778,N_33796,N_32970);
and U35779 (N_35779,N_33354,N_34405);
or U35780 (N_35780,N_33332,N_33181);
and U35781 (N_35781,N_32610,N_33936);
and U35782 (N_35782,N_34069,N_32905);
and U35783 (N_35783,N_34408,N_33205);
nor U35784 (N_35784,N_34691,N_34241);
nand U35785 (N_35785,N_33592,N_34573);
or U35786 (N_35786,N_34048,N_33008);
or U35787 (N_35787,N_33950,N_32536);
or U35788 (N_35788,N_34590,N_32874);
and U35789 (N_35789,N_33963,N_33452);
or U35790 (N_35790,N_33169,N_34265);
nor U35791 (N_35791,N_33910,N_34659);
nor U35792 (N_35792,N_34277,N_34191);
nor U35793 (N_35793,N_33525,N_32933);
and U35794 (N_35794,N_34952,N_32514);
nand U35795 (N_35795,N_33182,N_32720);
and U35796 (N_35796,N_33282,N_33293);
nand U35797 (N_35797,N_33613,N_34171);
or U35798 (N_35798,N_33146,N_33378);
or U35799 (N_35799,N_32799,N_34708);
and U35800 (N_35800,N_33695,N_34436);
nor U35801 (N_35801,N_34393,N_32881);
xor U35802 (N_35802,N_33534,N_32678);
or U35803 (N_35803,N_33723,N_33040);
nor U35804 (N_35804,N_34403,N_34920);
nor U35805 (N_35805,N_34831,N_32951);
xor U35806 (N_35806,N_33916,N_34734);
nand U35807 (N_35807,N_32952,N_32665);
xor U35808 (N_35808,N_33823,N_34997);
nand U35809 (N_35809,N_33727,N_34373);
nor U35810 (N_35810,N_33698,N_33943);
xnor U35811 (N_35811,N_34718,N_34703);
xor U35812 (N_35812,N_32562,N_33928);
xnor U35813 (N_35813,N_34977,N_34578);
nand U35814 (N_35814,N_33662,N_34012);
or U35815 (N_35815,N_34430,N_33853);
xor U35816 (N_35816,N_33140,N_33116);
nor U35817 (N_35817,N_34180,N_33602);
or U35818 (N_35818,N_34895,N_34490);
or U35819 (N_35819,N_33567,N_33132);
and U35820 (N_35820,N_33405,N_34762);
nand U35821 (N_35821,N_34474,N_33412);
or U35822 (N_35822,N_32721,N_33769);
or U35823 (N_35823,N_32841,N_33144);
nand U35824 (N_35824,N_33179,N_34081);
and U35825 (N_35825,N_34881,N_34203);
and U35826 (N_35826,N_34299,N_34821);
nor U35827 (N_35827,N_34066,N_33262);
or U35828 (N_35828,N_34515,N_33728);
xnor U35829 (N_35829,N_32617,N_33538);
nand U35830 (N_35830,N_34664,N_34884);
or U35831 (N_35831,N_34309,N_34273);
or U35832 (N_35832,N_33964,N_33870);
xnor U35833 (N_35833,N_34972,N_34266);
or U35834 (N_35834,N_33020,N_32700);
xor U35835 (N_35835,N_34903,N_34705);
or U35836 (N_35836,N_33673,N_34121);
xor U35837 (N_35837,N_34930,N_32923);
nand U35838 (N_35838,N_32676,N_33741);
xor U35839 (N_35839,N_33942,N_33649);
nor U35840 (N_35840,N_32748,N_33856);
nor U35841 (N_35841,N_34844,N_34085);
or U35842 (N_35842,N_34767,N_33951);
or U35843 (N_35843,N_33654,N_34056);
nor U35844 (N_35844,N_33987,N_32855);
or U35845 (N_35845,N_33343,N_33056);
and U35846 (N_35846,N_33639,N_34733);
nor U35847 (N_35847,N_34876,N_33501);
nand U35848 (N_35848,N_34092,N_34828);
xnor U35849 (N_35849,N_34830,N_32906);
and U35850 (N_35850,N_34356,N_33762);
or U35851 (N_35851,N_33317,N_34146);
or U35852 (N_35852,N_33482,N_34210);
or U35853 (N_35853,N_33138,N_34334);
nand U35854 (N_35854,N_34296,N_33240);
and U35855 (N_35855,N_33621,N_33330);
and U35856 (N_35856,N_32546,N_34181);
xnor U35857 (N_35857,N_34670,N_33165);
or U35858 (N_35858,N_34699,N_33861);
xnor U35859 (N_35859,N_33938,N_34414);
or U35860 (N_35860,N_34377,N_33209);
or U35861 (N_35861,N_33235,N_33821);
and U35862 (N_35862,N_34292,N_34917);
nor U35863 (N_35863,N_32824,N_33211);
xnor U35864 (N_35864,N_34851,N_33458);
nor U35865 (N_35865,N_33737,N_33283);
xor U35866 (N_35866,N_33830,N_33840);
or U35867 (N_35867,N_34756,N_33151);
nand U35868 (N_35868,N_34324,N_34646);
or U35869 (N_35869,N_33267,N_33519);
xnor U35870 (N_35870,N_33721,N_32839);
and U35871 (N_35871,N_33308,N_33591);
xor U35872 (N_35872,N_32551,N_33940);
and U35873 (N_35873,N_34224,N_34386);
xor U35874 (N_35874,N_32823,N_33980);
xnor U35875 (N_35875,N_34019,N_34285);
and U35876 (N_35876,N_34043,N_33507);
or U35877 (N_35877,N_33509,N_33549);
nand U35878 (N_35878,N_33478,N_32539);
nor U35879 (N_35879,N_33407,N_32662);
or U35880 (N_35880,N_34110,N_32541);
or U35881 (N_35881,N_34960,N_34835);
nand U35882 (N_35882,N_34519,N_33121);
xnor U35883 (N_35883,N_33888,N_34080);
nor U35884 (N_35884,N_32880,N_33258);
and U35885 (N_35885,N_32653,N_34537);
xor U35886 (N_35886,N_33115,N_34246);
and U35887 (N_35887,N_34577,N_32781);
and U35888 (N_35888,N_33589,N_33974);
and U35889 (N_35889,N_34088,N_34257);
nand U35890 (N_35890,N_34232,N_34409);
or U35891 (N_35891,N_33280,N_34097);
nor U35892 (N_35892,N_34962,N_34605);
xnor U35893 (N_35893,N_34242,N_32699);
nand U35894 (N_35894,N_33914,N_33242);
nor U35895 (N_35895,N_34520,N_34198);
or U35896 (N_35896,N_32512,N_34569);
xor U35897 (N_35897,N_33999,N_34321);
or U35898 (N_35898,N_33899,N_33543);
nand U35899 (N_35899,N_33383,N_33113);
and U35900 (N_35900,N_33859,N_33778);
nand U35901 (N_35901,N_32511,N_34745);
and U35902 (N_35902,N_32886,N_33284);
nor U35903 (N_35903,N_33874,N_34611);
nor U35904 (N_35904,N_34894,N_32765);
nor U35905 (N_35905,N_34270,N_34298);
nor U35906 (N_35906,N_32821,N_32707);
and U35907 (N_35907,N_32949,N_32776);
xor U35908 (N_35908,N_34022,N_33425);
and U35909 (N_35909,N_32966,N_33279);
nand U35910 (N_35910,N_33989,N_34557);
nand U35911 (N_35911,N_34550,N_34877);
and U35912 (N_35912,N_32633,N_32647);
xor U35913 (N_35913,N_33919,N_34372);
or U35914 (N_35914,N_32564,N_32649);
nor U35915 (N_35915,N_32925,N_34501);
xor U35916 (N_35916,N_34843,N_34809);
xnor U35917 (N_35917,N_34222,N_32805);
nand U35918 (N_35918,N_33528,N_34060);
or U35919 (N_35919,N_33799,N_33586);
xor U35920 (N_35920,N_33324,N_32663);
xor U35921 (N_35921,N_34114,N_34177);
and U35922 (N_35922,N_33060,N_34124);
xnor U35923 (N_35923,N_33521,N_33447);
or U35924 (N_35924,N_33993,N_33883);
nand U35925 (N_35925,N_33092,N_33788);
xnor U35926 (N_35926,N_34271,N_34093);
nor U35927 (N_35927,N_33510,N_33735);
nor U35928 (N_35928,N_34613,N_33476);
xor U35929 (N_35929,N_33598,N_32566);
and U35930 (N_35930,N_34428,N_32809);
xor U35931 (N_35931,N_32669,N_32592);
and U35932 (N_35932,N_33120,N_34953);
xnor U35933 (N_35933,N_33954,N_34507);
xnor U35934 (N_35934,N_33851,N_34351);
xnor U35935 (N_35935,N_33664,N_32714);
nand U35936 (N_35936,N_34591,N_34540);
xnor U35937 (N_35937,N_32978,N_34940);
nor U35938 (N_35938,N_32629,N_32547);
and U35939 (N_35939,N_34026,N_32540);
and U35940 (N_35940,N_33265,N_32997);
nand U35941 (N_35941,N_34483,N_32615);
nand U35942 (N_35942,N_33243,N_34402);
or U35943 (N_35943,N_34148,N_32935);
nand U35944 (N_35944,N_33985,N_33109);
xor U35945 (N_35945,N_34150,N_33620);
nand U35946 (N_35946,N_34432,N_34706);
or U35947 (N_35947,N_34197,N_34221);
nor U35948 (N_35948,N_34685,N_34264);
xnor U35949 (N_35949,N_33436,N_32943);
or U35950 (N_35950,N_34853,N_34499);
nand U35951 (N_35951,N_33818,N_33815);
or U35952 (N_35952,N_34013,N_33061);
xnor U35953 (N_35953,N_32887,N_33348);
nand U35954 (N_35954,N_33108,N_32670);
or U35955 (N_35955,N_33643,N_33922);
or U35956 (N_35956,N_34082,N_34986);
or U35957 (N_35957,N_33504,N_33552);
nor U35958 (N_35958,N_34846,N_34795);
or U35959 (N_35959,N_33274,N_34127);
nand U35960 (N_35960,N_33780,N_34849);
or U35961 (N_35961,N_32998,N_33204);
xnor U35962 (N_35962,N_33634,N_33522);
nand U35963 (N_35963,N_34448,N_34716);
or U35964 (N_35964,N_34753,N_33338);
nand U35965 (N_35965,N_33387,N_34267);
and U35966 (N_35966,N_33699,N_33886);
nand U35967 (N_35967,N_33333,N_32574);
and U35968 (N_35968,N_33033,N_32912);
xnor U35969 (N_35969,N_33712,N_33253);
or U35970 (N_35970,N_33296,N_33441);
nand U35971 (N_35971,N_34594,N_33863);
and U35972 (N_35972,N_34536,N_34445);
nor U35973 (N_35973,N_32842,N_32867);
or U35974 (N_35974,N_32708,N_34554);
nand U35975 (N_35975,N_34875,N_34250);
and U35976 (N_35976,N_32959,N_33462);
nor U35977 (N_35977,N_34120,N_32791);
xnor U35978 (N_35978,N_34838,N_33955);
nand U35979 (N_35979,N_32756,N_33518);
nor U35980 (N_35980,N_33537,N_33897);
and U35981 (N_35981,N_33248,N_33878);
and U35982 (N_35982,N_34498,N_34518);
xor U35983 (N_35983,N_33364,N_33771);
nand U35984 (N_35984,N_33848,N_33640);
nand U35985 (N_35985,N_32940,N_32939);
xor U35986 (N_35986,N_34565,N_34727);
nand U35987 (N_35987,N_32833,N_33373);
nor U35988 (N_35988,N_34200,N_34887);
and U35989 (N_35989,N_34649,N_32554);
and U35990 (N_35990,N_32894,N_32870);
and U35991 (N_35991,N_33677,N_32873);
nor U35992 (N_35992,N_33063,N_33081);
nand U35993 (N_35993,N_33117,N_34008);
or U35994 (N_35994,N_33037,N_33088);
xor U35995 (N_35995,N_33290,N_33612);
nor U35996 (N_35996,N_33341,N_33548);
or U35997 (N_35997,N_33754,N_32938);
xor U35998 (N_35998,N_34194,N_33836);
xnor U35999 (N_35999,N_34002,N_32928);
and U36000 (N_36000,N_32980,N_33036);
nor U36001 (N_36001,N_34359,N_33857);
or U36002 (N_36002,N_34786,N_33716);
xor U36003 (N_36003,N_34744,N_33231);
nor U36004 (N_36004,N_33390,N_32946);
nor U36005 (N_36005,N_33004,N_33163);
nand U36006 (N_36006,N_34228,N_33198);
or U36007 (N_36007,N_33309,N_33923);
xor U36008 (N_36008,N_33774,N_33783);
or U36009 (N_36009,N_34743,N_33607);
nor U36010 (N_36010,N_34842,N_33523);
or U36011 (N_36011,N_34804,N_33576);
nand U36012 (N_36012,N_33803,N_33715);
or U36013 (N_36013,N_34626,N_33082);
and U36014 (N_36014,N_33214,N_34343);
xor U36015 (N_36015,N_34237,N_34401);
and U36016 (N_36016,N_34885,N_34566);
xnor U36017 (N_36017,N_33882,N_33423);
or U36018 (N_36018,N_34771,N_34169);
xnor U36019 (N_36019,N_34496,N_34772);
nand U36020 (N_36020,N_34354,N_34145);
xnor U36021 (N_36021,N_34376,N_34089);
nor U36022 (N_36022,N_34162,N_33381);
nand U36023 (N_36023,N_34971,N_33089);
xor U36024 (N_36024,N_32589,N_32641);
xnor U36025 (N_36025,N_34510,N_34583);
or U36026 (N_36026,N_33772,N_34503);
xnor U36027 (N_36027,N_33763,N_34506);
nor U36028 (N_36028,N_34164,N_33746);
nor U36029 (N_36029,N_33697,N_33134);
xnor U36030 (N_36030,N_34235,N_32613);
or U36031 (N_36031,N_34388,N_34654);
xnor U36032 (N_36032,N_33862,N_34680);
nand U36033 (N_36033,N_32518,N_32605);
xnor U36034 (N_36034,N_33416,N_33512);
and U36035 (N_36035,N_34961,N_33358);
nor U36036 (N_36036,N_33396,N_33199);
and U36037 (N_36037,N_32521,N_32509);
nor U36038 (N_36038,N_33139,N_34634);
or U36039 (N_36039,N_34535,N_33709);
or U36040 (N_36040,N_34185,N_34812);
nand U36041 (N_36041,N_32810,N_32755);
or U36042 (N_36042,N_34326,N_34274);
xor U36043 (N_36043,N_34037,N_34925);
nand U36044 (N_36044,N_33765,N_32985);
nor U36045 (N_36045,N_32921,N_34452);
xnor U36046 (N_36046,N_33850,N_33758);
xnor U36047 (N_36047,N_34459,N_32797);
nor U36048 (N_36048,N_34438,N_33917);
or U36049 (N_36049,N_34945,N_33292);
nand U36050 (N_36050,N_32519,N_32986);
nor U36051 (N_36051,N_34389,N_34293);
and U36052 (N_36052,N_32581,N_34017);
or U36053 (N_36053,N_33415,N_33834);
nor U36054 (N_36054,N_34542,N_32875);
and U36055 (N_36055,N_33657,N_32834);
xnor U36056 (N_36056,N_33775,N_33095);
xnor U36057 (N_36057,N_33370,N_32927);
nor U36058 (N_36058,N_32694,N_34548);
and U36059 (N_36059,N_34482,N_32725);
nand U36060 (N_36060,N_34178,N_34485);
nor U36061 (N_36061,N_32936,N_32763);
nand U36062 (N_36062,N_33080,N_34580);
xnor U36063 (N_36063,N_33670,N_32818);
or U36064 (N_36064,N_33719,N_33362);
xnor U36065 (N_36065,N_34761,N_33767);
nand U36066 (N_36066,N_33911,N_34173);
or U36067 (N_36067,N_33885,N_34574);
and U36068 (N_36068,N_34544,N_34158);
nand U36069 (N_36069,N_34597,N_34308);
and U36070 (N_36070,N_32759,N_33550);
or U36071 (N_36071,N_32782,N_33369);
nor U36072 (N_36072,N_34883,N_33892);
nand U36073 (N_36073,N_32501,N_34684);
or U36074 (N_36074,N_33814,N_32544);
nand U36075 (N_36075,N_32517,N_34469);
nand U36076 (N_36076,N_33766,N_34370);
and U36077 (N_36077,N_34160,N_33263);
or U36078 (N_36078,N_32825,N_33189);
and U36079 (N_36079,N_33271,N_33024);
nand U36080 (N_36080,N_34375,N_33641);
nand U36081 (N_36081,N_33359,N_33872);
nand U36082 (N_36082,N_34787,N_32911);
nor U36083 (N_36083,N_33825,N_34065);
and U36084 (N_36084,N_32689,N_33481);
or U36085 (N_36085,N_33018,N_34766);
and U36086 (N_36086,N_32508,N_32990);
or U36087 (N_36087,N_32994,N_32510);
xnor U36088 (N_36088,N_34063,N_34101);
or U36089 (N_36089,N_32862,N_33325);
xnor U36090 (N_36090,N_34218,N_32624);
and U36091 (N_36091,N_34307,N_32968);
nand U36092 (N_36092,N_33837,N_34990);
nor U36093 (N_36093,N_34543,N_34451);
nor U36094 (N_36094,N_33562,N_33571);
xnor U36095 (N_36095,N_34865,N_34807);
or U36096 (N_36096,N_34007,N_33172);
or U36097 (N_36097,N_34425,N_34549);
nor U36098 (N_36098,N_34058,N_32941);
or U36099 (N_36099,N_34306,N_33101);
xnor U36100 (N_36100,N_33321,N_32637);
nand U36101 (N_36101,N_32977,N_33722);
nor U36102 (N_36102,N_33445,N_32648);
and U36103 (N_36103,N_34193,N_34287);
and U36104 (N_36104,N_32754,N_33801);
nor U36105 (N_36105,N_34395,N_33969);
nor U36106 (N_36106,N_34371,N_33449);
xor U36107 (N_36107,N_34551,N_34589);
xor U36108 (N_36108,N_34959,N_33067);
or U36109 (N_36109,N_33014,N_34163);
and U36110 (N_36110,N_34165,N_34526);
nor U36111 (N_36111,N_34102,N_33645);
and U36112 (N_36112,N_33414,N_32962);
nor U36113 (N_36113,N_34024,N_34564);
nand U36114 (N_36114,N_33511,N_32773);
and U36115 (N_36115,N_33162,N_33255);
or U36116 (N_36116,N_33422,N_34329);
or U36117 (N_36117,N_33962,N_34283);
or U36118 (N_36118,N_34712,N_34912);
nand U36119 (N_36119,N_34286,N_33517);
xnor U36120 (N_36120,N_34337,N_34132);
xnor U36121 (N_36121,N_34099,N_33471);
or U36122 (N_36122,N_34261,N_34004);
and U36123 (N_36123,N_32569,N_33459);
nor U36124 (N_36124,N_32947,N_34983);
or U36125 (N_36125,N_33474,N_33675);
nand U36126 (N_36126,N_34032,N_34802);
or U36127 (N_36127,N_34486,N_33408);
nand U36128 (N_36128,N_34281,N_33960);
and U36129 (N_36129,N_33889,N_34775);
nor U36130 (N_36130,N_34617,N_33773);
nand U36131 (N_36131,N_34435,N_34650);
nor U36132 (N_36132,N_33238,N_34478);
xor U36133 (N_36133,N_34263,N_33866);
nand U36134 (N_36134,N_34805,N_32907);
or U36135 (N_36135,N_32811,N_34166);
or U36136 (N_36136,N_33226,N_32877);
nand U36137 (N_36137,N_34103,N_34822);
nand U36138 (N_36138,N_34361,N_34645);
xor U36139 (N_36139,N_34531,N_32553);
nor U36140 (N_36140,N_32916,N_32829);
nor U36141 (N_36141,N_32819,N_32757);
xor U36142 (N_36142,N_34576,N_33401);
or U36143 (N_36143,N_33579,N_34642);
or U36144 (N_36144,N_33306,N_34638);
xnor U36145 (N_36145,N_34119,N_33062);
nor U36146 (N_36146,N_32552,N_34111);
or U36147 (N_36147,N_33404,N_34135);
or U36148 (N_36148,N_33239,N_33692);
xor U36149 (N_36149,N_32929,N_33155);
or U36150 (N_36150,N_34245,N_34968);
xor U36151 (N_36151,N_33130,N_33782);
or U36152 (N_36152,N_33277,N_33786);
or U36153 (N_36153,N_33533,N_33355);
nand U36154 (N_36154,N_33802,N_34852);
xor U36155 (N_36155,N_34473,N_33973);
xnor U36156 (N_36156,N_32871,N_32914);
nor U36157 (N_36157,N_34508,N_33463);
nor U36158 (N_36158,N_33027,N_32973);
or U36159 (N_36159,N_33264,N_33957);
and U36160 (N_36160,N_33218,N_33342);
nand U36161 (N_36161,N_34860,N_33514);
xnor U36162 (N_36162,N_33346,N_33527);
and U36163 (N_36163,N_32762,N_32889);
and U36164 (N_36164,N_32798,N_34834);
nand U36165 (N_36165,N_33291,N_34949);
xor U36166 (N_36166,N_34915,N_32775);
nor U36167 (N_36167,N_33222,N_33729);
xnor U36168 (N_36168,N_34154,N_32542);
and U36169 (N_36169,N_34303,N_33367);
xnor U36170 (N_36170,N_33768,N_33114);
nor U36171 (N_36171,N_33038,N_33072);
nand U36172 (N_36172,N_33966,N_33058);
xor U36173 (N_36173,N_34233,N_34906);
and U36174 (N_36174,N_33302,N_34896);
and U36175 (N_36175,N_34696,N_32785);
nand U36176 (N_36176,N_32538,N_33322);
and U36177 (N_36177,N_32890,N_33749);
nor U36178 (N_36178,N_34423,N_34190);
nor U36179 (N_36179,N_32531,N_34871);
and U36180 (N_36180,N_34790,N_34737);
nand U36181 (N_36181,N_33564,N_33789);
or U36182 (N_36182,N_34406,N_33580);
nor U36183 (N_36183,N_33584,N_34141);
nor U36184 (N_36184,N_33213,N_34601);
nand U36185 (N_36185,N_33581,N_34909);
nand U36186 (N_36186,N_34999,N_34357);
or U36187 (N_36187,N_34196,N_33046);
and U36188 (N_36188,N_32808,N_32957);
and U36189 (N_36189,N_33220,N_34929);
or U36190 (N_36190,N_33094,N_34516);
xnor U36191 (N_36191,N_34662,N_33759);
nor U36192 (N_36192,N_34675,N_33353);
or U36193 (N_36193,N_33502,N_33393);
and U36194 (N_36194,N_34892,N_32522);
nand U36195 (N_36195,N_33905,N_34392);
and U36196 (N_36196,N_33453,N_33939);
or U36197 (N_36197,N_32903,N_34470);
and U36198 (N_36198,N_33485,N_33472);
or U36199 (N_36199,N_34927,N_32856);
xor U36200 (N_36200,N_34533,N_34399);
nor U36201 (N_36201,N_32585,N_33438);
nand U36202 (N_36202,N_34976,N_34768);
nand U36203 (N_36203,N_33817,N_33952);
and U36204 (N_36204,N_34770,N_33596);
nor U36205 (N_36205,N_32560,N_33386);
and U36206 (N_36206,N_32932,N_33929);
or U36207 (N_36207,N_33924,N_34981);
nand U36208 (N_36208,N_32816,N_32848);
and U36209 (N_36209,N_32858,N_33937);
nor U36210 (N_36210,N_33996,N_34707);
nand U36211 (N_36211,N_33219,N_32644);
nand U36212 (N_36212,N_32576,N_33900);
xnor U36213 (N_36213,N_34491,N_33555);
xor U36214 (N_36214,N_34965,N_33319);
nand U36215 (N_36215,N_34336,N_34621);
nor U36216 (N_36216,N_34511,N_34117);
xor U36217 (N_36217,N_34175,N_33110);
and U36218 (N_36218,N_34234,N_32558);
or U36219 (N_36219,N_34094,N_33069);
and U36220 (N_36220,N_32761,N_32988);
nor U36221 (N_36221,N_33832,N_34118);
nand U36222 (N_36222,N_34776,N_32500);
nor U36223 (N_36223,N_34847,N_34053);
and U36224 (N_36224,N_33465,N_33287);
or U36225 (N_36225,N_33273,N_34211);
and U36226 (N_36226,N_33587,N_34051);
or U36227 (N_36227,N_33927,N_32920);
nor U36228 (N_36228,N_34623,N_33526);
xnor U36229 (N_36229,N_34870,N_34128);
nand U36230 (N_36230,N_34468,N_34969);
nor U36231 (N_36231,N_34552,N_33276);
nor U36232 (N_36232,N_33532,N_34873);
or U36233 (N_36233,N_34545,N_32723);
nor U36234 (N_36234,N_32752,N_34061);
and U36235 (N_36235,N_34814,N_33648);
nand U36236 (N_36236,N_34527,N_33506);
or U36237 (N_36237,N_34268,N_34368);
or U36238 (N_36238,N_33971,N_34748);
nand U36239 (N_36239,N_34910,N_32744);
nand U36240 (N_36240,N_33009,N_33334);
and U36241 (N_36241,N_33912,N_32563);
nor U36242 (N_36242,N_32630,N_33846);
or U36243 (N_36243,N_34176,N_33495);
nand U36244 (N_36244,N_32845,N_32618);
xor U36245 (N_36245,N_33984,N_33259);
nor U36246 (N_36246,N_32795,N_34741);
nor U36247 (N_36247,N_33932,N_34188);
and U36248 (N_36248,N_33616,N_33377);
nand U36249 (N_36249,N_33880,N_32556);
or U36250 (N_36250,N_33662,N_33965);
and U36251 (N_36251,N_32647,N_33529);
nand U36252 (N_36252,N_32781,N_33857);
nor U36253 (N_36253,N_33749,N_33213);
nor U36254 (N_36254,N_33282,N_33130);
nand U36255 (N_36255,N_34220,N_32674);
xor U36256 (N_36256,N_34227,N_32865);
xnor U36257 (N_36257,N_34906,N_33403);
xor U36258 (N_36258,N_33655,N_34026);
and U36259 (N_36259,N_33508,N_34288);
and U36260 (N_36260,N_34529,N_34863);
xor U36261 (N_36261,N_32728,N_33721);
nor U36262 (N_36262,N_33713,N_33308);
nand U36263 (N_36263,N_34111,N_32917);
and U36264 (N_36264,N_33098,N_33911);
or U36265 (N_36265,N_33866,N_34364);
and U36266 (N_36266,N_34060,N_34700);
and U36267 (N_36267,N_33684,N_33439);
nor U36268 (N_36268,N_33434,N_32519);
nor U36269 (N_36269,N_34720,N_34124);
xor U36270 (N_36270,N_34677,N_33417);
nand U36271 (N_36271,N_33400,N_34703);
nand U36272 (N_36272,N_34811,N_33137);
and U36273 (N_36273,N_34469,N_33900);
and U36274 (N_36274,N_34627,N_32511);
xnor U36275 (N_36275,N_32860,N_33615);
xor U36276 (N_36276,N_34158,N_33764);
or U36277 (N_36277,N_33213,N_33371);
nor U36278 (N_36278,N_33721,N_33727);
and U36279 (N_36279,N_34086,N_33865);
nand U36280 (N_36280,N_33882,N_34335);
nand U36281 (N_36281,N_34656,N_32598);
or U36282 (N_36282,N_32783,N_34420);
nand U36283 (N_36283,N_33823,N_32980);
or U36284 (N_36284,N_32937,N_33836);
nor U36285 (N_36285,N_34398,N_33298);
nand U36286 (N_36286,N_33307,N_34281);
or U36287 (N_36287,N_34586,N_33834);
and U36288 (N_36288,N_32776,N_33478);
nor U36289 (N_36289,N_34338,N_33646);
and U36290 (N_36290,N_33446,N_34873);
and U36291 (N_36291,N_34213,N_33916);
xor U36292 (N_36292,N_34414,N_34116);
xor U36293 (N_36293,N_34474,N_33664);
or U36294 (N_36294,N_32973,N_32582);
and U36295 (N_36295,N_33152,N_33074);
nand U36296 (N_36296,N_34885,N_34827);
nor U36297 (N_36297,N_33319,N_33193);
xor U36298 (N_36298,N_34164,N_33013);
and U36299 (N_36299,N_33063,N_34376);
or U36300 (N_36300,N_32572,N_34453);
xor U36301 (N_36301,N_33636,N_34862);
xnor U36302 (N_36302,N_34990,N_33175);
nand U36303 (N_36303,N_34908,N_32849);
nor U36304 (N_36304,N_33366,N_34778);
or U36305 (N_36305,N_32678,N_34561);
and U36306 (N_36306,N_33720,N_33704);
or U36307 (N_36307,N_33415,N_32787);
or U36308 (N_36308,N_33038,N_34486);
nor U36309 (N_36309,N_32724,N_33460);
xnor U36310 (N_36310,N_32749,N_34806);
xor U36311 (N_36311,N_33534,N_34557);
nor U36312 (N_36312,N_32825,N_32854);
nand U36313 (N_36313,N_34515,N_33195);
xnor U36314 (N_36314,N_33977,N_33455);
xnor U36315 (N_36315,N_33682,N_34739);
nand U36316 (N_36316,N_32534,N_33629);
and U36317 (N_36317,N_34430,N_33603);
nand U36318 (N_36318,N_34169,N_34278);
nor U36319 (N_36319,N_32701,N_34269);
nor U36320 (N_36320,N_33378,N_34448);
nor U36321 (N_36321,N_32625,N_33361);
or U36322 (N_36322,N_34163,N_32823);
and U36323 (N_36323,N_32767,N_33683);
or U36324 (N_36324,N_34812,N_34557);
nor U36325 (N_36325,N_33347,N_32858);
nor U36326 (N_36326,N_33983,N_33169);
and U36327 (N_36327,N_33896,N_32670);
xnor U36328 (N_36328,N_33823,N_33292);
nand U36329 (N_36329,N_34594,N_32729);
nand U36330 (N_36330,N_32602,N_33851);
and U36331 (N_36331,N_34314,N_34475);
nand U36332 (N_36332,N_33198,N_32564);
and U36333 (N_36333,N_34976,N_33557);
nand U36334 (N_36334,N_33809,N_32723);
nand U36335 (N_36335,N_32811,N_34634);
nand U36336 (N_36336,N_34931,N_34929);
nand U36337 (N_36337,N_33372,N_34767);
and U36338 (N_36338,N_34197,N_32782);
nor U36339 (N_36339,N_33971,N_34359);
and U36340 (N_36340,N_33684,N_33947);
or U36341 (N_36341,N_32815,N_34865);
or U36342 (N_36342,N_32749,N_33372);
and U36343 (N_36343,N_32911,N_33588);
nor U36344 (N_36344,N_32675,N_32597);
nand U36345 (N_36345,N_34548,N_32726);
or U36346 (N_36346,N_34048,N_34015);
or U36347 (N_36347,N_33897,N_33485);
xor U36348 (N_36348,N_33607,N_32685);
and U36349 (N_36349,N_33091,N_33281);
nand U36350 (N_36350,N_33692,N_33416);
xor U36351 (N_36351,N_33917,N_33515);
xor U36352 (N_36352,N_34467,N_33272);
or U36353 (N_36353,N_33377,N_32857);
and U36354 (N_36354,N_32980,N_32570);
nand U36355 (N_36355,N_32857,N_34861);
or U36356 (N_36356,N_32786,N_34632);
and U36357 (N_36357,N_33984,N_34602);
nor U36358 (N_36358,N_33439,N_32755);
nand U36359 (N_36359,N_32717,N_34526);
nor U36360 (N_36360,N_34537,N_32700);
or U36361 (N_36361,N_33079,N_32665);
nor U36362 (N_36362,N_34160,N_34373);
xor U36363 (N_36363,N_34489,N_34321);
nand U36364 (N_36364,N_32995,N_34100);
nand U36365 (N_36365,N_33917,N_34410);
xor U36366 (N_36366,N_33203,N_34423);
xnor U36367 (N_36367,N_32538,N_32993);
nand U36368 (N_36368,N_34819,N_34189);
or U36369 (N_36369,N_34783,N_33170);
xnor U36370 (N_36370,N_33221,N_32752);
nor U36371 (N_36371,N_34093,N_34350);
xnor U36372 (N_36372,N_32852,N_33426);
xnor U36373 (N_36373,N_32680,N_34478);
xor U36374 (N_36374,N_34316,N_33822);
nor U36375 (N_36375,N_34011,N_34032);
and U36376 (N_36376,N_32511,N_34458);
xnor U36377 (N_36377,N_33471,N_34165);
nand U36378 (N_36378,N_33879,N_33568);
or U36379 (N_36379,N_32814,N_34260);
and U36380 (N_36380,N_32591,N_34947);
or U36381 (N_36381,N_34632,N_34988);
nor U36382 (N_36382,N_33992,N_34214);
or U36383 (N_36383,N_33527,N_33606);
or U36384 (N_36384,N_33276,N_33272);
nor U36385 (N_36385,N_34864,N_33621);
or U36386 (N_36386,N_33418,N_33717);
or U36387 (N_36387,N_33911,N_33157);
and U36388 (N_36388,N_33760,N_33603);
xnor U36389 (N_36389,N_33149,N_34701);
xnor U36390 (N_36390,N_33423,N_32780);
xnor U36391 (N_36391,N_34263,N_33856);
and U36392 (N_36392,N_32785,N_34104);
xnor U36393 (N_36393,N_33685,N_32619);
or U36394 (N_36394,N_33010,N_33155);
and U36395 (N_36395,N_34451,N_33810);
xor U36396 (N_36396,N_33371,N_33135);
or U36397 (N_36397,N_34126,N_33475);
nand U36398 (N_36398,N_33874,N_34267);
or U36399 (N_36399,N_32509,N_33654);
nand U36400 (N_36400,N_32608,N_34511);
or U36401 (N_36401,N_33327,N_34528);
nand U36402 (N_36402,N_34260,N_33227);
xor U36403 (N_36403,N_34317,N_32628);
and U36404 (N_36404,N_34466,N_33543);
and U36405 (N_36405,N_33009,N_34306);
and U36406 (N_36406,N_32725,N_32788);
nor U36407 (N_36407,N_34393,N_32989);
or U36408 (N_36408,N_34092,N_33455);
xor U36409 (N_36409,N_32721,N_34782);
xnor U36410 (N_36410,N_33228,N_32785);
nand U36411 (N_36411,N_33500,N_34900);
nor U36412 (N_36412,N_33175,N_32503);
xnor U36413 (N_36413,N_34138,N_33202);
nand U36414 (N_36414,N_34023,N_34984);
or U36415 (N_36415,N_32541,N_34310);
and U36416 (N_36416,N_33401,N_34382);
nor U36417 (N_36417,N_32867,N_34918);
xor U36418 (N_36418,N_32568,N_34022);
and U36419 (N_36419,N_34240,N_33199);
nand U36420 (N_36420,N_33585,N_33813);
xnor U36421 (N_36421,N_33678,N_33631);
and U36422 (N_36422,N_34641,N_34403);
or U36423 (N_36423,N_34712,N_34665);
and U36424 (N_36424,N_32924,N_34585);
xor U36425 (N_36425,N_34039,N_34308);
nor U36426 (N_36426,N_34175,N_32543);
nand U36427 (N_36427,N_32899,N_34604);
xnor U36428 (N_36428,N_33443,N_33263);
and U36429 (N_36429,N_33968,N_34819);
nand U36430 (N_36430,N_33597,N_34466);
nor U36431 (N_36431,N_34577,N_33083);
or U36432 (N_36432,N_34451,N_32881);
xor U36433 (N_36433,N_34530,N_33674);
nand U36434 (N_36434,N_33654,N_33032);
nor U36435 (N_36435,N_34399,N_32640);
or U36436 (N_36436,N_32968,N_34358);
and U36437 (N_36437,N_33522,N_34794);
or U36438 (N_36438,N_33529,N_34286);
and U36439 (N_36439,N_34640,N_33590);
and U36440 (N_36440,N_34298,N_32880);
nor U36441 (N_36441,N_32676,N_34868);
or U36442 (N_36442,N_32642,N_34892);
xnor U36443 (N_36443,N_32602,N_34230);
nor U36444 (N_36444,N_34784,N_34309);
and U36445 (N_36445,N_32684,N_33809);
and U36446 (N_36446,N_33287,N_34806);
xnor U36447 (N_36447,N_33321,N_33687);
or U36448 (N_36448,N_34676,N_34819);
xnor U36449 (N_36449,N_33340,N_34497);
nand U36450 (N_36450,N_32600,N_34012);
nor U36451 (N_36451,N_33932,N_33552);
and U36452 (N_36452,N_32714,N_33454);
nand U36453 (N_36453,N_34290,N_34615);
and U36454 (N_36454,N_32978,N_33343);
and U36455 (N_36455,N_34160,N_34620);
or U36456 (N_36456,N_34914,N_34137);
or U36457 (N_36457,N_34034,N_34485);
nand U36458 (N_36458,N_34677,N_33541);
nand U36459 (N_36459,N_34394,N_32823);
nand U36460 (N_36460,N_32906,N_34907);
or U36461 (N_36461,N_34482,N_33789);
nand U36462 (N_36462,N_34476,N_34916);
or U36463 (N_36463,N_32783,N_32577);
nor U36464 (N_36464,N_34833,N_34995);
nor U36465 (N_36465,N_32894,N_33431);
or U36466 (N_36466,N_32643,N_34156);
xnor U36467 (N_36467,N_34762,N_34946);
xnor U36468 (N_36468,N_33461,N_33574);
and U36469 (N_36469,N_33234,N_33990);
and U36470 (N_36470,N_33239,N_33947);
xnor U36471 (N_36471,N_34493,N_34558);
xor U36472 (N_36472,N_33909,N_34782);
xnor U36473 (N_36473,N_33183,N_33826);
xnor U36474 (N_36474,N_34438,N_34601);
nor U36475 (N_36475,N_34475,N_34682);
nand U36476 (N_36476,N_33700,N_33814);
nor U36477 (N_36477,N_33777,N_34086);
or U36478 (N_36478,N_34990,N_33938);
nand U36479 (N_36479,N_34996,N_34604);
nand U36480 (N_36480,N_32748,N_34613);
nor U36481 (N_36481,N_34353,N_34825);
nand U36482 (N_36482,N_34485,N_33330);
nor U36483 (N_36483,N_33006,N_32888);
nor U36484 (N_36484,N_33177,N_34493);
nor U36485 (N_36485,N_34172,N_33085);
xor U36486 (N_36486,N_33407,N_34646);
nor U36487 (N_36487,N_33174,N_34318);
and U36488 (N_36488,N_34826,N_33039);
or U36489 (N_36489,N_33617,N_33592);
xnor U36490 (N_36490,N_34941,N_33984);
nor U36491 (N_36491,N_33804,N_33852);
nand U36492 (N_36492,N_32527,N_32926);
or U36493 (N_36493,N_32867,N_33296);
nand U36494 (N_36494,N_34158,N_32978);
nor U36495 (N_36495,N_34306,N_32823);
nor U36496 (N_36496,N_33995,N_34745);
nand U36497 (N_36497,N_34613,N_32760);
nand U36498 (N_36498,N_33807,N_33590);
or U36499 (N_36499,N_34284,N_34164);
nand U36500 (N_36500,N_34142,N_34514);
and U36501 (N_36501,N_34073,N_34116);
xnor U36502 (N_36502,N_32896,N_33094);
or U36503 (N_36503,N_33612,N_33388);
and U36504 (N_36504,N_34229,N_32666);
nand U36505 (N_36505,N_34155,N_34628);
nand U36506 (N_36506,N_33763,N_34567);
nor U36507 (N_36507,N_32557,N_33138);
and U36508 (N_36508,N_34857,N_34937);
or U36509 (N_36509,N_33316,N_33367);
nand U36510 (N_36510,N_34136,N_34315);
nand U36511 (N_36511,N_32538,N_32772);
and U36512 (N_36512,N_34761,N_32565);
and U36513 (N_36513,N_34436,N_33723);
or U36514 (N_36514,N_33992,N_33678);
nor U36515 (N_36515,N_34821,N_33380);
nand U36516 (N_36516,N_32867,N_32930);
nand U36517 (N_36517,N_33166,N_34292);
or U36518 (N_36518,N_33885,N_33097);
or U36519 (N_36519,N_33620,N_33804);
xnor U36520 (N_36520,N_33201,N_33337);
nor U36521 (N_36521,N_34905,N_34432);
nor U36522 (N_36522,N_32799,N_32972);
xor U36523 (N_36523,N_34387,N_34970);
and U36524 (N_36524,N_34854,N_34920);
xor U36525 (N_36525,N_33027,N_32502);
and U36526 (N_36526,N_34184,N_33428);
xnor U36527 (N_36527,N_33454,N_33671);
xor U36528 (N_36528,N_33995,N_32803);
or U36529 (N_36529,N_34674,N_34136);
nor U36530 (N_36530,N_32894,N_33982);
or U36531 (N_36531,N_33396,N_34540);
and U36532 (N_36532,N_33585,N_33841);
nor U36533 (N_36533,N_34839,N_32514);
or U36534 (N_36534,N_32678,N_32584);
nor U36535 (N_36535,N_34132,N_33313);
nand U36536 (N_36536,N_34767,N_33816);
nand U36537 (N_36537,N_34547,N_34809);
or U36538 (N_36538,N_34112,N_32701);
or U36539 (N_36539,N_34923,N_34050);
xnor U36540 (N_36540,N_34792,N_33761);
nand U36541 (N_36541,N_33571,N_33494);
nand U36542 (N_36542,N_32570,N_32679);
and U36543 (N_36543,N_32672,N_33869);
nand U36544 (N_36544,N_32639,N_34316);
nand U36545 (N_36545,N_32787,N_33372);
or U36546 (N_36546,N_34099,N_33774);
nand U36547 (N_36547,N_34964,N_32868);
and U36548 (N_36548,N_32934,N_34772);
nand U36549 (N_36549,N_33227,N_33737);
nor U36550 (N_36550,N_34035,N_33438);
or U36551 (N_36551,N_33317,N_34106);
xnor U36552 (N_36552,N_33127,N_34957);
xor U36553 (N_36553,N_33094,N_33909);
or U36554 (N_36554,N_34384,N_34589);
and U36555 (N_36555,N_33056,N_34973);
nor U36556 (N_36556,N_34406,N_33410);
xor U36557 (N_36557,N_34841,N_34887);
and U36558 (N_36558,N_34155,N_34643);
xor U36559 (N_36559,N_33569,N_32823);
xor U36560 (N_36560,N_34485,N_34386);
nor U36561 (N_36561,N_32713,N_32793);
nand U36562 (N_36562,N_32766,N_33753);
or U36563 (N_36563,N_33891,N_34291);
xnor U36564 (N_36564,N_32709,N_32799);
xor U36565 (N_36565,N_33256,N_32521);
and U36566 (N_36566,N_34336,N_32643);
nand U36567 (N_36567,N_34390,N_33227);
nor U36568 (N_36568,N_34488,N_33095);
or U36569 (N_36569,N_34472,N_34586);
or U36570 (N_36570,N_32695,N_32628);
or U36571 (N_36571,N_34176,N_33785);
and U36572 (N_36572,N_34305,N_32867);
and U36573 (N_36573,N_33992,N_32768);
xor U36574 (N_36574,N_33233,N_33117);
or U36575 (N_36575,N_34795,N_33698);
xor U36576 (N_36576,N_32565,N_32510);
and U36577 (N_36577,N_32944,N_33594);
or U36578 (N_36578,N_33731,N_34009);
xnor U36579 (N_36579,N_33247,N_33344);
or U36580 (N_36580,N_33262,N_33806);
xor U36581 (N_36581,N_33596,N_32912);
and U36582 (N_36582,N_33155,N_32931);
or U36583 (N_36583,N_34559,N_33011);
and U36584 (N_36584,N_32776,N_33029);
xor U36585 (N_36585,N_34744,N_32846);
nand U36586 (N_36586,N_33085,N_34741);
xor U36587 (N_36587,N_32890,N_34054);
and U36588 (N_36588,N_34674,N_33563);
xnor U36589 (N_36589,N_34808,N_34040);
xnor U36590 (N_36590,N_32946,N_33665);
nor U36591 (N_36591,N_33710,N_33787);
nor U36592 (N_36592,N_33427,N_33789);
and U36593 (N_36593,N_34639,N_33435);
nand U36594 (N_36594,N_34749,N_34214);
or U36595 (N_36595,N_34478,N_34447);
and U36596 (N_36596,N_33709,N_34248);
and U36597 (N_36597,N_32728,N_33608);
and U36598 (N_36598,N_32689,N_34164);
xor U36599 (N_36599,N_32790,N_33093);
nand U36600 (N_36600,N_34948,N_33912);
or U36601 (N_36601,N_33636,N_33194);
and U36602 (N_36602,N_33815,N_33233);
xor U36603 (N_36603,N_32916,N_33140);
and U36604 (N_36604,N_33951,N_34152);
xnor U36605 (N_36605,N_32641,N_32987);
xnor U36606 (N_36606,N_34428,N_34665);
nand U36607 (N_36607,N_32873,N_34389);
or U36608 (N_36608,N_34246,N_34202);
and U36609 (N_36609,N_33431,N_33300);
nand U36610 (N_36610,N_33718,N_34656);
and U36611 (N_36611,N_33896,N_33029);
nand U36612 (N_36612,N_34340,N_34182);
nor U36613 (N_36613,N_32544,N_33473);
xor U36614 (N_36614,N_33408,N_34656);
and U36615 (N_36615,N_34935,N_34973);
xnor U36616 (N_36616,N_33618,N_34039);
and U36617 (N_36617,N_33889,N_34576);
xor U36618 (N_36618,N_33345,N_33052);
and U36619 (N_36619,N_34188,N_34111);
or U36620 (N_36620,N_33793,N_34161);
nand U36621 (N_36621,N_32813,N_33831);
nand U36622 (N_36622,N_33914,N_34002);
nand U36623 (N_36623,N_34447,N_34127);
nor U36624 (N_36624,N_34612,N_33302);
and U36625 (N_36625,N_33337,N_34090);
xor U36626 (N_36626,N_34436,N_34255);
and U36627 (N_36627,N_33421,N_33666);
nor U36628 (N_36628,N_32532,N_33567);
nand U36629 (N_36629,N_34200,N_34282);
nand U36630 (N_36630,N_33777,N_34746);
nand U36631 (N_36631,N_33939,N_34166);
nor U36632 (N_36632,N_32875,N_33245);
xor U36633 (N_36633,N_34082,N_32867);
xor U36634 (N_36634,N_33488,N_32727);
nand U36635 (N_36635,N_33241,N_34065);
xor U36636 (N_36636,N_34686,N_33473);
or U36637 (N_36637,N_33923,N_33549);
or U36638 (N_36638,N_33484,N_32732);
and U36639 (N_36639,N_34132,N_34167);
and U36640 (N_36640,N_32996,N_33662);
or U36641 (N_36641,N_33104,N_33661);
nor U36642 (N_36642,N_33534,N_32668);
and U36643 (N_36643,N_34875,N_32675);
nor U36644 (N_36644,N_34139,N_33540);
and U36645 (N_36645,N_34913,N_34030);
and U36646 (N_36646,N_34250,N_33652);
and U36647 (N_36647,N_34306,N_34420);
nor U36648 (N_36648,N_34217,N_33480);
or U36649 (N_36649,N_33631,N_33753);
nor U36650 (N_36650,N_32812,N_32827);
nand U36651 (N_36651,N_33660,N_34354);
nand U36652 (N_36652,N_34301,N_34709);
nand U36653 (N_36653,N_33736,N_34280);
nand U36654 (N_36654,N_33107,N_32873);
and U36655 (N_36655,N_32699,N_33443);
and U36656 (N_36656,N_34007,N_33963);
nor U36657 (N_36657,N_34426,N_32506);
xor U36658 (N_36658,N_33136,N_32896);
or U36659 (N_36659,N_32737,N_34747);
xnor U36660 (N_36660,N_33852,N_33327);
xnor U36661 (N_36661,N_32752,N_34352);
or U36662 (N_36662,N_34216,N_34486);
and U36663 (N_36663,N_34901,N_33835);
or U36664 (N_36664,N_32543,N_33826);
and U36665 (N_36665,N_33292,N_33593);
and U36666 (N_36666,N_34134,N_33769);
nor U36667 (N_36667,N_32863,N_32858);
nor U36668 (N_36668,N_34925,N_34848);
xnor U36669 (N_36669,N_33996,N_33925);
or U36670 (N_36670,N_33051,N_33722);
or U36671 (N_36671,N_33004,N_34098);
and U36672 (N_36672,N_33813,N_34526);
and U36673 (N_36673,N_33254,N_34662);
nand U36674 (N_36674,N_34356,N_34838);
xor U36675 (N_36675,N_33167,N_32533);
xor U36676 (N_36676,N_34812,N_34342);
or U36677 (N_36677,N_34389,N_32799);
or U36678 (N_36678,N_33208,N_32727);
nand U36679 (N_36679,N_33952,N_34963);
nand U36680 (N_36680,N_33088,N_34261);
xnor U36681 (N_36681,N_33405,N_34901);
nand U36682 (N_36682,N_32922,N_34381);
nor U36683 (N_36683,N_33083,N_33369);
or U36684 (N_36684,N_33876,N_32766);
or U36685 (N_36685,N_32592,N_32997);
nor U36686 (N_36686,N_34785,N_32990);
or U36687 (N_36687,N_34533,N_34363);
xnor U36688 (N_36688,N_34196,N_34191);
or U36689 (N_36689,N_33165,N_34131);
or U36690 (N_36690,N_34830,N_33023);
nand U36691 (N_36691,N_33699,N_33184);
or U36692 (N_36692,N_32976,N_33838);
or U36693 (N_36693,N_34602,N_33336);
and U36694 (N_36694,N_33200,N_34154);
nand U36695 (N_36695,N_32970,N_32981);
xor U36696 (N_36696,N_32713,N_33022);
nand U36697 (N_36697,N_33862,N_32910);
or U36698 (N_36698,N_32830,N_33122);
nor U36699 (N_36699,N_34740,N_33394);
and U36700 (N_36700,N_32969,N_33465);
or U36701 (N_36701,N_32892,N_33814);
and U36702 (N_36702,N_34963,N_33279);
xnor U36703 (N_36703,N_34201,N_32651);
nand U36704 (N_36704,N_34277,N_33770);
xnor U36705 (N_36705,N_34362,N_33405);
nand U36706 (N_36706,N_34977,N_33026);
and U36707 (N_36707,N_32939,N_34338);
xor U36708 (N_36708,N_34304,N_34805);
nand U36709 (N_36709,N_34589,N_34120);
nand U36710 (N_36710,N_34104,N_33791);
nor U36711 (N_36711,N_34818,N_33829);
or U36712 (N_36712,N_34602,N_34951);
nor U36713 (N_36713,N_33031,N_34338);
and U36714 (N_36714,N_33377,N_34964);
nand U36715 (N_36715,N_34119,N_32542);
nor U36716 (N_36716,N_32608,N_33032);
nand U36717 (N_36717,N_33972,N_34432);
and U36718 (N_36718,N_33691,N_33972);
or U36719 (N_36719,N_33377,N_34879);
xnor U36720 (N_36720,N_33397,N_34870);
and U36721 (N_36721,N_34893,N_32658);
or U36722 (N_36722,N_34761,N_34593);
nor U36723 (N_36723,N_32734,N_34827);
xnor U36724 (N_36724,N_33216,N_33641);
and U36725 (N_36725,N_33014,N_33226);
and U36726 (N_36726,N_33960,N_33220);
nand U36727 (N_36727,N_34977,N_34629);
or U36728 (N_36728,N_32828,N_34357);
and U36729 (N_36729,N_33397,N_33019);
nor U36730 (N_36730,N_34414,N_33417);
xor U36731 (N_36731,N_34897,N_32744);
or U36732 (N_36732,N_32617,N_33184);
xnor U36733 (N_36733,N_34396,N_34529);
nor U36734 (N_36734,N_34536,N_34342);
nor U36735 (N_36735,N_34812,N_34958);
or U36736 (N_36736,N_34755,N_33233);
xor U36737 (N_36737,N_34337,N_34791);
and U36738 (N_36738,N_32797,N_34012);
nand U36739 (N_36739,N_32700,N_32750);
and U36740 (N_36740,N_32707,N_32950);
or U36741 (N_36741,N_34216,N_33219);
nor U36742 (N_36742,N_34485,N_32877);
nor U36743 (N_36743,N_33968,N_34258);
nand U36744 (N_36744,N_34354,N_33156);
xor U36745 (N_36745,N_34533,N_32950);
or U36746 (N_36746,N_34959,N_32763);
or U36747 (N_36747,N_34393,N_33572);
or U36748 (N_36748,N_34670,N_34322);
nand U36749 (N_36749,N_34414,N_34719);
or U36750 (N_36750,N_33579,N_32796);
nor U36751 (N_36751,N_33779,N_33224);
nand U36752 (N_36752,N_33590,N_34324);
and U36753 (N_36753,N_33767,N_34516);
nor U36754 (N_36754,N_32545,N_33996);
nand U36755 (N_36755,N_33776,N_34331);
nand U36756 (N_36756,N_32975,N_32658);
and U36757 (N_36757,N_33213,N_34692);
nand U36758 (N_36758,N_34993,N_32670);
nand U36759 (N_36759,N_34758,N_34227);
nand U36760 (N_36760,N_32990,N_34853);
nand U36761 (N_36761,N_34711,N_34610);
xnor U36762 (N_36762,N_34272,N_33353);
and U36763 (N_36763,N_33849,N_34496);
xnor U36764 (N_36764,N_34080,N_33316);
nand U36765 (N_36765,N_33903,N_34108);
or U36766 (N_36766,N_32906,N_33814);
nor U36767 (N_36767,N_34322,N_33920);
or U36768 (N_36768,N_34870,N_33483);
and U36769 (N_36769,N_32602,N_32710);
xnor U36770 (N_36770,N_34376,N_34717);
xor U36771 (N_36771,N_34303,N_32851);
nand U36772 (N_36772,N_33038,N_34930);
nor U36773 (N_36773,N_34276,N_32525);
or U36774 (N_36774,N_34850,N_34246);
nand U36775 (N_36775,N_33987,N_33657);
and U36776 (N_36776,N_33907,N_34961);
nand U36777 (N_36777,N_32702,N_32698);
xnor U36778 (N_36778,N_34869,N_34352);
and U36779 (N_36779,N_32818,N_32615);
or U36780 (N_36780,N_33563,N_34096);
or U36781 (N_36781,N_34115,N_34808);
and U36782 (N_36782,N_34804,N_33720);
nor U36783 (N_36783,N_32768,N_32576);
xnor U36784 (N_36784,N_32736,N_34141);
xor U36785 (N_36785,N_32887,N_34224);
xor U36786 (N_36786,N_34706,N_33503);
and U36787 (N_36787,N_32820,N_34244);
and U36788 (N_36788,N_33666,N_34339);
xnor U36789 (N_36789,N_32669,N_33556);
or U36790 (N_36790,N_33108,N_34144);
or U36791 (N_36791,N_34986,N_32634);
and U36792 (N_36792,N_33659,N_34372);
nand U36793 (N_36793,N_34495,N_34138);
nand U36794 (N_36794,N_33946,N_33420);
or U36795 (N_36795,N_33775,N_32588);
nand U36796 (N_36796,N_33701,N_34105);
xnor U36797 (N_36797,N_33954,N_34694);
or U36798 (N_36798,N_34518,N_34751);
nor U36799 (N_36799,N_33111,N_33120);
and U36800 (N_36800,N_33000,N_34386);
xor U36801 (N_36801,N_32779,N_34221);
and U36802 (N_36802,N_32654,N_32666);
or U36803 (N_36803,N_33693,N_34116);
nand U36804 (N_36804,N_33484,N_34970);
xnor U36805 (N_36805,N_33985,N_34821);
nor U36806 (N_36806,N_32786,N_34377);
xor U36807 (N_36807,N_34391,N_33428);
and U36808 (N_36808,N_34506,N_34172);
or U36809 (N_36809,N_34928,N_34717);
or U36810 (N_36810,N_34002,N_32890);
nor U36811 (N_36811,N_33186,N_32953);
nand U36812 (N_36812,N_33026,N_34134);
nor U36813 (N_36813,N_33391,N_32781);
or U36814 (N_36814,N_33634,N_33142);
xor U36815 (N_36815,N_32942,N_34668);
nor U36816 (N_36816,N_33072,N_33946);
or U36817 (N_36817,N_33926,N_33533);
nand U36818 (N_36818,N_33994,N_34825);
nor U36819 (N_36819,N_33674,N_33722);
nand U36820 (N_36820,N_33843,N_33942);
nand U36821 (N_36821,N_34347,N_34376);
nor U36822 (N_36822,N_33303,N_34370);
and U36823 (N_36823,N_33262,N_32628);
and U36824 (N_36824,N_34974,N_34655);
nand U36825 (N_36825,N_34395,N_34104);
nand U36826 (N_36826,N_33723,N_34080);
or U36827 (N_36827,N_34071,N_33254);
xnor U36828 (N_36828,N_34937,N_33532);
and U36829 (N_36829,N_32620,N_33543);
nand U36830 (N_36830,N_33891,N_33067);
nor U36831 (N_36831,N_33553,N_33871);
nand U36832 (N_36832,N_32663,N_32585);
nor U36833 (N_36833,N_32876,N_34502);
nor U36834 (N_36834,N_34746,N_34067);
nand U36835 (N_36835,N_34633,N_34056);
and U36836 (N_36836,N_32551,N_32699);
xor U36837 (N_36837,N_33660,N_33584);
nand U36838 (N_36838,N_34497,N_33839);
and U36839 (N_36839,N_32978,N_34418);
and U36840 (N_36840,N_32946,N_33463);
nor U36841 (N_36841,N_32564,N_34849);
nor U36842 (N_36842,N_34976,N_33684);
xnor U36843 (N_36843,N_34240,N_33947);
or U36844 (N_36844,N_34992,N_34837);
and U36845 (N_36845,N_33932,N_33205);
and U36846 (N_36846,N_34982,N_32676);
xor U36847 (N_36847,N_34339,N_32749);
nand U36848 (N_36848,N_34243,N_32845);
nor U36849 (N_36849,N_34536,N_33590);
xnor U36850 (N_36850,N_34189,N_34254);
and U36851 (N_36851,N_34508,N_33013);
nor U36852 (N_36852,N_33282,N_33926);
and U36853 (N_36853,N_34870,N_33117);
or U36854 (N_36854,N_32747,N_34190);
or U36855 (N_36855,N_33340,N_32566);
nor U36856 (N_36856,N_34375,N_32575);
nand U36857 (N_36857,N_33762,N_33617);
nor U36858 (N_36858,N_32711,N_34103);
nand U36859 (N_36859,N_32788,N_32636);
and U36860 (N_36860,N_34792,N_32797);
nor U36861 (N_36861,N_33906,N_34878);
xnor U36862 (N_36862,N_34574,N_33455);
or U36863 (N_36863,N_32692,N_34155);
nand U36864 (N_36864,N_33460,N_34167);
or U36865 (N_36865,N_32507,N_33361);
xnor U36866 (N_36866,N_32648,N_33666);
xnor U36867 (N_36867,N_32910,N_33130);
nor U36868 (N_36868,N_32801,N_33295);
or U36869 (N_36869,N_33119,N_32708);
xor U36870 (N_36870,N_32899,N_34655);
and U36871 (N_36871,N_33772,N_32758);
nor U36872 (N_36872,N_34173,N_32828);
and U36873 (N_36873,N_33503,N_33901);
xnor U36874 (N_36874,N_34806,N_32948);
xor U36875 (N_36875,N_34860,N_33579);
nand U36876 (N_36876,N_33478,N_33458);
or U36877 (N_36877,N_33975,N_33735);
xnor U36878 (N_36878,N_34685,N_32937);
xnor U36879 (N_36879,N_34145,N_34540);
or U36880 (N_36880,N_33130,N_33818);
nand U36881 (N_36881,N_33430,N_34810);
nand U36882 (N_36882,N_32687,N_32596);
nand U36883 (N_36883,N_32798,N_33896);
nand U36884 (N_36884,N_34720,N_34682);
nand U36885 (N_36885,N_34523,N_34487);
or U36886 (N_36886,N_33211,N_32551);
or U36887 (N_36887,N_32584,N_34713);
and U36888 (N_36888,N_34484,N_32819);
or U36889 (N_36889,N_34044,N_34312);
nor U36890 (N_36890,N_34512,N_34077);
xnor U36891 (N_36891,N_34277,N_34339);
nor U36892 (N_36892,N_32688,N_33535);
nor U36893 (N_36893,N_32703,N_34742);
or U36894 (N_36894,N_34038,N_32718);
nand U36895 (N_36895,N_32614,N_32827);
or U36896 (N_36896,N_34609,N_34317);
or U36897 (N_36897,N_33198,N_34168);
xor U36898 (N_36898,N_34658,N_33825);
xnor U36899 (N_36899,N_34319,N_33798);
xor U36900 (N_36900,N_33965,N_32723);
nand U36901 (N_36901,N_33691,N_33867);
and U36902 (N_36902,N_33793,N_34669);
or U36903 (N_36903,N_34308,N_34903);
xor U36904 (N_36904,N_34566,N_33812);
nand U36905 (N_36905,N_32917,N_34079);
and U36906 (N_36906,N_34803,N_33026);
and U36907 (N_36907,N_34975,N_32984);
or U36908 (N_36908,N_32885,N_33918);
xor U36909 (N_36909,N_34137,N_34901);
nor U36910 (N_36910,N_34370,N_34219);
nor U36911 (N_36911,N_34194,N_34748);
xnor U36912 (N_36912,N_33439,N_34705);
nor U36913 (N_36913,N_33212,N_32691);
xnor U36914 (N_36914,N_32997,N_32622);
and U36915 (N_36915,N_33941,N_32506);
xnor U36916 (N_36916,N_34574,N_34053);
nand U36917 (N_36917,N_33804,N_33737);
nand U36918 (N_36918,N_32705,N_33374);
xnor U36919 (N_36919,N_33884,N_34885);
nand U36920 (N_36920,N_34939,N_32605);
xnor U36921 (N_36921,N_33497,N_34819);
xnor U36922 (N_36922,N_33620,N_34079);
xnor U36923 (N_36923,N_32785,N_33581);
and U36924 (N_36924,N_34170,N_34709);
nor U36925 (N_36925,N_34181,N_34998);
and U36926 (N_36926,N_32829,N_33317);
xor U36927 (N_36927,N_33768,N_34893);
xor U36928 (N_36928,N_34411,N_32674);
or U36929 (N_36929,N_34272,N_32685);
xor U36930 (N_36930,N_34319,N_32976);
nand U36931 (N_36931,N_34421,N_34360);
or U36932 (N_36932,N_33457,N_34320);
nor U36933 (N_36933,N_33680,N_34183);
xor U36934 (N_36934,N_32804,N_33696);
nor U36935 (N_36935,N_34985,N_33056);
and U36936 (N_36936,N_34388,N_32895);
nor U36937 (N_36937,N_34417,N_33894);
and U36938 (N_36938,N_34040,N_34968);
nand U36939 (N_36939,N_34131,N_33509);
xnor U36940 (N_36940,N_32526,N_32535);
or U36941 (N_36941,N_34313,N_32947);
nand U36942 (N_36942,N_33092,N_33833);
and U36943 (N_36943,N_34193,N_33704);
nand U36944 (N_36944,N_32616,N_33863);
or U36945 (N_36945,N_33078,N_32848);
nor U36946 (N_36946,N_34229,N_34869);
nor U36947 (N_36947,N_33803,N_33059);
or U36948 (N_36948,N_32701,N_33514);
and U36949 (N_36949,N_33132,N_34004);
nand U36950 (N_36950,N_33845,N_33471);
nor U36951 (N_36951,N_32592,N_33017);
or U36952 (N_36952,N_34738,N_33737);
or U36953 (N_36953,N_33686,N_34624);
nand U36954 (N_36954,N_32965,N_32869);
nand U36955 (N_36955,N_33431,N_34761);
or U36956 (N_36956,N_32784,N_33667);
nand U36957 (N_36957,N_34105,N_34773);
xnor U36958 (N_36958,N_33252,N_34314);
nand U36959 (N_36959,N_33070,N_34285);
and U36960 (N_36960,N_34086,N_33134);
nor U36961 (N_36961,N_33933,N_32597);
xnor U36962 (N_36962,N_34654,N_33720);
nor U36963 (N_36963,N_34181,N_34843);
nor U36964 (N_36964,N_33889,N_33214);
or U36965 (N_36965,N_34746,N_34244);
nand U36966 (N_36966,N_33087,N_33362);
xor U36967 (N_36967,N_33717,N_34211);
nand U36968 (N_36968,N_33309,N_33183);
or U36969 (N_36969,N_33656,N_34308);
nor U36970 (N_36970,N_34962,N_32510);
and U36971 (N_36971,N_34237,N_34999);
nor U36972 (N_36972,N_34445,N_34677);
and U36973 (N_36973,N_32610,N_34485);
xor U36974 (N_36974,N_33167,N_33555);
nand U36975 (N_36975,N_33274,N_34113);
and U36976 (N_36976,N_33978,N_32669);
nand U36977 (N_36977,N_32673,N_33634);
or U36978 (N_36978,N_33679,N_34554);
or U36979 (N_36979,N_34528,N_34131);
xor U36980 (N_36980,N_34155,N_32508);
and U36981 (N_36981,N_33730,N_33190);
and U36982 (N_36982,N_34077,N_32678);
or U36983 (N_36983,N_33127,N_32870);
xor U36984 (N_36984,N_32987,N_34418);
nor U36985 (N_36985,N_34462,N_33095);
nand U36986 (N_36986,N_33327,N_33663);
or U36987 (N_36987,N_34322,N_33294);
xnor U36988 (N_36988,N_34915,N_33179);
nor U36989 (N_36989,N_32733,N_32991);
and U36990 (N_36990,N_34059,N_34388);
xnor U36991 (N_36991,N_32568,N_34370);
nor U36992 (N_36992,N_34504,N_34974);
nand U36993 (N_36993,N_32716,N_32907);
nor U36994 (N_36994,N_33410,N_32673);
nand U36995 (N_36995,N_33928,N_34093);
or U36996 (N_36996,N_33478,N_34937);
nor U36997 (N_36997,N_32878,N_34903);
and U36998 (N_36998,N_32608,N_34224);
nand U36999 (N_36999,N_34589,N_34433);
or U37000 (N_37000,N_33628,N_34624);
nor U37001 (N_37001,N_34009,N_33286);
and U37002 (N_37002,N_33464,N_34515);
nor U37003 (N_37003,N_34639,N_33675);
xor U37004 (N_37004,N_32513,N_32532);
or U37005 (N_37005,N_33426,N_34086);
xnor U37006 (N_37006,N_33513,N_33661);
xnor U37007 (N_37007,N_33983,N_33282);
and U37008 (N_37008,N_32559,N_33428);
and U37009 (N_37009,N_33013,N_33815);
nand U37010 (N_37010,N_32860,N_33974);
and U37011 (N_37011,N_34623,N_34056);
xnor U37012 (N_37012,N_33568,N_33876);
xnor U37013 (N_37013,N_34544,N_34670);
nor U37014 (N_37014,N_34960,N_34447);
nor U37015 (N_37015,N_33138,N_33937);
xor U37016 (N_37016,N_33560,N_34783);
nand U37017 (N_37017,N_33318,N_33255);
xor U37018 (N_37018,N_33566,N_34406);
or U37019 (N_37019,N_34356,N_33017);
and U37020 (N_37020,N_34373,N_34171);
xnor U37021 (N_37021,N_34471,N_33344);
nand U37022 (N_37022,N_33631,N_34070);
or U37023 (N_37023,N_32635,N_32571);
xnor U37024 (N_37024,N_33165,N_34895);
nor U37025 (N_37025,N_32803,N_34318);
nand U37026 (N_37026,N_34882,N_33426);
nand U37027 (N_37027,N_33076,N_34779);
and U37028 (N_37028,N_34862,N_33303);
or U37029 (N_37029,N_32811,N_33289);
and U37030 (N_37030,N_34105,N_34328);
or U37031 (N_37031,N_32561,N_32824);
and U37032 (N_37032,N_33522,N_34126);
and U37033 (N_37033,N_33945,N_33244);
or U37034 (N_37034,N_32951,N_33226);
and U37035 (N_37035,N_33395,N_33614);
and U37036 (N_37036,N_34902,N_34214);
nor U37037 (N_37037,N_32717,N_34060);
nand U37038 (N_37038,N_32985,N_34383);
xnor U37039 (N_37039,N_34298,N_33289);
nand U37040 (N_37040,N_34839,N_33563);
nand U37041 (N_37041,N_33090,N_34869);
xor U37042 (N_37042,N_34538,N_34259);
xnor U37043 (N_37043,N_33194,N_33467);
xnor U37044 (N_37044,N_34837,N_34620);
nor U37045 (N_37045,N_33447,N_34958);
nand U37046 (N_37046,N_34827,N_33446);
nand U37047 (N_37047,N_33186,N_33121);
xnor U37048 (N_37048,N_34416,N_33012);
xnor U37049 (N_37049,N_33006,N_33073);
and U37050 (N_37050,N_32553,N_33517);
nor U37051 (N_37051,N_34763,N_33548);
or U37052 (N_37052,N_33355,N_33082);
and U37053 (N_37053,N_33770,N_33125);
and U37054 (N_37054,N_34266,N_34664);
nand U37055 (N_37055,N_34423,N_32508);
xnor U37056 (N_37056,N_34251,N_34121);
nand U37057 (N_37057,N_32649,N_32795);
nand U37058 (N_37058,N_34082,N_34804);
nand U37059 (N_37059,N_33752,N_32735);
nor U37060 (N_37060,N_32533,N_33272);
and U37061 (N_37061,N_34289,N_32841);
xor U37062 (N_37062,N_34815,N_32874);
and U37063 (N_37063,N_32754,N_34055);
or U37064 (N_37064,N_32585,N_33513);
nand U37065 (N_37065,N_34207,N_33155);
nor U37066 (N_37066,N_33946,N_33546);
and U37067 (N_37067,N_34008,N_32566);
nand U37068 (N_37068,N_34612,N_32970);
nor U37069 (N_37069,N_34965,N_33991);
or U37070 (N_37070,N_33497,N_34037);
or U37071 (N_37071,N_33761,N_33896);
or U37072 (N_37072,N_33657,N_33414);
nand U37073 (N_37073,N_34816,N_34093);
or U37074 (N_37074,N_33710,N_33091);
nand U37075 (N_37075,N_34280,N_33615);
or U37076 (N_37076,N_33919,N_34302);
nand U37077 (N_37077,N_33124,N_33235);
xor U37078 (N_37078,N_32563,N_34947);
nand U37079 (N_37079,N_32845,N_34067);
or U37080 (N_37080,N_33390,N_33173);
or U37081 (N_37081,N_34245,N_32876);
nand U37082 (N_37082,N_33645,N_32895);
xor U37083 (N_37083,N_32625,N_32840);
nor U37084 (N_37084,N_34128,N_33245);
and U37085 (N_37085,N_33304,N_34731);
xor U37086 (N_37086,N_33004,N_33444);
or U37087 (N_37087,N_32685,N_34457);
xnor U37088 (N_37088,N_32825,N_34871);
and U37089 (N_37089,N_33297,N_33403);
nor U37090 (N_37090,N_34493,N_34648);
or U37091 (N_37091,N_34888,N_34074);
nand U37092 (N_37092,N_34979,N_33118);
nor U37093 (N_37093,N_34387,N_33655);
and U37094 (N_37094,N_33472,N_34220);
nand U37095 (N_37095,N_34861,N_34634);
nor U37096 (N_37096,N_32697,N_34921);
xnor U37097 (N_37097,N_33495,N_34619);
or U37098 (N_37098,N_34835,N_33372);
nand U37099 (N_37099,N_32581,N_33921);
or U37100 (N_37100,N_33332,N_33073);
and U37101 (N_37101,N_34007,N_32999);
and U37102 (N_37102,N_32837,N_32519);
nor U37103 (N_37103,N_33499,N_34356);
or U37104 (N_37104,N_34841,N_32611);
xor U37105 (N_37105,N_33834,N_32842);
or U37106 (N_37106,N_32782,N_33194);
xor U37107 (N_37107,N_33481,N_32516);
or U37108 (N_37108,N_33004,N_34073);
or U37109 (N_37109,N_34319,N_34716);
or U37110 (N_37110,N_34637,N_32873);
nand U37111 (N_37111,N_34248,N_34047);
xnor U37112 (N_37112,N_34527,N_32854);
nand U37113 (N_37113,N_33232,N_32715);
and U37114 (N_37114,N_32683,N_32567);
nor U37115 (N_37115,N_32567,N_33471);
or U37116 (N_37116,N_33988,N_34864);
and U37117 (N_37117,N_34578,N_32543);
xor U37118 (N_37118,N_34328,N_34405);
xor U37119 (N_37119,N_33604,N_33252);
or U37120 (N_37120,N_34171,N_34588);
nor U37121 (N_37121,N_33980,N_33634);
or U37122 (N_37122,N_32571,N_33384);
nor U37123 (N_37123,N_33654,N_34347);
and U37124 (N_37124,N_34991,N_33606);
xnor U37125 (N_37125,N_34275,N_34320);
or U37126 (N_37126,N_33894,N_33742);
nor U37127 (N_37127,N_33753,N_32946);
or U37128 (N_37128,N_33942,N_33587);
or U37129 (N_37129,N_34058,N_33919);
nor U37130 (N_37130,N_33899,N_34264);
xnor U37131 (N_37131,N_34379,N_33127);
and U37132 (N_37132,N_33355,N_34111);
and U37133 (N_37133,N_34330,N_34250);
nor U37134 (N_37134,N_34345,N_34831);
xnor U37135 (N_37135,N_32850,N_34360);
or U37136 (N_37136,N_33381,N_32931);
xor U37137 (N_37137,N_33488,N_32997);
nor U37138 (N_37138,N_33112,N_33809);
nor U37139 (N_37139,N_34830,N_33770);
nand U37140 (N_37140,N_33038,N_33411);
xnor U37141 (N_37141,N_33241,N_33334);
and U37142 (N_37142,N_34361,N_34188);
xor U37143 (N_37143,N_33337,N_34774);
xnor U37144 (N_37144,N_32886,N_32697);
or U37145 (N_37145,N_34762,N_34613);
xor U37146 (N_37146,N_34939,N_33402);
or U37147 (N_37147,N_33932,N_32677);
and U37148 (N_37148,N_33772,N_33365);
or U37149 (N_37149,N_32847,N_33267);
nand U37150 (N_37150,N_32661,N_33857);
xor U37151 (N_37151,N_33490,N_34582);
xnor U37152 (N_37152,N_34859,N_34955);
and U37153 (N_37153,N_32712,N_34225);
or U37154 (N_37154,N_34568,N_33693);
nand U37155 (N_37155,N_33722,N_32715);
xor U37156 (N_37156,N_33778,N_34791);
xor U37157 (N_37157,N_34623,N_34823);
xor U37158 (N_37158,N_33768,N_33420);
nand U37159 (N_37159,N_34610,N_33471);
or U37160 (N_37160,N_34018,N_34307);
and U37161 (N_37161,N_34818,N_33276);
nor U37162 (N_37162,N_33387,N_34318);
and U37163 (N_37163,N_33394,N_33642);
xnor U37164 (N_37164,N_32950,N_33087);
and U37165 (N_37165,N_34250,N_34101);
nor U37166 (N_37166,N_34206,N_33287);
nor U37167 (N_37167,N_33886,N_34772);
nand U37168 (N_37168,N_32674,N_32977);
nand U37169 (N_37169,N_32674,N_32838);
nand U37170 (N_37170,N_33138,N_34678);
xnor U37171 (N_37171,N_33982,N_34683);
or U37172 (N_37172,N_32626,N_32830);
and U37173 (N_37173,N_34190,N_34403);
nor U37174 (N_37174,N_34572,N_34951);
and U37175 (N_37175,N_32892,N_34633);
nand U37176 (N_37176,N_33593,N_34969);
nand U37177 (N_37177,N_34749,N_34082);
xnor U37178 (N_37178,N_32666,N_33343);
xor U37179 (N_37179,N_33279,N_34811);
nor U37180 (N_37180,N_34929,N_34876);
xor U37181 (N_37181,N_32694,N_33426);
nand U37182 (N_37182,N_34117,N_32580);
or U37183 (N_37183,N_34099,N_33189);
nor U37184 (N_37184,N_32889,N_33855);
nor U37185 (N_37185,N_34282,N_32668);
nor U37186 (N_37186,N_33129,N_33367);
nor U37187 (N_37187,N_32504,N_34833);
nor U37188 (N_37188,N_34477,N_34848);
and U37189 (N_37189,N_34838,N_33423);
xor U37190 (N_37190,N_33364,N_32595);
and U37191 (N_37191,N_34519,N_33307);
and U37192 (N_37192,N_33916,N_34097);
nand U37193 (N_37193,N_34450,N_32999);
nand U37194 (N_37194,N_33033,N_32561);
or U37195 (N_37195,N_32861,N_34507);
or U37196 (N_37196,N_33496,N_33607);
and U37197 (N_37197,N_32836,N_34017);
nor U37198 (N_37198,N_34011,N_34825);
xnor U37199 (N_37199,N_33692,N_34881);
or U37200 (N_37200,N_33212,N_33041);
xor U37201 (N_37201,N_33243,N_33815);
and U37202 (N_37202,N_33408,N_33108);
or U37203 (N_37203,N_33064,N_33526);
nor U37204 (N_37204,N_33964,N_33256);
nand U37205 (N_37205,N_32762,N_32631);
or U37206 (N_37206,N_34724,N_34903);
and U37207 (N_37207,N_34254,N_33471);
nand U37208 (N_37208,N_32873,N_32850);
nor U37209 (N_37209,N_34627,N_33151);
xor U37210 (N_37210,N_34444,N_33763);
xnor U37211 (N_37211,N_33842,N_33161);
nand U37212 (N_37212,N_32617,N_34806);
xor U37213 (N_37213,N_33091,N_34031);
and U37214 (N_37214,N_33044,N_34633);
nand U37215 (N_37215,N_33760,N_34587);
or U37216 (N_37216,N_33408,N_34290);
nand U37217 (N_37217,N_34889,N_34425);
nor U37218 (N_37218,N_33622,N_34641);
or U37219 (N_37219,N_34766,N_33572);
xnor U37220 (N_37220,N_34695,N_33308);
nor U37221 (N_37221,N_32567,N_34131);
and U37222 (N_37222,N_32648,N_34289);
nand U37223 (N_37223,N_32865,N_33814);
nand U37224 (N_37224,N_32861,N_32804);
and U37225 (N_37225,N_33850,N_32804);
or U37226 (N_37226,N_32757,N_32710);
nand U37227 (N_37227,N_34447,N_33288);
and U37228 (N_37228,N_34097,N_32845);
or U37229 (N_37229,N_34288,N_34238);
xor U37230 (N_37230,N_34768,N_34850);
xor U37231 (N_37231,N_33039,N_33852);
nor U37232 (N_37232,N_34873,N_34021);
and U37233 (N_37233,N_33864,N_34233);
nand U37234 (N_37234,N_34927,N_33489);
xor U37235 (N_37235,N_32579,N_32952);
nor U37236 (N_37236,N_34248,N_34289);
nor U37237 (N_37237,N_32972,N_34494);
nand U37238 (N_37238,N_34786,N_34028);
or U37239 (N_37239,N_33850,N_33208);
xnor U37240 (N_37240,N_34981,N_33850);
xor U37241 (N_37241,N_34313,N_34006);
nand U37242 (N_37242,N_32769,N_33448);
or U37243 (N_37243,N_32545,N_34486);
nand U37244 (N_37244,N_33839,N_33274);
and U37245 (N_37245,N_34629,N_32679);
nand U37246 (N_37246,N_33301,N_32782);
nand U37247 (N_37247,N_33702,N_34626);
xor U37248 (N_37248,N_34795,N_34192);
xnor U37249 (N_37249,N_33106,N_33710);
xnor U37250 (N_37250,N_34743,N_34057);
nor U37251 (N_37251,N_34225,N_34923);
xnor U37252 (N_37252,N_32874,N_33807);
nand U37253 (N_37253,N_33695,N_34787);
xnor U37254 (N_37254,N_34881,N_32916);
nor U37255 (N_37255,N_34421,N_32957);
xnor U37256 (N_37256,N_32782,N_34781);
or U37257 (N_37257,N_32975,N_33132);
nand U37258 (N_37258,N_34954,N_34539);
or U37259 (N_37259,N_33130,N_33825);
xor U37260 (N_37260,N_34792,N_32535);
nor U37261 (N_37261,N_34002,N_33252);
or U37262 (N_37262,N_33631,N_32669);
nand U37263 (N_37263,N_34487,N_34158);
xnor U37264 (N_37264,N_34585,N_33738);
and U37265 (N_37265,N_33728,N_34305);
xnor U37266 (N_37266,N_33356,N_34117);
nor U37267 (N_37267,N_34775,N_34372);
nand U37268 (N_37268,N_34558,N_34533);
nor U37269 (N_37269,N_34496,N_34654);
or U37270 (N_37270,N_33271,N_34617);
nor U37271 (N_37271,N_34797,N_33466);
or U37272 (N_37272,N_33027,N_33489);
and U37273 (N_37273,N_34605,N_33857);
nand U37274 (N_37274,N_34214,N_32896);
and U37275 (N_37275,N_33943,N_32701);
or U37276 (N_37276,N_33189,N_33734);
and U37277 (N_37277,N_32697,N_33526);
xnor U37278 (N_37278,N_33340,N_32551);
or U37279 (N_37279,N_34860,N_33366);
nor U37280 (N_37280,N_33182,N_32608);
xnor U37281 (N_37281,N_34898,N_33167);
nor U37282 (N_37282,N_33226,N_34314);
or U37283 (N_37283,N_32537,N_33646);
or U37284 (N_37284,N_34745,N_34958);
nor U37285 (N_37285,N_32756,N_33553);
and U37286 (N_37286,N_34664,N_34044);
or U37287 (N_37287,N_33821,N_33513);
xor U37288 (N_37288,N_34497,N_33881);
xor U37289 (N_37289,N_33944,N_32846);
xnor U37290 (N_37290,N_32623,N_34097);
or U37291 (N_37291,N_33826,N_33317);
nor U37292 (N_37292,N_34761,N_34830);
and U37293 (N_37293,N_33054,N_32635);
or U37294 (N_37294,N_33670,N_34880);
or U37295 (N_37295,N_34405,N_33519);
or U37296 (N_37296,N_33533,N_32779);
nand U37297 (N_37297,N_34439,N_32919);
or U37298 (N_37298,N_34028,N_34434);
xnor U37299 (N_37299,N_32576,N_33272);
nor U37300 (N_37300,N_33167,N_33469);
nand U37301 (N_37301,N_33038,N_33212);
and U37302 (N_37302,N_32814,N_32950);
or U37303 (N_37303,N_33912,N_34345);
and U37304 (N_37304,N_32699,N_32864);
nand U37305 (N_37305,N_34485,N_33441);
or U37306 (N_37306,N_33407,N_33691);
nor U37307 (N_37307,N_33825,N_32925);
nor U37308 (N_37308,N_34312,N_34098);
and U37309 (N_37309,N_33974,N_32852);
or U37310 (N_37310,N_34045,N_33883);
or U37311 (N_37311,N_33203,N_33238);
nor U37312 (N_37312,N_34432,N_34098);
nand U37313 (N_37313,N_32766,N_32824);
xor U37314 (N_37314,N_33395,N_33261);
nor U37315 (N_37315,N_33949,N_32807);
or U37316 (N_37316,N_34580,N_34309);
nor U37317 (N_37317,N_34573,N_33216);
nor U37318 (N_37318,N_33892,N_33005);
nand U37319 (N_37319,N_33807,N_33497);
or U37320 (N_37320,N_32910,N_33080);
nand U37321 (N_37321,N_33707,N_33044);
xor U37322 (N_37322,N_34926,N_33939);
xor U37323 (N_37323,N_34866,N_34287);
or U37324 (N_37324,N_34327,N_33168);
or U37325 (N_37325,N_34850,N_34106);
nor U37326 (N_37326,N_32788,N_33212);
xnor U37327 (N_37327,N_33526,N_32878);
xor U37328 (N_37328,N_33048,N_32935);
or U37329 (N_37329,N_34961,N_32957);
nor U37330 (N_37330,N_33729,N_33389);
or U37331 (N_37331,N_33447,N_33556);
or U37332 (N_37332,N_32613,N_34404);
nand U37333 (N_37333,N_34641,N_33694);
nand U37334 (N_37334,N_32539,N_33030);
and U37335 (N_37335,N_33584,N_34826);
and U37336 (N_37336,N_32542,N_32916);
or U37337 (N_37337,N_33171,N_34354);
nor U37338 (N_37338,N_32926,N_34650);
or U37339 (N_37339,N_32788,N_33222);
and U37340 (N_37340,N_34110,N_34150);
nor U37341 (N_37341,N_34235,N_34617);
nor U37342 (N_37342,N_34555,N_34401);
and U37343 (N_37343,N_33556,N_33950);
nor U37344 (N_37344,N_32501,N_34678);
xor U37345 (N_37345,N_34274,N_34591);
or U37346 (N_37346,N_34217,N_32957);
xor U37347 (N_37347,N_33715,N_34566);
nor U37348 (N_37348,N_33410,N_33937);
nor U37349 (N_37349,N_33677,N_33632);
xnor U37350 (N_37350,N_32538,N_33205);
nand U37351 (N_37351,N_33316,N_32780);
or U37352 (N_37352,N_34516,N_34181);
and U37353 (N_37353,N_34511,N_34796);
nand U37354 (N_37354,N_34484,N_33655);
and U37355 (N_37355,N_34453,N_34348);
xnor U37356 (N_37356,N_32616,N_33666);
nor U37357 (N_37357,N_32563,N_33642);
xnor U37358 (N_37358,N_32539,N_34888);
or U37359 (N_37359,N_33324,N_32606);
xor U37360 (N_37360,N_32853,N_34220);
xor U37361 (N_37361,N_34210,N_32572);
xor U37362 (N_37362,N_32503,N_33341);
and U37363 (N_37363,N_34777,N_33763);
or U37364 (N_37364,N_33014,N_34580);
or U37365 (N_37365,N_34344,N_33168);
or U37366 (N_37366,N_33095,N_34164);
and U37367 (N_37367,N_33698,N_33779);
and U37368 (N_37368,N_33081,N_33214);
and U37369 (N_37369,N_33188,N_34754);
or U37370 (N_37370,N_33064,N_33642);
or U37371 (N_37371,N_34776,N_34586);
or U37372 (N_37372,N_34325,N_33063);
and U37373 (N_37373,N_34591,N_34908);
or U37374 (N_37374,N_32568,N_34603);
xor U37375 (N_37375,N_34629,N_34197);
nand U37376 (N_37376,N_34507,N_33971);
nor U37377 (N_37377,N_34675,N_34507);
and U37378 (N_37378,N_33104,N_33658);
and U37379 (N_37379,N_32741,N_33846);
nand U37380 (N_37380,N_32631,N_32998);
or U37381 (N_37381,N_34928,N_34988);
xnor U37382 (N_37382,N_34144,N_34012);
nand U37383 (N_37383,N_34079,N_34727);
and U37384 (N_37384,N_34531,N_33374);
xor U37385 (N_37385,N_32689,N_33501);
nand U37386 (N_37386,N_33684,N_33256);
xor U37387 (N_37387,N_34202,N_34998);
or U37388 (N_37388,N_34946,N_33861);
or U37389 (N_37389,N_33177,N_34870);
xor U37390 (N_37390,N_34083,N_32616);
nor U37391 (N_37391,N_33846,N_34899);
nand U37392 (N_37392,N_32545,N_34649);
and U37393 (N_37393,N_34329,N_34054);
and U37394 (N_37394,N_34814,N_33612);
or U37395 (N_37395,N_34277,N_33379);
nor U37396 (N_37396,N_33583,N_33959);
and U37397 (N_37397,N_32984,N_34664);
xnor U37398 (N_37398,N_33049,N_33158);
nor U37399 (N_37399,N_34934,N_34617);
and U37400 (N_37400,N_33336,N_33850);
xnor U37401 (N_37401,N_33244,N_32755);
nor U37402 (N_37402,N_33684,N_33647);
or U37403 (N_37403,N_33495,N_34804);
xor U37404 (N_37404,N_34731,N_34611);
xor U37405 (N_37405,N_33873,N_34735);
nor U37406 (N_37406,N_33632,N_34616);
or U37407 (N_37407,N_34554,N_33617);
and U37408 (N_37408,N_34375,N_34633);
or U37409 (N_37409,N_34017,N_33805);
nand U37410 (N_37410,N_33246,N_33225);
and U37411 (N_37411,N_32556,N_32792);
nand U37412 (N_37412,N_32856,N_32507);
nor U37413 (N_37413,N_34140,N_33385);
or U37414 (N_37414,N_33001,N_34943);
or U37415 (N_37415,N_33284,N_33724);
nand U37416 (N_37416,N_33291,N_34520);
or U37417 (N_37417,N_33179,N_32804);
and U37418 (N_37418,N_33494,N_32540);
or U37419 (N_37419,N_32642,N_33985);
or U37420 (N_37420,N_34742,N_32634);
xnor U37421 (N_37421,N_33289,N_34035);
xnor U37422 (N_37422,N_34774,N_34295);
nand U37423 (N_37423,N_33964,N_34322);
nor U37424 (N_37424,N_33430,N_34575);
xnor U37425 (N_37425,N_33402,N_34807);
nor U37426 (N_37426,N_33862,N_34841);
nor U37427 (N_37427,N_32937,N_34395);
xnor U37428 (N_37428,N_32852,N_34987);
nor U37429 (N_37429,N_34264,N_33375);
and U37430 (N_37430,N_33631,N_33037);
or U37431 (N_37431,N_34478,N_32969);
and U37432 (N_37432,N_32650,N_33964);
xnor U37433 (N_37433,N_33630,N_32511);
nor U37434 (N_37434,N_34567,N_33668);
or U37435 (N_37435,N_34264,N_34084);
and U37436 (N_37436,N_33093,N_32722);
nor U37437 (N_37437,N_34780,N_34094);
xor U37438 (N_37438,N_32608,N_34454);
nand U37439 (N_37439,N_34079,N_34378);
and U37440 (N_37440,N_34965,N_33836);
or U37441 (N_37441,N_34188,N_34809);
and U37442 (N_37442,N_32991,N_34677);
xnor U37443 (N_37443,N_34924,N_34026);
nand U37444 (N_37444,N_33306,N_33113);
xnor U37445 (N_37445,N_34108,N_34602);
and U37446 (N_37446,N_33921,N_33712);
or U37447 (N_37447,N_32621,N_34217);
nand U37448 (N_37448,N_34117,N_33331);
nor U37449 (N_37449,N_33660,N_34144);
or U37450 (N_37450,N_34878,N_33322);
and U37451 (N_37451,N_34285,N_34063);
nor U37452 (N_37452,N_34471,N_34174);
nand U37453 (N_37453,N_34204,N_34829);
xor U37454 (N_37454,N_34295,N_33457);
nor U37455 (N_37455,N_34549,N_33606);
nor U37456 (N_37456,N_34852,N_33247);
or U37457 (N_37457,N_33786,N_33784);
nand U37458 (N_37458,N_32673,N_32922);
or U37459 (N_37459,N_34341,N_32678);
nand U37460 (N_37460,N_33418,N_33648);
nand U37461 (N_37461,N_32754,N_34564);
xor U37462 (N_37462,N_34206,N_32575);
nor U37463 (N_37463,N_33371,N_32554);
nand U37464 (N_37464,N_34431,N_34882);
nor U37465 (N_37465,N_34699,N_34728);
xor U37466 (N_37466,N_33003,N_33624);
xnor U37467 (N_37467,N_32999,N_32998);
nand U37468 (N_37468,N_33007,N_32772);
nand U37469 (N_37469,N_33140,N_34107);
nand U37470 (N_37470,N_34492,N_34431);
and U37471 (N_37471,N_34525,N_34376);
nor U37472 (N_37472,N_33668,N_34035);
nor U37473 (N_37473,N_34916,N_33166);
xnor U37474 (N_37474,N_33106,N_34821);
and U37475 (N_37475,N_33822,N_33452);
nor U37476 (N_37476,N_34238,N_32953);
or U37477 (N_37477,N_33651,N_33904);
nand U37478 (N_37478,N_34502,N_32694);
and U37479 (N_37479,N_33853,N_33554);
and U37480 (N_37480,N_33393,N_33242);
nand U37481 (N_37481,N_34972,N_32944);
xnor U37482 (N_37482,N_34661,N_34066);
xor U37483 (N_37483,N_34468,N_32947);
or U37484 (N_37484,N_34560,N_33114);
xor U37485 (N_37485,N_34013,N_34405);
or U37486 (N_37486,N_33175,N_33982);
nor U37487 (N_37487,N_34716,N_33009);
and U37488 (N_37488,N_34112,N_33737);
or U37489 (N_37489,N_34510,N_33779);
or U37490 (N_37490,N_33503,N_34767);
or U37491 (N_37491,N_33273,N_34524);
and U37492 (N_37492,N_34429,N_32569);
and U37493 (N_37493,N_34616,N_34852);
nand U37494 (N_37494,N_33457,N_34442);
nor U37495 (N_37495,N_32812,N_33260);
xor U37496 (N_37496,N_34615,N_33707);
nor U37497 (N_37497,N_34499,N_34949);
nand U37498 (N_37498,N_33725,N_33798);
xor U37499 (N_37499,N_33517,N_33455);
xor U37500 (N_37500,N_37187,N_36323);
or U37501 (N_37501,N_35514,N_35354);
and U37502 (N_37502,N_36898,N_37360);
or U37503 (N_37503,N_35383,N_35673);
or U37504 (N_37504,N_35830,N_37154);
xor U37505 (N_37505,N_36132,N_36689);
nand U37506 (N_37506,N_35305,N_36589);
xor U37507 (N_37507,N_36933,N_35298);
and U37508 (N_37508,N_35567,N_35303);
or U37509 (N_37509,N_36914,N_36722);
and U37510 (N_37510,N_35572,N_36265);
nand U37511 (N_37511,N_35777,N_36764);
nor U37512 (N_37512,N_36171,N_35621);
nand U37513 (N_37513,N_36170,N_35637);
nor U37514 (N_37514,N_35711,N_35481);
nand U37515 (N_37515,N_37025,N_35594);
or U37516 (N_37516,N_37388,N_36311);
nor U37517 (N_37517,N_36198,N_35047);
nor U37518 (N_37518,N_35728,N_35304);
nor U37519 (N_37519,N_36231,N_36945);
or U37520 (N_37520,N_35401,N_35242);
or U37521 (N_37521,N_36013,N_37250);
or U37522 (N_37522,N_35645,N_36820);
and U37523 (N_37523,N_37036,N_37459);
nor U37524 (N_37524,N_35036,N_36921);
and U37525 (N_37525,N_35456,N_36291);
and U37526 (N_37526,N_35244,N_36612);
xor U37527 (N_37527,N_36906,N_35694);
nand U37528 (N_37528,N_36672,N_37491);
nor U37529 (N_37529,N_36570,N_36919);
or U37530 (N_37530,N_36254,N_35863);
and U37531 (N_37531,N_37478,N_35628);
or U37532 (N_37532,N_35794,N_36294);
or U37533 (N_37533,N_35617,N_36189);
xor U37534 (N_37534,N_37055,N_37394);
or U37535 (N_37535,N_36536,N_36687);
nor U37536 (N_37536,N_36033,N_36610);
or U37537 (N_37537,N_36923,N_35730);
xor U37538 (N_37538,N_36724,N_36809);
nand U37539 (N_37539,N_37012,N_35018);
nand U37540 (N_37540,N_37209,N_35806);
nand U37541 (N_37541,N_35565,N_35760);
nor U37542 (N_37542,N_35425,N_35165);
and U37543 (N_37543,N_35926,N_36212);
xor U37544 (N_37544,N_35353,N_35738);
and U37545 (N_37545,N_35992,N_37447);
nand U37546 (N_37546,N_35217,N_35721);
or U37547 (N_37547,N_37110,N_35624);
nand U37548 (N_37548,N_35124,N_35143);
or U37549 (N_37549,N_35345,N_35319);
nand U37550 (N_37550,N_36204,N_36194);
or U37551 (N_37551,N_36550,N_37128);
nor U37552 (N_37552,N_35449,N_37008);
and U37553 (N_37553,N_36941,N_35037);
nand U37554 (N_37554,N_37014,N_35857);
or U37555 (N_37555,N_36356,N_35526);
or U37556 (N_37556,N_35381,N_35856);
nor U37557 (N_37557,N_36258,N_35224);
nor U37558 (N_37558,N_35220,N_36917);
nand U37559 (N_37559,N_35487,N_36414);
and U37560 (N_37560,N_36025,N_36325);
or U37561 (N_37561,N_35897,N_37069);
nor U37562 (N_37562,N_36327,N_36837);
nand U37563 (N_37563,N_37100,N_37442);
or U37564 (N_37564,N_35291,N_36275);
nor U37565 (N_37565,N_37386,N_37161);
nor U37566 (N_37566,N_35392,N_36515);
or U37567 (N_37567,N_36293,N_36752);
or U37568 (N_37568,N_35137,N_35558);
xor U37569 (N_37569,N_37169,N_37392);
xnor U37570 (N_37570,N_36247,N_35840);
and U37571 (N_37571,N_36065,N_35971);
and U37572 (N_37572,N_35468,N_37125);
nor U37573 (N_37573,N_36700,N_35619);
and U37574 (N_37574,N_35498,N_35632);
nor U37575 (N_37575,N_37301,N_36116);
or U37576 (N_37576,N_35564,N_35774);
or U37577 (N_37577,N_36238,N_35104);
or U37578 (N_37578,N_37051,N_35180);
and U37579 (N_37579,N_37197,N_35876);
xnor U37580 (N_37580,N_35816,N_36813);
nor U37581 (N_37581,N_36250,N_36931);
nand U37582 (N_37582,N_35732,N_35512);
or U37583 (N_37583,N_36779,N_35791);
nand U37584 (N_37584,N_36645,N_35672);
nor U37585 (N_37585,N_35663,N_37264);
and U37586 (N_37586,N_35973,N_36426);
and U37587 (N_37587,N_35548,N_35459);
and U37588 (N_37588,N_35804,N_37200);
nand U37589 (N_37589,N_36774,N_35636);
xnor U37590 (N_37590,N_37319,N_35823);
and U37591 (N_37591,N_35397,N_36101);
and U37592 (N_37592,N_37257,N_36856);
nand U37593 (N_37593,N_36241,N_35301);
and U37594 (N_37594,N_36805,N_36948);
xor U37595 (N_37595,N_37380,N_36090);
nor U37596 (N_37596,N_36347,N_35315);
and U37597 (N_37597,N_36737,N_35693);
nor U37598 (N_37598,N_37099,N_35908);
xnor U37599 (N_37599,N_36218,N_36835);
or U37600 (N_37600,N_35890,N_37406);
nand U37601 (N_37601,N_35972,N_35350);
nor U37602 (N_37602,N_37498,N_37061);
nand U37603 (N_37603,N_35284,N_37040);
nor U37604 (N_37604,N_35440,N_35019);
xor U37605 (N_37605,N_36169,N_37371);
and U37606 (N_37606,N_35348,N_35287);
nor U37607 (N_37607,N_36015,N_37103);
and U37608 (N_37608,N_36709,N_37087);
nor U37609 (N_37609,N_36979,N_37033);
xor U37610 (N_37610,N_35706,N_35595);
nor U37611 (N_37611,N_36380,N_36843);
or U37612 (N_37612,N_36904,N_37156);
xnor U37613 (N_37613,N_35753,N_36901);
or U37614 (N_37614,N_36011,N_35403);
nor U37615 (N_37615,N_37046,N_36188);
or U37616 (N_37616,N_36242,N_36609);
nand U37617 (N_37617,N_35030,N_35824);
xor U37618 (N_37618,N_36100,N_36374);
xor U37619 (N_37619,N_36431,N_35333);
or U37620 (N_37620,N_36335,N_35592);
nor U37621 (N_37621,N_36699,N_36145);
or U37622 (N_37622,N_35409,N_36838);
xnor U37623 (N_37623,N_36074,N_37080);
and U37624 (N_37624,N_35915,N_36817);
or U37625 (N_37625,N_36759,N_37149);
nor U37626 (N_37626,N_36551,N_36583);
nand U37627 (N_37627,N_35480,N_36987);
and U37628 (N_37628,N_36746,N_36739);
or U37629 (N_37629,N_37353,N_37283);
or U37630 (N_37630,N_36996,N_35455);
nand U37631 (N_37631,N_37453,N_36423);
and U37632 (N_37632,N_35911,N_37031);
and U37633 (N_37633,N_35067,N_36306);
and U37634 (N_37634,N_36346,N_36590);
and U37635 (N_37635,N_36442,N_35292);
xnor U37636 (N_37636,N_36045,N_35610);
and U37637 (N_37637,N_36519,N_36326);
and U37638 (N_37638,N_36539,N_35923);
nand U37639 (N_37639,N_35399,N_37321);
nor U37640 (N_37640,N_37372,N_36602);
or U37641 (N_37641,N_36888,N_36775);
or U37642 (N_37642,N_35574,N_36468);
nor U37643 (N_37643,N_36117,N_36027);
xor U37644 (N_37644,N_36989,N_35518);
xnor U37645 (N_37645,N_36109,N_36521);
and U37646 (N_37646,N_36394,N_35331);
and U37647 (N_37647,N_36929,N_36041);
xor U37648 (N_37648,N_36190,N_36295);
and U37649 (N_37649,N_37456,N_37436);
xor U37650 (N_37650,N_35070,N_36068);
xor U37651 (N_37651,N_35695,N_37071);
or U37652 (N_37652,N_35937,N_36371);
xnor U37653 (N_37653,N_36344,N_37193);
or U37654 (N_37654,N_37235,N_35611);
nor U37655 (N_37655,N_36851,N_36760);
nor U37656 (N_37656,N_36220,N_36088);
or U37657 (N_37657,N_36062,N_36611);
and U37658 (N_37658,N_35761,N_35547);
xnor U37659 (N_37659,N_36897,N_35068);
nand U37660 (N_37660,N_36582,N_35144);
nand U37661 (N_37661,N_37349,N_36039);
and U37662 (N_37662,N_35552,N_36451);
nor U37663 (N_37663,N_36186,N_36164);
nand U37664 (N_37664,N_36177,N_36822);
xnor U37665 (N_37665,N_37047,N_36260);
or U37666 (N_37666,N_37278,N_35054);
nor U37667 (N_37667,N_37252,N_35269);
nor U37668 (N_37668,N_35077,N_37146);
nor U37669 (N_37669,N_35869,N_36997);
and U37670 (N_37670,N_36466,N_35546);
xor U37671 (N_37671,N_35934,N_37496);
and U37672 (N_37672,N_35274,N_35898);
xnor U37673 (N_37673,N_35275,N_35531);
nand U37674 (N_37674,N_36797,N_37077);
and U37675 (N_37675,N_35846,N_35789);
xnor U37676 (N_37676,N_36653,N_37310);
nand U37677 (N_37677,N_37366,N_36905);
nor U37678 (N_37678,N_35961,N_36391);
and U37679 (N_37679,N_36530,N_36318);
and U37680 (N_37680,N_36690,N_37243);
nor U37681 (N_37681,N_36926,N_36044);
xnor U37682 (N_37682,N_35423,N_35211);
xor U37683 (N_37683,N_36865,N_35262);
xnor U37684 (N_37684,N_37309,N_35559);
xor U37685 (N_37685,N_36879,N_36078);
and U37686 (N_37686,N_37056,N_35888);
nand U37687 (N_37687,N_37236,N_35776);
nand U37688 (N_37688,N_35589,N_35079);
nand U37689 (N_37689,N_36955,N_36581);
nor U37690 (N_37690,N_36518,N_35767);
and U37691 (N_37691,N_35346,N_36962);
nand U37692 (N_37692,N_35190,N_36930);
or U37693 (N_37693,N_35954,N_35667);
and U37694 (N_37694,N_35475,N_36184);
nor U37695 (N_37695,N_35379,N_35635);
and U37696 (N_37696,N_36385,N_37297);
and U37697 (N_37697,N_35873,N_36704);
and U37698 (N_37698,N_36034,N_35603);
xnor U37699 (N_37699,N_35545,N_36122);
and U37700 (N_37700,N_35110,N_35225);
nor U37701 (N_37701,N_35807,N_36556);
nor U37702 (N_37702,N_35085,N_37094);
nor U37703 (N_37703,N_35763,N_36368);
xor U37704 (N_37704,N_36280,N_35729);
nor U37705 (N_37705,N_35839,N_35527);
or U37706 (N_37706,N_36830,N_35832);
xnor U37707 (N_37707,N_36532,N_37145);
and U37708 (N_37708,N_36983,N_35090);
nand U37709 (N_37709,N_36743,N_35543);
xor U37710 (N_37710,N_35720,N_37162);
and U37711 (N_37711,N_37472,N_37376);
xnor U37712 (N_37712,N_36036,N_36854);
nor U37713 (N_37713,N_35162,N_37488);
or U37714 (N_37714,N_36113,N_36751);
nor U37715 (N_37715,N_37474,N_36691);
or U37716 (N_37716,N_36562,N_36787);
xor U37717 (N_37717,N_36205,N_35207);
xor U37718 (N_37718,N_35272,N_36299);
or U37719 (N_37719,N_35587,N_36428);
nor U37720 (N_37720,N_36961,N_37095);
xor U37721 (N_37721,N_36453,N_36975);
and U37722 (N_37722,N_35618,N_35172);
or U37723 (N_37723,N_35302,N_37318);
and U37724 (N_37724,N_35115,N_35445);
or U37725 (N_37725,N_37433,N_36988);
or U37726 (N_37726,N_36440,N_35058);
xnor U37727 (N_37727,N_35447,N_36083);
nand U37728 (N_37728,N_35450,N_36175);
or U37729 (N_37729,N_36781,N_35845);
or U37730 (N_37730,N_35792,N_35002);
and U37731 (N_37731,N_36492,N_36663);
xor U37732 (N_37732,N_36496,N_35435);
nor U37733 (N_37733,N_35553,N_36899);
and U37734 (N_37734,N_37176,N_35192);
nor U37735 (N_37735,N_37052,N_35411);
nor U37736 (N_37736,N_36567,N_35271);
xor U37737 (N_37737,N_37242,N_37163);
and U37738 (N_37738,N_35679,N_37228);
or U37739 (N_37739,N_35772,N_37013);
and U37740 (N_37740,N_36810,N_35142);
nand U37741 (N_37741,N_35363,N_36107);
nand U37742 (N_37742,N_35247,N_35529);
nand U37743 (N_37743,N_36136,N_36892);
nor U37744 (N_37744,N_37091,N_36907);
or U37745 (N_37745,N_35560,N_37473);
and U37746 (N_37746,N_37195,N_36232);
xor U37747 (N_37747,N_37059,N_37284);
and U37748 (N_37748,N_35286,N_35834);
or U37749 (N_37749,N_36730,N_35669);
nand U37750 (N_37750,N_37454,N_37221);
nor U37751 (N_37751,N_36922,N_35027);
xor U37752 (N_37752,N_36890,N_36985);
nand U37753 (N_37753,N_36364,N_36939);
or U37754 (N_37754,N_36097,N_35283);
and U37755 (N_37755,N_35835,N_36072);
xnor U37756 (N_37756,N_36566,N_35135);
xnor U37757 (N_37757,N_36008,N_35474);
nand U37758 (N_37758,N_36460,N_35735);
nand U37759 (N_37759,N_36370,N_35386);
nor U37760 (N_37760,N_37455,N_36412);
nor U37761 (N_37761,N_35203,N_35001);
xnor U37762 (N_37762,N_36677,N_36869);
xnor U37763 (N_37763,N_35365,N_36725);
nand U37764 (N_37764,N_36447,N_36698);
nor U37765 (N_37765,N_36464,N_37305);
nor U37766 (N_37766,N_35650,N_36173);
nand U37767 (N_37767,N_36719,N_35389);
and U37768 (N_37768,N_36614,N_36417);
or U37769 (N_37769,N_35402,N_35431);
xnor U37770 (N_37770,N_36285,N_36833);
and U37771 (N_37771,N_36655,N_35842);
and U37772 (N_37772,N_36284,N_35415);
and U37773 (N_37773,N_35372,N_36971);
nor U37774 (N_37774,N_36674,N_35179);
or U37775 (N_37775,N_37212,N_35182);
or U37776 (N_37776,N_36341,N_37089);
and U37777 (N_37777,N_36425,N_36219);
and U37778 (N_37778,N_35899,N_36266);
xor U37779 (N_37779,N_35928,N_35183);
nand U37780 (N_37780,N_35096,N_37030);
and U37781 (N_37781,N_35657,N_35751);
nor U37782 (N_37782,N_36824,N_37097);
nand U37783 (N_37783,N_35727,N_35576);
nor U37784 (N_37784,N_36501,N_35341);
nor U37785 (N_37785,N_36030,N_35483);
nor U37786 (N_37786,N_37494,N_35375);
or U37787 (N_37787,N_35544,N_35975);
and U37788 (N_37788,N_35434,N_36469);
or U37789 (N_37789,N_36383,N_36007);
nand U37790 (N_37790,N_35311,N_36729);
nor U37791 (N_37791,N_35599,N_36046);
nand U37792 (N_37792,N_36659,N_36728);
xnor U37793 (N_37793,N_36375,N_37460);
xor U37794 (N_37794,N_37111,N_36421);
nand U37795 (N_37795,N_36165,N_36222);
nand U37796 (N_37796,N_35871,N_36935);
nor U37797 (N_37797,N_35590,N_35245);
or U37798 (N_37798,N_35197,N_36757);
nand U37799 (N_37799,N_35979,N_36320);
nor U37800 (N_37800,N_35836,N_35627);
nand U37801 (N_37801,N_35356,N_35974);
and U37802 (N_37802,N_36552,N_36849);
or U37803 (N_37803,N_37397,N_35081);
nor U37804 (N_37804,N_36508,N_36744);
nor U37805 (N_37805,N_36353,N_35034);
nor U37806 (N_37806,N_36801,N_35781);
xnor U37807 (N_37807,N_37035,N_37352);
and U37808 (N_37808,N_37441,N_35660);
nor U37809 (N_37809,N_37357,N_36727);
and U37810 (N_37810,N_36471,N_36620);
xnor U37811 (N_37811,N_37377,N_35532);
or U37812 (N_37812,N_35882,N_37331);
nand U37813 (N_37813,N_36628,N_37464);
nand U37814 (N_37814,N_35317,N_36883);
and U37815 (N_37815,N_36489,N_35990);
nand U37816 (N_37816,N_35583,N_37470);
and U37817 (N_37817,N_36287,N_35510);
nand U37818 (N_37818,N_36348,N_37079);
or U37819 (N_37819,N_36016,N_35308);
nor U37820 (N_37820,N_35458,N_35596);
xor U37821 (N_37821,N_36951,N_35243);
nand U37822 (N_37822,N_37107,N_36130);
or U37823 (N_37823,N_36367,N_35766);
xor U37824 (N_37824,N_36404,N_35230);
nand U37825 (N_37825,N_37115,N_35579);
nand U37826 (N_37826,N_35361,N_36494);
nor U37827 (N_37827,N_37203,N_37304);
nor U37828 (N_37828,N_37275,N_36847);
or U37829 (N_37829,N_37373,N_35102);
nor U37830 (N_37830,N_37188,N_36497);
or U37831 (N_37831,N_35360,N_35819);
and U37832 (N_37832,N_36026,N_35578);
or U37833 (N_37833,N_35511,N_36507);
and U37834 (N_37834,N_36276,N_35848);
or U37835 (N_37835,N_35654,N_37244);
xnor U37836 (N_37836,N_36599,N_36203);
nand U37837 (N_37837,N_36511,N_36063);
nand U37838 (N_37838,N_37015,N_35795);
and U37839 (N_37839,N_35404,N_35612);
nor U37840 (N_37840,N_37322,N_37292);
xor U37841 (N_37841,N_37152,N_35091);
xnor U37842 (N_37842,N_35801,N_37237);
nand U37843 (N_37843,N_36671,N_37281);
nand U37844 (N_37844,N_37072,N_36191);
nand U37845 (N_37845,N_35370,N_35408);
and U37846 (N_37846,N_36210,N_37348);
nand U37847 (N_37847,N_37417,N_35050);
or U37848 (N_37848,N_36111,N_35593);
and U37849 (N_37849,N_35537,N_35955);
nand U37850 (N_37850,N_35670,N_36139);
and U37851 (N_37851,N_36185,N_36120);
nor U37852 (N_37852,N_36243,N_37458);
and U37853 (N_37853,N_35380,N_36778);
xnor U37854 (N_37854,N_36777,N_36178);
nand U37855 (N_37855,N_35384,N_35555);
nor U37856 (N_37856,N_37326,N_37120);
and U37857 (N_37857,N_36946,N_35563);
nand U37858 (N_37858,N_37337,N_35521);
xnor U37859 (N_37859,N_37375,N_35613);
nand U37860 (N_37860,N_35206,N_37182);
or U37861 (N_37861,N_36502,N_35336);
or U37862 (N_37862,N_35833,N_35259);
xnor U37863 (N_37863,N_37101,N_35038);
nand U37864 (N_37864,N_36605,N_35860);
or U37865 (N_37865,N_36694,N_35949);
and U37866 (N_37866,N_35905,N_36732);
or U37867 (N_37867,N_36903,N_37183);
nand U37868 (N_37868,N_36487,N_37363);
nand U37869 (N_37869,N_35134,N_35719);
or U37870 (N_37870,N_36340,N_35111);
and U37871 (N_37871,N_35894,N_36754);
or U37872 (N_37872,N_36850,N_36211);
nand U37873 (N_37873,N_37190,N_36234);
nor U37874 (N_37874,N_35277,N_37016);
nand U37875 (N_37875,N_37409,N_36156);
nand U37876 (N_37876,N_37286,N_36253);
nand U37877 (N_37877,N_37159,N_36439);
and U37878 (N_37878,N_36315,N_36522);
nand U37879 (N_37879,N_35364,N_36182);
and U37880 (N_37880,N_36312,N_35234);
nand U37881 (N_37881,N_36862,N_36932);
xor U37882 (N_37882,N_37285,N_36223);
xnor U37883 (N_37883,N_36475,N_37475);
nor U37884 (N_37884,N_35062,N_36334);
nand U37885 (N_37885,N_35813,N_36540);
nor U37886 (N_37886,N_36576,N_37076);
or U37887 (N_37887,N_36429,N_36245);
xnor U37888 (N_37888,N_37266,N_35122);
nand U37889 (N_37889,N_37206,N_36493);
nor U37890 (N_37890,N_36328,N_35322);
nor U37891 (N_37891,N_36043,N_35820);
or U37892 (N_37892,N_37450,N_36119);
and U37893 (N_37893,N_36525,N_36531);
nand U37894 (N_37894,N_36573,N_36118);
nor U37895 (N_37895,N_35200,N_36816);
xnor U37896 (N_37896,N_36267,N_37290);
or U37897 (N_37897,N_35764,N_36443);
or U37898 (N_37898,N_37062,N_35205);
nor U37899 (N_37899,N_36998,N_36594);
or U37900 (N_37900,N_36350,N_35889);
and U37901 (N_37901,N_37256,N_37383);
or U37902 (N_37902,N_35467,N_35011);
or U37903 (N_37903,N_35265,N_37302);
xnor U37904 (N_37904,N_35128,N_35718);
nor U37905 (N_37905,N_35466,N_36162);
nand U37906 (N_37906,N_37452,N_36924);
nor U37907 (N_37907,N_35157,N_37437);
xor U37908 (N_37908,N_37350,N_36142);
nand U37909 (N_37909,N_35734,N_35708);
nand U37910 (N_37910,N_36791,N_35492);
nand U37911 (N_37911,N_36361,N_35022);
nand U37912 (N_37912,N_37265,N_35999);
or U37913 (N_37913,N_37023,N_37117);
xor U37914 (N_37914,N_36051,N_37178);
nand U37915 (N_37915,N_36982,N_36372);
nand U37916 (N_37916,N_36802,N_37446);
xnor U37917 (N_37917,N_35138,N_36121);
or U37918 (N_37918,N_36057,N_36112);
or U37919 (N_37919,N_37045,N_35060);
or U37920 (N_37920,N_36304,N_36456);
and U37921 (N_37921,N_35094,N_35649);
nand U37922 (N_37922,N_35051,N_37413);
or U37923 (N_37923,N_37004,N_35799);
and U37924 (N_37924,N_36235,N_36174);
nor U37925 (N_37925,N_35496,N_35290);
nand U37926 (N_37926,N_36715,N_35859);
nand U37927 (N_37927,N_37142,N_36419);
or U37928 (N_37928,N_36363,N_35585);
xnor U37929 (N_37929,N_35503,N_35000);
nor U37930 (N_37930,N_35198,N_37484);
or U37931 (N_37931,N_35917,N_36049);
nor U37932 (N_37932,N_36852,N_36548);
or U37933 (N_37933,N_35131,N_35698);
xnor U37934 (N_37934,N_35687,N_35705);
and U37935 (N_37935,N_36969,N_35248);
nor U37936 (N_37936,N_35261,N_36916);
nand U37937 (N_37937,N_35398,N_36619);
nor U37938 (N_37938,N_35754,N_37037);
nor U37939 (N_37939,N_36277,N_35378);
and U37940 (N_37940,N_37430,N_35844);
nor U37941 (N_37941,N_36894,N_35214);
and U37942 (N_37942,N_36673,N_36633);
nand U37943 (N_37943,N_35658,N_37485);
and U37944 (N_37944,N_37368,N_36472);
or U37945 (N_37945,N_37065,N_36129);
nand U37946 (N_37946,N_36938,N_37216);
and U37947 (N_37947,N_37499,N_37407);
nand U37948 (N_37948,N_35043,N_37053);
and U37949 (N_37949,N_36131,N_35114);
and U37950 (N_37950,N_36829,N_35166);
nand U37951 (N_37951,N_35817,N_35802);
and U37952 (N_37952,N_36703,N_36427);
xor U37953 (N_37953,N_35053,N_35268);
nor U37954 (N_37954,N_36152,N_37401);
xor U37955 (N_37955,N_35021,N_35638);
and U37956 (N_37956,N_35215,N_37253);
xor U37957 (N_37957,N_35089,N_36669);
and U37958 (N_37958,N_37020,N_35504);
xnor U37959 (N_37959,N_36362,N_37300);
and U37960 (N_37960,N_36031,N_37044);
nand U37961 (N_37961,N_36240,N_36541);
or U37962 (N_37962,N_35607,N_35530);
nand U37963 (N_37963,N_35195,N_36085);
nand U37964 (N_37964,N_36402,N_36138);
xnor U37965 (N_37965,N_35749,N_36651);
and U37966 (N_37966,N_36753,N_35906);
xor U37967 (N_37967,N_35469,N_35864);
or U37968 (N_37968,N_36076,N_36547);
or U37969 (N_37969,N_36504,N_35861);
or U37970 (N_37970,N_36839,N_37355);
or U37971 (N_37971,N_36289,N_35522);
and U37972 (N_37972,N_36734,N_37421);
or U37973 (N_37973,N_36106,N_35310);
xor U37974 (N_37974,N_36920,N_35520);
nor U37975 (N_37975,N_36200,N_35965);
nand U37976 (N_37976,N_35995,N_35812);
xor U37977 (N_37977,N_37431,N_37445);
nand U37978 (N_37978,N_36512,N_35251);
and U37979 (N_37979,N_35441,N_35991);
or U37980 (N_37980,N_37075,N_35156);
or U37981 (N_37981,N_36546,N_36643);
and U37982 (N_37982,N_35938,N_36405);
or U37983 (N_37983,N_36006,N_37308);
xnor U37984 (N_37984,N_36832,N_36861);
nor U37985 (N_37985,N_37070,N_35099);
nand U37986 (N_37986,N_36403,N_36390);
nor U37987 (N_37987,N_36735,N_35313);
nand U37988 (N_37988,N_37261,N_35723);
xor U37989 (N_37989,N_36600,N_36064);
xor U37990 (N_37990,N_35178,N_36141);
nor U37991 (N_37991,N_36143,N_36825);
or U37992 (N_37992,N_35228,N_36798);
nor U37993 (N_37993,N_35454,N_35069);
xnor U37994 (N_37994,N_37404,N_36554);
and U37995 (N_37995,N_37127,N_35410);
or U37996 (N_37996,N_36317,N_35373);
or U37997 (N_37997,N_36526,N_36668);
and U37998 (N_37998,N_36792,N_36596);
nor U37999 (N_37999,N_37288,N_35193);
xnor U38000 (N_38000,N_35289,N_35154);
nor U38001 (N_38001,N_35895,N_35463);
xnor U38002 (N_38002,N_36964,N_35968);
or U38003 (N_38003,N_35575,N_36571);
and U38004 (N_38004,N_36108,N_36351);
nor U38005 (N_38005,N_35647,N_35396);
and U38006 (N_38006,N_35351,N_35107);
nor U38007 (N_38007,N_36230,N_36410);
nor U38008 (N_38008,N_36061,N_35780);
or U38009 (N_38009,N_37440,N_36936);
and U38010 (N_38010,N_36538,N_35014);
nand U38011 (N_38011,N_36199,N_37057);
nand U38012 (N_38012,N_35023,N_35707);
nand U38013 (N_38013,N_37429,N_35235);
or U38014 (N_38014,N_36401,N_35258);
or U38015 (N_38015,N_36593,N_36314);
nand U38016 (N_38016,N_35850,N_36995);
or U38017 (N_38017,N_35473,N_36054);
nand U38018 (N_38018,N_36058,N_35981);
nand U38019 (N_38019,N_35872,N_36826);
nand U38020 (N_38020,N_35597,N_36217);
nand U38021 (N_38021,N_36776,N_35347);
and U38022 (N_38022,N_37327,N_35071);
and U38023 (N_38023,N_35394,N_35163);
nor U38024 (N_38024,N_35083,N_37425);
xnor U38025 (N_38025,N_36382,N_36823);
and U38026 (N_38026,N_36695,N_36168);
or U38027 (N_38027,N_37391,N_36248);
or U38028 (N_38028,N_36741,N_35927);
nand U38029 (N_38029,N_35338,N_36733);
xnor U38030 (N_38030,N_35256,N_36092);
and U38031 (N_38031,N_35641,N_36692);
and U38032 (N_38032,N_35750,N_35428);
and U38033 (N_38033,N_36081,N_35479);
or U38034 (N_38034,N_37258,N_37449);
or U38035 (N_38035,N_37272,N_36020);
and U38036 (N_38036,N_36179,N_35907);
nor U38037 (N_38037,N_37066,N_37096);
nand U38038 (N_38038,N_36731,N_35216);
or U38039 (N_38039,N_35909,N_37239);
nand U38040 (N_38040,N_35329,N_35212);
nor U38041 (N_38041,N_36283,N_35334);
nor U38042 (N_38042,N_36069,N_36855);
nand U38043 (N_38043,N_36876,N_36202);
or U38044 (N_38044,N_35987,N_35159);
or U38045 (N_38045,N_37314,N_35421);
nor U38046 (N_38046,N_36214,N_35847);
or U38047 (N_38047,N_36667,N_35790);
nand U38048 (N_38048,N_35983,N_36229);
nand U38049 (N_38049,N_35039,N_36192);
and U38050 (N_38050,N_37294,N_35901);
or U38051 (N_38051,N_36070,N_36681);
xnor U38052 (N_38052,N_35939,N_35952);
xor U38053 (N_38053,N_36696,N_36435);
nor U38054 (N_38054,N_37019,N_37427);
and U38055 (N_38055,N_35945,N_35914);
nand U38056 (N_38056,N_36569,N_36079);
or U38057 (N_38057,N_35238,N_36377);
nand U38058 (N_38058,N_37005,N_36622);
xnor U38059 (N_38059,N_35008,N_36711);
or U38060 (N_38060,N_36316,N_36766);
nor U38061 (N_38061,N_36448,N_37296);
xor U38062 (N_38062,N_35606,N_35095);
nor U38063 (N_38063,N_35841,N_35139);
or U38064 (N_38064,N_37268,N_37027);
or U38065 (N_38065,N_36846,N_37315);
nand U38066 (N_38066,N_35699,N_36398);
or U38067 (N_38067,N_35484,N_35616);
and U38068 (N_38068,N_36355,N_35340);
nand U38069 (N_38069,N_36127,N_36208);
nor U38070 (N_38070,N_35132,N_35229);
xor U38071 (N_38071,N_37365,N_35222);
xnor U38072 (N_38072,N_35352,N_36246);
nand U38073 (N_38073,N_35690,N_35035);
nor U38074 (N_38074,N_35885,N_36767);
nand U38075 (N_38075,N_36953,N_35644);
or U38076 (N_38076,N_36761,N_35488);
nand U38077 (N_38077,N_35282,N_37426);
and U38078 (N_38078,N_35685,N_36607);
nor U38079 (N_38079,N_35202,N_36154);
and U38080 (N_38080,N_36524,N_36868);
xor U38081 (N_38081,N_35826,N_36454);
and U38082 (N_38082,N_35838,N_36572);
and U38083 (N_38083,N_37420,N_35739);
nor U38084 (N_38084,N_35867,N_37487);
and U38085 (N_38085,N_35443,N_35395);
nand U38086 (N_38086,N_35634,N_37137);
or U38087 (N_38087,N_36708,N_35024);
and U38088 (N_38088,N_36296,N_36913);
nand U38089 (N_38089,N_35541,N_36424);
or U38090 (N_38090,N_37400,N_35293);
or U38091 (N_38091,N_36999,N_35491);
nand U38092 (N_38092,N_36226,N_36080);
or U38093 (N_38093,N_35884,N_36577);
xnor U38094 (N_38094,N_36662,N_37153);
nand U38095 (N_38095,N_36652,N_37260);
or U38096 (N_38096,N_36249,N_36972);
nand U38097 (N_38097,N_36279,N_36514);
and U38098 (N_38098,N_37254,N_35032);
or U38099 (N_38099,N_37387,N_35296);
nand U38100 (N_38100,N_37259,N_36588);
and U38101 (N_38101,N_35745,N_37359);
or U38102 (N_38102,N_35254,N_37274);
or U38103 (N_38103,N_37121,N_36038);
nor U38104 (N_38104,N_35084,N_35601);
and U38105 (N_38105,N_37241,N_36882);
nand U38106 (N_38106,N_37382,N_35285);
nor U38107 (N_38107,N_35219,N_37138);
xnor U38108 (N_38108,N_36543,N_36087);
nand U38109 (N_38109,N_35921,N_37358);
nand U38110 (N_38110,N_35337,N_36957);
nand U38111 (N_38111,N_36149,N_35571);
or U38112 (N_38112,N_36912,N_37038);
xnor U38113 (N_38113,N_35448,N_36842);
nor U38114 (N_38114,N_35600,N_36153);
xor U38115 (N_38115,N_35862,N_36345);
nor U38116 (N_38116,N_35117,N_37010);
or U38117 (N_38117,N_35877,N_36360);
nand U38118 (N_38118,N_35168,N_37245);
or U38119 (N_38119,N_36990,N_35316);
nand U38120 (N_38120,N_36915,N_36018);
xnor U38121 (N_38121,N_36252,N_35540);
or U38122 (N_38122,N_36161,N_35233);
and U38123 (N_38123,N_37050,N_35515);
or U38124 (N_38124,N_37282,N_35874);
and U38125 (N_38125,N_35295,N_36392);
or U38126 (N_38126,N_36629,N_37220);
nor U38127 (N_38127,N_36298,N_36873);
xnor U38128 (N_38128,N_35460,N_35717);
xnor U38129 (N_38129,N_37098,N_35920);
nand U38130 (N_38130,N_36886,N_35101);
nand U38131 (N_38131,N_35825,N_35539);
and U38132 (N_38132,N_36216,N_35056);
nand U38133 (N_38133,N_35940,N_36896);
nor U38134 (N_38134,N_36591,N_36771);
and U38135 (N_38135,N_37280,N_35811);
xor U38136 (N_38136,N_35536,N_37007);
nor U38137 (N_38137,N_36155,N_36597);
nor U38138 (N_38138,N_35809,N_35327);
and U38139 (N_38139,N_35005,N_36834);
and U38140 (N_38140,N_36270,N_37299);
nand U38141 (N_38141,N_37133,N_35556);
or U38142 (N_38142,N_36408,N_36866);
xnor U38143 (N_38143,N_37328,N_35609);
nor U38144 (N_38144,N_36658,N_35849);
nand U38145 (N_38145,N_37108,N_36053);
and U38146 (N_38146,N_36221,N_35958);
nor U38147 (N_38147,N_35478,N_36561);
nand U38148 (N_38148,N_35605,N_36706);
and U38149 (N_38149,N_35201,N_35470);
and U38150 (N_38150,N_37028,N_36444);
or U38151 (N_38151,N_36828,N_37122);
or U38152 (N_38152,N_35436,N_36840);
nor U38153 (N_38153,N_36970,N_35976);
nand U38154 (N_38154,N_35342,N_37333);
and U38155 (N_38155,N_36386,N_36397);
nor U38156 (N_38156,N_35726,N_36959);
or U38157 (N_38157,N_35012,N_36499);
nand U38158 (N_38158,N_35710,N_37289);
xnor U38159 (N_38159,N_36804,N_35088);
nor U38160 (N_38160,N_35957,N_35080);
nand U38161 (N_38161,N_36399,N_36215);
xor U38162 (N_38162,N_37490,N_37114);
xor U38163 (N_38163,N_36263,N_36366);
and U38164 (N_38164,N_36678,N_36467);
nand U38165 (N_38165,N_36480,N_37438);
and U38166 (N_38166,N_35167,N_35189);
or U38167 (N_38167,N_37344,N_36624);
xnor U38168 (N_38168,N_35267,N_36770);
nand U38169 (N_38169,N_37324,N_36613);
or U38170 (N_38170,N_37262,N_35509);
xnor U38171 (N_38171,N_37342,N_36172);
xor U38172 (N_38172,N_36307,N_35253);
or U38173 (N_38173,N_36559,N_35371);
xor U38174 (N_38174,N_35808,N_36578);
and U38175 (N_38175,N_36942,N_35788);
nor U38176 (N_38176,N_35922,N_35471);
and U38177 (N_38177,N_35815,N_37049);
nand U38178 (N_38178,N_37354,N_35614);
nor U38179 (N_38179,N_35343,N_37148);
nor U38180 (N_38180,N_36003,N_35306);
nand U38181 (N_38181,N_35980,N_35500);
nor U38182 (N_38182,N_36048,N_36763);
or U38183 (N_38183,N_37341,N_36373);
nor U38184 (N_38184,N_37060,N_36535);
and U38185 (N_38185,N_36877,N_37312);
and U38186 (N_38186,N_37480,N_37408);
nor U38187 (N_38187,N_35046,N_35903);
xor U38188 (N_38188,N_36393,N_37029);
or U38189 (N_38189,N_36047,N_36818);
and U38190 (N_38190,N_37227,N_35146);
nand U38191 (N_38191,N_35086,N_35701);
or U38192 (N_38192,N_35947,N_35309);
nor U38193 (N_38193,N_36365,N_36302);
xor U38194 (N_38194,N_36649,N_35608);
or U38195 (N_38195,N_36244,N_35963);
and U38196 (N_38196,N_37223,N_35577);
and U38197 (N_38197,N_37090,N_37054);
or U38198 (N_38198,N_36274,N_37444);
or U38199 (N_38199,N_35925,N_35887);
and U38200 (N_38200,N_36748,N_36617);
or U38201 (N_38201,N_35643,N_36349);
or U38202 (N_38202,N_35300,N_36473);
xor U38203 (N_38203,N_36021,N_35943);
nor U38204 (N_38204,N_36024,N_35472);
nand U38205 (N_38205,N_36657,N_35742);
and U38206 (N_38206,N_35507,N_36369);
nand U38207 (N_38207,N_36028,N_35800);
nand U38208 (N_38208,N_35074,N_36498);
xnor U38209 (N_38209,N_35551,N_37181);
or U38210 (N_38210,N_37412,N_37381);
xor U38211 (N_38211,N_35418,N_37230);
xnor U38212 (N_38212,N_37043,N_36563);
and U38213 (N_38213,N_37067,N_35762);
and U38214 (N_38214,N_37002,N_36720);
nand U38215 (N_38215,N_35376,N_35956);
and U38216 (N_38216,N_37334,N_35076);
nor U38217 (N_38217,N_37240,N_35013);
xor U38218 (N_38218,N_37419,N_35765);
nand U38219 (N_38219,N_35969,N_37347);
xnor U38220 (N_38220,N_36621,N_37384);
nor U38221 (N_38221,N_35489,N_35713);
or U38222 (N_38222,N_36745,N_36157);
and U38223 (N_38223,N_36806,N_35916);
or U38224 (N_38224,N_37074,N_36650);
nor U38225 (N_38225,N_36636,N_35513);
nand U38226 (N_38226,N_37210,N_35006);
nand U38227 (N_38227,N_35640,N_36750);
xor U38228 (N_38228,N_35218,N_37039);
nand U38229 (N_38229,N_36096,N_36413);
nand U38230 (N_38230,N_37385,N_36799);
or U38231 (N_38231,N_35175,N_36615);
nor U38232 (N_38232,N_36814,N_35822);
nor U38233 (N_38233,N_35953,N_36352);
nor U38234 (N_38234,N_37196,N_36803);
xnor U38235 (N_38235,N_35892,N_35582);
nor U38236 (N_38236,N_35049,N_35756);
nand U38237 (N_38237,N_35367,N_37422);
nor U38238 (N_38238,N_36808,N_35424);
xor U38239 (N_38239,N_35246,N_35164);
nand U38240 (N_38240,N_36196,N_35858);
xor U38241 (N_38241,N_36513,N_37224);
or U38242 (N_38242,N_35072,N_36415);
xor U38243 (N_38243,N_35103,N_36251);
nand U38244 (N_38244,N_36584,N_37234);
or U38245 (N_38245,N_35681,N_36261);
xor U38246 (N_38246,N_37451,N_35692);
xnor U38247 (N_38247,N_36262,N_35573);
and U38248 (N_38248,N_36844,N_36705);
nand U38249 (N_38249,N_36411,N_36795);
and U38250 (N_38250,N_36321,N_35516);
xnor U38251 (N_38251,N_37270,N_35988);
nand U38252 (N_38252,N_36432,N_35325);
or U38253 (N_38253,N_37477,N_35941);
nand U38254 (N_38254,N_36984,N_35998);
or U38255 (N_38255,N_36910,N_37104);
nand U38256 (N_38256,N_36269,N_35683);
and U38257 (N_38257,N_35227,N_36292);
xor U38258 (N_38258,N_37000,N_37064);
nor U38259 (N_38259,N_36864,N_36965);
nand U38260 (N_38260,N_35896,N_36575);
or U38261 (N_38261,N_36807,N_36960);
or U38262 (N_38262,N_37463,N_37248);
nor U38263 (N_38263,N_35664,N_35109);
nor U38264 (N_38264,N_36012,N_36474);
and U38265 (N_38265,N_36272,N_37293);
nor U38266 (N_38266,N_36565,N_36384);
and U38267 (N_38267,N_35486,N_36968);
or U38268 (N_38268,N_37298,N_35075);
xor U38269 (N_38269,N_36322,N_35620);
and U38270 (N_38270,N_35320,N_36004);
and U38271 (N_38271,N_36845,N_36158);
xor U38272 (N_38272,N_36793,N_35731);
nor U38273 (N_38273,N_35413,N_36313);
or U38274 (N_38274,N_36137,N_35902);
xor U38275 (N_38275,N_35240,N_35147);
nor U38276 (N_38276,N_35913,N_36585);
nand U38277 (N_38277,N_35188,N_36836);
or U38278 (N_38278,N_35063,N_35312);
or U38279 (N_38279,N_36301,N_36701);
or U38280 (N_38280,N_37112,N_36005);
and U38281 (N_38281,N_36680,N_36376);
nor U38282 (N_38282,N_37317,N_37144);
nand U38283 (N_38283,N_35580,N_37448);
xor U38284 (N_38284,N_37116,N_35204);
and U38285 (N_38285,N_36603,N_35160);
nor U38286 (N_38286,N_35570,N_35855);
and U38287 (N_38287,N_35810,N_36050);
nand U38288 (N_38288,N_36660,N_35199);
xor U38289 (N_38289,N_37058,N_36902);
xor U38290 (N_38290,N_35149,N_36490);
xor U38291 (N_38291,N_37263,N_36510);
nor U38292 (N_38292,N_35535,N_36239);
nor U38293 (N_38293,N_37231,N_36135);
xnor U38294 (N_38294,N_35659,N_35827);
and U38295 (N_38295,N_36863,N_37136);
or U38296 (N_38296,N_35561,N_36934);
nand U38297 (N_38297,N_36627,N_36150);
or U38298 (N_38298,N_36994,N_36874);
or U38299 (N_38299,N_36717,N_37147);
or U38300 (N_38300,N_36528,N_36387);
and U38301 (N_38301,N_37157,N_37246);
or U38302 (N_38302,N_35680,N_36331);
or U38303 (N_38303,N_36870,N_36201);
nand U38304 (N_38304,N_36022,N_35653);
and U38305 (N_38305,N_36553,N_35931);
nand U38306 (N_38306,N_35651,N_37106);
nor U38307 (N_38307,N_35959,N_36640);
nand U38308 (N_38308,N_37174,N_36433);
xnor U38309 (N_38309,N_35665,N_35755);
or U38310 (N_38310,N_37011,N_37194);
xor U38311 (N_38311,N_36032,N_35323);
or U38312 (N_38312,N_36723,N_35773);
nor U38313 (N_38313,N_36140,N_36986);
xnor U38314 (N_38314,N_36319,N_35031);
nand U38315 (N_38315,N_35678,N_35538);
xnor U38316 (N_38316,N_36441,N_36716);
nand U38317 (N_38317,N_35533,N_37389);
or U38318 (N_38318,N_37339,N_37222);
and U38319 (N_38319,N_36002,N_35629);
xor U38320 (N_38320,N_36981,N_35092);
nor U38321 (N_38321,N_36305,N_35505);
or U38322 (N_38322,N_36950,N_35831);
and U38323 (N_38323,N_35055,N_36486);
nor U38324 (N_38324,N_35549,N_37177);
and U38325 (N_38325,N_35112,N_36925);
and U38326 (N_38326,N_35688,N_37180);
and U38327 (N_38327,N_35697,N_37362);
nor U38328 (N_38328,N_35779,N_37215);
nor U38329 (N_38329,N_37130,N_35153);
nor U38330 (N_38330,N_36963,N_36071);
xor U38331 (N_38331,N_37217,N_35740);
and U38332 (N_38332,N_36872,N_37179);
xor U38333 (N_38333,N_35209,N_35758);
or U38334 (N_38334,N_36488,N_37139);
or U38335 (N_38335,N_36909,N_36000);
nand U38336 (N_38336,N_35769,N_36476);
xnor U38337 (N_38337,N_37102,N_35508);
and U38338 (N_38338,N_36449,N_36434);
nor U38339 (N_38339,N_36089,N_36455);
and U38340 (N_38340,N_37443,N_35982);
or U38341 (N_38341,N_36308,N_36009);
nor U38342 (N_38342,N_35078,N_36648);
xor U38343 (N_38343,N_37462,N_37432);
or U38344 (N_38344,N_36227,N_36773);
xnor U38345 (N_38345,N_37423,N_37414);
nand U38346 (N_38346,N_36646,N_36477);
or U38347 (N_38347,N_36407,N_35446);
and U38348 (N_38348,N_36166,N_36452);
nor U38349 (N_38349,N_35064,N_35432);
nand U38350 (N_38350,N_37323,N_36059);
xor U38351 (N_38351,N_36181,N_37479);
or U38352 (N_38352,N_35960,N_36437);
and U38353 (N_38353,N_35173,N_36358);
nand U38354 (N_38354,N_36871,N_37084);
or U38355 (N_38355,N_35042,N_35231);
xor U38356 (N_38356,N_36601,N_35082);
nor U38357 (N_38357,N_36282,N_36450);
xnor U38358 (N_38358,N_36891,N_37082);
nor U38359 (N_38359,N_36623,N_36714);
nand U38360 (N_38360,N_35339,N_36974);
and U38361 (N_38361,N_36483,N_35385);
or U38362 (N_38362,N_37396,N_35633);
nor U38363 (N_38363,N_36207,N_37201);
xnor U38364 (N_38364,N_36290,N_35281);
xnor U38365 (N_38365,N_36647,N_36271);
or U38366 (N_38366,N_37021,N_35004);
and U38367 (N_38367,N_36557,N_36324);
or U38368 (N_38368,N_35948,N_36400);
nand U38369 (N_38369,N_35422,N_35686);
and U38370 (N_38370,N_35052,N_37164);
and U38371 (N_38371,N_37495,N_35878);
or U38372 (N_38372,N_35935,N_36579);
or U38373 (N_38373,N_37307,N_37086);
and U38374 (N_38374,N_35725,N_35962);
or U38375 (N_38375,N_35566,N_36359);
and U38376 (N_38376,N_35747,N_36023);
xor U38377 (N_38377,N_36631,N_36756);
nand U38378 (N_38378,N_35676,N_35796);
or U38379 (N_38379,N_35208,N_35451);
and U38380 (N_38380,N_36592,N_36782);
and U38381 (N_38381,N_37186,N_35785);
nor U38382 (N_38382,N_36688,N_37118);
nor U38383 (N_38383,N_36197,N_35133);
nand U38384 (N_38384,N_36418,N_35097);
nand U38385 (N_38385,N_36675,N_35523);
xor U38386 (N_38386,N_35407,N_35462);
nor U38387 (N_38387,N_36762,N_36568);
and U38388 (N_38388,N_37461,N_35866);
nand U38389 (N_38389,N_37415,N_35733);
nand U38390 (N_38390,N_36718,N_37279);
xnor U38391 (N_38391,N_36430,N_36618);
nor U38392 (N_38392,N_36259,N_37205);
and U38393 (N_38393,N_35554,N_35196);
or U38394 (N_38394,N_35984,N_36634);
and U38395 (N_38395,N_35502,N_35737);
nand U38396 (N_38396,N_37219,N_35715);
nand U38397 (N_38397,N_36052,N_37113);
nor U38398 (N_38398,N_37172,N_35716);
nor U38399 (N_38399,N_35299,N_36895);
or U38400 (N_38400,N_37022,N_36209);
xor U38401 (N_38401,N_36500,N_36911);
xor U38402 (N_38402,N_35388,N_37457);
or U38403 (N_38403,N_35989,N_35026);
and U38404 (N_38404,N_35045,N_35374);
xor U38405 (N_38405,N_36110,N_35623);
nor U38406 (N_38406,N_35433,N_36608);
nor U38407 (N_38407,N_36056,N_36257);
and U38408 (N_38408,N_36713,N_36516);
nor U38409 (N_38409,N_35118,N_36014);
nor U38410 (N_38410,N_35145,N_35668);
and U38411 (N_38411,N_37313,N_37405);
or U38412 (N_38412,N_36768,N_35865);
and U38413 (N_38413,N_36859,N_35986);
xor U38414 (N_38414,N_36707,N_35757);
and U38415 (N_38415,N_36815,N_35724);
xnor U38416 (N_38416,N_36148,N_35252);
and U38417 (N_38417,N_37199,N_35924);
xor U38418 (N_38418,N_36329,N_37269);
xnor U38419 (N_38419,N_36338,N_35677);
nand U38420 (N_38420,N_35040,N_35318);
or U38421 (N_38421,N_35630,N_35170);
nor U38422 (N_38422,N_35752,N_37369);
nor U38423 (N_38423,N_35714,N_35266);
or U38424 (N_38424,N_35420,N_35438);
or U38425 (N_38425,N_35997,N_36664);
and U38426 (N_38426,N_36993,N_36193);
nor U38427 (N_38427,N_37175,N_35648);
xor U38428 (N_38428,N_37123,N_36503);
xor U38429 (N_38429,N_35506,N_37255);
and U38430 (N_38430,N_37338,N_37378);
nor U38431 (N_38431,N_37273,N_35497);
or U38432 (N_38432,N_35349,N_37119);
and U38433 (N_38433,N_36104,N_35517);
xor U38434 (N_38434,N_36884,N_35263);
or U38435 (N_38435,N_36574,N_35591);
nor U38436 (N_38436,N_36697,N_35519);
and U38437 (N_38437,N_35324,N_35951);
nand U38438 (N_38438,N_36509,N_36580);
nand U38439 (N_38439,N_36067,N_36586);
or U38440 (N_38440,N_36183,N_36747);
nor U38441 (N_38441,N_37251,N_35391);
and U38442 (N_38442,N_37218,N_35465);
and U38443 (N_38443,N_37329,N_35598);
nand U38444 (N_38444,N_35007,N_37325);
xor U38445 (N_38445,N_37208,N_37158);
or U38446 (N_38446,N_35452,N_35406);
or U38447 (N_38447,N_37083,N_36176);
and U38448 (N_38448,N_36465,N_35586);
xor U38449 (N_38449,N_35626,N_36780);
nor U38450 (N_38450,N_37467,N_37063);
and U38451 (N_38451,N_37171,N_35891);
nor U38452 (N_38452,N_35652,N_36992);
xnor U38453 (N_38453,N_35116,N_37402);
nand U38454 (N_38454,N_35400,N_37189);
and U38455 (N_38455,N_35970,N_35270);
and U38456 (N_38456,N_37143,N_37003);
or U38457 (N_38457,N_37068,N_36144);
or U38458 (N_38458,N_37134,N_35696);
nor U38459 (N_38459,N_37277,N_36310);
xor U38460 (N_38460,N_36755,N_35994);
nand U38461 (N_38461,N_36928,N_36388);
xnor U38462 (N_38462,N_37497,N_35978);
and U38463 (N_38463,N_35029,N_36693);
or U38464 (N_38464,N_37345,N_36381);
nor U38465 (N_38465,N_35087,N_35743);
xor U38466 (N_38466,N_37073,N_37006);
xor U38467 (N_38467,N_35239,N_35655);
nor U38468 (N_38468,N_36860,N_37471);
xor U38469 (N_38469,N_35712,N_35525);
nor U38470 (N_38470,N_36542,N_35430);
xor U38471 (N_38471,N_36564,N_36286);
and U38472 (N_38472,N_36679,N_36598);
xnor U38473 (N_38473,N_35426,N_36042);
xor U38474 (N_38474,N_35881,N_35783);
nor U38475 (N_38475,N_35457,N_36479);
and U38476 (N_38476,N_36943,N_35656);
nand U38477 (N_38477,N_36604,N_35569);
nor U38478 (N_38478,N_35288,N_35028);
and U38479 (N_38479,N_36019,N_37465);
xnor U38480 (N_38480,N_35942,N_35439);
nand U38481 (N_38481,N_36463,N_35119);
or U38482 (N_38482,N_37191,N_36060);
nand U38483 (N_38483,N_35919,N_36880);
nand U38484 (N_38484,N_35369,N_35335);
nor U38485 (N_38485,N_35414,N_35344);
and U38486 (N_38486,N_37041,N_37018);
xnor U38487 (N_38487,N_35359,N_37192);
and U38488 (N_38488,N_37185,N_36422);
or U38489 (N_38489,N_35048,N_37416);
or U38490 (N_38490,N_35358,N_35155);
nand U38491 (N_38491,N_37173,N_35893);
nand U38492 (N_38492,N_37287,N_35416);
xor U38493 (N_38493,N_35477,N_36103);
and U38494 (N_38494,N_36459,N_35542);
or U38495 (N_38495,N_37466,N_35184);
nand U38496 (N_38496,N_36606,N_35944);
or U38497 (N_38497,N_37489,N_36066);
nand U38498 (N_38498,N_36991,N_36710);
or U38499 (N_38499,N_35223,N_36683);
nand U38500 (N_38500,N_36520,N_35744);
xor U38501 (N_38501,N_35843,N_37001);
xnor U38502 (N_38502,N_36949,N_35332);
and U38503 (N_38503,N_37085,N_36811);
nand U38504 (N_38504,N_36666,N_36354);
nand U38505 (N_38505,N_35171,N_37428);
nand U38506 (N_38506,N_35853,N_36632);
xor U38507 (N_38507,N_36637,N_36937);
nand U38508 (N_38508,N_35588,N_37335);
nor U38509 (N_38509,N_35044,N_37361);
and U38510 (N_38510,N_35232,N_35464);
xnor U38511 (N_38511,N_35297,N_36167);
nor U38512 (N_38512,N_35113,N_36958);
nand U38513 (N_38513,N_37247,N_35821);
xor U38514 (N_38514,N_35770,N_36236);
or U38515 (N_38515,N_36330,N_35803);
and U38516 (N_38516,N_35482,N_35176);
or U38517 (N_38517,N_36740,N_36885);
or U38518 (N_38518,N_36676,N_35568);
nand U38519 (N_38519,N_36505,N_35025);
and U38520 (N_38520,N_36124,N_35187);
or U38521 (N_38521,N_36126,N_35020);
xnor U38522 (N_38522,N_36918,N_36084);
and U38523 (N_38523,N_36721,N_35562);
nor U38524 (N_38524,N_37167,N_35996);
nor U38525 (N_38525,N_35106,N_36395);
nor U38526 (N_38526,N_36264,N_36446);
nor U38527 (N_38527,N_37165,N_35368);
or U38528 (N_38528,N_36297,N_36180);
and U38529 (N_38529,N_36545,N_36379);
or U38530 (N_38530,N_37403,N_35797);
and U38531 (N_38531,N_36682,N_36789);
nor U38532 (N_38532,N_36123,N_36146);
or U38533 (N_38533,N_35009,N_35930);
and U38534 (N_38534,N_36555,N_37303);
and U38535 (N_38535,N_37393,N_36160);
xor U38536 (N_38536,N_36783,N_36134);
nand U38537 (N_38537,N_35280,N_36644);
or U38538 (N_38538,N_35151,N_35152);
or U38539 (N_38539,N_36954,N_35828);
and U38540 (N_38540,N_36927,N_35851);
xnor U38541 (N_38541,N_35883,N_36956);
nand U38542 (N_38542,N_35213,N_35524);
nand U38543 (N_38543,N_35485,N_35330);
and U38544 (N_38544,N_36256,N_36517);
nand U38545 (N_38545,N_35260,N_36409);
nor U38546 (N_38546,N_36765,N_35405);
nor U38547 (N_38547,N_35033,N_35273);
nand U38548 (N_38548,N_37493,N_36967);
or U38549 (N_38549,N_36827,N_36642);
nand U38550 (N_38550,N_36237,N_35814);
nor U38551 (N_38551,N_36233,N_35390);
and U38552 (N_38552,N_35490,N_37370);
nand U38553 (N_38553,N_35355,N_36095);
nor U38554 (N_38554,N_37078,N_36278);
and U38555 (N_38555,N_35264,N_36893);
nor U38556 (N_38556,N_36017,N_37140);
and U38557 (N_38557,N_35362,N_36635);
and U38558 (N_38558,N_36484,N_35127);
xnor U38559 (N_38559,N_35977,N_36529);
and U38560 (N_38560,N_35550,N_36273);
xor U38561 (N_38561,N_35017,N_35936);
nand U38562 (N_38562,N_36309,N_36670);
xnor U38563 (N_38563,N_37081,N_35700);
and U38564 (N_38564,N_37202,N_36300);
nor U38565 (N_38565,N_35691,N_37346);
nor U38566 (N_38566,N_35169,N_37306);
or U38567 (N_38567,N_37232,N_35377);
nand U38568 (N_38568,N_36686,N_37320);
and U38569 (N_38569,N_37214,N_36641);
and U38570 (N_38570,N_37395,N_36800);
nand U38571 (N_38571,N_35868,N_37332);
nor U38572 (N_38572,N_35557,N_36749);
or U38573 (N_38573,N_37410,N_36357);
xnor U38574 (N_38574,N_35140,N_35702);
xor U38575 (N_38575,N_36098,N_36420);
or U38576 (N_38576,N_35236,N_36001);
and U38577 (N_38577,N_36665,N_36281);
nand U38578 (N_38578,N_35125,N_35003);
xnor U38579 (N_38579,N_36337,N_35210);
nor U38580 (N_38580,N_35393,N_35778);
nor U38581 (N_38581,N_35784,N_36125);
or U38582 (N_38582,N_35880,N_35249);
nor U38583 (N_38583,N_36887,N_35041);
or U38584 (N_38584,N_37150,N_36977);
or U38585 (N_38585,N_37009,N_36086);
nand U38586 (N_38586,N_35100,N_36889);
or U38587 (N_38587,N_36857,N_35015);
xnor U38588 (N_38588,N_36029,N_36654);
nand U38589 (N_38589,N_35057,N_37170);
nand U38590 (N_38590,N_36094,N_36099);
nor U38591 (N_38591,N_35581,N_36533);
nand U38592 (N_38592,N_36952,N_36255);
nor U38593 (N_38593,N_37184,N_37469);
and U38594 (N_38594,N_37225,N_37271);
nand U38595 (N_38595,N_37024,N_37424);
nor U38596 (N_38596,N_35602,N_36853);
and U38597 (N_38597,N_37124,N_35798);
nand U38598 (N_38598,N_37093,N_37398);
or U38599 (N_38599,N_35495,N_35946);
xnor U38600 (N_38600,N_35120,N_36940);
nand U38601 (N_38601,N_36461,N_35684);
nor U38602 (N_38602,N_37291,N_36831);
xnor U38603 (N_38603,N_36900,N_35912);
nand U38604 (N_38604,N_35158,N_36980);
or U38605 (N_38605,N_37198,N_36187);
nand U38606 (N_38606,N_35279,N_37486);
xor U38607 (N_38607,N_35854,N_35250);
xnor U38608 (N_38608,N_36626,N_35357);
xnor U38609 (N_38609,N_36702,N_37048);
xor U38610 (N_38610,N_37168,N_36342);
xor U38611 (N_38611,N_36544,N_36639);
nand U38612 (N_38612,N_35237,N_36947);
xnor U38613 (N_38613,N_35501,N_36841);
nor U38614 (N_38614,N_37468,N_37229);
nor U38615 (N_38615,N_35061,N_35933);
nor U38616 (N_38616,N_36093,N_36973);
xor U38617 (N_38617,N_36819,N_35786);
and U38618 (N_38618,N_35759,N_35493);
and U38619 (N_38619,N_36616,N_35499);
and U38620 (N_38620,N_36506,N_35741);
nor U38621 (N_38621,N_36944,N_37226);
nand U38622 (N_38622,N_36128,N_36812);
nand U38623 (N_38623,N_36788,N_35615);
nand U38624 (N_38624,N_36333,N_35307);
or U38625 (N_38625,N_37141,N_36147);
xor U38626 (N_38626,N_35121,N_36436);
xor U38627 (N_38627,N_37207,N_35278);
and U38628 (N_38628,N_35775,N_37135);
or U38629 (N_38629,N_36470,N_35429);
xor U38630 (N_38630,N_35771,N_36055);
or U38631 (N_38631,N_35161,N_36661);
or U38632 (N_38632,N_36481,N_35852);
and U38633 (N_38633,N_35129,N_35010);
nand U38634 (N_38634,N_36881,N_37126);
xor U38635 (N_38635,N_36712,N_35703);
xnor U38636 (N_38636,N_35709,N_35226);
xor U38637 (N_38637,N_36458,N_35674);
or U38638 (N_38638,N_37211,N_36534);
xor U38639 (N_38639,N_35964,N_35257);
nor U38640 (N_38640,N_36638,N_35148);
or U38641 (N_38641,N_35417,N_35093);
xnor U38642 (N_38642,N_35904,N_36684);
nor U38643 (N_38643,N_35444,N_35646);
nor U38644 (N_38644,N_35108,N_36549);
xor U38645 (N_38645,N_36336,N_37481);
nor U38646 (N_38646,N_36040,N_35631);
and U38647 (N_38647,N_36495,N_37160);
nor U38648 (N_38648,N_36821,N_35639);
or U38649 (N_38649,N_35967,N_35314);
nand U38650 (N_38650,N_35255,N_36560);
nor U38651 (N_38651,N_35412,N_35382);
and U38652 (N_38652,N_36091,N_36225);
or U38653 (N_38653,N_37343,N_36133);
and U38654 (N_38654,N_36105,N_36288);
xnor U38655 (N_38655,N_35671,N_35437);
nor U38656 (N_38656,N_36656,N_36796);
xnor U38657 (N_38657,N_36738,N_37351);
and U38658 (N_38658,N_37131,N_35059);
and U38659 (N_38659,N_36978,N_36858);
xnor U38660 (N_38660,N_35736,N_36976);
xor U38661 (N_38661,N_36037,N_37295);
xor U38662 (N_38662,N_36736,N_37166);
xor U38663 (N_38663,N_35126,N_36527);
nand U38664 (N_38664,N_35453,N_36790);
nor U38665 (N_38665,N_35662,N_35105);
nor U38666 (N_38666,N_35622,N_37026);
nor U38667 (N_38667,N_36848,N_36758);
or U38668 (N_38668,N_35185,N_35625);
xor U38669 (N_38669,N_37374,N_37418);
nor U38670 (N_38670,N_35829,N_35066);
xnor U38671 (N_38671,N_37105,N_35174);
nand U38672 (N_38672,N_35141,N_37238);
or U38673 (N_38673,N_36625,N_35419);
nor U38674 (N_38674,N_37434,N_36685);
xor U38675 (N_38675,N_36445,N_35746);
nand U38676 (N_38676,N_35689,N_35328);
nand U38677 (N_38677,N_36159,N_35186);
nand U38678 (N_38678,N_35065,N_35748);
nand U38679 (N_38679,N_36378,N_35787);
or U38680 (N_38680,N_35870,N_35150);
nand U38681 (N_38681,N_37109,N_36082);
and U38682 (N_38682,N_37151,N_35528);
and U38683 (N_38683,N_36228,N_35221);
xor U38684 (N_38684,N_35642,N_37476);
and U38685 (N_38685,N_35366,N_37316);
xnor U38686 (N_38686,N_35918,N_35427);
nand U38687 (N_38687,N_36457,N_37249);
and U38688 (N_38688,N_37492,N_37340);
nor U38689 (N_38689,N_37390,N_37032);
nor U38690 (N_38690,N_36406,N_36523);
and U38691 (N_38691,N_36794,N_37017);
nor U38692 (N_38692,N_36784,N_37129);
and U38693 (N_38693,N_36785,N_35722);
nand U38694 (N_38694,N_37233,N_37439);
xnor U38695 (N_38695,N_35910,N_37204);
nor U38696 (N_38696,N_36485,N_35966);
or U38697 (N_38697,N_35875,N_35704);
nor U38698 (N_38698,N_36878,N_36102);
xnor U38699 (N_38699,N_35098,N_36075);
and U38700 (N_38700,N_37411,N_35276);
nand U38701 (N_38701,N_35604,N_36115);
xor U38702 (N_38702,N_35929,N_37482);
nor U38703 (N_38703,N_36195,N_36482);
nand U38704 (N_38704,N_37336,N_35387);
or U38705 (N_38705,N_37330,N_36224);
and U38706 (N_38706,N_36163,N_37092);
and U38707 (N_38707,N_35682,N_36268);
xor U38708 (N_38708,N_37379,N_37276);
or U38709 (N_38709,N_35534,N_36114);
nor U38710 (N_38710,N_36206,N_37155);
nand U38711 (N_38711,N_36462,N_36726);
xnor U38712 (N_38712,N_37034,N_35879);
and U38713 (N_38713,N_37213,N_36742);
nor U38714 (N_38714,N_35136,N_35837);
nor U38715 (N_38715,N_35191,N_36966);
and U38716 (N_38716,N_35321,N_35442);
xor U38717 (N_38717,N_36587,N_35985);
xor U38718 (N_38718,N_36213,N_35016);
nand U38719 (N_38719,N_36343,N_35194);
and U38720 (N_38720,N_36867,N_36077);
nand U38721 (N_38721,N_36389,N_35805);
and U38722 (N_38722,N_37399,N_36073);
xor U38723 (N_38723,N_36908,N_35461);
xnor U38724 (N_38724,N_35661,N_35584);
nor U38725 (N_38725,N_36010,N_35675);
nand U38726 (N_38726,N_35181,N_35241);
xnor U38727 (N_38727,N_37435,N_36491);
and U38728 (N_38728,N_35073,N_36035);
or U38729 (N_38729,N_36478,N_37367);
or U38730 (N_38730,N_37267,N_35666);
xor U38731 (N_38731,N_36396,N_37483);
and U38732 (N_38732,N_37311,N_35818);
and U38733 (N_38733,N_36151,N_37132);
xor U38734 (N_38734,N_35886,N_35326);
or U38735 (N_38735,N_35993,N_37356);
xor U38736 (N_38736,N_36786,N_36772);
or U38737 (N_38737,N_35130,N_35294);
or U38738 (N_38738,N_35476,N_36416);
nor U38739 (N_38739,N_36303,N_35932);
nand U38740 (N_38740,N_35177,N_35494);
and U38741 (N_38741,N_36558,N_36339);
nor U38742 (N_38742,N_35793,N_35768);
nand U38743 (N_38743,N_36537,N_37088);
or U38744 (N_38744,N_35782,N_35950);
or U38745 (N_38745,N_36769,N_36630);
nand U38746 (N_38746,N_37364,N_35123);
and U38747 (N_38747,N_36875,N_37042);
or U38748 (N_38748,N_36595,N_36438);
or U38749 (N_38749,N_35900,N_36332);
nor U38750 (N_38750,N_36853,N_35506);
nor U38751 (N_38751,N_35796,N_35448);
or U38752 (N_38752,N_35374,N_35091);
nor U38753 (N_38753,N_35771,N_36763);
nand U38754 (N_38754,N_37048,N_36108);
nor U38755 (N_38755,N_35214,N_36642);
xor U38756 (N_38756,N_36094,N_35108);
xnor U38757 (N_38757,N_35180,N_35736);
and U38758 (N_38758,N_37050,N_37412);
nand U38759 (N_38759,N_36574,N_36794);
and U38760 (N_38760,N_35058,N_35907);
or U38761 (N_38761,N_36927,N_36142);
and U38762 (N_38762,N_35644,N_35643);
or U38763 (N_38763,N_35814,N_35635);
or U38764 (N_38764,N_36312,N_35724);
or U38765 (N_38765,N_36147,N_35249);
nor U38766 (N_38766,N_36907,N_36174);
and U38767 (N_38767,N_37355,N_35037);
nor U38768 (N_38768,N_36314,N_36419);
and U38769 (N_38769,N_35225,N_35875);
nor U38770 (N_38770,N_36654,N_36593);
or U38771 (N_38771,N_36817,N_36911);
nor U38772 (N_38772,N_35014,N_35925);
xnor U38773 (N_38773,N_36794,N_36402);
nor U38774 (N_38774,N_35698,N_36614);
and U38775 (N_38775,N_35131,N_37307);
and U38776 (N_38776,N_36065,N_35896);
xnor U38777 (N_38777,N_36391,N_37257);
nand U38778 (N_38778,N_35449,N_36529);
xor U38779 (N_38779,N_37406,N_37476);
or U38780 (N_38780,N_35256,N_35426);
xnor U38781 (N_38781,N_35680,N_36327);
nor U38782 (N_38782,N_37256,N_35104);
or U38783 (N_38783,N_36654,N_35956);
or U38784 (N_38784,N_36559,N_35252);
or U38785 (N_38785,N_36517,N_36089);
nand U38786 (N_38786,N_35129,N_35372);
nor U38787 (N_38787,N_35432,N_35068);
xor U38788 (N_38788,N_35175,N_35733);
nand U38789 (N_38789,N_37343,N_36426);
nor U38790 (N_38790,N_35339,N_37163);
nand U38791 (N_38791,N_36897,N_36683);
nand U38792 (N_38792,N_36834,N_35755);
nor U38793 (N_38793,N_36494,N_35619);
nor U38794 (N_38794,N_36450,N_36779);
xnor U38795 (N_38795,N_35164,N_36169);
nor U38796 (N_38796,N_35665,N_35997);
or U38797 (N_38797,N_36231,N_36669);
or U38798 (N_38798,N_36696,N_36707);
nor U38799 (N_38799,N_37227,N_37021);
xor U38800 (N_38800,N_35965,N_35438);
and U38801 (N_38801,N_36243,N_36127);
and U38802 (N_38802,N_37184,N_35869);
xnor U38803 (N_38803,N_37067,N_35722);
nand U38804 (N_38804,N_37219,N_35671);
nand U38805 (N_38805,N_36420,N_36837);
and U38806 (N_38806,N_37411,N_35846);
xor U38807 (N_38807,N_37040,N_37135);
or U38808 (N_38808,N_36575,N_36525);
nor U38809 (N_38809,N_35261,N_35089);
nor U38810 (N_38810,N_36905,N_35955);
nand U38811 (N_38811,N_35062,N_37307);
and U38812 (N_38812,N_36267,N_35771);
or U38813 (N_38813,N_37296,N_36726);
xnor U38814 (N_38814,N_35458,N_36650);
nand U38815 (N_38815,N_35106,N_36660);
and U38816 (N_38816,N_35003,N_36606);
nand U38817 (N_38817,N_37476,N_36808);
nor U38818 (N_38818,N_36964,N_36429);
xor U38819 (N_38819,N_37019,N_37300);
nand U38820 (N_38820,N_35611,N_35022);
nand U38821 (N_38821,N_36115,N_35690);
xor U38822 (N_38822,N_36768,N_37251);
xnor U38823 (N_38823,N_36628,N_36736);
nor U38824 (N_38824,N_35968,N_36868);
and U38825 (N_38825,N_37308,N_36343);
or U38826 (N_38826,N_37006,N_36115);
and U38827 (N_38827,N_36135,N_36142);
xnor U38828 (N_38828,N_35770,N_36217);
and U38829 (N_38829,N_37087,N_36157);
and U38830 (N_38830,N_35607,N_35491);
nor U38831 (N_38831,N_36309,N_36902);
and U38832 (N_38832,N_35823,N_35603);
nor U38833 (N_38833,N_37387,N_37315);
and U38834 (N_38834,N_35448,N_35417);
nor U38835 (N_38835,N_35873,N_35937);
and U38836 (N_38836,N_35166,N_36887);
xor U38837 (N_38837,N_35957,N_36684);
xnor U38838 (N_38838,N_35223,N_37253);
or U38839 (N_38839,N_36669,N_36832);
or U38840 (N_38840,N_37228,N_37415);
nor U38841 (N_38841,N_35231,N_35177);
or U38842 (N_38842,N_36053,N_36511);
xor U38843 (N_38843,N_35223,N_35073);
xor U38844 (N_38844,N_36238,N_35369);
nor U38845 (N_38845,N_35205,N_35442);
nor U38846 (N_38846,N_37386,N_35393);
or U38847 (N_38847,N_37345,N_36934);
nand U38848 (N_38848,N_37015,N_37358);
or U38849 (N_38849,N_36236,N_36268);
or U38850 (N_38850,N_35378,N_37109);
nand U38851 (N_38851,N_35963,N_36544);
or U38852 (N_38852,N_37423,N_36348);
or U38853 (N_38853,N_37050,N_37475);
or U38854 (N_38854,N_37177,N_37017);
and U38855 (N_38855,N_35010,N_36085);
nor U38856 (N_38856,N_35837,N_35512);
nand U38857 (N_38857,N_36025,N_35014);
nand U38858 (N_38858,N_36352,N_35430);
nand U38859 (N_38859,N_37403,N_35561);
and U38860 (N_38860,N_35707,N_37100);
nor U38861 (N_38861,N_35936,N_35526);
and U38862 (N_38862,N_35124,N_35976);
and U38863 (N_38863,N_36537,N_35630);
nand U38864 (N_38864,N_36721,N_35822);
nand U38865 (N_38865,N_35044,N_35021);
and U38866 (N_38866,N_37071,N_35238);
nand U38867 (N_38867,N_36332,N_35565);
nand U38868 (N_38868,N_37169,N_35764);
xor U38869 (N_38869,N_36839,N_37348);
or U38870 (N_38870,N_35389,N_37137);
and U38871 (N_38871,N_35346,N_36315);
nand U38872 (N_38872,N_36387,N_35550);
or U38873 (N_38873,N_35361,N_35616);
nand U38874 (N_38874,N_37154,N_37142);
nand U38875 (N_38875,N_36592,N_35562);
and U38876 (N_38876,N_35122,N_36833);
xor U38877 (N_38877,N_35386,N_36306);
and U38878 (N_38878,N_36428,N_35517);
nor U38879 (N_38879,N_37057,N_36327);
and U38880 (N_38880,N_35192,N_35777);
nand U38881 (N_38881,N_36162,N_35338);
nor U38882 (N_38882,N_37217,N_35608);
and U38883 (N_38883,N_36718,N_35788);
and U38884 (N_38884,N_35577,N_37208);
and U38885 (N_38885,N_35475,N_35189);
and U38886 (N_38886,N_36126,N_35425);
nor U38887 (N_38887,N_37145,N_36003);
xor U38888 (N_38888,N_37058,N_35015);
and U38889 (N_38889,N_36393,N_37363);
nor U38890 (N_38890,N_37012,N_35483);
nand U38891 (N_38891,N_36334,N_35182);
or U38892 (N_38892,N_35981,N_35896);
or U38893 (N_38893,N_35369,N_36093);
nor U38894 (N_38894,N_35768,N_37074);
and U38895 (N_38895,N_35532,N_35674);
and U38896 (N_38896,N_35726,N_37261);
nand U38897 (N_38897,N_36059,N_36434);
nand U38898 (N_38898,N_36998,N_37269);
or U38899 (N_38899,N_37172,N_36236);
nor U38900 (N_38900,N_37373,N_37034);
xor U38901 (N_38901,N_35423,N_35196);
and U38902 (N_38902,N_36643,N_35045);
nor U38903 (N_38903,N_37476,N_36956);
nand U38904 (N_38904,N_36990,N_36440);
or U38905 (N_38905,N_37305,N_36286);
or U38906 (N_38906,N_35549,N_36206);
or U38907 (N_38907,N_35563,N_37343);
nand U38908 (N_38908,N_36838,N_35552);
xor U38909 (N_38909,N_37386,N_35716);
nor U38910 (N_38910,N_35795,N_37250);
xnor U38911 (N_38911,N_35702,N_35082);
and U38912 (N_38912,N_37183,N_36994);
nor U38913 (N_38913,N_35394,N_35072);
or U38914 (N_38914,N_35675,N_35866);
nand U38915 (N_38915,N_36365,N_36053);
nor U38916 (N_38916,N_36238,N_36378);
xnor U38917 (N_38917,N_35803,N_36569);
and U38918 (N_38918,N_35742,N_36906);
nand U38919 (N_38919,N_35483,N_35631);
and U38920 (N_38920,N_35053,N_36224);
nor U38921 (N_38921,N_37037,N_35748);
and U38922 (N_38922,N_35045,N_36838);
nor U38923 (N_38923,N_36484,N_36383);
nand U38924 (N_38924,N_35711,N_36822);
or U38925 (N_38925,N_36735,N_36648);
xor U38926 (N_38926,N_35853,N_37090);
nand U38927 (N_38927,N_35529,N_35701);
nand U38928 (N_38928,N_35971,N_37238);
xnor U38929 (N_38929,N_35663,N_35353);
nor U38930 (N_38930,N_37128,N_36018);
nor U38931 (N_38931,N_35802,N_36037);
nand U38932 (N_38932,N_36991,N_35858);
nor U38933 (N_38933,N_37074,N_35391);
and U38934 (N_38934,N_35694,N_36170);
xor U38935 (N_38935,N_37423,N_35095);
or U38936 (N_38936,N_35519,N_36992);
nand U38937 (N_38937,N_36011,N_35196);
xor U38938 (N_38938,N_36774,N_37397);
or U38939 (N_38939,N_36378,N_37304);
and U38940 (N_38940,N_37004,N_35655);
xor U38941 (N_38941,N_37305,N_36331);
nand U38942 (N_38942,N_35143,N_35745);
nand U38943 (N_38943,N_35582,N_36974);
or U38944 (N_38944,N_36501,N_35180);
or U38945 (N_38945,N_35284,N_36615);
and U38946 (N_38946,N_35713,N_35749);
xnor U38947 (N_38947,N_35788,N_35554);
or U38948 (N_38948,N_36691,N_36203);
nor U38949 (N_38949,N_35475,N_36589);
and U38950 (N_38950,N_35780,N_36901);
nor U38951 (N_38951,N_36711,N_35083);
nand U38952 (N_38952,N_35130,N_35961);
nand U38953 (N_38953,N_36192,N_36264);
or U38954 (N_38954,N_37292,N_35234);
nand U38955 (N_38955,N_35901,N_35042);
and U38956 (N_38956,N_35754,N_36952);
nor U38957 (N_38957,N_36645,N_37175);
xor U38958 (N_38958,N_35957,N_36630);
and U38959 (N_38959,N_35854,N_37460);
or U38960 (N_38960,N_35927,N_36034);
and U38961 (N_38961,N_36952,N_35767);
nand U38962 (N_38962,N_35693,N_35422);
or U38963 (N_38963,N_36746,N_36780);
and U38964 (N_38964,N_36323,N_36759);
or U38965 (N_38965,N_36173,N_36437);
xnor U38966 (N_38966,N_35135,N_35890);
nor U38967 (N_38967,N_36623,N_35497);
nand U38968 (N_38968,N_35848,N_37150);
nor U38969 (N_38969,N_35685,N_35797);
and U38970 (N_38970,N_36253,N_36654);
and U38971 (N_38971,N_36032,N_36691);
nor U38972 (N_38972,N_35302,N_35433);
and U38973 (N_38973,N_36696,N_37458);
and U38974 (N_38974,N_37367,N_35172);
nand U38975 (N_38975,N_37170,N_36936);
and U38976 (N_38976,N_37294,N_37409);
and U38977 (N_38977,N_36577,N_35790);
nor U38978 (N_38978,N_36397,N_36541);
xor U38979 (N_38979,N_35722,N_36606);
nand U38980 (N_38980,N_35463,N_36210);
and U38981 (N_38981,N_37241,N_35269);
or U38982 (N_38982,N_35927,N_36009);
or U38983 (N_38983,N_37392,N_35610);
nand U38984 (N_38984,N_35212,N_36780);
or U38985 (N_38985,N_35612,N_35800);
xor U38986 (N_38986,N_35714,N_35255);
nor U38987 (N_38987,N_35310,N_35398);
nor U38988 (N_38988,N_35682,N_36684);
nor U38989 (N_38989,N_35090,N_35424);
nor U38990 (N_38990,N_35557,N_36260);
and U38991 (N_38991,N_36167,N_35836);
or U38992 (N_38992,N_35792,N_37321);
nor U38993 (N_38993,N_35351,N_36524);
or U38994 (N_38994,N_35069,N_37154);
nor U38995 (N_38995,N_36770,N_36444);
or U38996 (N_38996,N_36104,N_35746);
nand U38997 (N_38997,N_35856,N_35062);
or U38998 (N_38998,N_35055,N_36879);
nor U38999 (N_38999,N_35764,N_37092);
xor U39000 (N_39000,N_35224,N_36862);
or U39001 (N_39001,N_35380,N_36766);
and U39002 (N_39002,N_36371,N_36044);
nor U39003 (N_39003,N_37113,N_37270);
and U39004 (N_39004,N_37354,N_37172);
xnor U39005 (N_39005,N_35375,N_35737);
and U39006 (N_39006,N_35803,N_36712);
and U39007 (N_39007,N_36038,N_37197);
nand U39008 (N_39008,N_35655,N_35200);
or U39009 (N_39009,N_35985,N_35830);
xor U39010 (N_39010,N_35985,N_35848);
xnor U39011 (N_39011,N_36862,N_36318);
xor U39012 (N_39012,N_36255,N_36515);
nor U39013 (N_39013,N_35425,N_37497);
nand U39014 (N_39014,N_35006,N_36737);
nor U39015 (N_39015,N_35018,N_36011);
xor U39016 (N_39016,N_36577,N_35330);
nor U39017 (N_39017,N_37480,N_37323);
nor U39018 (N_39018,N_36661,N_35041);
nor U39019 (N_39019,N_35601,N_35487);
or U39020 (N_39020,N_35423,N_36061);
and U39021 (N_39021,N_36581,N_36749);
and U39022 (N_39022,N_35645,N_36069);
nand U39023 (N_39023,N_35648,N_36723);
nor U39024 (N_39024,N_36394,N_35493);
and U39025 (N_39025,N_36346,N_37113);
and U39026 (N_39026,N_35432,N_36803);
nor U39027 (N_39027,N_35780,N_36860);
nor U39028 (N_39028,N_36885,N_37308);
xnor U39029 (N_39029,N_36988,N_36696);
xnor U39030 (N_39030,N_36487,N_37217);
nor U39031 (N_39031,N_36617,N_37062);
nand U39032 (N_39032,N_36788,N_36849);
or U39033 (N_39033,N_37004,N_36537);
nor U39034 (N_39034,N_36313,N_36250);
or U39035 (N_39035,N_37307,N_35867);
or U39036 (N_39036,N_36569,N_35868);
nor U39037 (N_39037,N_36953,N_35047);
or U39038 (N_39038,N_36296,N_35616);
xor U39039 (N_39039,N_37159,N_35919);
or U39040 (N_39040,N_36243,N_35701);
and U39041 (N_39041,N_36311,N_35961);
nor U39042 (N_39042,N_35195,N_36178);
nor U39043 (N_39043,N_35622,N_35399);
or U39044 (N_39044,N_37394,N_36161);
nand U39045 (N_39045,N_37185,N_35577);
and U39046 (N_39046,N_35770,N_35743);
and U39047 (N_39047,N_35276,N_36743);
or U39048 (N_39048,N_36187,N_35616);
nor U39049 (N_39049,N_36691,N_36587);
and U39050 (N_39050,N_35778,N_36247);
nand U39051 (N_39051,N_35496,N_35674);
and U39052 (N_39052,N_35440,N_36628);
nor U39053 (N_39053,N_35698,N_35211);
and U39054 (N_39054,N_36822,N_35844);
and U39055 (N_39055,N_35570,N_37404);
xor U39056 (N_39056,N_36785,N_37462);
or U39057 (N_39057,N_36362,N_36883);
and U39058 (N_39058,N_35668,N_37287);
xnor U39059 (N_39059,N_36081,N_35398);
nor U39060 (N_39060,N_35426,N_36223);
or U39061 (N_39061,N_36131,N_36099);
nor U39062 (N_39062,N_37318,N_36545);
xor U39063 (N_39063,N_36026,N_36210);
or U39064 (N_39064,N_36247,N_36887);
and U39065 (N_39065,N_36879,N_35182);
nand U39066 (N_39066,N_35355,N_37398);
nand U39067 (N_39067,N_35583,N_36285);
nor U39068 (N_39068,N_35496,N_35657);
xnor U39069 (N_39069,N_35019,N_35450);
or U39070 (N_39070,N_35767,N_37177);
nand U39071 (N_39071,N_35533,N_35789);
and U39072 (N_39072,N_36165,N_36238);
nand U39073 (N_39073,N_35505,N_35551);
xnor U39074 (N_39074,N_37245,N_35759);
and U39075 (N_39075,N_35661,N_35263);
xnor U39076 (N_39076,N_35314,N_36663);
and U39077 (N_39077,N_37243,N_37391);
and U39078 (N_39078,N_36920,N_36930);
xnor U39079 (N_39079,N_35104,N_35250);
and U39080 (N_39080,N_35245,N_37150);
xnor U39081 (N_39081,N_35777,N_35933);
and U39082 (N_39082,N_35849,N_35203);
nor U39083 (N_39083,N_36094,N_36658);
nand U39084 (N_39084,N_36325,N_36452);
xnor U39085 (N_39085,N_36855,N_35826);
xnor U39086 (N_39086,N_35881,N_35173);
or U39087 (N_39087,N_36670,N_36807);
xor U39088 (N_39088,N_35321,N_37206);
nand U39089 (N_39089,N_36843,N_35556);
nor U39090 (N_39090,N_35290,N_35528);
nand U39091 (N_39091,N_36783,N_36148);
nand U39092 (N_39092,N_37193,N_35640);
and U39093 (N_39093,N_35009,N_36902);
or U39094 (N_39094,N_36050,N_37293);
xnor U39095 (N_39095,N_36370,N_36377);
nand U39096 (N_39096,N_36255,N_37446);
xnor U39097 (N_39097,N_35767,N_36384);
nand U39098 (N_39098,N_36040,N_36808);
or U39099 (N_39099,N_35673,N_36832);
nand U39100 (N_39100,N_36834,N_36629);
nor U39101 (N_39101,N_35985,N_36340);
or U39102 (N_39102,N_35048,N_36995);
xor U39103 (N_39103,N_36634,N_37345);
and U39104 (N_39104,N_35414,N_36244);
nor U39105 (N_39105,N_35574,N_35946);
xor U39106 (N_39106,N_36860,N_37210);
xnor U39107 (N_39107,N_35851,N_35949);
nand U39108 (N_39108,N_35293,N_35194);
xor U39109 (N_39109,N_36671,N_36250);
and U39110 (N_39110,N_35538,N_36780);
and U39111 (N_39111,N_35223,N_35791);
or U39112 (N_39112,N_35842,N_35460);
nor U39113 (N_39113,N_37049,N_37102);
nand U39114 (N_39114,N_37290,N_36613);
or U39115 (N_39115,N_37110,N_35173);
nor U39116 (N_39116,N_36656,N_37120);
or U39117 (N_39117,N_37000,N_35172);
nand U39118 (N_39118,N_35703,N_36124);
nor U39119 (N_39119,N_35261,N_36437);
or U39120 (N_39120,N_36773,N_35828);
xnor U39121 (N_39121,N_36454,N_35282);
and U39122 (N_39122,N_35274,N_37046);
xor U39123 (N_39123,N_36489,N_35681);
nor U39124 (N_39124,N_36854,N_35568);
or U39125 (N_39125,N_35118,N_36289);
or U39126 (N_39126,N_35786,N_35689);
nor U39127 (N_39127,N_35567,N_36560);
xnor U39128 (N_39128,N_35426,N_36766);
xnor U39129 (N_39129,N_35580,N_35799);
or U39130 (N_39130,N_37307,N_35917);
and U39131 (N_39131,N_35735,N_37211);
or U39132 (N_39132,N_36574,N_36665);
nor U39133 (N_39133,N_35837,N_36925);
and U39134 (N_39134,N_35908,N_36543);
nand U39135 (N_39135,N_35200,N_35818);
or U39136 (N_39136,N_36470,N_35188);
nand U39137 (N_39137,N_36719,N_35731);
and U39138 (N_39138,N_36696,N_36371);
or U39139 (N_39139,N_35747,N_37102);
nor U39140 (N_39140,N_36912,N_36058);
or U39141 (N_39141,N_37082,N_36287);
nand U39142 (N_39142,N_36799,N_36403);
and U39143 (N_39143,N_36734,N_37342);
and U39144 (N_39144,N_35152,N_36085);
and U39145 (N_39145,N_35609,N_37029);
and U39146 (N_39146,N_37241,N_35838);
nor U39147 (N_39147,N_36430,N_36425);
nand U39148 (N_39148,N_36185,N_36152);
xnor U39149 (N_39149,N_36300,N_35720);
nand U39150 (N_39150,N_35797,N_35743);
and U39151 (N_39151,N_36561,N_35563);
nor U39152 (N_39152,N_36051,N_36456);
nor U39153 (N_39153,N_35430,N_35325);
nor U39154 (N_39154,N_37015,N_35313);
and U39155 (N_39155,N_35934,N_36103);
nand U39156 (N_39156,N_37210,N_36808);
nor U39157 (N_39157,N_36447,N_35602);
or U39158 (N_39158,N_36417,N_35388);
nor U39159 (N_39159,N_35811,N_35138);
or U39160 (N_39160,N_36957,N_35508);
or U39161 (N_39161,N_35266,N_36252);
nand U39162 (N_39162,N_36314,N_36953);
xnor U39163 (N_39163,N_35897,N_35720);
nor U39164 (N_39164,N_37092,N_36959);
nor U39165 (N_39165,N_37261,N_35227);
xor U39166 (N_39166,N_36965,N_35705);
and U39167 (N_39167,N_37328,N_36809);
nor U39168 (N_39168,N_37238,N_36428);
or U39169 (N_39169,N_35444,N_36133);
and U39170 (N_39170,N_37425,N_35410);
xor U39171 (N_39171,N_35705,N_35903);
nor U39172 (N_39172,N_36028,N_35242);
xor U39173 (N_39173,N_35713,N_36984);
nand U39174 (N_39174,N_35464,N_37399);
nor U39175 (N_39175,N_35676,N_35545);
nor U39176 (N_39176,N_37326,N_35525);
or U39177 (N_39177,N_37038,N_36366);
nor U39178 (N_39178,N_36748,N_37014);
and U39179 (N_39179,N_35399,N_35290);
nor U39180 (N_39180,N_37204,N_36317);
or U39181 (N_39181,N_35391,N_37020);
nor U39182 (N_39182,N_36052,N_37161);
and U39183 (N_39183,N_36945,N_35330);
or U39184 (N_39184,N_35855,N_36814);
and U39185 (N_39185,N_36013,N_35610);
xnor U39186 (N_39186,N_35904,N_35471);
nor U39187 (N_39187,N_36310,N_35467);
nand U39188 (N_39188,N_37119,N_35541);
or U39189 (N_39189,N_37207,N_35116);
nor U39190 (N_39190,N_36135,N_35926);
or U39191 (N_39191,N_37403,N_35545);
xor U39192 (N_39192,N_35567,N_35424);
nand U39193 (N_39193,N_35139,N_35629);
nand U39194 (N_39194,N_36387,N_35816);
xnor U39195 (N_39195,N_35851,N_35835);
xor U39196 (N_39196,N_37364,N_37149);
and U39197 (N_39197,N_35472,N_35209);
nand U39198 (N_39198,N_36174,N_36089);
or U39199 (N_39199,N_36557,N_37345);
nand U39200 (N_39200,N_36271,N_35219);
nor U39201 (N_39201,N_35647,N_35222);
xor U39202 (N_39202,N_35438,N_37479);
and U39203 (N_39203,N_35101,N_37298);
and U39204 (N_39204,N_36221,N_37014);
nand U39205 (N_39205,N_35319,N_35429);
and U39206 (N_39206,N_35868,N_35110);
nand U39207 (N_39207,N_35108,N_36099);
nor U39208 (N_39208,N_36365,N_37498);
nor U39209 (N_39209,N_35259,N_36315);
nor U39210 (N_39210,N_37105,N_35758);
nand U39211 (N_39211,N_37361,N_36409);
nor U39212 (N_39212,N_36379,N_37032);
or U39213 (N_39213,N_35391,N_37481);
nand U39214 (N_39214,N_37298,N_35283);
nand U39215 (N_39215,N_35620,N_36014);
nand U39216 (N_39216,N_36846,N_37256);
nand U39217 (N_39217,N_36914,N_35735);
nor U39218 (N_39218,N_35368,N_37235);
nor U39219 (N_39219,N_35302,N_35636);
nand U39220 (N_39220,N_35220,N_35501);
nand U39221 (N_39221,N_36045,N_36173);
and U39222 (N_39222,N_37372,N_36807);
xor U39223 (N_39223,N_35581,N_37084);
nor U39224 (N_39224,N_36916,N_35161);
and U39225 (N_39225,N_36116,N_36393);
nor U39226 (N_39226,N_36347,N_36914);
nor U39227 (N_39227,N_36979,N_37019);
xor U39228 (N_39228,N_35047,N_36318);
or U39229 (N_39229,N_36502,N_35025);
or U39230 (N_39230,N_37478,N_36381);
xnor U39231 (N_39231,N_36809,N_36091);
nand U39232 (N_39232,N_35861,N_35199);
nand U39233 (N_39233,N_36822,N_37150);
nor U39234 (N_39234,N_36663,N_35473);
and U39235 (N_39235,N_35466,N_37203);
xnor U39236 (N_39236,N_35013,N_36232);
xor U39237 (N_39237,N_37483,N_36386);
and U39238 (N_39238,N_35482,N_37351);
nand U39239 (N_39239,N_35374,N_36372);
and U39240 (N_39240,N_35737,N_36041);
xnor U39241 (N_39241,N_36955,N_36415);
and U39242 (N_39242,N_36099,N_35929);
nor U39243 (N_39243,N_36938,N_36930);
nand U39244 (N_39244,N_37374,N_37478);
nand U39245 (N_39245,N_36767,N_35263);
nor U39246 (N_39246,N_36169,N_35004);
or U39247 (N_39247,N_35540,N_35431);
and U39248 (N_39248,N_35433,N_36210);
nand U39249 (N_39249,N_36778,N_36526);
nand U39250 (N_39250,N_35924,N_37277);
or U39251 (N_39251,N_35835,N_35409);
or U39252 (N_39252,N_35143,N_36579);
or U39253 (N_39253,N_35740,N_36874);
nor U39254 (N_39254,N_35336,N_36094);
nand U39255 (N_39255,N_36076,N_35969);
xor U39256 (N_39256,N_35190,N_36465);
or U39257 (N_39257,N_36605,N_36662);
or U39258 (N_39258,N_36769,N_35748);
and U39259 (N_39259,N_35367,N_35580);
nor U39260 (N_39260,N_37433,N_35394);
nor U39261 (N_39261,N_37028,N_35149);
nor U39262 (N_39262,N_36118,N_36688);
or U39263 (N_39263,N_35737,N_35649);
and U39264 (N_39264,N_36356,N_35518);
xnor U39265 (N_39265,N_35172,N_35622);
xnor U39266 (N_39266,N_35179,N_36921);
and U39267 (N_39267,N_36974,N_36102);
nand U39268 (N_39268,N_35068,N_35327);
nand U39269 (N_39269,N_35207,N_35526);
and U39270 (N_39270,N_36292,N_36566);
xor U39271 (N_39271,N_35206,N_37494);
or U39272 (N_39272,N_36601,N_35367);
nor U39273 (N_39273,N_35973,N_35415);
xnor U39274 (N_39274,N_35064,N_35223);
xnor U39275 (N_39275,N_35920,N_35173);
nand U39276 (N_39276,N_36836,N_37402);
nor U39277 (N_39277,N_37211,N_36074);
nand U39278 (N_39278,N_35141,N_36467);
or U39279 (N_39279,N_35706,N_37059);
or U39280 (N_39280,N_37341,N_35352);
and U39281 (N_39281,N_37380,N_35383);
or U39282 (N_39282,N_35849,N_35768);
xnor U39283 (N_39283,N_36815,N_37150);
or U39284 (N_39284,N_36696,N_35901);
and U39285 (N_39285,N_36507,N_37234);
nor U39286 (N_39286,N_35132,N_35901);
or U39287 (N_39287,N_35903,N_36667);
nor U39288 (N_39288,N_36778,N_36060);
nor U39289 (N_39289,N_37038,N_36597);
or U39290 (N_39290,N_36544,N_35322);
and U39291 (N_39291,N_37175,N_37168);
and U39292 (N_39292,N_36468,N_36337);
and U39293 (N_39293,N_35078,N_37295);
or U39294 (N_39294,N_37359,N_35454);
xnor U39295 (N_39295,N_35152,N_35844);
or U39296 (N_39296,N_35341,N_36301);
xor U39297 (N_39297,N_35336,N_35818);
or U39298 (N_39298,N_35238,N_36884);
nor U39299 (N_39299,N_37069,N_35135);
or U39300 (N_39300,N_35064,N_36001);
or U39301 (N_39301,N_35217,N_35222);
nor U39302 (N_39302,N_35505,N_35185);
xor U39303 (N_39303,N_36349,N_35278);
xor U39304 (N_39304,N_37127,N_35081);
nand U39305 (N_39305,N_36503,N_35595);
and U39306 (N_39306,N_35267,N_36036);
and U39307 (N_39307,N_36452,N_36623);
nand U39308 (N_39308,N_36884,N_35074);
nor U39309 (N_39309,N_36792,N_35005);
xor U39310 (N_39310,N_35208,N_37051);
and U39311 (N_39311,N_36263,N_36285);
or U39312 (N_39312,N_35690,N_37357);
or U39313 (N_39313,N_36575,N_37144);
nand U39314 (N_39314,N_35808,N_35861);
nand U39315 (N_39315,N_37313,N_37242);
or U39316 (N_39316,N_36870,N_37013);
and U39317 (N_39317,N_37087,N_37162);
xnor U39318 (N_39318,N_35940,N_35466);
xor U39319 (N_39319,N_35302,N_37468);
xnor U39320 (N_39320,N_36446,N_35133);
nor U39321 (N_39321,N_36465,N_36168);
or U39322 (N_39322,N_35905,N_35179);
nor U39323 (N_39323,N_35413,N_35366);
and U39324 (N_39324,N_36765,N_35326);
and U39325 (N_39325,N_35534,N_35611);
and U39326 (N_39326,N_36517,N_36309);
or U39327 (N_39327,N_35177,N_36187);
nor U39328 (N_39328,N_35982,N_36263);
xnor U39329 (N_39329,N_36329,N_35528);
nor U39330 (N_39330,N_35383,N_36992);
or U39331 (N_39331,N_35200,N_36730);
or U39332 (N_39332,N_35150,N_36418);
nand U39333 (N_39333,N_35345,N_37190);
nand U39334 (N_39334,N_36612,N_36897);
or U39335 (N_39335,N_35498,N_37193);
or U39336 (N_39336,N_35689,N_37367);
or U39337 (N_39337,N_36479,N_37009);
nor U39338 (N_39338,N_35092,N_36841);
nor U39339 (N_39339,N_35027,N_35764);
nor U39340 (N_39340,N_35307,N_35682);
and U39341 (N_39341,N_35976,N_35168);
xnor U39342 (N_39342,N_36952,N_35493);
nand U39343 (N_39343,N_35900,N_36680);
nor U39344 (N_39344,N_35303,N_35058);
xor U39345 (N_39345,N_35025,N_36187);
xnor U39346 (N_39346,N_36974,N_35305);
xor U39347 (N_39347,N_36162,N_37430);
xor U39348 (N_39348,N_35860,N_37119);
or U39349 (N_39349,N_35211,N_35822);
xnor U39350 (N_39350,N_35921,N_36785);
and U39351 (N_39351,N_35833,N_36030);
nor U39352 (N_39352,N_36056,N_36963);
nor U39353 (N_39353,N_37116,N_36970);
nor U39354 (N_39354,N_37333,N_35857);
and U39355 (N_39355,N_37337,N_35750);
xor U39356 (N_39356,N_35599,N_35758);
and U39357 (N_39357,N_36248,N_35240);
xor U39358 (N_39358,N_37010,N_37141);
and U39359 (N_39359,N_35138,N_37106);
or U39360 (N_39360,N_37213,N_37174);
nor U39361 (N_39361,N_36741,N_35740);
and U39362 (N_39362,N_35560,N_37091);
and U39363 (N_39363,N_36147,N_37243);
and U39364 (N_39364,N_35368,N_35005);
nand U39365 (N_39365,N_37194,N_37083);
xnor U39366 (N_39366,N_36178,N_37440);
nand U39367 (N_39367,N_36901,N_36553);
or U39368 (N_39368,N_36212,N_36283);
xnor U39369 (N_39369,N_36134,N_36538);
nand U39370 (N_39370,N_35352,N_36180);
and U39371 (N_39371,N_35555,N_35820);
and U39372 (N_39372,N_36133,N_35536);
or U39373 (N_39373,N_35566,N_37399);
and U39374 (N_39374,N_36423,N_35325);
nor U39375 (N_39375,N_36212,N_35454);
nand U39376 (N_39376,N_35520,N_36010);
nor U39377 (N_39377,N_35366,N_35058);
nand U39378 (N_39378,N_35661,N_35623);
or U39379 (N_39379,N_36191,N_36600);
nand U39380 (N_39380,N_37242,N_35994);
or U39381 (N_39381,N_35879,N_35651);
nor U39382 (N_39382,N_35445,N_35683);
or U39383 (N_39383,N_37439,N_36611);
and U39384 (N_39384,N_37092,N_35423);
nor U39385 (N_39385,N_36713,N_36178);
nand U39386 (N_39386,N_35138,N_35697);
xnor U39387 (N_39387,N_36463,N_36357);
nand U39388 (N_39388,N_35353,N_35098);
nand U39389 (N_39389,N_37397,N_36220);
and U39390 (N_39390,N_35795,N_37281);
nor U39391 (N_39391,N_35251,N_36676);
and U39392 (N_39392,N_35534,N_37108);
nor U39393 (N_39393,N_37312,N_36285);
xor U39394 (N_39394,N_35536,N_35871);
nor U39395 (N_39395,N_35076,N_36367);
nor U39396 (N_39396,N_36602,N_37276);
nand U39397 (N_39397,N_36353,N_37401);
nor U39398 (N_39398,N_36472,N_37184);
and U39399 (N_39399,N_37449,N_35943);
nor U39400 (N_39400,N_37294,N_37355);
nand U39401 (N_39401,N_37458,N_36718);
and U39402 (N_39402,N_36353,N_36818);
nand U39403 (N_39403,N_36080,N_37134);
nand U39404 (N_39404,N_36626,N_36926);
nor U39405 (N_39405,N_35155,N_35147);
and U39406 (N_39406,N_37111,N_37101);
nor U39407 (N_39407,N_37478,N_35215);
nor U39408 (N_39408,N_35984,N_35303);
or U39409 (N_39409,N_36320,N_35313);
xor U39410 (N_39410,N_35248,N_36600);
nand U39411 (N_39411,N_37325,N_36551);
xor U39412 (N_39412,N_35043,N_36133);
xnor U39413 (N_39413,N_35609,N_35006);
nor U39414 (N_39414,N_36366,N_35958);
nand U39415 (N_39415,N_36607,N_37395);
or U39416 (N_39416,N_35618,N_35564);
nand U39417 (N_39417,N_35015,N_36362);
or U39418 (N_39418,N_36779,N_36884);
nor U39419 (N_39419,N_37266,N_36660);
or U39420 (N_39420,N_36500,N_35908);
and U39421 (N_39421,N_36217,N_36646);
or U39422 (N_39422,N_36054,N_37397);
or U39423 (N_39423,N_35579,N_37428);
nor U39424 (N_39424,N_37392,N_35644);
xor U39425 (N_39425,N_37348,N_35309);
nor U39426 (N_39426,N_36500,N_37116);
xor U39427 (N_39427,N_35332,N_36762);
or U39428 (N_39428,N_37152,N_37111);
nand U39429 (N_39429,N_36936,N_35199);
nand U39430 (N_39430,N_36656,N_36782);
or U39431 (N_39431,N_36490,N_36967);
nor U39432 (N_39432,N_36093,N_37493);
nand U39433 (N_39433,N_36338,N_35943);
nand U39434 (N_39434,N_36887,N_35978);
and U39435 (N_39435,N_36072,N_37045);
or U39436 (N_39436,N_37380,N_35949);
or U39437 (N_39437,N_36325,N_37431);
and U39438 (N_39438,N_36441,N_37045);
or U39439 (N_39439,N_35658,N_35707);
and U39440 (N_39440,N_35578,N_36833);
and U39441 (N_39441,N_37385,N_35632);
xor U39442 (N_39442,N_36289,N_36849);
and U39443 (N_39443,N_35291,N_36099);
and U39444 (N_39444,N_35865,N_35662);
and U39445 (N_39445,N_37385,N_35240);
nand U39446 (N_39446,N_36902,N_35664);
nand U39447 (N_39447,N_36171,N_35879);
nor U39448 (N_39448,N_36474,N_36560);
nor U39449 (N_39449,N_36012,N_36517);
or U39450 (N_39450,N_37142,N_35273);
nand U39451 (N_39451,N_37268,N_36991);
nor U39452 (N_39452,N_36345,N_35504);
xnor U39453 (N_39453,N_36316,N_36576);
xor U39454 (N_39454,N_37229,N_35052);
nor U39455 (N_39455,N_36151,N_35342);
and U39456 (N_39456,N_35767,N_35272);
and U39457 (N_39457,N_35537,N_35909);
or U39458 (N_39458,N_36523,N_36087);
xor U39459 (N_39459,N_35295,N_36180);
nand U39460 (N_39460,N_35887,N_36694);
and U39461 (N_39461,N_36857,N_35357);
and U39462 (N_39462,N_36303,N_37055);
nor U39463 (N_39463,N_35228,N_36026);
nor U39464 (N_39464,N_36315,N_36038);
or U39465 (N_39465,N_35007,N_37016);
nand U39466 (N_39466,N_36648,N_35409);
and U39467 (N_39467,N_36457,N_37373);
or U39468 (N_39468,N_36611,N_37108);
and U39469 (N_39469,N_36484,N_35143);
or U39470 (N_39470,N_36169,N_35801);
nand U39471 (N_39471,N_35135,N_36640);
nand U39472 (N_39472,N_37237,N_35444);
nand U39473 (N_39473,N_35131,N_36954);
nand U39474 (N_39474,N_35441,N_37227);
nand U39475 (N_39475,N_36498,N_36737);
and U39476 (N_39476,N_37048,N_35705);
nor U39477 (N_39477,N_36477,N_35553);
and U39478 (N_39478,N_35550,N_36435);
and U39479 (N_39479,N_37173,N_36944);
and U39480 (N_39480,N_36666,N_36768);
or U39481 (N_39481,N_36728,N_37325);
and U39482 (N_39482,N_36815,N_36488);
nand U39483 (N_39483,N_35862,N_35902);
and U39484 (N_39484,N_36773,N_36747);
or U39485 (N_39485,N_36563,N_35662);
nor U39486 (N_39486,N_35058,N_35038);
nand U39487 (N_39487,N_35225,N_37113);
and U39488 (N_39488,N_37266,N_36307);
nor U39489 (N_39489,N_36123,N_35505);
and U39490 (N_39490,N_36285,N_37139);
xnor U39491 (N_39491,N_36580,N_36678);
or U39492 (N_39492,N_36315,N_36986);
nand U39493 (N_39493,N_36598,N_35267);
xnor U39494 (N_39494,N_36481,N_35978);
nor U39495 (N_39495,N_35015,N_36517);
xor U39496 (N_39496,N_36159,N_36033);
and U39497 (N_39497,N_35676,N_36619);
nor U39498 (N_39498,N_36887,N_35802);
nor U39499 (N_39499,N_36362,N_35020);
or U39500 (N_39500,N_37071,N_36935);
nand U39501 (N_39501,N_36924,N_36710);
nand U39502 (N_39502,N_36412,N_35094);
or U39503 (N_39503,N_35116,N_36839);
and U39504 (N_39504,N_37453,N_36702);
nand U39505 (N_39505,N_35845,N_36164);
nand U39506 (N_39506,N_35012,N_35854);
nand U39507 (N_39507,N_35881,N_37201);
nand U39508 (N_39508,N_37256,N_37080);
nand U39509 (N_39509,N_35198,N_36881);
xor U39510 (N_39510,N_37085,N_35567);
or U39511 (N_39511,N_36745,N_35609);
nand U39512 (N_39512,N_36200,N_35117);
nor U39513 (N_39513,N_35392,N_36865);
or U39514 (N_39514,N_36669,N_35819);
nand U39515 (N_39515,N_37039,N_37397);
xor U39516 (N_39516,N_36895,N_35584);
nand U39517 (N_39517,N_35080,N_36090);
nor U39518 (N_39518,N_36943,N_35116);
and U39519 (N_39519,N_36927,N_36775);
xnor U39520 (N_39520,N_37154,N_37223);
nand U39521 (N_39521,N_36866,N_36811);
nor U39522 (N_39522,N_36383,N_35478);
xor U39523 (N_39523,N_36384,N_35415);
nand U39524 (N_39524,N_36876,N_36538);
xnor U39525 (N_39525,N_35785,N_36227);
or U39526 (N_39526,N_36887,N_35607);
or U39527 (N_39527,N_35305,N_37013);
xor U39528 (N_39528,N_37358,N_37248);
nor U39529 (N_39529,N_36876,N_36581);
and U39530 (N_39530,N_37154,N_37474);
and U39531 (N_39531,N_36351,N_36754);
or U39532 (N_39532,N_37093,N_35509);
xnor U39533 (N_39533,N_36965,N_35156);
and U39534 (N_39534,N_37477,N_36189);
and U39535 (N_39535,N_36581,N_35147);
or U39536 (N_39536,N_35419,N_35614);
nand U39537 (N_39537,N_36214,N_37087);
nor U39538 (N_39538,N_36975,N_35684);
nor U39539 (N_39539,N_35738,N_36589);
nor U39540 (N_39540,N_36820,N_35022);
or U39541 (N_39541,N_37145,N_35193);
nor U39542 (N_39542,N_35058,N_35133);
or U39543 (N_39543,N_36704,N_37025);
or U39544 (N_39544,N_35975,N_36911);
nand U39545 (N_39545,N_37213,N_35764);
and U39546 (N_39546,N_36191,N_37119);
or U39547 (N_39547,N_35648,N_35255);
xor U39548 (N_39548,N_36890,N_36308);
xnor U39549 (N_39549,N_36593,N_35825);
and U39550 (N_39550,N_36773,N_37211);
xor U39551 (N_39551,N_36959,N_37152);
and U39552 (N_39552,N_35668,N_37268);
xor U39553 (N_39553,N_37396,N_37012);
or U39554 (N_39554,N_37451,N_36366);
nand U39555 (N_39555,N_37209,N_36885);
nand U39556 (N_39556,N_36854,N_35464);
nand U39557 (N_39557,N_37404,N_37428);
nand U39558 (N_39558,N_35102,N_37330);
or U39559 (N_39559,N_35355,N_35102);
or U39560 (N_39560,N_36409,N_35393);
and U39561 (N_39561,N_36028,N_35872);
and U39562 (N_39562,N_35223,N_36618);
nor U39563 (N_39563,N_37065,N_35579);
or U39564 (N_39564,N_36725,N_36245);
or U39565 (N_39565,N_37411,N_37436);
nor U39566 (N_39566,N_36462,N_37488);
nor U39567 (N_39567,N_35026,N_36204);
nand U39568 (N_39568,N_35789,N_35908);
nor U39569 (N_39569,N_36984,N_36631);
xor U39570 (N_39570,N_35376,N_36707);
nor U39571 (N_39571,N_36329,N_36249);
or U39572 (N_39572,N_36334,N_37029);
and U39573 (N_39573,N_35176,N_35752);
and U39574 (N_39574,N_36238,N_35003);
nor U39575 (N_39575,N_36635,N_36573);
or U39576 (N_39576,N_35180,N_37450);
xor U39577 (N_39577,N_35645,N_37400);
xnor U39578 (N_39578,N_36337,N_35421);
xor U39579 (N_39579,N_35592,N_36533);
nor U39580 (N_39580,N_36703,N_35333);
nor U39581 (N_39581,N_36429,N_35931);
or U39582 (N_39582,N_36599,N_35962);
nor U39583 (N_39583,N_36397,N_35748);
nor U39584 (N_39584,N_36255,N_36001);
xnor U39585 (N_39585,N_35380,N_36367);
nand U39586 (N_39586,N_36966,N_36388);
nor U39587 (N_39587,N_37387,N_37108);
or U39588 (N_39588,N_37234,N_36728);
nand U39589 (N_39589,N_36322,N_35110);
nand U39590 (N_39590,N_35423,N_37181);
xor U39591 (N_39591,N_36153,N_37065);
xnor U39592 (N_39592,N_36344,N_37257);
nand U39593 (N_39593,N_35541,N_36929);
xor U39594 (N_39594,N_35318,N_36769);
or U39595 (N_39595,N_37445,N_36850);
or U39596 (N_39596,N_37465,N_36334);
nand U39597 (N_39597,N_35026,N_36351);
xor U39598 (N_39598,N_36560,N_36041);
and U39599 (N_39599,N_35429,N_37265);
nand U39600 (N_39600,N_36482,N_36605);
xnor U39601 (N_39601,N_35292,N_36641);
nand U39602 (N_39602,N_35894,N_37317);
xnor U39603 (N_39603,N_36076,N_35931);
nand U39604 (N_39604,N_36942,N_37267);
nand U39605 (N_39605,N_36543,N_37330);
xor U39606 (N_39606,N_35685,N_37260);
and U39607 (N_39607,N_37359,N_35974);
nand U39608 (N_39608,N_37093,N_36268);
xor U39609 (N_39609,N_35561,N_37174);
or U39610 (N_39610,N_35999,N_36684);
xnor U39611 (N_39611,N_35504,N_36022);
or U39612 (N_39612,N_37124,N_36792);
or U39613 (N_39613,N_35222,N_35170);
xnor U39614 (N_39614,N_35630,N_36085);
and U39615 (N_39615,N_36027,N_35778);
nand U39616 (N_39616,N_36196,N_36707);
nand U39617 (N_39617,N_35908,N_35478);
nor U39618 (N_39618,N_37462,N_36222);
nand U39619 (N_39619,N_35837,N_35321);
xnor U39620 (N_39620,N_37228,N_36773);
xnor U39621 (N_39621,N_37321,N_37018);
or U39622 (N_39622,N_36137,N_35278);
nand U39623 (N_39623,N_36167,N_36144);
nor U39624 (N_39624,N_35069,N_35967);
nor U39625 (N_39625,N_36916,N_35313);
xnor U39626 (N_39626,N_35695,N_36488);
nor U39627 (N_39627,N_35707,N_36064);
or U39628 (N_39628,N_36763,N_35490);
or U39629 (N_39629,N_36446,N_35025);
and U39630 (N_39630,N_36190,N_37173);
nor U39631 (N_39631,N_37301,N_37210);
xnor U39632 (N_39632,N_36013,N_36905);
nand U39633 (N_39633,N_35255,N_35189);
nor U39634 (N_39634,N_35127,N_37071);
xor U39635 (N_39635,N_36906,N_37214);
nand U39636 (N_39636,N_35587,N_36461);
nand U39637 (N_39637,N_36493,N_35422);
xor U39638 (N_39638,N_36008,N_36998);
nand U39639 (N_39639,N_35081,N_37262);
xnor U39640 (N_39640,N_35453,N_36306);
and U39641 (N_39641,N_37054,N_36010);
nor U39642 (N_39642,N_36349,N_37042);
nand U39643 (N_39643,N_36608,N_35563);
and U39644 (N_39644,N_35517,N_36429);
xor U39645 (N_39645,N_35325,N_35031);
xnor U39646 (N_39646,N_36241,N_36854);
nand U39647 (N_39647,N_36208,N_37363);
or U39648 (N_39648,N_35073,N_35511);
or U39649 (N_39649,N_37008,N_36834);
nor U39650 (N_39650,N_35380,N_37461);
xor U39651 (N_39651,N_36450,N_35895);
and U39652 (N_39652,N_37498,N_37327);
xor U39653 (N_39653,N_37110,N_35395);
xor U39654 (N_39654,N_35423,N_35955);
nor U39655 (N_39655,N_35899,N_35665);
nand U39656 (N_39656,N_36687,N_36738);
nor U39657 (N_39657,N_35837,N_36210);
or U39658 (N_39658,N_35243,N_35300);
or U39659 (N_39659,N_35574,N_37073);
nand U39660 (N_39660,N_37302,N_36579);
or U39661 (N_39661,N_37414,N_35560);
nor U39662 (N_39662,N_36149,N_35265);
and U39663 (N_39663,N_35161,N_35431);
xnor U39664 (N_39664,N_36550,N_35457);
xor U39665 (N_39665,N_35921,N_36521);
nand U39666 (N_39666,N_35523,N_35140);
nand U39667 (N_39667,N_35663,N_36176);
and U39668 (N_39668,N_35069,N_36460);
and U39669 (N_39669,N_36073,N_36795);
xnor U39670 (N_39670,N_37369,N_35609);
nor U39671 (N_39671,N_36779,N_36515);
xor U39672 (N_39672,N_36823,N_35754);
or U39673 (N_39673,N_35469,N_35185);
xnor U39674 (N_39674,N_35131,N_35429);
or U39675 (N_39675,N_36485,N_36585);
xnor U39676 (N_39676,N_36009,N_35971);
and U39677 (N_39677,N_35894,N_36149);
and U39678 (N_39678,N_36700,N_37004);
or U39679 (N_39679,N_36530,N_36637);
nand U39680 (N_39680,N_35216,N_36580);
xor U39681 (N_39681,N_35430,N_35098);
and U39682 (N_39682,N_36726,N_36717);
and U39683 (N_39683,N_35640,N_36017);
or U39684 (N_39684,N_35448,N_35906);
xor U39685 (N_39685,N_36415,N_37427);
nor U39686 (N_39686,N_35013,N_35158);
xor U39687 (N_39687,N_35115,N_36885);
and U39688 (N_39688,N_35966,N_36121);
xnor U39689 (N_39689,N_35679,N_37456);
nor U39690 (N_39690,N_37213,N_36704);
or U39691 (N_39691,N_35941,N_35215);
nand U39692 (N_39692,N_35735,N_36353);
nor U39693 (N_39693,N_35795,N_37237);
nor U39694 (N_39694,N_36460,N_36749);
and U39695 (N_39695,N_36183,N_35194);
or U39696 (N_39696,N_35709,N_35765);
and U39697 (N_39697,N_37241,N_35297);
xor U39698 (N_39698,N_35404,N_35357);
nor U39699 (N_39699,N_36178,N_36175);
or U39700 (N_39700,N_35872,N_35301);
nor U39701 (N_39701,N_36415,N_36356);
nor U39702 (N_39702,N_35847,N_35537);
xnor U39703 (N_39703,N_37455,N_35482);
nor U39704 (N_39704,N_36811,N_35221);
nor U39705 (N_39705,N_35028,N_37321);
and U39706 (N_39706,N_37472,N_36068);
nand U39707 (N_39707,N_37324,N_37225);
and U39708 (N_39708,N_35378,N_36693);
xnor U39709 (N_39709,N_35475,N_35599);
xor U39710 (N_39710,N_36353,N_36336);
xor U39711 (N_39711,N_35102,N_36415);
xnor U39712 (N_39712,N_36196,N_37010);
xnor U39713 (N_39713,N_36184,N_35671);
nor U39714 (N_39714,N_35079,N_35331);
nand U39715 (N_39715,N_35460,N_35787);
nor U39716 (N_39716,N_36368,N_36261);
xnor U39717 (N_39717,N_36379,N_36633);
nor U39718 (N_39718,N_36150,N_36268);
or U39719 (N_39719,N_35516,N_36637);
xnor U39720 (N_39720,N_36538,N_36148);
nand U39721 (N_39721,N_36243,N_35717);
and U39722 (N_39722,N_36689,N_36603);
xnor U39723 (N_39723,N_35434,N_36167);
xnor U39724 (N_39724,N_36207,N_35566);
nor U39725 (N_39725,N_35618,N_35797);
xor U39726 (N_39726,N_37498,N_35115);
nor U39727 (N_39727,N_35794,N_35763);
and U39728 (N_39728,N_35943,N_36003);
nor U39729 (N_39729,N_36387,N_36113);
and U39730 (N_39730,N_35380,N_35839);
nor U39731 (N_39731,N_37035,N_36211);
nor U39732 (N_39732,N_36261,N_36561);
and U39733 (N_39733,N_35398,N_35719);
xnor U39734 (N_39734,N_36687,N_36147);
or U39735 (N_39735,N_36891,N_36582);
xnor U39736 (N_39736,N_36497,N_37240);
and U39737 (N_39737,N_36109,N_36803);
and U39738 (N_39738,N_36862,N_35301);
or U39739 (N_39739,N_35562,N_35000);
and U39740 (N_39740,N_36952,N_35066);
xnor U39741 (N_39741,N_35030,N_37302);
nor U39742 (N_39742,N_35259,N_35386);
nor U39743 (N_39743,N_35398,N_36066);
or U39744 (N_39744,N_35015,N_35939);
nand U39745 (N_39745,N_36687,N_35382);
nor U39746 (N_39746,N_36226,N_36070);
xor U39747 (N_39747,N_37132,N_35649);
or U39748 (N_39748,N_36151,N_35334);
xor U39749 (N_39749,N_35814,N_37096);
or U39750 (N_39750,N_37243,N_36500);
or U39751 (N_39751,N_35767,N_37250);
nor U39752 (N_39752,N_36467,N_36782);
xor U39753 (N_39753,N_36466,N_35377);
nand U39754 (N_39754,N_35334,N_36449);
or U39755 (N_39755,N_36527,N_35140);
xnor U39756 (N_39756,N_37334,N_36297);
and U39757 (N_39757,N_37449,N_36437);
or U39758 (N_39758,N_36905,N_37093);
and U39759 (N_39759,N_36858,N_37395);
xor U39760 (N_39760,N_35540,N_35514);
or U39761 (N_39761,N_37419,N_37216);
nand U39762 (N_39762,N_37007,N_36642);
nor U39763 (N_39763,N_35439,N_35237);
nand U39764 (N_39764,N_36052,N_37416);
xor U39765 (N_39765,N_36108,N_37066);
or U39766 (N_39766,N_36525,N_37072);
and U39767 (N_39767,N_35266,N_35873);
nand U39768 (N_39768,N_37267,N_35686);
and U39769 (N_39769,N_36334,N_37080);
and U39770 (N_39770,N_37048,N_36911);
nand U39771 (N_39771,N_36922,N_36363);
and U39772 (N_39772,N_36781,N_36276);
xor U39773 (N_39773,N_37313,N_36096);
or U39774 (N_39774,N_37098,N_36129);
or U39775 (N_39775,N_36498,N_36590);
nor U39776 (N_39776,N_36098,N_36200);
and U39777 (N_39777,N_36699,N_37065);
xor U39778 (N_39778,N_37369,N_35909);
or U39779 (N_39779,N_36488,N_35694);
or U39780 (N_39780,N_35532,N_35264);
xnor U39781 (N_39781,N_35335,N_35993);
xor U39782 (N_39782,N_35426,N_35263);
or U39783 (N_39783,N_35108,N_37438);
and U39784 (N_39784,N_36026,N_35600);
or U39785 (N_39785,N_35814,N_36335);
or U39786 (N_39786,N_35457,N_36038);
and U39787 (N_39787,N_35702,N_35843);
nor U39788 (N_39788,N_37476,N_36313);
xor U39789 (N_39789,N_36146,N_35188);
nand U39790 (N_39790,N_37289,N_36493);
xor U39791 (N_39791,N_37136,N_36529);
nand U39792 (N_39792,N_36590,N_35338);
xnor U39793 (N_39793,N_36039,N_36424);
nor U39794 (N_39794,N_37308,N_36440);
or U39795 (N_39795,N_35068,N_35946);
nand U39796 (N_39796,N_35895,N_35849);
nor U39797 (N_39797,N_36880,N_37438);
or U39798 (N_39798,N_35756,N_36906);
nor U39799 (N_39799,N_36315,N_35104);
xnor U39800 (N_39800,N_36221,N_36851);
nor U39801 (N_39801,N_35439,N_37465);
xor U39802 (N_39802,N_36779,N_36626);
nand U39803 (N_39803,N_35827,N_35059);
or U39804 (N_39804,N_35893,N_35139);
xnor U39805 (N_39805,N_36986,N_36191);
nor U39806 (N_39806,N_35659,N_36035);
nand U39807 (N_39807,N_37103,N_35456);
nand U39808 (N_39808,N_35422,N_35596);
and U39809 (N_39809,N_36501,N_37322);
nand U39810 (N_39810,N_35622,N_36113);
xor U39811 (N_39811,N_36183,N_35683);
nand U39812 (N_39812,N_36007,N_36543);
nand U39813 (N_39813,N_37415,N_35380);
or U39814 (N_39814,N_36763,N_35697);
xor U39815 (N_39815,N_36779,N_36529);
and U39816 (N_39816,N_35646,N_37492);
nor U39817 (N_39817,N_37433,N_35357);
nor U39818 (N_39818,N_36442,N_37166);
xor U39819 (N_39819,N_36994,N_36828);
nor U39820 (N_39820,N_36536,N_35428);
nand U39821 (N_39821,N_36323,N_35305);
nor U39822 (N_39822,N_36437,N_36014);
nor U39823 (N_39823,N_36651,N_36894);
or U39824 (N_39824,N_36408,N_37298);
nor U39825 (N_39825,N_36844,N_35460);
xor U39826 (N_39826,N_36323,N_37483);
nor U39827 (N_39827,N_37471,N_35106);
nor U39828 (N_39828,N_37217,N_36356);
and U39829 (N_39829,N_36174,N_37076);
nor U39830 (N_39830,N_37416,N_35898);
and U39831 (N_39831,N_35977,N_36015);
and U39832 (N_39832,N_35142,N_36848);
or U39833 (N_39833,N_35084,N_35505);
xor U39834 (N_39834,N_36098,N_36981);
or U39835 (N_39835,N_36763,N_35388);
xor U39836 (N_39836,N_37436,N_36801);
or U39837 (N_39837,N_35754,N_35318);
xor U39838 (N_39838,N_36739,N_37046);
and U39839 (N_39839,N_37330,N_36529);
and U39840 (N_39840,N_35360,N_36870);
and U39841 (N_39841,N_37092,N_35866);
nand U39842 (N_39842,N_35036,N_36332);
nand U39843 (N_39843,N_36213,N_36350);
nand U39844 (N_39844,N_36372,N_36334);
and U39845 (N_39845,N_36393,N_36444);
or U39846 (N_39846,N_36077,N_36358);
and U39847 (N_39847,N_36158,N_36502);
and U39848 (N_39848,N_36803,N_36604);
nand U39849 (N_39849,N_35706,N_37208);
and U39850 (N_39850,N_36515,N_37109);
or U39851 (N_39851,N_36807,N_35295);
xnor U39852 (N_39852,N_35106,N_37331);
nand U39853 (N_39853,N_37433,N_37002);
xnor U39854 (N_39854,N_36748,N_35245);
or U39855 (N_39855,N_35080,N_35943);
nor U39856 (N_39856,N_35565,N_35456);
nor U39857 (N_39857,N_36140,N_35385);
xor U39858 (N_39858,N_35201,N_36381);
nand U39859 (N_39859,N_35855,N_35395);
xor U39860 (N_39860,N_36926,N_35645);
xor U39861 (N_39861,N_35547,N_35025);
and U39862 (N_39862,N_36502,N_37488);
nand U39863 (N_39863,N_37360,N_35362);
xor U39864 (N_39864,N_36496,N_37296);
nand U39865 (N_39865,N_35502,N_37008);
or U39866 (N_39866,N_37033,N_36319);
and U39867 (N_39867,N_36445,N_36816);
and U39868 (N_39868,N_36820,N_35084);
nor U39869 (N_39869,N_35636,N_35473);
and U39870 (N_39870,N_36362,N_37073);
nand U39871 (N_39871,N_36448,N_37186);
xor U39872 (N_39872,N_35891,N_37422);
and U39873 (N_39873,N_36485,N_37179);
nand U39874 (N_39874,N_37167,N_37031);
nor U39875 (N_39875,N_37070,N_35813);
or U39876 (N_39876,N_36706,N_36926);
nor U39877 (N_39877,N_35180,N_35134);
nand U39878 (N_39878,N_35771,N_36974);
nand U39879 (N_39879,N_35781,N_36485);
or U39880 (N_39880,N_36377,N_36732);
or U39881 (N_39881,N_36210,N_35670);
xnor U39882 (N_39882,N_36592,N_37229);
or U39883 (N_39883,N_36152,N_37210);
or U39884 (N_39884,N_36756,N_35606);
nor U39885 (N_39885,N_35842,N_37054);
nand U39886 (N_39886,N_36879,N_36683);
nand U39887 (N_39887,N_35700,N_37450);
or U39888 (N_39888,N_36902,N_35554);
or U39889 (N_39889,N_37069,N_36334);
nor U39890 (N_39890,N_35740,N_37456);
or U39891 (N_39891,N_36394,N_37271);
nand U39892 (N_39892,N_36686,N_36243);
or U39893 (N_39893,N_36029,N_35175);
and U39894 (N_39894,N_36869,N_36730);
xnor U39895 (N_39895,N_37185,N_37352);
nand U39896 (N_39896,N_36468,N_37044);
and U39897 (N_39897,N_37350,N_35528);
and U39898 (N_39898,N_36370,N_35345);
xnor U39899 (N_39899,N_36083,N_35126);
or U39900 (N_39900,N_35270,N_36414);
nor U39901 (N_39901,N_36287,N_36107);
nand U39902 (N_39902,N_36189,N_35889);
or U39903 (N_39903,N_35929,N_35700);
and U39904 (N_39904,N_37276,N_36501);
or U39905 (N_39905,N_36384,N_36208);
nand U39906 (N_39906,N_35059,N_35828);
or U39907 (N_39907,N_35286,N_36252);
and U39908 (N_39908,N_37338,N_35231);
and U39909 (N_39909,N_37161,N_35836);
nor U39910 (N_39910,N_35938,N_36870);
and U39911 (N_39911,N_36949,N_36065);
nor U39912 (N_39912,N_36132,N_35059);
xor U39913 (N_39913,N_35629,N_35020);
nand U39914 (N_39914,N_37300,N_35900);
and U39915 (N_39915,N_36799,N_37138);
or U39916 (N_39916,N_35428,N_36026);
nand U39917 (N_39917,N_35836,N_37396);
or U39918 (N_39918,N_35074,N_36615);
nand U39919 (N_39919,N_35369,N_36561);
or U39920 (N_39920,N_35858,N_36132);
or U39921 (N_39921,N_36583,N_36981);
and U39922 (N_39922,N_36484,N_37040);
and U39923 (N_39923,N_36755,N_35941);
and U39924 (N_39924,N_35668,N_36670);
nand U39925 (N_39925,N_37245,N_35579);
or U39926 (N_39926,N_35757,N_37132);
and U39927 (N_39927,N_35813,N_35766);
and U39928 (N_39928,N_37180,N_35153);
and U39929 (N_39929,N_36350,N_36485);
xnor U39930 (N_39930,N_35122,N_37465);
nor U39931 (N_39931,N_36316,N_37319);
nor U39932 (N_39932,N_35191,N_36651);
and U39933 (N_39933,N_37024,N_37265);
xor U39934 (N_39934,N_35185,N_36828);
and U39935 (N_39935,N_36899,N_36179);
or U39936 (N_39936,N_37423,N_37213);
and U39937 (N_39937,N_36233,N_35955);
and U39938 (N_39938,N_36277,N_36448);
nand U39939 (N_39939,N_36481,N_36168);
nand U39940 (N_39940,N_37326,N_35968);
nor U39941 (N_39941,N_35811,N_36672);
nand U39942 (N_39942,N_35569,N_36558);
and U39943 (N_39943,N_35621,N_36034);
and U39944 (N_39944,N_35240,N_35471);
or U39945 (N_39945,N_35818,N_37258);
nand U39946 (N_39946,N_36353,N_36937);
nor U39947 (N_39947,N_35526,N_37046);
and U39948 (N_39948,N_36254,N_35993);
nor U39949 (N_39949,N_36478,N_35650);
and U39950 (N_39950,N_36981,N_36059);
nor U39951 (N_39951,N_36874,N_36018);
and U39952 (N_39952,N_35781,N_36134);
and U39953 (N_39953,N_35539,N_37370);
and U39954 (N_39954,N_36851,N_36264);
nor U39955 (N_39955,N_36571,N_35336);
xor U39956 (N_39956,N_36560,N_35150);
and U39957 (N_39957,N_37041,N_37374);
nand U39958 (N_39958,N_35307,N_36799);
xor U39959 (N_39959,N_36020,N_36448);
or U39960 (N_39960,N_37033,N_35007);
or U39961 (N_39961,N_36866,N_37238);
xnor U39962 (N_39962,N_36992,N_36454);
xnor U39963 (N_39963,N_35715,N_35228);
or U39964 (N_39964,N_37134,N_36954);
or U39965 (N_39965,N_37347,N_35385);
xnor U39966 (N_39966,N_36897,N_37196);
xor U39967 (N_39967,N_37107,N_37379);
xor U39968 (N_39968,N_36226,N_36799);
nand U39969 (N_39969,N_36928,N_36878);
nand U39970 (N_39970,N_35076,N_37469);
nand U39971 (N_39971,N_35132,N_37119);
or U39972 (N_39972,N_36738,N_36993);
and U39973 (N_39973,N_36983,N_36914);
nor U39974 (N_39974,N_36742,N_36544);
xor U39975 (N_39975,N_35787,N_36381);
nor U39976 (N_39976,N_35043,N_36290);
nor U39977 (N_39977,N_37488,N_35322);
nand U39978 (N_39978,N_36616,N_37416);
xor U39979 (N_39979,N_35709,N_37277);
or U39980 (N_39980,N_36331,N_35100);
or U39981 (N_39981,N_35259,N_35380);
and U39982 (N_39982,N_36345,N_37370);
or U39983 (N_39983,N_35409,N_37199);
nor U39984 (N_39984,N_35670,N_36857);
or U39985 (N_39985,N_35958,N_35612);
nand U39986 (N_39986,N_35438,N_35477);
nand U39987 (N_39987,N_36435,N_36279);
or U39988 (N_39988,N_36372,N_35976);
nor U39989 (N_39989,N_35856,N_36507);
nand U39990 (N_39990,N_37117,N_36803);
or U39991 (N_39991,N_37318,N_36607);
and U39992 (N_39992,N_36917,N_35206);
xnor U39993 (N_39993,N_36827,N_36217);
nand U39994 (N_39994,N_36793,N_35446);
or U39995 (N_39995,N_36026,N_35333);
or U39996 (N_39996,N_35199,N_37130);
or U39997 (N_39997,N_35265,N_37212);
nand U39998 (N_39998,N_35063,N_35252);
nand U39999 (N_39999,N_37333,N_35679);
and U40000 (N_40000,N_39371,N_39171);
xnor U40001 (N_40001,N_38499,N_39783);
or U40002 (N_40002,N_37696,N_38878);
nand U40003 (N_40003,N_37671,N_39958);
nand U40004 (N_40004,N_39681,N_38573);
nand U40005 (N_40005,N_38233,N_39427);
and U40006 (N_40006,N_39178,N_39538);
xor U40007 (N_40007,N_38191,N_39658);
xor U40008 (N_40008,N_38046,N_39084);
nor U40009 (N_40009,N_38894,N_39484);
xor U40010 (N_40010,N_38348,N_39109);
nand U40011 (N_40011,N_38908,N_39527);
nor U40012 (N_40012,N_38879,N_38565);
and U40013 (N_40013,N_39587,N_39065);
nor U40014 (N_40014,N_37712,N_37779);
or U40015 (N_40015,N_38958,N_38359);
or U40016 (N_40016,N_38783,N_39684);
xnor U40017 (N_40017,N_38396,N_39468);
nor U40018 (N_40018,N_38987,N_39829);
nand U40019 (N_40019,N_37832,N_38409);
or U40020 (N_40020,N_39889,N_37957);
nor U40021 (N_40021,N_37670,N_39475);
nand U40022 (N_40022,N_39387,N_37730);
nand U40023 (N_40023,N_37871,N_39888);
and U40024 (N_40024,N_38655,N_39942);
xor U40025 (N_40025,N_39792,N_39754);
xnor U40026 (N_40026,N_38229,N_39214);
or U40027 (N_40027,N_39460,N_37778);
nor U40028 (N_40028,N_38781,N_39983);
and U40029 (N_40029,N_38403,N_39859);
xnor U40030 (N_40030,N_39014,N_39010);
or U40031 (N_40031,N_37714,N_37589);
and U40032 (N_40032,N_38757,N_39169);
or U40033 (N_40033,N_37815,N_38373);
xor U40034 (N_40034,N_38462,N_37812);
and U40035 (N_40035,N_39858,N_39261);
nor U40036 (N_40036,N_37943,N_37662);
nor U40037 (N_40037,N_38004,N_39221);
nor U40038 (N_40038,N_38181,N_39087);
nand U40039 (N_40039,N_38684,N_38604);
nor U40040 (N_40040,N_38401,N_37822);
or U40041 (N_40041,N_37993,N_39588);
xor U40042 (N_40042,N_39059,N_39631);
nor U40043 (N_40043,N_39762,N_38135);
nand U40044 (N_40044,N_37776,N_39710);
or U40045 (N_40045,N_39630,N_39943);
nand U40046 (N_40046,N_38612,N_37583);
or U40047 (N_40047,N_39477,N_39976);
nor U40048 (N_40048,N_39691,N_39993);
nand U40049 (N_40049,N_37699,N_37795);
or U40050 (N_40050,N_38389,N_39434);
and U40051 (N_40051,N_39713,N_38753);
or U40052 (N_40052,N_39351,N_39112);
or U40053 (N_40053,N_38444,N_38982);
xnor U40054 (N_40054,N_38569,N_38416);
nand U40055 (N_40055,N_37571,N_38308);
nand U40056 (N_40056,N_39992,N_39760);
or U40057 (N_40057,N_38095,N_39313);
and U40058 (N_40058,N_37676,N_37992);
nand U40059 (N_40059,N_37572,N_38548);
nor U40060 (N_40060,N_39865,N_37614);
nor U40061 (N_40061,N_37680,N_38797);
xor U40062 (N_40062,N_38697,N_39137);
or U40063 (N_40063,N_37690,N_38588);
and U40064 (N_40064,N_39503,N_38031);
or U40065 (N_40065,N_37538,N_38966);
nand U40066 (N_40066,N_39322,N_37843);
and U40067 (N_40067,N_39046,N_39105);
xnor U40068 (N_40068,N_38848,N_38353);
or U40069 (N_40069,N_39330,N_37539);
nand U40070 (N_40070,N_37942,N_39800);
or U40071 (N_40071,N_39959,N_38550);
nor U40072 (N_40072,N_38645,N_38463);
nand U40073 (N_40073,N_38841,N_38286);
nand U40074 (N_40074,N_39396,N_38405);
and U40075 (N_40075,N_39148,N_39608);
nor U40076 (N_40076,N_39664,N_39880);
and U40077 (N_40077,N_38429,N_39439);
and U40078 (N_40078,N_39676,N_38376);
or U40079 (N_40079,N_39197,N_39416);
nor U40080 (N_40080,N_39817,N_37526);
and U40081 (N_40081,N_38424,N_38358);
nand U40082 (N_40082,N_38025,N_39055);
nor U40083 (N_40083,N_39687,N_39256);
nand U40084 (N_40084,N_39181,N_39293);
and U40085 (N_40085,N_38452,N_39053);
and U40086 (N_40086,N_37711,N_38541);
xor U40087 (N_40087,N_38754,N_39209);
nor U40088 (N_40088,N_38602,N_38108);
or U40089 (N_40089,N_39575,N_37541);
nand U40090 (N_40090,N_39867,N_39671);
or U40091 (N_40091,N_39906,N_39541);
or U40092 (N_40092,N_39271,N_39624);
nand U40093 (N_40093,N_37665,N_39894);
xor U40094 (N_40094,N_38702,N_39830);
nand U40095 (N_40095,N_37978,N_37713);
or U40096 (N_40096,N_39868,N_38070);
xnor U40097 (N_40097,N_37753,N_37727);
and U40098 (N_40098,N_39043,N_39781);
and U40099 (N_40099,N_37648,N_38110);
nor U40100 (N_40100,N_38605,N_38498);
or U40101 (N_40101,N_39599,N_38460);
xor U40102 (N_40102,N_39950,N_39977);
nor U40103 (N_40103,N_38009,N_38137);
or U40104 (N_40104,N_38941,N_38384);
nand U40105 (N_40105,N_39998,N_39405);
nand U40106 (N_40106,N_39196,N_38562);
or U40107 (N_40107,N_37846,N_38397);
or U40108 (N_40108,N_38053,N_38242);
nand U40109 (N_40109,N_39091,N_37724);
nor U40110 (N_40110,N_38810,N_39714);
nand U40111 (N_40111,N_38954,N_39431);
nand U40112 (N_40112,N_38472,N_37792);
nor U40113 (N_40113,N_38622,N_37827);
or U40114 (N_40114,N_39081,N_39450);
nand U40115 (N_40115,N_38129,N_39912);
and U40116 (N_40116,N_38974,N_37718);
or U40117 (N_40117,N_39544,N_39827);
or U40118 (N_40118,N_39886,N_37944);
and U40119 (N_40119,N_37950,N_38372);
and U40120 (N_40120,N_38903,N_38620);
or U40121 (N_40121,N_38634,N_39839);
nand U40122 (N_40122,N_37903,N_39025);
or U40123 (N_40123,N_37899,N_39884);
and U40124 (N_40124,N_38625,N_39307);
nand U40125 (N_40125,N_37577,N_38496);
nor U40126 (N_40126,N_39097,N_39455);
and U40127 (N_40127,N_37986,N_38193);
and U40128 (N_40128,N_38784,N_39409);
xor U40129 (N_40129,N_38259,N_39147);
and U40130 (N_40130,N_37601,N_38709);
nor U40131 (N_40131,N_39142,N_38114);
xnor U40132 (N_40132,N_39364,N_37698);
xor U40133 (N_40133,N_37945,N_37655);
nand U40134 (N_40134,N_37856,N_39502);
nand U40135 (N_40135,N_39806,N_38207);
or U40136 (N_40136,N_38212,N_38247);
and U40137 (N_40137,N_38189,N_38935);
and U40138 (N_40138,N_38663,N_38329);
or U40139 (N_40139,N_39339,N_37606);
and U40140 (N_40140,N_39188,N_38050);
and U40141 (N_40141,N_39149,N_38079);
nor U40142 (N_40142,N_38724,N_39238);
nor U40143 (N_40143,N_37552,N_39236);
nor U40144 (N_40144,N_37576,N_39936);
xor U40145 (N_40145,N_39838,N_38598);
xor U40146 (N_40146,N_39642,N_38426);
or U40147 (N_40147,N_39410,N_38431);
nand U40148 (N_40148,N_38607,N_39465);
and U40149 (N_40149,N_37729,N_38725);
and U40150 (N_40150,N_38327,N_37531);
or U40151 (N_40151,N_38458,N_38186);
nor U40152 (N_40152,N_39385,N_38871);
xnor U40153 (N_40153,N_39769,N_39433);
and U40154 (N_40154,N_38280,N_39739);
nand U40155 (N_40155,N_37567,N_39733);
xor U40156 (N_40156,N_38807,N_39015);
xor U40157 (N_40157,N_39907,N_39116);
nand U40158 (N_40158,N_37656,N_39517);
nand U40159 (N_40159,N_37635,N_38309);
and U40160 (N_40160,N_38703,N_38323);
xor U40161 (N_40161,N_39489,N_38410);
and U40162 (N_40162,N_39776,N_38494);
xor U40163 (N_40163,N_38872,N_39359);
or U40164 (N_40164,N_37824,N_37609);
or U40165 (N_40165,N_38098,N_39741);
and U40166 (N_40166,N_39613,N_37761);
or U40167 (N_40167,N_37592,N_39951);
nor U40168 (N_40168,N_37633,N_37748);
xor U40169 (N_40169,N_39117,N_39301);
nand U40170 (N_40170,N_38707,N_38819);
nor U40171 (N_40171,N_38511,N_39303);
nor U40172 (N_40172,N_39625,N_39216);
nand U40173 (N_40173,N_37514,N_38084);
nor U40174 (N_40174,N_39798,N_38934);
and U40175 (N_40175,N_39737,N_38537);
nor U40176 (N_40176,N_38271,N_39092);
or U40177 (N_40177,N_38115,N_38970);
xnor U40178 (N_40178,N_38613,N_39047);
nor U40179 (N_40179,N_38255,N_38282);
and U40180 (N_40180,N_38912,N_37627);
or U40181 (N_40181,N_39824,N_37762);
and U40182 (N_40182,N_38322,N_38669);
or U40183 (N_40183,N_37743,N_37508);
xor U40184 (N_40184,N_39758,N_38930);
nor U40185 (N_40185,N_38274,N_39444);
xor U40186 (N_40186,N_38777,N_38172);
xnor U40187 (N_40187,N_39241,N_39481);
nand U40188 (N_40188,N_38928,N_38469);
or U40189 (N_40189,N_39571,N_38342);
nor U40190 (N_40190,N_39278,N_37891);
nor U40191 (N_40191,N_39164,N_38619);
nor U40192 (N_40192,N_37869,N_37533);
and U40193 (N_40193,N_39296,N_39660);
nor U40194 (N_40194,N_38354,N_39374);
nor U40195 (N_40195,N_38069,N_38347);
nand U40196 (N_40196,N_37784,N_39856);
and U40197 (N_40197,N_37506,N_38853);
nand U40198 (N_40198,N_38262,N_37968);
or U40199 (N_40199,N_38532,N_37740);
and U40200 (N_40200,N_39060,N_38759);
xor U40201 (N_40201,N_39228,N_39677);
nand U40202 (N_40202,N_38951,N_39258);
and U40203 (N_40203,N_38026,N_37825);
xnor U40204 (N_40204,N_38988,N_37930);
nor U40205 (N_40205,N_37675,N_38226);
xor U40206 (N_40206,N_38836,N_38385);
nor U40207 (N_40207,N_39380,N_37878);
or U40208 (N_40208,N_38720,N_38874);
and U40209 (N_40209,N_38546,N_38977);
xnor U40210 (N_40210,N_38307,N_38438);
or U40211 (N_40211,N_38028,N_39008);
and U40212 (N_40212,N_38060,N_39213);
or U40213 (N_40213,N_39414,N_38782);
and U40214 (N_40214,N_38592,N_38746);
or U40215 (N_40215,N_38361,N_38177);
nand U40216 (N_40216,N_39350,N_39659);
or U40217 (N_40217,N_37616,N_38545);
xnor U40218 (N_40218,N_39173,N_38317);
or U40219 (N_40219,N_39735,N_38006);
xor U40220 (N_40220,N_39666,N_38459);
and U40221 (N_40221,N_39392,N_37587);
or U40222 (N_40222,N_37672,N_37604);
nor U40223 (N_40223,N_38464,N_39198);
and U40224 (N_40224,N_39230,N_39694);
and U40225 (N_40225,N_37769,N_39985);
or U40226 (N_40226,N_39842,N_39143);
and U40227 (N_40227,N_38497,N_38632);
xnor U40228 (N_40228,N_39127,N_38370);
and U40229 (N_40229,N_37892,N_37782);
nand U40230 (N_40230,N_38117,N_38611);
nand U40231 (N_40231,N_38556,N_38804);
nand U40232 (N_40232,N_39500,N_37537);
nand U40233 (N_40233,N_39609,N_39832);
xnor U40234 (N_40234,N_39021,N_39504);
nand U40235 (N_40235,N_38980,N_38743);
or U40236 (N_40236,N_37852,N_39333);
or U40237 (N_40237,N_39354,N_39882);
nand U40238 (N_40238,N_39336,N_39962);
and U40239 (N_40239,N_38440,N_39550);
or U40240 (N_40240,N_38363,N_39222);
or U40241 (N_40241,N_38895,N_37980);
xnor U40242 (N_40242,N_38811,N_38456);
xor U40243 (N_40243,N_38946,N_38378);
nand U40244 (N_40244,N_39342,N_39376);
nand U40245 (N_40245,N_39534,N_39501);
xor U40246 (N_40246,N_38855,N_37835);
nand U40247 (N_40247,N_39286,N_39125);
xnor U40248 (N_40248,N_39218,N_37598);
xnor U40249 (N_40249,N_38767,N_38633);
or U40250 (N_40250,N_39123,N_39509);
and U40251 (N_40251,N_38981,N_37688);
xnor U40252 (N_40252,N_38395,N_37553);
xnor U40253 (N_40253,N_38953,N_39411);
or U40254 (N_40254,N_39399,N_38577);
nand U40255 (N_40255,N_37826,N_39761);
nor U40256 (N_40256,N_37544,N_39352);
or U40257 (N_40257,N_37600,N_38715);
or U40258 (N_40258,N_39203,N_39182);
and U40259 (N_40259,N_38517,N_39417);
and U40260 (N_40260,N_37912,N_37591);
nor U40261 (N_40261,N_39172,N_38963);
xnor U40262 (N_40262,N_37501,N_37739);
nor U40263 (N_40263,N_39548,N_37535);
xnor U40264 (N_40264,N_38995,N_39346);
nand U40265 (N_40265,N_39662,N_38744);
xnor U40266 (N_40266,N_38300,N_38507);
and U40267 (N_40267,N_37750,N_39855);
or U40268 (N_40268,N_38333,N_37645);
xnor U40269 (N_40269,N_39802,N_38735);
nor U40270 (N_40270,N_38991,N_37906);
nor U40271 (N_40271,N_38106,N_39833);
and U40272 (N_40272,N_37954,N_38586);
nor U40273 (N_40273,N_38869,N_38552);
xor U40274 (N_40274,N_39646,N_37654);
nor U40275 (N_40275,N_37678,N_37908);
or U40276 (N_40276,N_38814,N_37643);
xor U40277 (N_40277,N_38943,N_37578);
nor U40278 (N_40278,N_38156,N_37580);
and U40279 (N_40279,N_39554,N_38480);
nor U40280 (N_40280,N_37517,N_39004);
or U40281 (N_40281,N_37709,N_38474);
or U40282 (N_40282,N_39701,N_37594);
nand U40283 (N_40283,N_39030,N_37816);
or U40284 (N_40284,N_39239,N_38430);
nor U40285 (N_40285,N_37859,N_38606);
xor U40286 (N_40286,N_37525,N_39140);
and U40287 (N_40287,N_37518,N_38231);
or U40288 (N_40288,N_38829,N_39177);
and U40289 (N_40289,N_39639,N_39215);
nor U40290 (N_40290,N_39315,N_37926);
nand U40291 (N_40291,N_39299,N_38230);
xnor U40292 (N_40292,N_38194,N_37702);
or U40293 (N_40293,N_39133,N_39514);
nor U40294 (N_40294,N_39184,N_39996);
nand U40295 (N_40295,N_37689,N_39837);
nor U40296 (N_40296,N_38876,N_38867);
nand U40297 (N_40297,N_39049,N_37962);
or U40298 (N_40298,N_38017,N_38983);
nor U40299 (N_40299,N_39029,N_39873);
or U40300 (N_40300,N_37925,N_38325);
nand U40301 (N_40301,N_37998,N_39079);
or U40302 (N_40302,N_37911,N_39668);
xnor U40303 (N_40303,N_37624,N_37575);
and U40304 (N_40304,N_38332,N_39745);
or U40305 (N_40305,N_39864,N_37660);
nor U40306 (N_40306,N_38791,N_39821);
xnor U40307 (N_40307,N_37854,N_37934);
or U40308 (N_40308,N_38644,N_38523);
xnor U40309 (N_40309,N_37733,N_37877);
and U40310 (N_40310,N_39227,N_39327);
nor U40311 (N_40311,N_39765,N_38938);
or U40312 (N_40312,N_39893,N_39237);
and U40313 (N_40313,N_39045,N_39887);
nor U40314 (N_40314,N_37639,N_38778);
nand U40315 (N_40315,N_37540,N_38649);
or U40316 (N_40316,N_39488,N_37651);
xor U40317 (N_40317,N_37982,N_39853);
and U40318 (N_40318,N_38176,N_38614);
or U40319 (N_40319,N_38630,N_38399);
or U40320 (N_40320,N_38875,N_38412);
and U40321 (N_40321,N_38553,N_38790);
nor U40322 (N_40322,N_39064,N_38445);
or U40323 (N_40323,N_38989,N_38432);
xnor U40324 (N_40324,N_38057,N_37707);
and U40325 (N_40325,N_37500,N_39332);
xnor U40326 (N_40326,N_38926,N_38400);
nor U40327 (N_40327,N_37933,N_37811);
nand U40328 (N_40328,N_39009,N_39193);
and U40329 (N_40329,N_39077,N_38566);
nor U40330 (N_40330,N_39102,N_37565);
xnor U40331 (N_40331,N_37916,N_38145);
nand U40332 (N_40332,N_39418,N_39695);
nand U40333 (N_40333,N_38243,N_37728);
nor U40334 (N_40334,N_38727,N_37617);
nor U40335 (N_40335,N_39016,N_37631);
xnor U40336 (N_40336,N_38221,N_38011);
nand U40337 (N_40337,N_38138,N_38623);
and U40338 (N_40338,N_39018,N_38199);
or U40339 (N_40339,N_39712,N_38330);
and U40340 (N_40340,N_38123,N_38774);
and U40341 (N_40341,N_38683,N_38688);
xnor U40342 (N_40342,N_38020,N_39778);
or U40343 (N_40343,N_39020,N_38232);
and U40344 (N_40344,N_37967,N_39369);
nand U40345 (N_40345,N_39643,N_39426);
and U40346 (N_40346,N_38419,N_39814);
xor U40347 (N_40347,N_38341,N_37649);
or U40348 (N_40348,N_39686,N_38955);
or U40349 (N_40349,N_38275,N_39306);
and U40350 (N_40350,N_37788,N_38408);
nand U40351 (N_40351,N_38040,N_39185);
nand U40352 (N_40352,N_38650,N_38719);
nand U40353 (N_40353,N_39999,N_39076);
xnor U40354 (N_40354,N_38956,N_39933);
nand U40355 (N_40355,N_38847,N_39437);
xor U40356 (N_40356,N_38336,N_39101);
xnor U40357 (N_40357,N_38473,N_38487);
xor U40358 (N_40358,N_38415,N_37994);
nand U40359 (N_40359,N_37701,N_37973);
or U40360 (N_40360,N_38937,N_39809);
or U40361 (N_40361,N_39606,N_38491);
or U40362 (N_40362,N_39982,N_39131);
xor U40363 (N_40363,N_39786,N_38215);
and U40364 (N_40364,N_37807,N_37618);
nor U40365 (N_40365,N_39493,N_39566);
and U40366 (N_40366,N_39152,N_39577);
and U40367 (N_40367,N_38014,N_39471);
nand U40368 (N_40368,N_38292,N_38418);
and U40369 (N_40369,N_38269,N_39860);
nand U40370 (N_40370,N_38975,N_39905);
nor U40371 (N_40371,N_37747,N_37974);
xor U40372 (N_40372,N_37918,N_39304);
nor U40373 (N_40373,N_39129,N_38466);
xor U40374 (N_40374,N_39083,N_38568);
nand U40375 (N_40375,N_39082,N_39452);
nand U40376 (N_40376,N_38856,N_37513);
or U40377 (N_40377,N_38706,N_39875);
xnor U40378 (N_40378,N_38299,N_38326);
nor U40379 (N_40379,N_37855,N_39913);
and U40380 (N_40380,N_37521,N_38152);
and U40381 (N_40381,N_38978,N_38227);
nor U40382 (N_40382,N_39300,N_39357);
nor U40383 (N_40383,N_38411,N_39024);
nand U40384 (N_40384,N_38355,N_39485);
or U40385 (N_40385,N_39779,N_38792);
nand U40386 (N_40386,N_38224,N_39526);
or U40387 (N_40387,N_38572,N_39945);
and U40388 (N_40388,N_37612,N_37751);
nor U40389 (N_40389,N_39528,N_39520);
xor U40390 (N_40390,N_38173,N_38167);
and U40391 (N_40391,N_38640,N_37781);
nor U40392 (N_40392,N_38621,N_39805);
or U40393 (N_40393,N_39547,N_39965);
xor U40394 (N_40394,N_39590,N_37504);
or U40395 (N_40395,N_38865,N_39498);
and U40396 (N_40396,N_37677,N_39954);
or U40397 (N_40397,N_38443,N_39449);
or U40398 (N_40398,N_37817,N_39916);
xnor U40399 (N_40399,N_37597,N_39629);
xnor U40400 (N_40400,N_38171,N_39784);
xnor U40401 (N_40401,N_38428,N_38099);
and U40402 (N_40402,N_38515,N_38001);
nand U40403 (N_40403,N_39289,N_37708);
nand U40404 (N_40404,N_38478,N_38997);
nand U40405 (N_40405,N_39665,N_39720);
xnor U40406 (N_40406,N_39937,N_38843);
nand U40407 (N_40407,N_38732,N_39326);
xor U40408 (N_40408,N_39755,N_38404);
nand U40409 (N_40409,N_37808,N_38907);
and U40410 (N_40410,N_38627,N_39930);
nand U40411 (N_40411,N_39287,N_39007);
xnor U40412 (N_40412,N_37622,N_39106);
xor U40413 (N_40413,N_39986,N_37510);
or U40414 (N_40414,N_38256,N_39707);
nand U40415 (N_40415,N_38858,N_38506);
xor U40416 (N_40416,N_38092,N_39750);
or U40417 (N_40417,N_39494,N_38039);
nand U40418 (N_40418,N_37684,N_38745);
nor U40419 (N_40419,N_38390,N_39787);
or U40420 (N_40420,N_39974,N_39028);
nor U40421 (N_40421,N_39206,N_38624);
nand U40422 (N_40422,N_38860,N_38344);
nor U40423 (N_40423,N_38125,N_37610);
or U40424 (N_40424,N_39308,N_38866);
xor U40425 (N_40425,N_37981,N_39562);
and U40426 (N_40426,N_39233,N_38524);
nor U40427 (N_40427,N_39358,N_37902);
nand U40428 (N_40428,N_39274,N_37704);
xnor U40429 (N_40429,N_39978,N_38514);
or U40430 (N_40430,N_37754,N_39461);
xnor U40431 (N_40431,N_37686,N_38136);
nor U40432 (N_40432,N_38334,N_38180);
and U40433 (N_40433,N_39096,N_37797);
xor U40434 (N_40434,N_39641,N_38849);
xnor U40435 (N_40435,N_37574,N_39220);
nand U40436 (N_40436,N_39085,N_38128);
nor U40437 (N_40437,N_39229,N_39251);
nor U40438 (N_40438,N_37775,N_37715);
and U40439 (N_40439,N_38162,N_38512);
nor U40440 (N_40440,N_37885,N_37806);
xnor U40441 (N_40441,N_39584,N_37872);
nand U40442 (N_40442,N_38818,N_38488);
nand U40443 (N_40443,N_39531,N_38100);
xnor U40444 (N_40444,N_38468,N_38713);
nand U40445 (N_40445,N_38339,N_38187);
nor U40446 (N_40446,N_39726,N_38711);
nor U40447 (N_40447,N_38324,N_39108);
or U40448 (N_40448,N_38113,N_39738);
nand U40449 (N_40449,N_38251,N_39883);
xor U40450 (N_40450,N_37849,N_39770);
nor U40451 (N_40451,N_38648,N_39589);
nor U40452 (N_40452,N_37726,N_39661);
nand U40453 (N_40453,N_39801,N_38660);
and U40454 (N_40454,N_38490,N_37858);
or U40455 (N_40455,N_39003,N_39089);
and U40456 (N_40456,N_39924,N_39199);
or U40457 (N_40457,N_39309,N_39176);
or U40458 (N_40458,N_37963,N_39652);
xnor U40459 (N_40459,N_38345,N_39247);
or U40460 (N_40460,N_39580,N_39277);
and U40461 (N_40461,N_38661,N_39161);
nor U40462 (N_40462,N_38758,N_39623);
nand U40463 (N_40463,N_38112,N_38285);
nor U40464 (N_40464,N_39191,N_39902);
nand U40465 (N_40465,N_37758,N_38571);
xor U40466 (N_40466,N_39632,N_39777);
or U40467 (N_40467,N_37886,N_39647);
and U40468 (N_40468,N_39255,N_38880);
xnor U40469 (N_40469,N_37995,N_38318);
nor U40470 (N_40470,N_38809,N_38842);
nor U40471 (N_40471,N_38971,N_39276);
and U40472 (N_40472,N_39675,N_39412);
or U40473 (N_40473,N_38658,N_38673);
or U40474 (N_40474,N_39651,N_39885);
and U40475 (N_40475,N_39944,N_39457);
or U40476 (N_40476,N_38529,N_39482);
and U40477 (N_40477,N_38337,N_39808);
and U40478 (N_40478,N_37771,N_38107);
nand U40479 (N_40479,N_38425,N_38219);
or U40480 (N_40480,N_38626,N_39037);
nand U40481 (N_40481,N_37697,N_38522);
xnor U40482 (N_40482,N_38051,N_39403);
and U40483 (N_40483,N_37809,N_39719);
and U40484 (N_40484,N_39680,N_39058);
or U40485 (N_40485,N_39698,N_38044);
nor U40486 (N_40486,N_38768,N_38824);
or U40487 (N_40487,N_38222,N_37890);
nor U40488 (N_40488,N_39640,N_39861);
nor U40489 (N_40489,N_38610,N_38617);
nor U40490 (N_40490,N_38766,N_37971);
or U40491 (N_40491,N_37532,N_39280);
nand U40492 (N_40492,N_38451,N_39929);
or U40493 (N_40493,N_39568,N_38615);
or U40494 (N_40494,N_37783,N_38276);
xnor U40495 (N_40495,N_37935,N_38760);
xor U40496 (N_40496,N_38692,N_39622);
xor U40497 (N_40497,N_38685,N_38901);
nor U40498 (N_40498,N_39166,N_38862);
and U40499 (N_40499,N_39711,N_37904);
nor U40500 (N_40500,N_38067,N_38969);
or U40501 (N_40501,N_39790,N_38296);
nand U40502 (N_40502,N_39476,N_39967);
nand U40503 (N_40503,N_38816,N_38539);
nor U40504 (N_40504,N_38197,N_37984);
nor U40505 (N_40505,N_39159,N_37907);
nor U40506 (N_40506,N_38513,N_38560);
nor U40507 (N_40507,N_39190,N_38839);
and U40508 (N_40508,N_39932,N_39334);
nor U40509 (N_40509,N_39969,N_37522);
xnor U40510 (N_40510,N_38942,N_39732);
nor U40511 (N_40511,N_39495,N_38749);
and U40512 (N_40512,N_39552,N_38543);
nand U40513 (N_40513,N_37634,N_39682);
and U40514 (N_40514,N_37620,N_38833);
and U40515 (N_40515,N_39766,N_39212);
xor U40516 (N_40516,N_37932,N_37985);
nor U40517 (N_40517,N_39920,N_39406);
nand U40518 (N_40518,N_39649,N_37595);
xor U40519 (N_40519,N_39845,N_38303);
and U40520 (N_40520,N_39823,N_38973);
xor U40521 (N_40521,N_37928,N_39282);
or U40522 (N_40522,N_38435,N_37650);
nand U40523 (N_40523,N_38712,N_38896);
and U40524 (N_40524,N_39540,N_37519);
nand U40525 (N_40525,N_39253,N_37823);
or U40526 (N_40526,N_38482,N_38321);
nand U40527 (N_40527,N_39593,N_38558);
xor U40528 (N_40528,N_39508,N_37923);
xor U40529 (N_40529,N_37719,N_38087);
nor U40530 (N_40530,N_39492,N_37529);
and U40531 (N_40531,N_37608,N_39210);
or U40532 (N_40532,N_37641,N_38828);
xnor U40533 (N_40533,N_38787,N_39831);
or U40534 (N_40534,N_37874,N_39960);
and U40535 (N_40535,N_39725,N_37927);
nor U40536 (N_40536,N_38141,N_38518);
nand U40537 (N_40537,N_39565,N_38146);
nand U40538 (N_40538,N_38691,N_38369);
or U40539 (N_40539,N_39926,N_38651);
nand U40540 (N_40540,N_37770,N_38155);
nor U40541 (N_40541,N_37922,N_38892);
nand U40542 (N_40542,N_37920,N_37759);
xnor U40543 (N_40543,N_39252,N_38055);
nor U40544 (N_40544,N_37585,N_37948);
xnor U40545 (N_40545,N_38105,N_39567);
nand U40546 (N_40546,N_38904,N_38889);
and U40547 (N_40547,N_39470,N_38350);
and U40548 (N_40548,N_38950,N_39231);
nor U40549 (N_40549,N_38398,N_38631);
and U40550 (N_40550,N_39355,N_38639);
or U40551 (N_40551,N_37611,N_39871);
and U40552 (N_40552,N_39219,N_38030);
xor U40553 (N_40553,N_38439,N_38019);
xor U40554 (N_40554,N_38674,N_37851);
nand U40555 (N_40555,N_39098,N_38433);
and U40556 (N_40556,N_38080,N_38047);
nor U40557 (N_40557,N_37693,N_39056);
nor U40558 (N_40558,N_38885,N_38593);
xnor U40559 (N_40559,N_38290,N_38228);
or U40560 (N_40560,N_38423,N_39442);
nor U40561 (N_40561,N_39595,N_37768);
nor U40562 (N_40562,N_38825,N_38690);
or U40563 (N_40563,N_38582,N_37710);
or U40564 (N_40564,N_38096,N_38919);
nand U40565 (N_40565,N_39292,N_39348);
xnor U40566 (N_40566,N_38748,N_38945);
and U40567 (N_40567,N_38461,N_38179);
nand U40568 (N_40568,N_38504,N_39126);
nand U40569 (N_40569,N_39591,N_39408);
xor U40570 (N_40570,N_39249,N_39722);
nor U40571 (N_40571,N_39425,N_38089);
nand U40572 (N_40572,N_38281,N_39421);
or U40573 (N_40573,N_39654,N_38591);
xor U40574 (N_40574,N_38881,N_38609);
and U40575 (N_40575,N_38716,N_38131);
nor U40576 (N_40576,N_37850,N_37683);
nor U40577 (N_40577,N_37725,N_38150);
nor U40578 (N_40578,N_39748,N_38122);
or U40579 (N_40579,N_39626,N_39044);
or U40580 (N_40580,N_39272,N_38705);
and U40581 (N_40581,N_39088,N_38704);
nor U40582 (N_40582,N_38457,N_39035);
or U40583 (N_40583,N_38003,N_38195);
nor U40584 (N_40584,N_39389,N_39156);
or U40585 (N_40585,N_38815,N_38618);
nor U40586 (N_40586,N_39440,N_39851);
and U40587 (N_40587,N_39435,N_39979);
or U40588 (N_40588,N_38086,N_39094);
and U40589 (N_40589,N_39155,N_39539);
nor U40590 (N_40590,N_39909,N_39794);
or U40591 (N_40591,N_38984,N_39115);
xor U40592 (N_40592,N_38252,N_39645);
and U40593 (N_40593,N_39242,N_38600);
or U40594 (N_40594,N_38273,N_39834);
nand U40595 (N_40595,N_39195,N_37734);
nand U40596 (N_40596,N_39795,N_38148);
nand U40597 (N_40597,N_38994,N_38202);
or U40598 (N_40598,N_38812,N_38267);
and U40599 (N_40599,N_39715,N_38111);
and U40600 (N_40600,N_39650,N_38023);
nor U40601 (N_40601,N_38139,N_38883);
and U40602 (N_40602,N_37602,N_38575);
or U40603 (N_40603,N_39343,N_37774);
xor U40604 (N_40604,N_39167,N_39881);
and U40605 (N_40605,N_37663,N_38035);
nor U40606 (N_40606,N_38864,N_39483);
and U40607 (N_40607,N_39914,N_39100);
xnor U40608 (N_40608,N_37559,N_39621);
nor U40609 (N_40609,N_38010,N_37528);
xnor U40610 (N_40610,N_38338,N_38542);
or U40611 (N_40611,N_38346,N_37703);
nor U40612 (N_40612,N_39507,N_37801);
xnor U40613 (N_40613,N_38312,N_38751);
xor U40614 (N_40614,N_38218,N_37556);
xnor U40615 (N_40615,N_37560,N_39697);
and U40616 (N_40616,N_39729,N_39878);
nor U40617 (N_40617,N_38489,N_39145);
nand U40618 (N_40618,N_38449,N_39573);
nor U40619 (N_40619,N_38701,N_38434);
nor U40620 (N_40620,N_37563,N_37605);
xnor U40621 (N_40621,N_39636,N_38109);
nor U40622 (N_40622,N_37901,N_37584);
nor U40623 (N_40623,N_39061,N_39451);
and U40624 (N_40624,N_38349,N_38185);
xor U40625 (N_40625,N_37630,N_39857);
and U40626 (N_40626,N_38121,N_39519);
and U40627 (N_40627,N_38447,N_38007);
and U40628 (N_40628,N_39723,N_39793);
and U40629 (N_40629,N_38154,N_38379);
and U40630 (N_40630,N_38104,N_39305);
and U40631 (N_40631,N_39560,N_39316);
xor U40632 (N_40632,N_39898,N_38520);
or U40633 (N_40633,N_37837,N_38929);
nand U40634 (N_40634,N_39340,N_38196);
or U40635 (N_40635,N_37969,N_39335);
and U40636 (N_40636,N_38840,N_38940);
nor U40637 (N_40637,N_37955,N_38964);
xor U40638 (N_40638,N_39260,N_38258);
nor U40639 (N_40639,N_38157,N_39223);
xnor U40640 (N_40640,N_38999,N_38647);
xor U40641 (N_40641,N_37561,N_39491);
xnor U40642 (N_40642,N_38266,N_39699);
nor U40643 (N_40643,N_37732,N_38140);
nand U40644 (N_40644,N_39708,N_37821);
xor U40645 (N_40645,N_38068,N_37936);
xor U40646 (N_40646,N_38960,N_38278);
or U40647 (N_40647,N_38846,N_38679);
nand U40648 (N_40648,N_38454,N_39653);
and U40649 (N_40649,N_38143,N_38959);
nand U40650 (N_40650,N_39522,N_38579);
and U40651 (N_40651,N_39964,N_39578);
nor U40652 (N_40652,N_39592,N_37786);
xnor U40653 (N_40653,N_39456,N_39462);
or U40654 (N_40654,N_39525,N_37810);
and U40655 (N_40655,N_39822,N_37542);
or U40656 (N_40656,N_39192,N_37705);
xor U40657 (N_40657,N_38158,N_39939);
nor U40658 (N_40658,N_38311,N_39702);
and U40659 (N_40659,N_38225,N_37642);
nor U40660 (N_40660,N_39521,N_39187);
nor U40661 (N_40661,N_38124,N_39611);
xor U40662 (N_40662,N_37880,N_38165);
or U40663 (N_40663,N_39103,N_39154);
xor U40664 (N_40664,N_39496,N_39120);
nand U40665 (N_40665,N_38775,N_39536);
nor U40666 (N_40666,N_39331,N_39782);
nor U40667 (N_40667,N_37813,N_39122);
nor U40668 (N_40668,N_38831,N_37638);
nor U40669 (N_40669,N_38772,N_39689);
nor U40670 (N_40670,N_39583,N_38750);
and U40671 (N_40671,N_38944,N_38913);
xor U40672 (N_40672,N_38694,N_38603);
nand U40673 (N_40673,N_39397,N_38240);
xnor U40674 (N_40674,N_39367,N_37549);
xnor U40675 (N_40675,N_37804,N_39789);
or U40676 (N_40676,N_39850,N_39872);
or U40677 (N_40677,N_38897,N_39341);
xnor U40678 (N_40678,N_38638,N_37744);
nand U40679 (N_40679,N_39717,N_38304);
or U40680 (N_40680,N_37887,N_38223);
nand U40681 (N_40681,N_39511,N_38799);
and U40682 (N_40682,N_38914,N_39533);
or U40683 (N_40683,N_37668,N_39516);
and U40684 (N_40684,N_39052,N_38305);
nor U40685 (N_40685,N_38120,N_38301);
or U40686 (N_40686,N_38533,N_38058);
nand U40687 (N_40687,N_39048,N_37599);
or U40688 (N_40688,N_39078,N_37905);
or U40689 (N_40689,N_39270,N_38710);
nor U40690 (N_40690,N_38295,N_38320);
nand U40691 (N_40691,N_38576,N_38470);
and U40692 (N_40692,N_38391,N_37796);
nor U40693 (N_40693,N_37863,N_38239);
or U40694 (N_40694,N_38134,N_39840);
xnor U40695 (N_40695,N_38298,N_39338);
or U40696 (N_40696,N_38877,N_38924);
and U40697 (N_40697,N_39057,N_38737);
or U40698 (N_40698,N_37745,N_38077);
or U40699 (N_40699,N_38728,N_38594);
nor U40700 (N_40700,N_38236,N_38779);
nand U40701 (N_40701,N_39585,N_38823);
and U40702 (N_40702,N_39935,N_39107);
nor U40703 (N_40703,N_38527,N_39811);
xnor U40704 (N_40704,N_39438,N_39721);
or U40705 (N_40705,N_38061,N_39564);
nand U40706 (N_40706,N_39803,N_38931);
xor U40707 (N_40707,N_39413,N_39011);
xnor U40708 (N_40708,N_39532,N_38835);
nand U40709 (N_40709,N_37946,N_39153);
and U40710 (N_40710,N_38448,N_37937);
or U40711 (N_40711,N_38268,N_39602);
and U40712 (N_40712,N_39730,N_37794);
or U40713 (N_40713,N_38965,N_39810);
and U40714 (N_40714,N_39472,N_38102);
nor U40715 (N_40715,N_38036,N_38992);
and U40716 (N_40716,N_39981,N_38371);
nor U40717 (N_40717,N_38563,N_37626);
or U40718 (N_40718,N_39572,N_38636);
and U40719 (N_40719,N_38288,N_39903);
or U40720 (N_40720,N_37958,N_38854);
xor U40721 (N_40721,N_39160,N_38248);
nor U40722 (N_40722,N_39012,N_39384);
and U40723 (N_40723,N_38918,N_39835);
xor U40724 (N_40724,N_37862,N_37791);
and U40725 (N_40725,N_37868,N_37951);
nand U40726 (N_40726,N_39473,N_39797);
nand U40727 (N_40727,N_39989,N_38643);
or U40728 (N_40728,N_38174,N_37961);
nand U40729 (N_40729,N_38037,N_38947);
nor U40730 (N_40730,N_38726,N_38996);
xor U40731 (N_40731,N_37593,N_38957);
nand U40732 (N_40732,N_39633,N_38073);
xor U40733 (N_40733,N_38731,N_39990);
xor U40734 (N_40734,N_39319,N_39144);
nor U40735 (N_40735,N_38005,N_38993);
or U40736 (N_40736,N_38211,N_37669);
and U40737 (N_40737,N_37658,N_39895);
nor U40738 (N_40738,N_39372,N_37896);
nand U40739 (N_40739,N_38045,N_37752);
nand U40740 (N_40740,N_39949,N_37716);
nor U40741 (N_40741,N_39246,N_38297);
nor U40742 (N_40742,N_39971,N_38083);
nand U40743 (N_40743,N_39486,N_38210);
nor U40744 (N_40744,N_39667,N_38420);
and U40745 (N_40745,N_39068,N_38769);
xor U40746 (N_40746,N_38319,N_38509);
xnor U40747 (N_40747,N_38949,N_38479);
nor U40748 (N_40748,N_39224,N_38314);
nand U40749 (N_40749,N_38733,N_39601);
xnor U40750 (N_40750,N_38021,N_39530);
nor U40751 (N_40751,N_39934,N_38851);
xor U40752 (N_40752,N_37509,N_37613);
or U40753 (N_40753,N_39474,N_37657);
nor U40754 (N_40754,N_39796,N_39419);
xnor U40755 (N_40755,N_37898,N_38362);
and U40756 (N_40756,N_38178,N_38421);
or U40757 (N_40757,N_37659,N_39535);
nor U40758 (N_40758,N_37691,N_38042);
xnor U40759 (N_40759,N_39463,N_38016);
or U40760 (N_40760,N_38161,N_39217);
nor U40761 (N_40761,N_39051,N_37834);
nand U40762 (N_40762,N_38902,N_38826);
xor U40763 (N_40763,N_37970,N_39607);
xor U40764 (N_40764,N_38596,N_39023);
and U40765 (N_40765,N_39031,N_39757);
or U40766 (N_40766,N_38531,N_39281);
nand U40767 (N_40767,N_39386,N_38920);
xnor U40768 (N_40768,N_38071,N_39013);
or U40769 (N_40769,N_38998,N_39050);
or U40770 (N_40770,N_38786,N_38821);
and U40771 (N_40771,N_38739,N_38075);
nor U40772 (N_40772,N_39373,N_39005);
nand U40773 (N_40773,N_37848,N_37581);
nand U40774 (N_40774,N_37550,N_38013);
nor U40775 (N_40775,N_38802,N_39731);
xor U40776 (N_40776,N_39362,N_38235);
and U40777 (N_40777,N_39398,N_38776);
xnor U40778 (N_40778,N_37505,N_37900);
nor U40779 (N_40779,N_39345,N_38773);
and U40780 (N_40780,N_38065,N_38056);
nand U40781 (N_40781,N_39813,N_38664);
xor U40782 (N_40782,N_39879,N_39728);
or U40783 (N_40783,N_37737,N_37562);
nand U40784 (N_40784,N_39204,N_39317);
or U40785 (N_40785,N_39407,N_37889);
nand U40786 (N_40786,N_39067,N_39648);
xor U40787 (N_40787,N_39542,N_39940);
nor U40788 (N_40788,N_38032,N_37915);
xnor U40789 (N_40789,N_37640,N_38310);
xor U40790 (N_40790,N_39370,N_37979);
and U40791 (N_40791,N_39353,N_37842);
nand U40792 (N_40792,N_38535,N_37664);
or U40793 (N_40793,N_39637,N_39266);
xor U40794 (N_40794,N_37749,N_37990);
or U40795 (N_40795,N_39320,N_38686);
nor U40796 (N_40796,N_38813,N_37590);
or U40797 (N_40797,N_38214,N_38936);
xnor U40798 (N_40798,N_39696,N_38291);
nor U40799 (N_40799,N_39961,N_38237);
nand U40800 (N_40800,N_38551,N_38365);
and U40801 (N_40801,N_39672,N_38817);
xnor U40802 (N_40802,N_38549,N_39443);
nor U40803 (N_40803,N_39163,N_38066);
xor U40804 (N_40804,N_38717,N_39957);
or U40805 (N_40805,N_39727,N_37685);
or U40806 (N_40806,N_37865,N_37819);
and U40807 (N_40807,N_39090,N_37674);
xnor U40808 (N_40808,N_39302,N_39870);
and U40809 (N_40809,N_37717,N_38608);
nand U40810 (N_40810,N_38962,N_39545);
and U40811 (N_40811,N_38335,N_38659);
xnor U40812 (N_40812,N_39458,N_38062);
xnor U40813 (N_40813,N_39825,N_39235);
or U40814 (N_40814,N_38857,N_38206);
xnor U40815 (N_40815,N_39054,N_37666);
nand U40816 (N_40816,N_39874,N_37636);
and U40817 (N_40817,N_39478,N_39852);
and U40818 (N_40818,N_38289,N_38534);
and U40819 (N_40819,N_38244,N_38381);
nand U40820 (N_40820,N_37845,N_38765);
nor U40821 (N_40821,N_38091,N_37520);
nand U40822 (N_40822,N_38900,N_37939);
and U40823 (N_40823,N_38861,N_39325);
or U40824 (N_40824,N_38386,N_39168);
or U40825 (N_40825,N_39688,N_39910);
or U40826 (N_40826,N_38933,N_39234);
or U40827 (N_40827,N_37570,N_37956);
nand U40828 (N_40828,N_38254,N_38590);
or U40829 (N_40829,N_37803,N_39297);
xor U40830 (N_40830,N_39284,N_38587);
and U40831 (N_40831,N_39749,N_39582);
nand U40832 (N_40832,N_37940,N_38601);
nand U40833 (N_40833,N_37952,N_39768);
nor U40834 (N_40834,N_39581,N_39614);
nor U40835 (N_40835,N_39579,N_37579);
or U40836 (N_40836,N_39170,N_38756);
or U40837 (N_40837,N_39877,N_39559);
xor U40838 (N_40838,N_37566,N_38101);
xnor U40839 (N_40839,N_39445,N_39165);
nand U40840 (N_40840,N_39378,N_39846);
nor U40841 (N_40841,N_38184,N_38838);
or U40842 (N_40842,N_39911,N_37881);
xor U40843 (N_40843,N_38921,N_37977);
or U40844 (N_40844,N_37515,N_38521);
nor U40845 (N_40845,N_39423,N_38175);
xor U40846 (N_40846,N_38736,N_39927);
and U40847 (N_40847,N_39901,N_37596);
or U40848 (N_40848,N_39424,N_39908);
and U40849 (N_40849,N_39480,N_38899);
nand U40850 (N_40850,N_38316,N_39430);
and U40851 (N_40851,N_39953,N_39063);
nor U40852 (N_40852,N_39311,N_38015);
or U40853 (N_40853,N_38911,N_37507);
nor U40854 (N_40854,N_38402,N_37847);
nand U40855 (N_40855,N_37966,N_39202);
nand U40856 (N_40856,N_38132,N_39616);
or U40857 (N_40857,N_39268,N_38064);
xnor U40858 (N_40858,N_37777,N_38343);
nand U40859 (N_40859,N_38976,N_38094);
and U40860 (N_40860,N_38652,N_37588);
nand U40861 (N_40861,N_39312,N_38806);
and U40862 (N_40862,N_38022,N_39896);
and U40863 (N_40863,N_39390,N_37564);
or U40864 (N_40864,N_39928,N_39464);
nand U40865 (N_40865,N_39447,N_38820);
xor U40866 (N_40866,N_38730,N_38203);
and U40867 (N_40867,N_37960,N_39970);
or U40868 (N_40868,N_37741,N_38505);
nand U40869 (N_40869,N_38407,N_37682);
or U40870 (N_40870,N_39890,N_39518);
and U40871 (N_40871,N_39995,N_38427);
nor U40872 (N_40872,N_39269,N_39179);
xnor U40873 (N_40873,N_39393,N_39062);
nor U40874 (N_40874,N_39618,N_37534);
and U40875 (N_40875,N_37953,N_38119);
xor U40876 (N_40876,N_39515,N_38486);
and U40877 (N_40877,N_37667,N_39892);
nor U40878 (N_40878,N_38740,N_39070);
and U40879 (N_40879,N_38525,N_37853);
or U40880 (N_40880,N_37722,N_39718);
nor U40881 (N_40881,N_39245,N_37831);
or U40882 (N_40882,N_38671,N_38169);
nand U40883 (N_40883,N_39617,N_37836);
nor U40884 (N_40884,N_38795,N_39854);
nand U40885 (N_40885,N_38803,N_37692);
or U40886 (N_40886,N_38763,N_38163);
nor U40887 (N_40887,N_38043,N_39288);
or U40888 (N_40888,N_39634,N_38249);
or U40889 (N_40889,N_37647,N_38850);
nor U40890 (N_40890,N_37895,N_39328);
and U40891 (N_40891,N_39700,N_38905);
xor U40892 (N_40892,N_37720,N_38351);
nand U40893 (N_40893,N_37516,N_37568);
xor U40894 (N_40894,N_38641,N_38844);
and U40895 (N_40895,N_38796,N_38642);
nand U40896 (N_40896,N_38264,N_39685);
nor U40897 (N_40897,N_38153,N_38510);
and U40898 (N_40898,N_38277,N_38722);
nand U40899 (N_40899,N_39074,N_38485);
and U40900 (N_40900,N_39273,N_38340);
xnor U40901 (N_40901,N_39963,N_39361);
nor U40902 (N_40902,N_38261,N_38059);
nand U40903 (N_40903,N_39764,N_38574);
nand U40904 (N_40904,N_38367,N_38762);
and U40905 (N_40905,N_38502,N_39040);
nand U40906 (N_40906,N_38771,N_37742);
nand U40907 (N_40907,N_37736,N_37621);
nand U40908 (N_40908,N_38103,N_39603);
or U40909 (N_40909,N_39138,N_37976);
and U40910 (N_40910,N_38698,N_39368);
xnor U40911 (N_40911,N_38088,N_39669);
xor U40912 (N_40912,N_37603,N_37873);
nand U40913 (N_40913,N_38082,N_37867);
or U40914 (N_40914,N_39774,N_37632);
and U40915 (N_40915,N_37888,N_39429);
or U40916 (N_40916,N_38682,N_39706);
or U40917 (N_40917,N_38217,N_38882);
and U40918 (N_40918,N_38967,N_39400);
and U40919 (N_40919,N_37829,N_39135);
xor U40920 (N_40920,N_39574,N_39975);
or U40921 (N_40921,N_38584,N_39436);
and U40922 (N_40922,N_39225,N_39972);
nand U40923 (N_40923,N_38374,N_39069);
nor U40924 (N_40924,N_37805,N_38360);
and U40925 (N_40925,N_38925,N_39263);
xnor U40926 (N_40926,N_39771,N_38368);
and U40927 (N_40927,N_38357,N_39828);
nand U40928 (N_40928,N_38681,N_39002);
nand U40929 (N_40929,N_39381,N_39968);
nand U40930 (N_40930,N_38700,N_39174);
xnor U40931 (N_40931,N_37909,N_37551);
nand U40932 (N_40932,N_37840,N_39124);
or U40933 (N_40933,N_39267,N_39673);
xor U40934 (N_40934,N_37828,N_38822);
or U40935 (N_40935,N_39324,N_39772);
nand U40936 (N_40936,N_39099,N_38417);
xnor U40937 (N_40937,N_38961,N_39988);
and U40938 (N_40938,N_39113,N_38041);
xnor U40939 (N_40939,N_39543,N_37694);
xor U40940 (N_40940,N_39919,N_37860);
and U40941 (N_40941,N_38500,N_39923);
nor U40942 (N_40942,N_39110,N_38008);
nand U40943 (N_40943,N_39298,N_39836);
or U40944 (N_40944,N_38406,N_39921);
nor U40945 (N_40945,N_39866,N_37838);
xor U40946 (N_40946,N_39506,N_39605);
or U40947 (N_40947,N_37767,N_39295);
and U40948 (N_40948,N_39692,N_38536);
xor U40949 (N_40949,N_39363,N_39360);
or U40950 (N_40950,N_37883,N_38182);
nand U40951 (N_40951,N_39841,N_39615);
nand U40952 (N_40952,N_37545,N_39594);
xnor U40953 (N_40953,N_38166,N_39162);
xor U40954 (N_40954,N_39186,N_39752);
and U40955 (N_40955,N_37637,N_39915);
and U40956 (N_40956,N_39490,N_39876);
nor U40957 (N_40957,N_39703,N_39984);
nor U40958 (N_40958,N_38708,N_38284);
and U40959 (N_40959,N_38693,N_39740);
nand U40960 (N_40960,N_38034,N_38837);
nand U40961 (N_40961,N_39746,N_38093);
nand U40962 (N_40962,N_38718,N_38201);
or U40963 (N_40963,N_39826,N_38677);
nand U40964 (N_40964,N_39257,N_38377);
or U40965 (N_40965,N_39264,N_38670);
or U40966 (N_40966,N_37839,N_39349);
and U40967 (N_40967,N_38597,N_38142);
and U40968 (N_40968,N_38678,N_39139);
or U40969 (N_40969,N_37546,N_37706);
and U40970 (N_40970,N_39446,N_38453);
xnor U40971 (N_40971,N_38554,N_39804);
nand U40972 (N_40972,N_38830,N_39036);
nand U40973 (N_40973,N_39404,N_39693);
nand U40974 (N_40974,N_38450,N_38738);
nand U40975 (N_40975,N_39922,N_38629);
xnor U40976 (N_40976,N_37949,N_39141);
or U40977 (N_40977,N_39812,N_37866);
nor U40978 (N_40978,N_39095,N_37628);
and U40979 (N_40979,N_39899,N_39775);
and U40980 (N_40980,N_39344,N_39254);
and U40981 (N_40981,N_38471,N_38761);
or U40982 (N_40982,N_38891,N_38909);
nand U40983 (N_40983,N_38250,N_38495);
nand U40984 (N_40984,N_39863,N_39948);
and U40985 (N_40985,N_38147,N_39743);
nor U40986 (N_40986,N_38886,N_38048);
xor U40987 (N_40987,N_38078,N_39466);
xnor U40988 (N_40988,N_37652,N_38805);
nor U40989 (N_40989,N_37653,N_39704);
and U40990 (N_40990,N_38130,N_38315);
and U40991 (N_40991,N_37924,N_39816);
or U40992 (N_40992,N_37723,N_38887);
and U40993 (N_40993,N_38972,N_38859);
and U40994 (N_40994,N_39980,N_39644);
or U40995 (N_40995,N_39756,N_38476);
xnor U40996 (N_40996,N_39310,N_39323);
nand U40997 (N_40997,N_38585,N_38910);
nand U40998 (N_40998,N_38437,N_39862);
and U40999 (N_40999,N_37919,N_37502);
nor U41000 (N_41000,N_38526,N_38986);
nand U41001 (N_41001,N_39285,N_38081);
nand U41002 (N_41002,N_37814,N_38968);
xor U41003 (N_41003,N_37536,N_38414);
or U41004 (N_41004,N_38952,N_39180);
xnor U41005 (N_41005,N_39111,N_38024);
and U41006 (N_41006,N_38559,N_37972);
or U41007 (N_41007,N_39157,N_39366);
and U41008 (N_41008,N_39275,N_38544);
nor U41009 (N_41009,N_37820,N_37629);
nand U41010 (N_41010,N_37623,N_38260);
nand U41011 (N_41011,N_39432,N_38793);
nor U41012 (N_41012,N_39952,N_38216);
or U41013 (N_41013,N_38246,N_38287);
nor U41014 (N_41014,N_39201,N_38493);
nand U41015 (N_41015,N_38755,N_37818);
nor U41016 (N_41016,N_38687,N_39788);
xor U41017 (N_41017,N_39093,N_38917);
and U41018 (N_41018,N_37772,N_39032);
or U41019 (N_41019,N_39034,N_38948);
nor U41020 (N_41020,N_38481,N_38653);
nor U41021 (N_41021,N_38635,N_38741);
nor U41022 (N_41022,N_39767,N_37615);
and U41023 (N_41023,N_37983,N_38027);
xor U41024 (N_41024,N_38366,N_39785);
or U41025 (N_41025,N_38063,N_38441);
and U41026 (N_41026,N_38788,N_38383);
or U41027 (N_41027,N_39897,N_38564);
and U41028 (N_41028,N_38000,N_39900);
or U41029 (N_41029,N_39576,N_37721);
nand U41030 (N_41030,N_38890,N_39973);
nor U41031 (N_41031,N_38672,N_39600);
or U41032 (N_41032,N_39947,N_39818);
and U41033 (N_41033,N_39819,N_39042);
nand U41034 (N_41034,N_38133,N_39388);
and U41035 (N_41035,N_39356,N_38666);
nand U41036 (N_41036,N_38118,N_38159);
or U41037 (N_41037,N_38002,N_39119);
xor U41038 (N_41038,N_39638,N_38168);
nor U41039 (N_41039,N_37790,N_39279);
nor U41040 (N_41040,N_39420,N_39556);
nor U41041 (N_41041,N_37503,N_38160);
xor U41042 (N_41042,N_39194,N_39402);
or U41043 (N_41043,N_37929,N_38873);
or U41044 (N_41044,N_39150,N_38516);
nand U41045 (N_41045,N_37527,N_38540);
nor U41046 (N_41046,N_38356,N_38801);
nand U41047 (N_41047,N_39994,N_37999);
xor U41048 (N_41048,N_37917,N_39679);
or U41049 (N_41049,N_38208,N_39848);
nor U41050 (N_41050,N_39946,N_38667);
or U41051 (N_41051,N_38446,N_37586);
nand U41052 (N_41052,N_38241,N_37787);
and U41053 (N_41053,N_39291,N_38393);
xnor U41054 (N_41054,N_38279,N_39931);
or U41055 (N_41055,N_39001,N_37763);
nor U41056 (N_41056,N_39265,N_39849);
or U41057 (N_41057,N_38637,N_38151);
nor U41058 (N_41058,N_37511,N_39017);
or U41059 (N_41059,N_38436,N_37844);
and U41060 (N_41060,N_38789,N_38742);
and U41061 (N_41061,N_39751,N_39244);
xnor U41062 (N_41062,N_39395,N_39175);
nor U41063 (N_41063,N_38721,N_38492);
nand U41064 (N_41064,N_38852,N_38665);
and U41065 (N_41065,N_37931,N_38798);
and U41066 (N_41066,N_38188,N_38192);
or U41067 (N_41067,N_39041,N_39454);
nand U41068 (N_41068,N_38049,N_37756);
nor U41069 (N_41069,N_39690,N_38581);
nor U41070 (N_41070,N_39596,N_37799);
and U41071 (N_41071,N_39917,N_39586);
xor U41072 (N_41072,N_37861,N_37687);
xor U41073 (N_41073,N_39513,N_38484);
xnor U41074 (N_41074,N_38072,N_38331);
or U41075 (N_41075,N_38680,N_39569);
nand U41076 (N_41076,N_37864,N_39627);
nand U41077 (N_41077,N_37569,N_38272);
xnor U41078 (N_41078,N_38413,N_39553);
nand U41079 (N_41079,N_38845,N_37938);
xor U41080 (N_41080,N_39628,N_38442);
xnor U41081 (N_41081,N_38979,N_39314);
and U41082 (N_41082,N_37910,N_37789);
nand U41083 (N_41083,N_38747,N_37988);
or U41084 (N_41084,N_37555,N_38808);
and U41085 (N_41085,N_38675,N_38097);
nand U41086 (N_41086,N_39132,N_39570);
nor U41087 (N_41087,N_39780,N_39610);
or U41088 (N_41088,N_39512,N_38939);
or U41089 (N_41089,N_38209,N_39211);
and U41090 (N_41090,N_39843,N_39537);
xnor U41091 (N_41091,N_39118,N_38646);
and U41092 (N_41092,N_39635,N_39558);
nor U41093 (N_41093,N_38090,N_38916);
xnor U41094 (N_41094,N_38263,N_39121);
or U41095 (N_41095,N_39337,N_39604);
xor U41096 (N_41096,N_38074,N_39448);
xnor U41097 (N_41097,N_39130,N_39391);
xor U41098 (N_41098,N_37557,N_39941);
xor U41099 (N_41099,N_38149,N_37673);
xor U41100 (N_41100,N_39487,N_39678);
nor U41101 (N_41101,N_38723,N_38567);
nand U41102 (N_41102,N_38387,N_38483);
or U41103 (N_41103,N_39987,N_37959);
xnor U41104 (N_41104,N_37989,N_38220);
xnor U41105 (N_41105,N_39071,N_38538);
or U41106 (N_41106,N_37547,N_38392);
nand U41107 (N_41107,N_38033,N_38475);
or U41108 (N_41108,N_38932,N_39529);
and U41109 (N_41109,N_38375,N_39189);
nor U41110 (N_41110,N_38302,N_38547);
nand U41111 (N_41111,N_37735,N_38734);
nand U41112 (N_41112,N_39027,N_39820);
and U41113 (N_41113,N_37554,N_38893);
and U41114 (N_41114,N_39136,N_38293);
nand U41115 (N_41115,N_38689,N_38530);
xnor U41116 (N_41116,N_37793,N_39955);
nor U41117 (N_41117,N_39469,N_39441);
nor U41118 (N_41118,N_38589,N_38029);
or U41119 (N_41119,N_38076,N_37870);
nor U41120 (N_41120,N_38465,N_37841);
nor U41121 (N_41121,N_37833,N_38729);
xor U41122 (N_41122,N_38190,N_37619);
nand U41123 (N_41123,N_37941,N_39250);
and U41124 (N_41124,N_38990,N_37524);
or U41125 (N_41125,N_39620,N_39597);
xor U41126 (N_41126,N_39799,N_37857);
nand U41127 (N_41127,N_38599,N_37543);
nand U41128 (N_41128,N_37975,N_37625);
nor U41129 (N_41129,N_39318,N_39208);
nor U41130 (N_41130,N_38578,N_37757);
nor U41131 (N_41131,N_38238,N_37921);
nand U41132 (N_41132,N_39382,N_39467);
nor U41133 (N_41133,N_38868,N_39997);
nand U41134 (N_41134,N_39026,N_39753);
or U41135 (N_41135,N_37876,N_37997);
nor U41136 (N_41136,N_38570,N_38985);
nand U41137 (N_41137,N_38922,N_39904);
nand U41138 (N_41138,N_39505,N_38205);
xnor U41139 (N_41139,N_39551,N_39619);
and U41140 (N_41140,N_38394,N_38313);
nor U41141 (N_41141,N_38764,N_39232);
and U41142 (N_41142,N_39709,N_38382);
nor U41143 (N_41143,N_39523,N_39563);
xnor U41144 (N_41144,N_37802,N_38923);
and U41145 (N_41145,N_39844,N_37695);
or U41146 (N_41146,N_38695,N_38245);
nor U41147 (N_41147,N_38662,N_37893);
and U41148 (N_41148,N_37800,N_39073);
xor U41149 (N_41149,N_38018,N_38422);
and U41150 (N_41150,N_39869,N_39151);
nor U41151 (N_41151,N_37913,N_37731);
nor U41152 (N_41152,N_39815,N_38676);
nor U41153 (N_41153,N_39734,N_38183);
or U41154 (N_41154,N_38213,N_37964);
nor U41155 (N_41155,N_38198,N_39248);
nand U41156 (N_41156,N_38380,N_37765);
nor U41157 (N_41157,N_39479,N_37661);
and U41158 (N_41158,N_39956,N_39401);
and U41159 (N_41159,N_39549,N_38116);
or U41160 (N_41160,N_37512,N_37766);
nor U41161 (N_41161,N_39670,N_39663);
xor U41162 (N_41162,N_39066,N_38528);
nand U41163 (N_41163,N_38870,N_39598);
and U41164 (N_41164,N_39080,N_39365);
nand U41165 (N_41165,N_39422,N_39006);
or U41166 (N_41166,N_38164,N_38770);
and U41167 (N_41167,N_38583,N_38834);
nand U41168 (N_41168,N_38503,N_38328);
xor U41169 (N_41169,N_37530,N_39243);
or U41170 (N_41170,N_39019,N_37681);
nand U41171 (N_41171,N_39991,N_39022);
nand U41172 (N_41172,N_39329,N_38654);
nor U41173 (N_41173,N_39321,N_38699);
and U41174 (N_41174,N_37646,N_38785);
or U41175 (N_41175,N_39674,N_38927);
nor U41176 (N_41176,N_38455,N_39000);
and U41177 (N_41177,N_38477,N_38580);
xnor U41178 (N_41178,N_39114,N_37746);
and U41179 (N_41179,N_39759,N_39226);
nand U41180 (N_41180,N_39524,N_39657);
and U41181 (N_41181,N_39966,N_38863);
and U41182 (N_41182,N_39656,N_39925);
nor U41183 (N_41183,N_37582,N_39104);
xnor U41184 (N_41184,N_38253,N_39459);
nor U41185 (N_41185,N_37738,N_39379);
nand U41186 (N_41186,N_38906,N_38257);
nand U41187 (N_41187,N_39262,N_38283);
and U41188 (N_41188,N_37679,N_37996);
or U41189 (N_41189,N_37700,N_38126);
nand U41190 (N_41190,N_38364,N_39158);
nor U41191 (N_41191,N_38595,N_37607);
or U41192 (N_41192,N_38832,N_37780);
or U41193 (N_41193,N_39072,N_38270);
nor U41194 (N_41194,N_37965,N_38555);
nand U41195 (N_41195,N_38888,N_37914);
and U41196 (N_41196,N_37523,N_37894);
nand U41197 (N_41197,N_39415,N_39763);
nand U41198 (N_41198,N_39428,N_38800);
or U41199 (N_41199,N_37558,N_39747);
nand U41200 (N_41200,N_39724,N_39546);
xnor U41201 (N_41201,N_38508,N_39205);
or U41202 (N_41202,N_38628,N_38714);
nor U41203 (N_41203,N_38794,N_38388);
nand U41204 (N_41204,N_39207,N_38294);
nand U41205 (N_41205,N_39612,N_37785);
nor U41206 (N_41206,N_39134,N_38519);
xnor U41207 (N_41207,N_38616,N_39294);
xnor U41208 (N_41208,N_39497,N_38696);
nand U41209 (N_41209,N_39555,N_37773);
nor U41210 (N_41210,N_39283,N_39510);
nand U41211 (N_41211,N_37830,N_39655);
nor U41212 (N_41212,N_37884,N_39744);
nand U41213 (N_41213,N_39200,N_39033);
nor U41214 (N_41214,N_38915,N_39847);
nor U41215 (N_41215,N_39086,N_39347);
nand U41216 (N_41216,N_38265,N_38052);
nand U41217 (N_41217,N_38501,N_39561);
or U41218 (N_41218,N_39377,N_39183);
nand U41219 (N_41219,N_38352,N_39742);
xor U41220 (N_41220,N_38898,N_37947);
and U41221 (N_41221,N_37764,N_39716);
and U41222 (N_41222,N_37897,N_39146);
nand U41223 (N_41223,N_39259,N_39038);
nand U41224 (N_41224,N_38204,N_37573);
nor U41225 (N_41225,N_37879,N_38657);
nand U41226 (N_41226,N_39375,N_38234);
nand U41227 (N_41227,N_39938,N_39453);
nand U41228 (N_41228,N_37798,N_38306);
nor U41229 (N_41229,N_38752,N_37755);
nand U41230 (N_41230,N_37991,N_38780);
or U41231 (N_41231,N_38170,N_39807);
or U41232 (N_41232,N_38656,N_38144);
or U41233 (N_41233,N_38827,N_39039);
nor U41234 (N_41234,N_38012,N_39891);
nor U41235 (N_41235,N_39290,N_38054);
or U41236 (N_41236,N_39557,N_38467);
and U41237 (N_41237,N_37644,N_37882);
nor U41238 (N_41238,N_39736,N_38884);
xor U41239 (N_41239,N_39683,N_38127);
nor U41240 (N_41240,N_38038,N_39075);
nor U41241 (N_41241,N_37875,N_37548);
nor U41242 (N_41242,N_37987,N_39705);
xnor U41243 (N_41243,N_39394,N_39773);
or U41244 (N_41244,N_37760,N_38668);
nand U41245 (N_41245,N_38085,N_39918);
or U41246 (N_41246,N_39383,N_38557);
nand U41247 (N_41247,N_39499,N_38200);
nor U41248 (N_41248,N_38561,N_39791);
nand U41249 (N_41249,N_39128,N_39240);
nor U41250 (N_41250,N_39201,N_39486);
and U41251 (N_41251,N_38070,N_39875);
nor U41252 (N_41252,N_38763,N_39552);
xor U41253 (N_41253,N_39309,N_39887);
and U41254 (N_41254,N_39343,N_39713);
xnor U41255 (N_41255,N_39767,N_39834);
nor U41256 (N_41256,N_38881,N_38307);
or U41257 (N_41257,N_39008,N_37675);
nand U41258 (N_41258,N_39143,N_38953);
and U41259 (N_41259,N_39061,N_38730);
nor U41260 (N_41260,N_39243,N_38042);
or U41261 (N_41261,N_39125,N_38244);
xnor U41262 (N_41262,N_39795,N_38153);
and U41263 (N_41263,N_39353,N_38261);
nand U41264 (N_41264,N_39723,N_39642);
xnor U41265 (N_41265,N_38191,N_38450);
xor U41266 (N_41266,N_39893,N_39024);
nand U41267 (N_41267,N_39012,N_37604);
xnor U41268 (N_41268,N_38027,N_38111);
xor U41269 (N_41269,N_38717,N_39069);
and U41270 (N_41270,N_38166,N_39648);
xnor U41271 (N_41271,N_38080,N_37532);
nand U41272 (N_41272,N_37827,N_39170);
nor U41273 (N_41273,N_39063,N_38305);
or U41274 (N_41274,N_39340,N_39292);
and U41275 (N_41275,N_37666,N_37904);
xnor U41276 (N_41276,N_38082,N_37640);
and U41277 (N_41277,N_37600,N_39981);
and U41278 (N_41278,N_38627,N_39546);
nor U41279 (N_41279,N_37520,N_37673);
and U41280 (N_41280,N_37641,N_38124);
xnor U41281 (N_41281,N_39004,N_39084);
nand U41282 (N_41282,N_39688,N_38918);
nor U41283 (N_41283,N_39359,N_39473);
xnor U41284 (N_41284,N_37507,N_38960);
and U41285 (N_41285,N_39068,N_37587);
nor U41286 (N_41286,N_39614,N_38908);
xnor U41287 (N_41287,N_38645,N_38724);
or U41288 (N_41288,N_39691,N_39903);
and U41289 (N_41289,N_38239,N_39435);
and U41290 (N_41290,N_38717,N_38445);
nor U41291 (N_41291,N_38944,N_38318);
nor U41292 (N_41292,N_37898,N_39025);
xor U41293 (N_41293,N_39980,N_39524);
xor U41294 (N_41294,N_38216,N_38018);
xor U41295 (N_41295,N_38394,N_39491);
nand U41296 (N_41296,N_38942,N_37803);
nor U41297 (N_41297,N_37922,N_38963);
nor U41298 (N_41298,N_37668,N_39838);
and U41299 (N_41299,N_38352,N_37630);
and U41300 (N_41300,N_39078,N_38893);
and U41301 (N_41301,N_39528,N_38139);
xnor U41302 (N_41302,N_38913,N_38406);
or U41303 (N_41303,N_39872,N_39566);
and U41304 (N_41304,N_39259,N_37820);
nor U41305 (N_41305,N_37598,N_38466);
or U41306 (N_41306,N_38755,N_38082);
nor U41307 (N_41307,N_38866,N_38841);
or U41308 (N_41308,N_39508,N_38075);
or U41309 (N_41309,N_39001,N_38048);
xnor U41310 (N_41310,N_39702,N_38162);
xnor U41311 (N_41311,N_37624,N_39044);
xnor U41312 (N_41312,N_38688,N_39517);
and U41313 (N_41313,N_38334,N_38746);
xor U41314 (N_41314,N_39701,N_39141);
xor U41315 (N_41315,N_39530,N_39611);
or U41316 (N_41316,N_39473,N_38251);
and U41317 (N_41317,N_39384,N_38593);
nor U41318 (N_41318,N_39398,N_38132);
nor U41319 (N_41319,N_38245,N_38084);
xor U41320 (N_41320,N_38992,N_39436);
nor U41321 (N_41321,N_38142,N_37692);
and U41322 (N_41322,N_38154,N_37954);
nand U41323 (N_41323,N_38509,N_38878);
or U41324 (N_41324,N_39204,N_39174);
and U41325 (N_41325,N_38501,N_39091);
nand U41326 (N_41326,N_38502,N_38840);
nor U41327 (N_41327,N_39879,N_39246);
xnor U41328 (N_41328,N_38924,N_37782);
and U41329 (N_41329,N_39956,N_38895);
nor U41330 (N_41330,N_38737,N_37999);
or U41331 (N_41331,N_37991,N_39970);
and U41332 (N_41332,N_38244,N_38986);
or U41333 (N_41333,N_39113,N_38724);
and U41334 (N_41334,N_37787,N_38193);
and U41335 (N_41335,N_38328,N_39845);
or U41336 (N_41336,N_38197,N_39184);
nand U41337 (N_41337,N_38030,N_39716);
or U41338 (N_41338,N_38952,N_37947);
nor U41339 (N_41339,N_38974,N_37924);
or U41340 (N_41340,N_38902,N_37615);
xor U41341 (N_41341,N_38865,N_39460);
nand U41342 (N_41342,N_38580,N_38768);
xor U41343 (N_41343,N_39808,N_39262);
or U41344 (N_41344,N_37810,N_39037);
or U41345 (N_41345,N_37980,N_38388);
nand U41346 (N_41346,N_39575,N_38357);
or U41347 (N_41347,N_39571,N_38132);
xnor U41348 (N_41348,N_39825,N_37512);
or U41349 (N_41349,N_39902,N_38208);
nand U41350 (N_41350,N_39461,N_39496);
or U41351 (N_41351,N_38264,N_38837);
nand U41352 (N_41352,N_39859,N_39855);
and U41353 (N_41353,N_38955,N_39797);
nand U41354 (N_41354,N_38014,N_38515);
nor U41355 (N_41355,N_39245,N_38844);
xnor U41356 (N_41356,N_38564,N_38151);
or U41357 (N_41357,N_37826,N_39248);
or U41358 (N_41358,N_37808,N_39017);
nand U41359 (N_41359,N_39360,N_39767);
xnor U41360 (N_41360,N_39708,N_38743);
nand U41361 (N_41361,N_38975,N_37939);
and U41362 (N_41362,N_39772,N_39576);
and U41363 (N_41363,N_37674,N_39861);
xor U41364 (N_41364,N_37635,N_38039);
or U41365 (N_41365,N_38923,N_38263);
nor U41366 (N_41366,N_38666,N_39128);
or U41367 (N_41367,N_38069,N_39420);
xor U41368 (N_41368,N_38303,N_38734);
nand U41369 (N_41369,N_38444,N_37819);
or U41370 (N_41370,N_38411,N_39837);
nor U41371 (N_41371,N_38002,N_37583);
nand U41372 (N_41372,N_38409,N_39975);
and U41373 (N_41373,N_38846,N_38770);
and U41374 (N_41374,N_38548,N_39436);
nand U41375 (N_41375,N_38100,N_38460);
xor U41376 (N_41376,N_38987,N_38788);
nor U41377 (N_41377,N_37694,N_38257);
and U41378 (N_41378,N_38016,N_39089);
nand U41379 (N_41379,N_39767,N_37632);
and U41380 (N_41380,N_39539,N_37801);
nor U41381 (N_41381,N_39931,N_37528);
xnor U41382 (N_41382,N_37742,N_38447);
nor U41383 (N_41383,N_39647,N_39732);
xnor U41384 (N_41384,N_38995,N_38410);
nor U41385 (N_41385,N_39297,N_37663);
nor U41386 (N_41386,N_37821,N_39827);
and U41387 (N_41387,N_39782,N_39153);
and U41388 (N_41388,N_39015,N_38760);
and U41389 (N_41389,N_39024,N_39471);
or U41390 (N_41390,N_39983,N_38851);
xor U41391 (N_41391,N_38603,N_39572);
nand U41392 (N_41392,N_38794,N_37795);
xnor U41393 (N_41393,N_39313,N_38084);
and U41394 (N_41394,N_37689,N_37770);
and U41395 (N_41395,N_38136,N_38663);
or U41396 (N_41396,N_38188,N_38108);
nor U41397 (N_41397,N_37563,N_39789);
nor U41398 (N_41398,N_39362,N_38443);
nor U41399 (N_41399,N_39713,N_38892);
nor U41400 (N_41400,N_38774,N_37567);
and U41401 (N_41401,N_37952,N_38969);
xnor U41402 (N_41402,N_38764,N_39354);
and U41403 (N_41403,N_39111,N_39683);
xnor U41404 (N_41404,N_39540,N_39228);
xnor U41405 (N_41405,N_39181,N_39272);
nor U41406 (N_41406,N_38449,N_37524);
xor U41407 (N_41407,N_39399,N_37816);
nand U41408 (N_41408,N_39804,N_39356);
xnor U41409 (N_41409,N_39344,N_37752);
xnor U41410 (N_41410,N_38044,N_39176);
or U41411 (N_41411,N_38405,N_39091);
xnor U41412 (N_41412,N_37511,N_39629);
nand U41413 (N_41413,N_38807,N_38289);
or U41414 (N_41414,N_39571,N_39810);
or U41415 (N_41415,N_39517,N_39584);
xnor U41416 (N_41416,N_37580,N_37919);
and U41417 (N_41417,N_38515,N_38672);
or U41418 (N_41418,N_39747,N_39562);
nor U41419 (N_41419,N_38675,N_37679);
and U41420 (N_41420,N_37764,N_39367);
xnor U41421 (N_41421,N_38795,N_38694);
nand U41422 (N_41422,N_39788,N_39520);
xnor U41423 (N_41423,N_38677,N_38077);
nand U41424 (N_41424,N_38162,N_37595);
nand U41425 (N_41425,N_38616,N_38505);
nand U41426 (N_41426,N_39807,N_39664);
nand U41427 (N_41427,N_38364,N_38115);
or U41428 (N_41428,N_39231,N_37574);
xnor U41429 (N_41429,N_38605,N_39914);
xnor U41430 (N_41430,N_38593,N_39576);
xor U41431 (N_41431,N_39837,N_39709);
nand U41432 (N_41432,N_37562,N_37893);
or U41433 (N_41433,N_38233,N_39307);
nor U41434 (N_41434,N_39144,N_37531);
nor U41435 (N_41435,N_37953,N_39530);
nand U41436 (N_41436,N_39366,N_38013);
and U41437 (N_41437,N_39725,N_37516);
xnor U41438 (N_41438,N_37811,N_39078);
and U41439 (N_41439,N_38683,N_39503);
nor U41440 (N_41440,N_39249,N_38013);
nor U41441 (N_41441,N_38526,N_39744);
or U41442 (N_41442,N_39783,N_38401);
xor U41443 (N_41443,N_39618,N_38970);
xor U41444 (N_41444,N_37550,N_39691);
nand U41445 (N_41445,N_39184,N_38536);
nor U41446 (N_41446,N_38691,N_37553);
or U41447 (N_41447,N_39572,N_38136);
nand U41448 (N_41448,N_39244,N_39656);
nand U41449 (N_41449,N_38251,N_38765);
nand U41450 (N_41450,N_39728,N_38176);
nand U41451 (N_41451,N_38809,N_37954);
xor U41452 (N_41452,N_39890,N_37694);
and U41453 (N_41453,N_38166,N_38531);
nand U41454 (N_41454,N_39080,N_37794);
nor U41455 (N_41455,N_38441,N_39531);
nor U41456 (N_41456,N_38019,N_38277);
or U41457 (N_41457,N_37615,N_39037);
or U41458 (N_41458,N_38618,N_38464);
xnor U41459 (N_41459,N_39367,N_38005);
or U41460 (N_41460,N_38378,N_38555);
nor U41461 (N_41461,N_38535,N_39100);
or U41462 (N_41462,N_38074,N_39233);
nand U41463 (N_41463,N_39815,N_37694);
and U41464 (N_41464,N_38494,N_38563);
and U41465 (N_41465,N_38078,N_38640);
xor U41466 (N_41466,N_39577,N_38500);
nand U41467 (N_41467,N_38264,N_37777);
xnor U41468 (N_41468,N_39585,N_38746);
or U41469 (N_41469,N_38920,N_38576);
and U41470 (N_41470,N_38146,N_38629);
nor U41471 (N_41471,N_38368,N_38354);
and U41472 (N_41472,N_37577,N_38284);
and U41473 (N_41473,N_39329,N_38831);
or U41474 (N_41474,N_38386,N_37552);
xor U41475 (N_41475,N_39831,N_38101);
nor U41476 (N_41476,N_39289,N_38857);
xor U41477 (N_41477,N_38632,N_39329);
and U41478 (N_41478,N_39330,N_39495);
or U41479 (N_41479,N_37728,N_37678);
xor U41480 (N_41480,N_37580,N_38456);
and U41481 (N_41481,N_38456,N_39641);
and U41482 (N_41482,N_38947,N_39310);
and U41483 (N_41483,N_37829,N_37938);
nor U41484 (N_41484,N_38278,N_39053);
xnor U41485 (N_41485,N_39738,N_38655);
nand U41486 (N_41486,N_38810,N_38526);
nor U41487 (N_41487,N_39771,N_38288);
or U41488 (N_41488,N_37700,N_39585);
and U41489 (N_41489,N_38940,N_39343);
and U41490 (N_41490,N_39933,N_39229);
nand U41491 (N_41491,N_38747,N_39599);
nand U41492 (N_41492,N_37546,N_38001);
nor U41493 (N_41493,N_39252,N_38522);
and U41494 (N_41494,N_38998,N_39352);
or U41495 (N_41495,N_39127,N_39389);
xor U41496 (N_41496,N_39883,N_39318);
xnor U41497 (N_41497,N_39512,N_38245);
and U41498 (N_41498,N_39691,N_39254);
or U41499 (N_41499,N_39569,N_39763);
xor U41500 (N_41500,N_38209,N_37532);
and U41501 (N_41501,N_37923,N_38060);
or U41502 (N_41502,N_37775,N_39595);
or U41503 (N_41503,N_39215,N_38903);
xnor U41504 (N_41504,N_39631,N_38924);
nor U41505 (N_41505,N_39577,N_39821);
nand U41506 (N_41506,N_38326,N_38342);
nand U41507 (N_41507,N_39874,N_39788);
nor U41508 (N_41508,N_38856,N_38666);
xnor U41509 (N_41509,N_38038,N_39178);
or U41510 (N_41510,N_39386,N_39839);
or U41511 (N_41511,N_39165,N_37949);
xnor U41512 (N_41512,N_37931,N_37896);
nand U41513 (N_41513,N_37680,N_39359);
nand U41514 (N_41514,N_39566,N_39284);
xor U41515 (N_41515,N_39394,N_38591);
nand U41516 (N_41516,N_39975,N_37700);
or U41517 (N_41517,N_39987,N_38647);
and U41518 (N_41518,N_37797,N_38350);
nor U41519 (N_41519,N_38435,N_39062);
xor U41520 (N_41520,N_39867,N_38710);
or U41521 (N_41521,N_39875,N_39945);
xor U41522 (N_41522,N_38570,N_39087);
nand U41523 (N_41523,N_38367,N_39043);
xor U41524 (N_41524,N_39045,N_38042);
nor U41525 (N_41525,N_38161,N_39791);
xor U41526 (N_41526,N_39610,N_37525);
xor U41527 (N_41527,N_38642,N_39688);
nor U41528 (N_41528,N_38882,N_38309);
and U41529 (N_41529,N_38017,N_39144);
nor U41530 (N_41530,N_38784,N_39513);
or U41531 (N_41531,N_37983,N_38661);
xor U41532 (N_41532,N_37954,N_38720);
xor U41533 (N_41533,N_39404,N_38288);
nor U41534 (N_41534,N_37802,N_39726);
or U41535 (N_41535,N_38013,N_39516);
nor U41536 (N_41536,N_38837,N_39249);
and U41537 (N_41537,N_38520,N_38079);
nor U41538 (N_41538,N_39608,N_38231);
nand U41539 (N_41539,N_38195,N_39547);
and U41540 (N_41540,N_39821,N_38190);
nand U41541 (N_41541,N_39735,N_39593);
or U41542 (N_41542,N_37862,N_39090);
or U41543 (N_41543,N_39188,N_38767);
nand U41544 (N_41544,N_39892,N_38354);
nor U41545 (N_41545,N_39746,N_38047);
xor U41546 (N_41546,N_39114,N_39224);
xnor U41547 (N_41547,N_38479,N_38597);
xor U41548 (N_41548,N_39580,N_38426);
nand U41549 (N_41549,N_38501,N_39034);
nor U41550 (N_41550,N_38266,N_39917);
nand U41551 (N_41551,N_39529,N_38810);
and U41552 (N_41552,N_39774,N_39222);
nand U41553 (N_41553,N_39321,N_39766);
and U41554 (N_41554,N_37693,N_39719);
nor U41555 (N_41555,N_37781,N_37814);
or U41556 (N_41556,N_38512,N_37569);
xor U41557 (N_41557,N_39132,N_39353);
or U41558 (N_41558,N_38510,N_37653);
nor U41559 (N_41559,N_38934,N_39556);
and U41560 (N_41560,N_39416,N_39470);
xor U41561 (N_41561,N_39103,N_38765);
nand U41562 (N_41562,N_39271,N_39408);
nor U41563 (N_41563,N_39753,N_38076);
nor U41564 (N_41564,N_39112,N_39731);
and U41565 (N_41565,N_38888,N_37623);
xnor U41566 (N_41566,N_39872,N_38141);
nor U41567 (N_41567,N_39187,N_39181);
nor U41568 (N_41568,N_38329,N_38715);
xor U41569 (N_41569,N_38153,N_39714);
and U41570 (N_41570,N_39325,N_38878);
or U41571 (N_41571,N_38731,N_37896);
nand U41572 (N_41572,N_37757,N_38728);
xnor U41573 (N_41573,N_37702,N_39271);
xor U41574 (N_41574,N_38444,N_39432);
nand U41575 (N_41575,N_38737,N_39681);
nor U41576 (N_41576,N_38913,N_39387);
nor U41577 (N_41577,N_39735,N_38413);
and U41578 (N_41578,N_37847,N_37614);
xnor U41579 (N_41579,N_39486,N_38787);
or U41580 (N_41580,N_38942,N_38492);
xor U41581 (N_41581,N_38792,N_37850);
nor U41582 (N_41582,N_37994,N_39834);
nor U41583 (N_41583,N_38154,N_38374);
or U41584 (N_41584,N_37662,N_37981);
or U41585 (N_41585,N_38771,N_39714);
nand U41586 (N_41586,N_38795,N_39495);
and U41587 (N_41587,N_38895,N_39293);
and U41588 (N_41588,N_37564,N_38134);
nor U41589 (N_41589,N_39147,N_37959);
xnor U41590 (N_41590,N_38710,N_37690);
nand U41591 (N_41591,N_39057,N_39315);
nor U41592 (N_41592,N_39686,N_38923);
or U41593 (N_41593,N_39414,N_37566);
nor U41594 (N_41594,N_38374,N_38637);
xor U41595 (N_41595,N_38358,N_39123);
xnor U41596 (N_41596,N_37911,N_38687);
or U41597 (N_41597,N_39761,N_39531);
nand U41598 (N_41598,N_39743,N_38989);
nand U41599 (N_41599,N_37596,N_37635);
xor U41600 (N_41600,N_38143,N_38345);
nand U41601 (N_41601,N_38616,N_39464);
and U41602 (N_41602,N_39304,N_37963);
xor U41603 (N_41603,N_39828,N_38505);
nor U41604 (N_41604,N_38380,N_39607);
and U41605 (N_41605,N_37550,N_37675);
and U41606 (N_41606,N_37518,N_37988);
and U41607 (N_41607,N_39273,N_38001);
or U41608 (N_41608,N_38056,N_39467);
or U41609 (N_41609,N_38013,N_39996);
and U41610 (N_41610,N_37743,N_37994);
nor U41611 (N_41611,N_38203,N_38282);
nand U41612 (N_41612,N_38390,N_38089);
nor U41613 (N_41613,N_37773,N_39307);
nand U41614 (N_41614,N_38114,N_37691);
and U41615 (N_41615,N_38589,N_38110);
nor U41616 (N_41616,N_39845,N_38292);
nand U41617 (N_41617,N_39355,N_38615);
nor U41618 (N_41618,N_39066,N_38382);
xnor U41619 (N_41619,N_38717,N_39542);
or U41620 (N_41620,N_39656,N_39716);
nor U41621 (N_41621,N_39958,N_38763);
and U41622 (N_41622,N_39101,N_39282);
xnor U41623 (N_41623,N_38915,N_39483);
nor U41624 (N_41624,N_37563,N_39051);
or U41625 (N_41625,N_38210,N_37987);
and U41626 (N_41626,N_38155,N_39693);
nor U41627 (N_41627,N_37606,N_39383);
or U41628 (N_41628,N_39884,N_38893);
and U41629 (N_41629,N_38960,N_39459);
or U41630 (N_41630,N_38122,N_37901);
nor U41631 (N_41631,N_39734,N_38644);
and U41632 (N_41632,N_38416,N_38428);
nor U41633 (N_41633,N_38579,N_39805);
nor U41634 (N_41634,N_38855,N_38335);
nand U41635 (N_41635,N_38425,N_39740);
and U41636 (N_41636,N_38658,N_38969);
nor U41637 (N_41637,N_38522,N_38118);
xor U41638 (N_41638,N_39374,N_37793);
xnor U41639 (N_41639,N_39076,N_39661);
xor U41640 (N_41640,N_38044,N_37940);
nand U41641 (N_41641,N_38703,N_39308);
and U41642 (N_41642,N_38204,N_38259);
and U41643 (N_41643,N_38388,N_38906);
nor U41644 (N_41644,N_38048,N_39962);
xor U41645 (N_41645,N_38388,N_38873);
xnor U41646 (N_41646,N_38370,N_39298);
nand U41647 (N_41647,N_38974,N_38753);
nand U41648 (N_41648,N_39343,N_37912);
xnor U41649 (N_41649,N_38513,N_39341);
nand U41650 (N_41650,N_38255,N_39956);
and U41651 (N_41651,N_39263,N_39545);
nand U41652 (N_41652,N_39659,N_37831);
or U41653 (N_41653,N_39802,N_38002);
or U41654 (N_41654,N_39993,N_37641);
xor U41655 (N_41655,N_39426,N_38137);
and U41656 (N_41656,N_38037,N_39883);
or U41657 (N_41657,N_39315,N_37530);
nor U41658 (N_41658,N_39740,N_38121);
and U41659 (N_41659,N_39685,N_39999);
xor U41660 (N_41660,N_39510,N_39215);
xnor U41661 (N_41661,N_38946,N_38084);
xnor U41662 (N_41662,N_38326,N_38412);
and U41663 (N_41663,N_37758,N_39761);
nand U41664 (N_41664,N_38373,N_39913);
nand U41665 (N_41665,N_38541,N_37854);
nor U41666 (N_41666,N_39033,N_38497);
nand U41667 (N_41667,N_39900,N_37756);
and U41668 (N_41668,N_38944,N_38395);
and U41669 (N_41669,N_38271,N_38301);
nand U41670 (N_41670,N_39205,N_38418);
or U41671 (N_41671,N_39214,N_37703);
and U41672 (N_41672,N_38122,N_39698);
xnor U41673 (N_41673,N_39638,N_39021);
nor U41674 (N_41674,N_39680,N_38415);
and U41675 (N_41675,N_39468,N_39555);
nor U41676 (N_41676,N_38313,N_38027);
or U41677 (N_41677,N_37857,N_37627);
nand U41678 (N_41678,N_39661,N_39277);
xnor U41679 (N_41679,N_38161,N_38419);
nor U41680 (N_41680,N_38448,N_37905);
and U41681 (N_41681,N_39906,N_39013);
or U41682 (N_41682,N_39032,N_38916);
or U41683 (N_41683,N_39147,N_38324);
and U41684 (N_41684,N_37662,N_39154);
and U41685 (N_41685,N_38228,N_39945);
or U41686 (N_41686,N_37584,N_38737);
nand U41687 (N_41687,N_39090,N_38385);
nor U41688 (N_41688,N_38421,N_38573);
and U41689 (N_41689,N_38674,N_37581);
nor U41690 (N_41690,N_38061,N_39332);
nor U41691 (N_41691,N_39242,N_39337);
xor U41692 (N_41692,N_38414,N_39186);
or U41693 (N_41693,N_39465,N_39358);
nor U41694 (N_41694,N_38230,N_38162);
or U41695 (N_41695,N_39770,N_39785);
xor U41696 (N_41696,N_39890,N_37825);
nand U41697 (N_41697,N_38655,N_37981);
and U41698 (N_41698,N_39895,N_38422);
nand U41699 (N_41699,N_39551,N_38103);
xnor U41700 (N_41700,N_37599,N_39823);
nand U41701 (N_41701,N_38366,N_38685);
nor U41702 (N_41702,N_39171,N_39097);
and U41703 (N_41703,N_39772,N_38254);
nand U41704 (N_41704,N_38811,N_37985);
xor U41705 (N_41705,N_37837,N_38993);
nand U41706 (N_41706,N_37771,N_39060);
nor U41707 (N_41707,N_37679,N_38192);
xnor U41708 (N_41708,N_37902,N_39048);
or U41709 (N_41709,N_38271,N_38455);
nand U41710 (N_41710,N_37898,N_37851);
nand U41711 (N_41711,N_38458,N_39777);
and U41712 (N_41712,N_37858,N_39506);
or U41713 (N_41713,N_38473,N_38978);
or U41714 (N_41714,N_38634,N_38233);
and U41715 (N_41715,N_38236,N_38789);
and U41716 (N_41716,N_39933,N_39261);
nand U41717 (N_41717,N_37792,N_37610);
nor U41718 (N_41718,N_39040,N_39298);
xor U41719 (N_41719,N_39552,N_38840);
and U41720 (N_41720,N_37843,N_37855);
nor U41721 (N_41721,N_39388,N_38595);
or U41722 (N_41722,N_39013,N_38198);
or U41723 (N_41723,N_37692,N_39359);
xor U41724 (N_41724,N_39779,N_39420);
nor U41725 (N_41725,N_39831,N_37500);
or U41726 (N_41726,N_39786,N_39774);
nor U41727 (N_41727,N_38180,N_39859);
and U41728 (N_41728,N_39069,N_39164);
nand U41729 (N_41729,N_38282,N_38689);
nand U41730 (N_41730,N_39345,N_39896);
nand U41731 (N_41731,N_38722,N_39194);
nand U41732 (N_41732,N_38226,N_38138);
or U41733 (N_41733,N_37934,N_39801);
xor U41734 (N_41734,N_39035,N_38122);
and U41735 (N_41735,N_39107,N_39181);
and U41736 (N_41736,N_37717,N_37596);
xor U41737 (N_41737,N_39416,N_39486);
nand U41738 (N_41738,N_38785,N_39024);
nand U41739 (N_41739,N_39631,N_37544);
nor U41740 (N_41740,N_39872,N_39056);
xnor U41741 (N_41741,N_38785,N_38930);
or U41742 (N_41742,N_39707,N_37771);
xor U41743 (N_41743,N_39687,N_38736);
nor U41744 (N_41744,N_37608,N_39841);
nand U41745 (N_41745,N_39451,N_37955);
or U41746 (N_41746,N_39552,N_39794);
and U41747 (N_41747,N_38348,N_39811);
or U41748 (N_41748,N_38409,N_39610);
nor U41749 (N_41749,N_38863,N_38001);
xnor U41750 (N_41750,N_39610,N_39240);
nor U41751 (N_41751,N_38561,N_38743);
nand U41752 (N_41752,N_38517,N_37675);
nand U41753 (N_41753,N_38554,N_39311);
and U41754 (N_41754,N_37949,N_37616);
nand U41755 (N_41755,N_39934,N_38412);
and U41756 (N_41756,N_39908,N_37562);
nand U41757 (N_41757,N_39021,N_37816);
xor U41758 (N_41758,N_37966,N_38282);
nand U41759 (N_41759,N_39609,N_38722);
or U41760 (N_41760,N_37783,N_38534);
nand U41761 (N_41761,N_39183,N_38035);
xor U41762 (N_41762,N_37677,N_38615);
and U41763 (N_41763,N_37792,N_38643);
nand U41764 (N_41764,N_38187,N_37882);
or U41765 (N_41765,N_39855,N_38269);
xor U41766 (N_41766,N_38957,N_39294);
or U41767 (N_41767,N_39379,N_38964);
nand U41768 (N_41768,N_38189,N_38539);
nor U41769 (N_41769,N_38302,N_39064);
or U41770 (N_41770,N_37669,N_39251);
and U41771 (N_41771,N_38018,N_38115);
or U41772 (N_41772,N_37784,N_37938);
nor U41773 (N_41773,N_37881,N_38907);
xor U41774 (N_41774,N_39778,N_39195);
xor U41775 (N_41775,N_38023,N_38770);
or U41776 (N_41776,N_39310,N_38032);
nand U41777 (N_41777,N_39281,N_37677);
or U41778 (N_41778,N_38735,N_39475);
and U41779 (N_41779,N_38530,N_39970);
nand U41780 (N_41780,N_38231,N_38166);
or U41781 (N_41781,N_39351,N_38740);
nand U41782 (N_41782,N_38208,N_37510);
nand U41783 (N_41783,N_38998,N_37976);
or U41784 (N_41784,N_38419,N_37688);
or U41785 (N_41785,N_38199,N_39137);
nand U41786 (N_41786,N_39996,N_39969);
xnor U41787 (N_41787,N_38553,N_39531);
nor U41788 (N_41788,N_39063,N_38636);
xnor U41789 (N_41789,N_38540,N_39588);
nand U41790 (N_41790,N_39560,N_38860);
xnor U41791 (N_41791,N_39108,N_38336);
xor U41792 (N_41792,N_37549,N_39431);
xor U41793 (N_41793,N_39235,N_39869);
xor U41794 (N_41794,N_38048,N_38176);
nand U41795 (N_41795,N_37680,N_38109);
or U41796 (N_41796,N_38715,N_39151);
or U41797 (N_41797,N_38748,N_39723);
nor U41798 (N_41798,N_39551,N_38619);
nor U41799 (N_41799,N_38437,N_39916);
nor U41800 (N_41800,N_38659,N_38689);
xor U41801 (N_41801,N_38342,N_39222);
and U41802 (N_41802,N_37763,N_38249);
nor U41803 (N_41803,N_38377,N_39861);
xnor U41804 (N_41804,N_38622,N_39382);
nor U41805 (N_41805,N_38489,N_39120);
xnor U41806 (N_41806,N_38239,N_38929);
nand U41807 (N_41807,N_37745,N_38056);
xor U41808 (N_41808,N_39645,N_38997);
or U41809 (N_41809,N_38000,N_37550);
and U41810 (N_41810,N_38279,N_38355);
xor U41811 (N_41811,N_39797,N_39280);
or U41812 (N_41812,N_39500,N_38504);
or U41813 (N_41813,N_39239,N_37947);
and U41814 (N_41814,N_37618,N_39800);
xor U41815 (N_41815,N_37692,N_37562);
nand U41816 (N_41816,N_39438,N_39179);
nand U41817 (N_41817,N_38609,N_38487);
nand U41818 (N_41818,N_38328,N_38776);
or U41819 (N_41819,N_38259,N_39524);
xor U41820 (N_41820,N_38209,N_38122);
or U41821 (N_41821,N_39361,N_38649);
nor U41822 (N_41822,N_38150,N_39285);
nand U41823 (N_41823,N_39439,N_39108);
nand U41824 (N_41824,N_38639,N_38270);
and U41825 (N_41825,N_38088,N_37955);
xnor U41826 (N_41826,N_38926,N_38022);
nand U41827 (N_41827,N_39284,N_39183);
nand U41828 (N_41828,N_38580,N_39417);
nand U41829 (N_41829,N_39150,N_39557);
nor U41830 (N_41830,N_37744,N_38740);
nand U41831 (N_41831,N_37749,N_38049);
nor U41832 (N_41832,N_37987,N_39445);
nor U41833 (N_41833,N_38212,N_39531);
nor U41834 (N_41834,N_39471,N_39964);
nor U41835 (N_41835,N_39437,N_38061);
xnor U41836 (N_41836,N_37957,N_38255);
nor U41837 (N_41837,N_37766,N_38188);
nor U41838 (N_41838,N_38963,N_38581);
nand U41839 (N_41839,N_39053,N_38683);
nand U41840 (N_41840,N_39246,N_38033);
xnor U41841 (N_41841,N_38269,N_39344);
xnor U41842 (N_41842,N_37540,N_39876);
xnor U41843 (N_41843,N_37697,N_38654);
nor U41844 (N_41844,N_39159,N_37862);
xor U41845 (N_41845,N_38706,N_38919);
nand U41846 (N_41846,N_37832,N_38793);
xor U41847 (N_41847,N_38773,N_37984);
nand U41848 (N_41848,N_37561,N_39732);
or U41849 (N_41849,N_39818,N_37711);
or U41850 (N_41850,N_38126,N_37562);
or U41851 (N_41851,N_38891,N_39614);
and U41852 (N_41852,N_39264,N_38413);
nor U41853 (N_41853,N_38235,N_38609);
or U41854 (N_41854,N_39379,N_38500);
xor U41855 (N_41855,N_38785,N_39794);
xnor U41856 (N_41856,N_37509,N_38031);
and U41857 (N_41857,N_39112,N_39153);
xnor U41858 (N_41858,N_39963,N_38942);
nand U41859 (N_41859,N_38753,N_37898);
and U41860 (N_41860,N_39239,N_38781);
nand U41861 (N_41861,N_39767,N_38890);
or U41862 (N_41862,N_38669,N_37954);
nor U41863 (N_41863,N_39669,N_39012);
nor U41864 (N_41864,N_39185,N_39511);
or U41865 (N_41865,N_39715,N_37562);
nand U41866 (N_41866,N_37899,N_38653);
nand U41867 (N_41867,N_38098,N_39178);
nand U41868 (N_41868,N_39428,N_39607);
or U41869 (N_41869,N_37699,N_37753);
or U41870 (N_41870,N_37908,N_39643);
xor U41871 (N_41871,N_37533,N_38472);
nor U41872 (N_41872,N_38168,N_37936);
xor U41873 (N_41873,N_39228,N_37508);
nand U41874 (N_41874,N_38217,N_38690);
nor U41875 (N_41875,N_38699,N_37973);
nand U41876 (N_41876,N_39060,N_38080);
and U41877 (N_41877,N_38654,N_37911);
or U41878 (N_41878,N_39670,N_38065);
nor U41879 (N_41879,N_38679,N_37635);
nand U41880 (N_41880,N_39440,N_39041);
nand U41881 (N_41881,N_39546,N_38774);
or U41882 (N_41882,N_37838,N_39202);
nor U41883 (N_41883,N_39296,N_37594);
xor U41884 (N_41884,N_39698,N_37925);
and U41885 (N_41885,N_37637,N_39032);
xor U41886 (N_41886,N_37590,N_38905);
nand U41887 (N_41887,N_37579,N_39680);
xor U41888 (N_41888,N_37905,N_38328);
nand U41889 (N_41889,N_39107,N_37993);
nand U41890 (N_41890,N_39841,N_39130);
or U41891 (N_41891,N_37866,N_37548);
and U41892 (N_41892,N_38853,N_38264);
xor U41893 (N_41893,N_39244,N_39599);
and U41894 (N_41894,N_39245,N_39066);
and U41895 (N_41895,N_38248,N_38898);
nand U41896 (N_41896,N_38056,N_38155);
or U41897 (N_41897,N_39660,N_38327);
and U41898 (N_41898,N_38029,N_39202);
or U41899 (N_41899,N_37875,N_37862);
and U41900 (N_41900,N_37788,N_38634);
and U41901 (N_41901,N_38683,N_37827);
nor U41902 (N_41902,N_38816,N_39356);
and U41903 (N_41903,N_37763,N_37910);
and U41904 (N_41904,N_38362,N_37521);
nand U41905 (N_41905,N_39033,N_38969);
nand U41906 (N_41906,N_38736,N_39287);
and U41907 (N_41907,N_38465,N_38090);
nor U41908 (N_41908,N_39636,N_38990);
and U41909 (N_41909,N_37771,N_37658);
nand U41910 (N_41910,N_39129,N_38237);
nor U41911 (N_41911,N_39182,N_38050);
and U41912 (N_41912,N_37775,N_39992);
nor U41913 (N_41913,N_37598,N_38286);
or U41914 (N_41914,N_37896,N_37802);
nor U41915 (N_41915,N_37735,N_39118);
and U41916 (N_41916,N_37524,N_39190);
nor U41917 (N_41917,N_39495,N_38072);
or U41918 (N_41918,N_38684,N_39947);
or U41919 (N_41919,N_38750,N_37795);
nor U41920 (N_41920,N_39599,N_38015);
nand U41921 (N_41921,N_39576,N_39581);
or U41922 (N_41922,N_39950,N_38664);
or U41923 (N_41923,N_37535,N_38132);
xnor U41924 (N_41924,N_39860,N_37823);
and U41925 (N_41925,N_38808,N_39742);
nor U41926 (N_41926,N_39677,N_37609);
or U41927 (N_41927,N_38085,N_39592);
and U41928 (N_41928,N_39867,N_37849);
nor U41929 (N_41929,N_39364,N_39063);
nor U41930 (N_41930,N_39332,N_38574);
or U41931 (N_41931,N_39366,N_38979);
xnor U41932 (N_41932,N_38370,N_37576);
or U41933 (N_41933,N_38825,N_38364);
or U41934 (N_41934,N_39702,N_39739);
xnor U41935 (N_41935,N_39404,N_37884);
nor U41936 (N_41936,N_39325,N_37665);
nand U41937 (N_41937,N_39890,N_39249);
nor U41938 (N_41938,N_39054,N_38044);
or U41939 (N_41939,N_37654,N_38156);
or U41940 (N_41940,N_39785,N_38894);
or U41941 (N_41941,N_38955,N_37532);
nand U41942 (N_41942,N_39460,N_39602);
and U41943 (N_41943,N_39657,N_37955);
xor U41944 (N_41944,N_38109,N_38410);
nor U41945 (N_41945,N_38250,N_39257);
or U41946 (N_41946,N_39546,N_37603);
nand U41947 (N_41947,N_38684,N_38445);
nand U41948 (N_41948,N_37808,N_38625);
and U41949 (N_41949,N_39029,N_38396);
nor U41950 (N_41950,N_38622,N_37971);
or U41951 (N_41951,N_37910,N_38308);
nand U41952 (N_41952,N_37587,N_39892);
xnor U41953 (N_41953,N_38014,N_39588);
or U41954 (N_41954,N_38921,N_38603);
nand U41955 (N_41955,N_39721,N_39988);
nand U41956 (N_41956,N_38802,N_38793);
or U41957 (N_41957,N_39098,N_37526);
and U41958 (N_41958,N_38860,N_37843);
and U41959 (N_41959,N_37984,N_39527);
or U41960 (N_41960,N_39885,N_38916);
and U41961 (N_41961,N_38314,N_39140);
nor U41962 (N_41962,N_38564,N_37741);
xnor U41963 (N_41963,N_39582,N_37624);
nor U41964 (N_41964,N_39178,N_38281);
nor U41965 (N_41965,N_38150,N_38660);
and U41966 (N_41966,N_38932,N_39962);
nand U41967 (N_41967,N_38264,N_39018);
or U41968 (N_41968,N_39803,N_39675);
and U41969 (N_41969,N_39409,N_39636);
nand U41970 (N_41970,N_39359,N_39498);
nor U41971 (N_41971,N_39652,N_39295);
and U41972 (N_41972,N_39325,N_37506);
xor U41973 (N_41973,N_39545,N_39214);
and U41974 (N_41974,N_39346,N_39125);
nor U41975 (N_41975,N_39803,N_37861);
nand U41976 (N_41976,N_39536,N_38504);
nand U41977 (N_41977,N_37566,N_39081);
or U41978 (N_41978,N_38909,N_38351);
nor U41979 (N_41979,N_39866,N_39795);
or U41980 (N_41980,N_38601,N_38117);
nor U41981 (N_41981,N_39853,N_37972);
or U41982 (N_41982,N_37717,N_39305);
xnor U41983 (N_41983,N_38519,N_38445);
nor U41984 (N_41984,N_39168,N_37889);
nand U41985 (N_41985,N_38193,N_38903);
nand U41986 (N_41986,N_39460,N_38505);
xor U41987 (N_41987,N_39836,N_37714);
or U41988 (N_41988,N_39126,N_39559);
xor U41989 (N_41989,N_39641,N_39217);
and U41990 (N_41990,N_39579,N_39456);
and U41991 (N_41991,N_39408,N_38598);
nand U41992 (N_41992,N_37924,N_37986);
nand U41993 (N_41993,N_37888,N_37648);
nand U41994 (N_41994,N_38642,N_38636);
nor U41995 (N_41995,N_39263,N_38307);
xor U41996 (N_41996,N_38951,N_38909);
or U41997 (N_41997,N_37715,N_37543);
nor U41998 (N_41998,N_38282,N_39786);
nand U41999 (N_41999,N_37800,N_37603);
nor U42000 (N_42000,N_37936,N_39293);
nand U42001 (N_42001,N_38627,N_37593);
or U42002 (N_42002,N_37720,N_39042);
and U42003 (N_42003,N_38183,N_39008);
nor U42004 (N_42004,N_38886,N_39215);
nor U42005 (N_42005,N_38190,N_38188);
xnor U42006 (N_42006,N_38656,N_38053);
nor U42007 (N_42007,N_37845,N_39964);
xnor U42008 (N_42008,N_39168,N_38566);
and U42009 (N_42009,N_39101,N_38987);
and U42010 (N_42010,N_38301,N_38203);
and U42011 (N_42011,N_38872,N_38303);
nand U42012 (N_42012,N_39848,N_38639);
nor U42013 (N_42013,N_38761,N_39054);
xnor U42014 (N_42014,N_38986,N_38264);
or U42015 (N_42015,N_38294,N_39195);
and U42016 (N_42016,N_39619,N_39909);
and U42017 (N_42017,N_39350,N_39529);
and U42018 (N_42018,N_37930,N_39048);
or U42019 (N_42019,N_39682,N_38773);
nand U42020 (N_42020,N_37869,N_39947);
nor U42021 (N_42021,N_37773,N_39397);
and U42022 (N_42022,N_39736,N_39983);
nand U42023 (N_42023,N_39645,N_38363);
and U42024 (N_42024,N_39133,N_39527);
and U42025 (N_42025,N_39189,N_37626);
xnor U42026 (N_42026,N_38180,N_38701);
nor U42027 (N_42027,N_39359,N_37817);
xor U42028 (N_42028,N_37604,N_39954);
nor U42029 (N_42029,N_38608,N_38827);
or U42030 (N_42030,N_37684,N_37784);
xor U42031 (N_42031,N_38772,N_37611);
and U42032 (N_42032,N_39928,N_38618);
nor U42033 (N_42033,N_39047,N_37928);
or U42034 (N_42034,N_37746,N_39844);
and U42035 (N_42035,N_38854,N_38672);
or U42036 (N_42036,N_38611,N_38560);
or U42037 (N_42037,N_38294,N_38232);
nor U42038 (N_42038,N_39714,N_39022);
or U42039 (N_42039,N_39370,N_39425);
nand U42040 (N_42040,N_39903,N_39016);
nand U42041 (N_42041,N_39513,N_37840);
or U42042 (N_42042,N_38749,N_39893);
and U42043 (N_42043,N_39931,N_39325);
xnor U42044 (N_42044,N_38064,N_38789);
and U42045 (N_42045,N_39184,N_39338);
nand U42046 (N_42046,N_39405,N_38311);
nand U42047 (N_42047,N_38292,N_38109);
xnor U42048 (N_42048,N_39449,N_38522);
xnor U42049 (N_42049,N_38435,N_38594);
xor U42050 (N_42050,N_38743,N_39028);
or U42051 (N_42051,N_39419,N_37773);
or U42052 (N_42052,N_38942,N_37968);
or U42053 (N_42053,N_37926,N_38166);
nor U42054 (N_42054,N_37506,N_38325);
xor U42055 (N_42055,N_39625,N_38690);
and U42056 (N_42056,N_39998,N_38451);
nor U42057 (N_42057,N_39410,N_39219);
xnor U42058 (N_42058,N_38552,N_39868);
nand U42059 (N_42059,N_37568,N_38325);
or U42060 (N_42060,N_39318,N_37866);
and U42061 (N_42061,N_38370,N_37642);
nor U42062 (N_42062,N_39944,N_39601);
or U42063 (N_42063,N_38589,N_38199);
or U42064 (N_42064,N_37805,N_38033);
xnor U42065 (N_42065,N_38148,N_39427);
nand U42066 (N_42066,N_39777,N_39955);
and U42067 (N_42067,N_38655,N_38644);
and U42068 (N_42068,N_37970,N_37810);
and U42069 (N_42069,N_37516,N_38002);
nor U42070 (N_42070,N_38548,N_38938);
xnor U42071 (N_42071,N_38486,N_39399);
or U42072 (N_42072,N_39829,N_39526);
and U42073 (N_42073,N_38793,N_38700);
nor U42074 (N_42074,N_39039,N_37862);
nor U42075 (N_42075,N_39531,N_38543);
xor U42076 (N_42076,N_38293,N_39622);
nand U42077 (N_42077,N_37722,N_38609);
xor U42078 (N_42078,N_39233,N_39306);
nand U42079 (N_42079,N_38029,N_39959);
or U42080 (N_42080,N_39115,N_38060);
and U42081 (N_42081,N_39765,N_39409);
nand U42082 (N_42082,N_37814,N_39694);
nor U42083 (N_42083,N_39418,N_37826);
and U42084 (N_42084,N_38734,N_38065);
or U42085 (N_42085,N_37820,N_39130);
and U42086 (N_42086,N_38831,N_39036);
and U42087 (N_42087,N_39484,N_39816);
xnor U42088 (N_42088,N_39360,N_39555);
or U42089 (N_42089,N_38812,N_39444);
nand U42090 (N_42090,N_39563,N_38026);
or U42091 (N_42091,N_38014,N_38202);
nand U42092 (N_42092,N_38032,N_38742);
and U42093 (N_42093,N_39257,N_37786);
nand U42094 (N_42094,N_39685,N_38777);
xor U42095 (N_42095,N_39039,N_38658);
or U42096 (N_42096,N_38896,N_37724);
and U42097 (N_42097,N_37898,N_37732);
or U42098 (N_42098,N_38061,N_39501);
xor U42099 (N_42099,N_38787,N_38224);
nor U42100 (N_42100,N_37618,N_38480);
and U42101 (N_42101,N_39023,N_37934);
and U42102 (N_42102,N_37960,N_39019);
nand U42103 (N_42103,N_38288,N_37874);
nor U42104 (N_42104,N_37765,N_39254);
xor U42105 (N_42105,N_38822,N_39853);
and U42106 (N_42106,N_39445,N_39719);
xor U42107 (N_42107,N_39345,N_39304);
xor U42108 (N_42108,N_38974,N_38711);
xnor U42109 (N_42109,N_38228,N_39250);
or U42110 (N_42110,N_39851,N_39091);
or U42111 (N_42111,N_38235,N_37623);
nand U42112 (N_42112,N_38925,N_38115);
nor U42113 (N_42113,N_38173,N_39002);
nor U42114 (N_42114,N_39632,N_38504);
and U42115 (N_42115,N_39941,N_38934);
nor U42116 (N_42116,N_39595,N_39417);
and U42117 (N_42117,N_38717,N_38361);
nand U42118 (N_42118,N_39695,N_38179);
or U42119 (N_42119,N_38886,N_38713);
or U42120 (N_42120,N_38622,N_37741);
nor U42121 (N_42121,N_39521,N_38110);
xnor U42122 (N_42122,N_39813,N_38637);
xor U42123 (N_42123,N_39251,N_39403);
nor U42124 (N_42124,N_38699,N_39733);
and U42125 (N_42125,N_39777,N_39182);
xnor U42126 (N_42126,N_39026,N_39483);
and U42127 (N_42127,N_39009,N_38345);
nor U42128 (N_42128,N_39691,N_37768);
nand U42129 (N_42129,N_38707,N_38475);
nor U42130 (N_42130,N_39944,N_39147);
and U42131 (N_42131,N_39877,N_39855);
xnor U42132 (N_42132,N_38080,N_39473);
nand U42133 (N_42133,N_38280,N_39404);
xnor U42134 (N_42134,N_39782,N_39806);
and U42135 (N_42135,N_37927,N_39049);
xor U42136 (N_42136,N_38360,N_37942);
xnor U42137 (N_42137,N_39534,N_39936);
or U42138 (N_42138,N_39946,N_37951);
or U42139 (N_42139,N_37756,N_38713);
nor U42140 (N_42140,N_38617,N_38207);
xnor U42141 (N_42141,N_37829,N_39331);
xnor U42142 (N_42142,N_39986,N_39156);
xnor U42143 (N_42143,N_39915,N_38311);
xnor U42144 (N_42144,N_37689,N_39613);
or U42145 (N_42145,N_38052,N_38586);
and U42146 (N_42146,N_39378,N_39836);
and U42147 (N_42147,N_38972,N_38181);
and U42148 (N_42148,N_39616,N_38606);
or U42149 (N_42149,N_38881,N_38907);
xor U42150 (N_42150,N_39176,N_37555);
xnor U42151 (N_42151,N_39884,N_39825);
and U42152 (N_42152,N_38092,N_39446);
xor U42153 (N_42153,N_38328,N_37684);
and U42154 (N_42154,N_39690,N_38420);
and U42155 (N_42155,N_39060,N_37844);
or U42156 (N_42156,N_39363,N_38702);
nor U42157 (N_42157,N_39773,N_38495);
nand U42158 (N_42158,N_38756,N_39421);
and U42159 (N_42159,N_39197,N_38906);
and U42160 (N_42160,N_39461,N_37666);
nand U42161 (N_42161,N_39011,N_38052);
nor U42162 (N_42162,N_39570,N_39381);
nor U42163 (N_42163,N_37603,N_39131);
or U42164 (N_42164,N_37712,N_39732);
xor U42165 (N_42165,N_39671,N_38315);
nand U42166 (N_42166,N_38883,N_39486);
nor U42167 (N_42167,N_39221,N_38041);
nor U42168 (N_42168,N_38879,N_39872);
and U42169 (N_42169,N_39218,N_38906);
nor U42170 (N_42170,N_39347,N_39503);
or U42171 (N_42171,N_38623,N_37857);
nand U42172 (N_42172,N_38062,N_38668);
xnor U42173 (N_42173,N_38147,N_38440);
xor U42174 (N_42174,N_38438,N_39547);
and U42175 (N_42175,N_39169,N_37663);
nor U42176 (N_42176,N_37791,N_38144);
xor U42177 (N_42177,N_37673,N_39377);
and U42178 (N_42178,N_38308,N_39751);
xor U42179 (N_42179,N_38777,N_38386);
nand U42180 (N_42180,N_38398,N_39456);
xor U42181 (N_42181,N_37557,N_39881);
nand U42182 (N_42182,N_39503,N_38523);
and U42183 (N_42183,N_38948,N_37886);
xnor U42184 (N_42184,N_38400,N_38259);
and U42185 (N_42185,N_39267,N_38835);
nor U42186 (N_42186,N_39539,N_39118);
or U42187 (N_42187,N_38232,N_38169);
nand U42188 (N_42188,N_37504,N_38649);
xnor U42189 (N_42189,N_37965,N_38464);
or U42190 (N_42190,N_38100,N_38846);
nor U42191 (N_42191,N_38230,N_37829);
or U42192 (N_42192,N_39251,N_39761);
and U42193 (N_42193,N_39003,N_37715);
and U42194 (N_42194,N_38683,N_38034);
or U42195 (N_42195,N_37947,N_37943);
nor U42196 (N_42196,N_39707,N_38320);
nand U42197 (N_42197,N_37555,N_38944);
nand U42198 (N_42198,N_39235,N_38792);
or U42199 (N_42199,N_39954,N_38136);
xor U42200 (N_42200,N_38464,N_37741);
nor U42201 (N_42201,N_39544,N_38484);
nand U42202 (N_42202,N_39347,N_37544);
xor U42203 (N_42203,N_38087,N_37990);
xor U42204 (N_42204,N_39503,N_37916);
nand U42205 (N_42205,N_39158,N_39498);
xor U42206 (N_42206,N_39801,N_39457);
nand U42207 (N_42207,N_38108,N_39144);
nand U42208 (N_42208,N_39728,N_39304);
nand U42209 (N_42209,N_37996,N_38345);
xnor U42210 (N_42210,N_39623,N_39246);
and U42211 (N_42211,N_37952,N_39704);
nor U42212 (N_42212,N_38873,N_37662);
xnor U42213 (N_42213,N_39532,N_39246);
nand U42214 (N_42214,N_37678,N_38197);
nor U42215 (N_42215,N_37589,N_39198);
xnor U42216 (N_42216,N_38810,N_39881);
or U42217 (N_42217,N_38018,N_37555);
and U42218 (N_42218,N_38345,N_38887);
nor U42219 (N_42219,N_39760,N_38035);
nand U42220 (N_42220,N_37760,N_39192);
nand U42221 (N_42221,N_39822,N_38066);
and U42222 (N_42222,N_37956,N_38809);
nand U42223 (N_42223,N_37621,N_38917);
or U42224 (N_42224,N_39703,N_39200);
nor U42225 (N_42225,N_38035,N_38412);
nand U42226 (N_42226,N_38611,N_38930);
xor U42227 (N_42227,N_37557,N_38950);
and U42228 (N_42228,N_39670,N_37994);
or U42229 (N_42229,N_39825,N_39028);
nor U42230 (N_42230,N_37622,N_37723);
nor U42231 (N_42231,N_38542,N_38150);
nand U42232 (N_42232,N_37517,N_39569);
xnor U42233 (N_42233,N_39132,N_38869);
nand U42234 (N_42234,N_39874,N_37820);
or U42235 (N_42235,N_38858,N_39945);
xor U42236 (N_42236,N_39030,N_38471);
nand U42237 (N_42237,N_39560,N_39881);
xnor U42238 (N_42238,N_39949,N_38954);
and U42239 (N_42239,N_38363,N_37517);
or U42240 (N_42240,N_39028,N_38067);
nand U42241 (N_42241,N_38988,N_39914);
xor U42242 (N_42242,N_38095,N_39122);
or U42243 (N_42243,N_38870,N_37960);
or U42244 (N_42244,N_39440,N_39821);
nand U42245 (N_42245,N_38293,N_38837);
and U42246 (N_42246,N_39171,N_39380);
xnor U42247 (N_42247,N_39729,N_38250);
and U42248 (N_42248,N_38197,N_38003);
nand U42249 (N_42249,N_37723,N_38474);
and U42250 (N_42250,N_39164,N_39259);
and U42251 (N_42251,N_39203,N_39188);
or U42252 (N_42252,N_37866,N_38107);
xor U42253 (N_42253,N_38316,N_37531);
nor U42254 (N_42254,N_38850,N_38607);
xnor U42255 (N_42255,N_38169,N_39554);
and U42256 (N_42256,N_38197,N_38486);
xor U42257 (N_42257,N_38056,N_37684);
xor U42258 (N_42258,N_37649,N_39634);
nor U42259 (N_42259,N_37740,N_38029);
nor U42260 (N_42260,N_39832,N_37697);
nand U42261 (N_42261,N_38859,N_37945);
and U42262 (N_42262,N_39501,N_39338);
and U42263 (N_42263,N_38511,N_37713);
nor U42264 (N_42264,N_38753,N_39622);
and U42265 (N_42265,N_38991,N_37992);
or U42266 (N_42266,N_38336,N_38189);
nand U42267 (N_42267,N_38641,N_39872);
nor U42268 (N_42268,N_39131,N_38314);
nor U42269 (N_42269,N_38630,N_37695);
or U42270 (N_42270,N_38913,N_38567);
and U42271 (N_42271,N_39090,N_38009);
nand U42272 (N_42272,N_37630,N_38913);
and U42273 (N_42273,N_38353,N_37926);
or U42274 (N_42274,N_38682,N_38446);
nand U42275 (N_42275,N_38314,N_38344);
or U42276 (N_42276,N_39406,N_38429);
xnor U42277 (N_42277,N_38188,N_38348);
nor U42278 (N_42278,N_39456,N_39924);
xor U42279 (N_42279,N_38555,N_38779);
or U42280 (N_42280,N_37664,N_38665);
or U42281 (N_42281,N_37955,N_38113);
nand U42282 (N_42282,N_37620,N_39180);
and U42283 (N_42283,N_39106,N_38889);
or U42284 (N_42284,N_39465,N_38597);
xor U42285 (N_42285,N_38142,N_38599);
nor U42286 (N_42286,N_39727,N_38337);
nand U42287 (N_42287,N_39393,N_38164);
or U42288 (N_42288,N_38290,N_38007);
nor U42289 (N_42289,N_39742,N_38910);
nor U42290 (N_42290,N_38984,N_38865);
nor U42291 (N_42291,N_39723,N_38209);
xnor U42292 (N_42292,N_39902,N_39188);
and U42293 (N_42293,N_38251,N_39407);
and U42294 (N_42294,N_39271,N_38044);
nand U42295 (N_42295,N_38088,N_37533);
and U42296 (N_42296,N_39650,N_38528);
xor U42297 (N_42297,N_38203,N_39763);
and U42298 (N_42298,N_39699,N_37653);
nor U42299 (N_42299,N_37614,N_37934);
nor U42300 (N_42300,N_39314,N_38266);
nand U42301 (N_42301,N_39717,N_38684);
or U42302 (N_42302,N_38438,N_39761);
nand U42303 (N_42303,N_38329,N_38424);
xnor U42304 (N_42304,N_38521,N_38057);
nor U42305 (N_42305,N_38058,N_38677);
and U42306 (N_42306,N_38019,N_39720);
or U42307 (N_42307,N_39665,N_38617);
xor U42308 (N_42308,N_39897,N_38374);
xnor U42309 (N_42309,N_38031,N_39208);
nor U42310 (N_42310,N_38258,N_39353);
nand U42311 (N_42311,N_38261,N_39190);
and U42312 (N_42312,N_39260,N_38046);
and U42313 (N_42313,N_39572,N_37591);
xor U42314 (N_42314,N_39569,N_37643);
nor U42315 (N_42315,N_39803,N_39120);
nor U42316 (N_42316,N_38504,N_38806);
and U42317 (N_42317,N_39159,N_39343);
xnor U42318 (N_42318,N_38119,N_38684);
nor U42319 (N_42319,N_38050,N_37872);
nor U42320 (N_42320,N_38065,N_38000);
nand U42321 (N_42321,N_39112,N_39121);
nor U42322 (N_42322,N_38823,N_39690);
nand U42323 (N_42323,N_39812,N_37765);
xnor U42324 (N_42324,N_38269,N_37530);
nor U42325 (N_42325,N_38459,N_39868);
nand U42326 (N_42326,N_39251,N_39664);
or U42327 (N_42327,N_38161,N_38633);
and U42328 (N_42328,N_38289,N_38398);
nand U42329 (N_42329,N_38163,N_38641);
or U42330 (N_42330,N_39149,N_38867);
xor U42331 (N_42331,N_38765,N_38957);
and U42332 (N_42332,N_38315,N_38215);
nand U42333 (N_42333,N_39368,N_39451);
nand U42334 (N_42334,N_39180,N_39484);
and U42335 (N_42335,N_39179,N_38404);
nor U42336 (N_42336,N_38353,N_38882);
nor U42337 (N_42337,N_38883,N_37934);
xor U42338 (N_42338,N_38131,N_37716);
nor U42339 (N_42339,N_38087,N_38513);
or U42340 (N_42340,N_39509,N_37537);
and U42341 (N_42341,N_39823,N_38484);
nand U42342 (N_42342,N_38106,N_39278);
nand U42343 (N_42343,N_39983,N_39688);
nand U42344 (N_42344,N_38362,N_38957);
nor U42345 (N_42345,N_37591,N_39426);
nor U42346 (N_42346,N_38918,N_39979);
xnor U42347 (N_42347,N_38243,N_39121);
and U42348 (N_42348,N_39769,N_37651);
nor U42349 (N_42349,N_38501,N_37572);
or U42350 (N_42350,N_38867,N_37712);
xor U42351 (N_42351,N_37943,N_39528);
xnor U42352 (N_42352,N_38169,N_39427);
and U42353 (N_42353,N_39579,N_38420);
nand U42354 (N_42354,N_39917,N_38707);
xor U42355 (N_42355,N_37930,N_38479);
nand U42356 (N_42356,N_39763,N_38082);
and U42357 (N_42357,N_39002,N_38013);
and U42358 (N_42358,N_39920,N_39094);
nor U42359 (N_42359,N_38209,N_38581);
nand U42360 (N_42360,N_37937,N_39690);
xnor U42361 (N_42361,N_38221,N_38605);
nor U42362 (N_42362,N_38678,N_39515);
xor U42363 (N_42363,N_38747,N_38727);
nand U42364 (N_42364,N_38836,N_37542);
and U42365 (N_42365,N_38268,N_38660);
and U42366 (N_42366,N_38599,N_38221);
nor U42367 (N_42367,N_37540,N_37597);
xnor U42368 (N_42368,N_38300,N_39096);
or U42369 (N_42369,N_38796,N_39507);
and U42370 (N_42370,N_38668,N_38506);
or U42371 (N_42371,N_38740,N_37805);
and U42372 (N_42372,N_39137,N_37614);
xnor U42373 (N_42373,N_38785,N_39733);
nand U42374 (N_42374,N_37969,N_39759);
xnor U42375 (N_42375,N_39654,N_39410);
or U42376 (N_42376,N_39869,N_38321);
or U42377 (N_42377,N_38988,N_39541);
nor U42378 (N_42378,N_39253,N_37571);
xnor U42379 (N_42379,N_39475,N_39626);
nand U42380 (N_42380,N_38403,N_38605);
xor U42381 (N_42381,N_37974,N_38645);
nand U42382 (N_42382,N_38701,N_39559);
nor U42383 (N_42383,N_38422,N_38987);
xnor U42384 (N_42384,N_37926,N_39080);
nand U42385 (N_42385,N_38763,N_37517);
nor U42386 (N_42386,N_39557,N_39889);
or U42387 (N_42387,N_38501,N_39115);
nor U42388 (N_42388,N_38158,N_39469);
nand U42389 (N_42389,N_37840,N_39745);
and U42390 (N_42390,N_38352,N_38728);
xor U42391 (N_42391,N_37584,N_38134);
and U42392 (N_42392,N_38774,N_37936);
xnor U42393 (N_42393,N_38762,N_37541);
nand U42394 (N_42394,N_39671,N_39964);
nand U42395 (N_42395,N_38726,N_38224);
and U42396 (N_42396,N_37917,N_39682);
xnor U42397 (N_42397,N_38988,N_39596);
xnor U42398 (N_42398,N_39297,N_38032);
or U42399 (N_42399,N_37566,N_38232);
nand U42400 (N_42400,N_37848,N_38080);
nand U42401 (N_42401,N_38287,N_39409);
xor U42402 (N_42402,N_39117,N_39730);
nand U42403 (N_42403,N_39298,N_39504);
or U42404 (N_42404,N_39160,N_39525);
nand U42405 (N_42405,N_38509,N_38834);
or U42406 (N_42406,N_38301,N_38882);
xnor U42407 (N_42407,N_37821,N_37600);
nand U42408 (N_42408,N_38475,N_39605);
nand U42409 (N_42409,N_38440,N_38824);
or U42410 (N_42410,N_39244,N_39145);
and U42411 (N_42411,N_39599,N_39144);
and U42412 (N_42412,N_38447,N_37506);
nor U42413 (N_42413,N_38082,N_39987);
or U42414 (N_42414,N_39600,N_37874);
nor U42415 (N_42415,N_38394,N_38905);
nor U42416 (N_42416,N_39723,N_38619);
nand U42417 (N_42417,N_39649,N_39993);
nor U42418 (N_42418,N_38590,N_39402);
nand U42419 (N_42419,N_39367,N_38726);
xor U42420 (N_42420,N_38743,N_39107);
and U42421 (N_42421,N_38132,N_39245);
nand U42422 (N_42422,N_39253,N_37657);
and U42423 (N_42423,N_38001,N_39413);
and U42424 (N_42424,N_38572,N_37501);
xor U42425 (N_42425,N_39916,N_39435);
nand U42426 (N_42426,N_37542,N_38646);
or U42427 (N_42427,N_39196,N_38204);
nand U42428 (N_42428,N_38912,N_38029);
and U42429 (N_42429,N_39922,N_39017);
or U42430 (N_42430,N_38392,N_38903);
or U42431 (N_42431,N_37607,N_39409);
xor U42432 (N_42432,N_37760,N_37997);
nand U42433 (N_42433,N_37975,N_39704);
nand U42434 (N_42434,N_39308,N_37813);
nand U42435 (N_42435,N_37512,N_39502);
xnor U42436 (N_42436,N_38243,N_38201);
nand U42437 (N_42437,N_37933,N_38361);
nand U42438 (N_42438,N_38383,N_39477);
nand U42439 (N_42439,N_37796,N_38856);
or U42440 (N_42440,N_38776,N_38019);
nand U42441 (N_42441,N_38957,N_37675);
nor U42442 (N_42442,N_38593,N_39657);
and U42443 (N_42443,N_38894,N_37767);
nand U42444 (N_42444,N_38086,N_38732);
and U42445 (N_42445,N_39646,N_38068);
or U42446 (N_42446,N_39551,N_38954);
and U42447 (N_42447,N_39767,N_37582);
nor U42448 (N_42448,N_38395,N_38566);
xnor U42449 (N_42449,N_37997,N_38301);
nor U42450 (N_42450,N_39244,N_39742);
or U42451 (N_42451,N_39192,N_39727);
xnor U42452 (N_42452,N_37844,N_37600);
nand U42453 (N_42453,N_37635,N_37830);
nor U42454 (N_42454,N_39506,N_39259);
nand U42455 (N_42455,N_37727,N_38741);
nor U42456 (N_42456,N_37909,N_38928);
nor U42457 (N_42457,N_38210,N_38216);
xnor U42458 (N_42458,N_38123,N_38328);
or U42459 (N_42459,N_38120,N_38254);
xnor U42460 (N_42460,N_38061,N_37655);
nor U42461 (N_42461,N_38729,N_39113);
nand U42462 (N_42462,N_38414,N_38598);
xor U42463 (N_42463,N_37589,N_37651);
nand U42464 (N_42464,N_39702,N_39219);
and U42465 (N_42465,N_38590,N_38237);
nand U42466 (N_42466,N_39476,N_38298);
nor U42467 (N_42467,N_39323,N_39780);
or U42468 (N_42468,N_38885,N_39680);
xor U42469 (N_42469,N_38045,N_38199);
or U42470 (N_42470,N_37553,N_38956);
and U42471 (N_42471,N_38113,N_37948);
nor U42472 (N_42472,N_38351,N_37584);
or U42473 (N_42473,N_37830,N_38866);
nand U42474 (N_42474,N_38140,N_38343);
and U42475 (N_42475,N_38908,N_39057);
and U42476 (N_42476,N_37501,N_38906);
xor U42477 (N_42477,N_38355,N_37536);
xnor U42478 (N_42478,N_37703,N_37700);
nor U42479 (N_42479,N_38502,N_39625);
and U42480 (N_42480,N_38031,N_39872);
or U42481 (N_42481,N_39002,N_39872);
or U42482 (N_42482,N_38912,N_38686);
xnor U42483 (N_42483,N_37714,N_37628);
xor U42484 (N_42484,N_39146,N_39904);
xnor U42485 (N_42485,N_38758,N_38505);
xor U42486 (N_42486,N_37867,N_38386);
xor U42487 (N_42487,N_38203,N_39626);
xor U42488 (N_42488,N_38708,N_38597);
nor U42489 (N_42489,N_38354,N_39296);
and U42490 (N_42490,N_39778,N_38862);
nand U42491 (N_42491,N_38873,N_37948);
nand U42492 (N_42492,N_39819,N_37518);
nor U42493 (N_42493,N_37686,N_39149);
xnor U42494 (N_42494,N_38656,N_38393);
nor U42495 (N_42495,N_38612,N_38031);
nor U42496 (N_42496,N_37643,N_39903);
and U42497 (N_42497,N_39060,N_38466);
nor U42498 (N_42498,N_37925,N_38939);
and U42499 (N_42499,N_37971,N_38722);
nor U42500 (N_42500,N_40251,N_41522);
nand U42501 (N_42501,N_41496,N_40878);
xnor U42502 (N_42502,N_40278,N_42397);
and U42503 (N_42503,N_42378,N_42466);
nand U42504 (N_42504,N_40308,N_41085);
nor U42505 (N_42505,N_40791,N_42388);
or U42506 (N_42506,N_42290,N_40919);
nand U42507 (N_42507,N_40794,N_41833);
nand U42508 (N_42508,N_41569,N_40509);
and U42509 (N_42509,N_41313,N_42447);
and U42510 (N_42510,N_40048,N_42228);
nor U42511 (N_42511,N_40062,N_40914);
nand U42512 (N_42512,N_40229,N_40266);
and U42513 (N_42513,N_40922,N_41612);
nor U42514 (N_42514,N_42385,N_40999);
nor U42515 (N_42515,N_42318,N_40905);
nand U42516 (N_42516,N_41451,N_41906);
nor U42517 (N_42517,N_40259,N_41784);
nand U42518 (N_42518,N_41865,N_41472);
nand U42519 (N_42519,N_41631,N_41221);
and U42520 (N_42520,N_40706,N_42138);
xor U42521 (N_42521,N_41911,N_42164);
and U42522 (N_42522,N_41386,N_40641);
nor U42523 (N_42523,N_40370,N_41940);
xnor U42524 (N_42524,N_41992,N_41859);
or U42525 (N_42525,N_40651,N_41072);
or U42526 (N_42526,N_40164,N_41203);
nor U42527 (N_42527,N_41069,N_40953);
xor U42528 (N_42528,N_41093,N_41272);
and U42529 (N_42529,N_41849,N_41256);
xnor U42530 (N_42530,N_41020,N_41573);
xor U42531 (N_42531,N_40753,N_40989);
nor U42532 (N_42532,N_41663,N_40979);
or U42533 (N_42533,N_42021,N_40193);
nand U42534 (N_42534,N_41922,N_41079);
and U42535 (N_42535,N_42023,N_41948);
xnor U42536 (N_42536,N_41314,N_41083);
or U42537 (N_42537,N_40392,N_41912);
and U42538 (N_42538,N_40369,N_42205);
nor U42539 (N_42539,N_41892,N_40085);
nand U42540 (N_42540,N_41581,N_41341);
or U42541 (N_42541,N_42077,N_42368);
xnor U42542 (N_42542,N_40961,N_42367);
and U42543 (N_42543,N_40937,N_40656);
and U42544 (N_42544,N_40262,N_40091);
nor U42545 (N_42545,N_40247,N_40415);
or U42546 (N_42546,N_42452,N_42090);
nor U42547 (N_42547,N_42065,N_41883);
and U42548 (N_42548,N_40783,N_41861);
and U42549 (N_42549,N_41009,N_41999);
and U42550 (N_42550,N_40101,N_40825);
and U42551 (N_42551,N_41866,N_40529);
and U42552 (N_42552,N_41116,N_40406);
xor U42553 (N_42553,N_40615,N_42297);
nor U42554 (N_42554,N_40993,N_42246);
xor U42555 (N_42555,N_42132,N_41404);
nor U42556 (N_42556,N_42155,N_41648);
nand U42557 (N_42557,N_40135,N_40936);
nand U42558 (N_42558,N_40560,N_41302);
or U42559 (N_42559,N_40359,N_41567);
nand U42560 (N_42560,N_40854,N_41145);
xnor U42561 (N_42561,N_41030,N_42232);
nand U42562 (N_42562,N_41794,N_40241);
nand U42563 (N_42563,N_40280,N_41413);
nor U42564 (N_42564,N_41089,N_40893);
or U42565 (N_42565,N_42028,N_40077);
nand U42566 (N_42566,N_42442,N_41381);
nand U42567 (N_42567,N_40918,N_41614);
and U42568 (N_42568,N_41147,N_42491);
or U42569 (N_42569,N_41936,N_41981);
nand U42570 (N_42570,N_40694,N_40442);
nand U42571 (N_42571,N_41318,N_40363);
nand U42572 (N_42572,N_40631,N_41260);
xor U42573 (N_42573,N_40899,N_42222);
xnor U42574 (N_42574,N_40632,N_41232);
xnor U42575 (N_42575,N_40365,N_42469);
or U42576 (N_42576,N_42443,N_42113);
nor U42577 (N_42577,N_41643,N_40527);
nand U42578 (N_42578,N_40648,N_40635);
and U42579 (N_42579,N_42371,N_41798);
and U42580 (N_42580,N_40441,N_41813);
xor U42581 (N_42581,N_41026,N_41852);
nor U42582 (N_42582,N_40029,N_40860);
or U42583 (N_42583,N_40275,N_40223);
nand U42584 (N_42584,N_41515,N_40831);
nand U42585 (N_42585,N_41641,N_40186);
or U42586 (N_42586,N_41476,N_41233);
or U42587 (N_42587,N_41727,N_40561);
xor U42588 (N_42588,N_40778,N_41445);
xnor U42589 (N_42589,N_41140,N_42172);
or U42590 (N_42590,N_41052,N_40121);
or U42591 (N_42591,N_41760,N_40707);
nand U42592 (N_42592,N_41745,N_42010);
nand U42593 (N_42593,N_40524,N_41755);
nand U42594 (N_42594,N_41566,N_42372);
nor U42595 (N_42595,N_41461,N_41730);
and U42596 (N_42596,N_41736,N_41667);
xor U42597 (N_42597,N_40986,N_41729);
or U42598 (N_42598,N_42379,N_41956);
and U42599 (N_42599,N_40337,N_42216);
or U42600 (N_42600,N_40735,N_40178);
and U42601 (N_42601,N_40503,N_42408);
nor U42602 (N_42602,N_40788,N_42067);
and U42603 (N_42603,N_40421,N_41795);
and U42604 (N_42604,N_41257,N_40996);
nand U42605 (N_42605,N_42211,N_42178);
or U42606 (N_42606,N_40440,N_41563);
xnor U42607 (N_42607,N_40790,N_42059);
and U42608 (N_42608,N_40254,N_41635);
nor U42609 (N_42609,N_42489,N_40130);
xnor U42610 (N_42610,N_41202,N_40469);
and U42611 (N_42611,N_41692,N_42152);
nor U42612 (N_42612,N_41489,N_42386);
xnor U42613 (N_42613,N_41903,N_41400);
xnor U42614 (N_42614,N_41128,N_41230);
nand U42615 (N_42615,N_41671,N_40901);
and U42616 (N_42616,N_40033,N_41562);
or U42617 (N_42617,N_41388,N_41756);
nand U42618 (N_42618,N_40722,N_41344);
and U42619 (N_42619,N_42061,N_42206);
and U42620 (N_42620,N_41226,N_42184);
nand U42621 (N_42621,N_40260,N_41923);
nor U42622 (N_42622,N_41448,N_42224);
or U42623 (N_42623,N_42012,N_40747);
nor U42624 (N_42624,N_41157,N_42374);
nand U42625 (N_42625,N_40611,N_41953);
nor U42626 (N_42626,N_40313,N_41991);
xor U42627 (N_42627,N_41066,N_41048);
xor U42628 (N_42628,N_41475,N_41658);
xnor U42629 (N_42629,N_40243,N_41190);
nand U42630 (N_42630,N_40506,N_40792);
or U42631 (N_42631,N_41686,N_42352);
and U42632 (N_42632,N_40328,N_40728);
nand U42633 (N_42633,N_40482,N_42230);
and U42634 (N_42634,N_40608,N_42338);
and U42635 (N_42635,N_41441,N_42497);
or U42636 (N_42636,N_40481,N_41076);
xor U42637 (N_42637,N_41354,N_41543);
or U42638 (N_42638,N_40143,N_42008);
or U42639 (N_42639,N_40207,N_41856);
and U42640 (N_42640,N_42045,N_41875);
xnor U42641 (N_42641,N_40601,N_42308);
nand U42642 (N_42642,N_41243,N_42042);
and U42643 (N_42643,N_40401,N_41882);
xor U42644 (N_42644,N_40677,N_42055);
nand U42645 (N_42645,N_40926,N_42109);
xor U42646 (N_42646,N_41575,N_41978);
xor U42647 (N_42647,N_42087,N_41169);
nand U42648 (N_42648,N_41674,N_41378);
or U42649 (N_42649,N_42175,N_41039);
and U42650 (N_42650,N_40981,N_40782);
and U42651 (N_42651,N_41802,N_42460);
xnor U42652 (N_42652,N_40625,N_41022);
nand U42653 (N_42653,N_40713,N_41787);
xnor U42654 (N_42654,N_41468,N_41974);
nand U42655 (N_42655,N_41278,N_41368);
xnor U42656 (N_42656,N_41086,N_41154);
xnor U42657 (N_42657,N_42248,N_41415);
and U42658 (N_42658,N_42085,N_40149);
xnor U42659 (N_42659,N_40938,N_41783);
nor U42660 (N_42660,N_41721,N_40940);
and U42661 (N_42661,N_41007,N_40110);
nand U42662 (N_42662,N_40982,N_40209);
nor U42663 (N_42663,N_40799,N_41121);
and U42664 (N_42664,N_42403,N_41160);
nor U42665 (N_42665,N_41764,N_40011);
xnor U42666 (N_42666,N_42270,N_41375);
and U42667 (N_42667,N_41768,N_41464);
and U42668 (N_42668,N_41509,N_40749);
or U42669 (N_42669,N_41073,N_41456);
or U42670 (N_42670,N_41176,N_40820);
xor U42671 (N_42671,N_42307,N_41336);
nor U42672 (N_42672,N_42160,N_42025);
xor U42673 (N_42673,N_42133,N_41952);
xor U42674 (N_42674,N_41210,N_40669);
nand U42675 (N_42675,N_40255,N_40589);
or U42676 (N_42676,N_42238,N_41239);
or U42677 (N_42677,N_41946,N_41327);
nor U42678 (N_42678,N_41251,N_41700);
or U42679 (N_42679,N_41647,N_40240);
or U42680 (N_42680,N_41850,N_40861);
nand U42681 (N_42681,N_40204,N_40472);
xor U42682 (N_42682,N_40386,N_40065);
nand U42683 (N_42683,N_42208,N_41961);
xor U42684 (N_42684,N_42425,N_40410);
or U42685 (N_42685,N_41045,N_40105);
xnor U42686 (N_42686,N_41574,N_41824);
and U42687 (N_42687,N_42310,N_41781);
xnor U42688 (N_42688,N_42415,N_41545);
xor U42689 (N_42689,N_40044,N_40023);
xor U42690 (N_42690,N_40134,N_41299);
nor U42691 (N_42691,N_42089,N_40590);
nor U42692 (N_42692,N_40807,N_40843);
nor U42693 (N_42693,N_40718,N_40063);
or U42694 (N_42694,N_41896,N_40715);
nor U42695 (N_42695,N_40984,N_41511);
xor U42696 (N_42696,N_40427,N_42414);
nand U42697 (N_42697,N_41062,N_41803);
xor U42698 (N_42698,N_42106,N_42038);
nand U42699 (N_42699,N_41238,N_41901);
or U42700 (N_42700,N_40086,N_40559);
xor U42701 (N_42701,N_41332,N_41786);
or U42702 (N_42702,N_42039,N_41275);
nor U42703 (N_42703,N_40092,N_40946);
nor U42704 (N_42704,N_41857,N_40399);
and U42705 (N_42705,N_41568,N_40955);
nor U42706 (N_42706,N_40903,N_40532);
and U42707 (N_42707,N_42462,N_41799);
and U42708 (N_42708,N_41293,N_41944);
xor U42709 (N_42709,N_41542,N_40881);
xor U42710 (N_42710,N_41735,N_40304);
nand U42711 (N_42711,N_42197,N_41357);
nand U42712 (N_42712,N_40634,N_41928);
nor U42713 (N_42713,N_41660,N_42110);
and U42714 (N_42714,N_40962,N_42080);
and U42715 (N_42715,N_41106,N_41038);
xnor U42716 (N_42716,N_41640,N_41159);
and U42717 (N_42717,N_41935,N_41317);
or U42718 (N_42718,N_41268,N_40617);
or U42719 (N_42719,N_42453,N_40423);
xnor U42720 (N_42720,N_41060,N_41576);
and U42721 (N_42721,N_40624,N_41312);
and U42722 (N_42722,N_42070,N_41077);
nand U42723 (N_42723,N_40281,N_40437);
or U42724 (N_42724,N_42467,N_41362);
and U42725 (N_42725,N_41734,N_41739);
xor U42726 (N_42726,N_40075,N_40991);
nand U42727 (N_42727,N_42114,N_40967);
nor U42728 (N_42728,N_40122,N_41891);
or U42729 (N_42729,N_40710,N_41544);
nor U42730 (N_42730,N_41138,N_41639);
and U42731 (N_42731,N_40521,N_41012);
xnor U42732 (N_42732,N_40570,N_40805);
nand U42733 (N_42733,N_41284,N_42141);
nand U42734 (N_42734,N_40599,N_42076);
or U42735 (N_42735,N_41282,N_41367);
xnor U42736 (N_42736,N_41831,N_41514);
and U42737 (N_42737,N_42422,N_41405);
nand U42738 (N_42738,N_41845,N_41333);
or U42739 (N_42739,N_40020,N_42487);
nand U42740 (N_42740,N_40815,N_41743);
or U42741 (N_42741,N_40238,N_41267);
nand U42742 (N_42742,N_40719,N_42325);
nor U42743 (N_42743,N_42256,N_41254);
or U42744 (N_42744,N_41290,N_41193);
and U42745 (N_42745,N_42103,N_40948);
or U42746 (N_42746,N_41494,N_41331);
nor U42747 (N_42747,N_41549,N_42366);
nor U42748 (N_42748,N_41876,N_42321);
xor U42749 (N_42749,N_41477,N_40541);
nor U42750 (N_42750,N_40496,N_40120);
xnor U42751 (N_42751,N_41701,N_41490);
and U42752 (N_42752,N_40975,N_40089);
or U42753 (N_42753,N_40580,N_41305);
xnor U42754 (N_42754,N_40419,N_41111);
and U42755 (N_42755,N_40612,N_41763);
xnor U42756 (N_42756,N_41123,N_41863);
nor U42757 (N_42757,N_40983,N_41538);
xor U42758 (N_42758,N_41589,N_41731);
nor U42759 (N_42759,N_41198,N_42468);
nand U42760 (N_42760,N_40428,N_40320);
or U42761 (N_42761,N_40454,N_40945);
nor U42762 (N_42762,N_41644,N_40483);
and U42763 (N_42763,N_40520,N_40236);
nor U42764 (N_42764,N_42476,N_41216);
xor U42765 (N_42765,N_40813,N_40555);
nand U42766 (N_42766,N_41450,N_41807);
nor U42767 (N_42767,N_40618,N_41829);
and U42768 (N_42768,N_41976,N_41526);
xnor U42769 (N_42769,N_41273,N_41291);
and U42770 (N_42770,N_41227,N_40663);
xnor U42771 (N_42771,N_41422,N_40645);
and U42772 (N_42772,N_40908,N_40097);
nand U42773 (N_42773,N_41791,N_42274);
nor U42774 (N_42774,N_41818,N_40675);
and U42775 (N_42775,N_40705,N_40367);
or U42776 (N_42776,N_40150,N_41929);
and U42777 (N_42777,N_41462,N_40154);
and U42778 (N_42778,N_42348,N_40330);
nand U42779 (N_42779,N_40581,N_41505);
nand U42780 (N_42780,N_40289,N_42299);
or U42781 (N_42781,N_42312,N_41682);
xor U42782 (N_42782,N_41200,N_41329);
xor U42783 (N_42783,N_41893,N_41649);
xor U42784 (N_42784,N_40391,N_41143);
or U42785 (N_42785,N_40679,N_41950);
nor U42786 (N_42786,N_40575,N_41114);
nor U42787 (N_42787,N_40144,N_41955);
nor U42788 (N_42788,N_41611,N_40334);
or U42789 (N_42789,N_42179,N_42236);
and U42790 (N_42790,N_40758,N_41155);
nand U42791 (N_42791,N_40389,N_42009);
nand U42792 (N_42792,N_41053,N_40119);
or U42793 (N_42793,N_42139,N_41390);
and U42794 (N_42794,N_42284,N_42257);
nor U42795 (N_42795,N_40864,N_40526);
or U42796 (N_42796,N_41192,N_40194);
or U42797 (N_42797,N_40851,N_41605);
and U42798 (N_42798,N_41555,N_41355);
xnor U42799 (N_42799,N_40818,N_41110);
or U42800 (N_42800,N_40080,N_41356);
or U42801 (N_42801,N_41826,N_40405);
or U42802 (N_42802,N_42041,N_42199);
nand U42803 (N_42803,N_40765,N_41492);
nor U42804 (N_42804,N_40510,N_42186);
nor U42805 (N_42805,N_42245,N_42212);
xnor U42806 (N_42806,N_40375,N_42051);
nor U42807 (N_42807,N_40809,N_41751);
or U42808 (N_42808,N_42354,N_40049);
or U42809 (N_42809,N_40803,N_41528);
or U42810 (N_42810,N_42240,N_42473);
or U42811 (N_42811,N_41161,N_40849);
xnor U42812 (N_42812,N_40358,N_41491);
or U42813 (N_42813,N_40569,N_41005);
nand U42814 (N_42814,N_40351,N_41100);
nor U42815 (N_42815,N_40733,N_42219);
nand U42816 (N_42816,N_40323,N_42389);
and U42817 (N_42817,N_41090,N_40286);
or U42818 (N_42818,N_41248,N_40219);
xnor U42819 (N_42819,N_41207,N_40288);
nand U42820 (N_42820,N_42235,N_40628);
nand U42821 (N_42821,N_41351,N_41015);
nand U42822 (N_42822,N_41990,N_40028);
nor U42823 (N_42823,N_41777,N_40811);
nand U42824 (N_42824,N_40103,N_40225);
or U42825 (N_42825,N_42081,N_41270);
and U42826 (N_42826,N_42058,N_40913);
nor U42827 (N_42827,N_40776,N_40264);
nor U42828 (N_42828,N_40703,N_42298);
nor U42829 (N_42829,N_41184,N_40959);
nand U42830 (N_42830,N_41889,N_42189);
nor U42831 (N_42831,N_40671,N_40489);
or U42832 (N_42832,N_41334,N_40382);
or U42833 (N_42833,N_40279,N_42084);
nand U42834 (N_42834,N_40468,N_40036);
nand U42835 (N_42835,N_40683,N_42401);
nand U42836 (N_42836,N_40342,N_40867);
nor U42837 (N_42837,N_42359,N_40587);
nand U42838 (N_42838,N_41792,N_41716);
nand U42839 (N_42839,N_42498,N_42183);
and U42840 (N_42840,N_42412,N_40923);
nor U42841 (N_42841,N_42158,N_41623);
nand U42842 (N_42842,N_41665,N_40514);
nor U42843 (N_42843,N_40985,N_42483);
and U42844 (N_42844,N_40270,N_40233);
nand U42845 (N_42845,N_41880,N_40252);
nor U42846 (N_42846,N_42168,N_42112);
and U42847 (N_42847,N_41151,N_40404);
and U42848 (N_42848,N_41695,N_40933);
nor U42849 (N_42849,N_41394,N_40630);
xor U42850 (N_42850,N_40015,N_42440);
xor U42851 (N_42851,N_40906,N_40109);
or U42852 (N_42852,N_40883,N_42022);
nor U42853 (N_42853,N_40868,N_42239);
nand U42854 (N_42854,N_41283,N_42384);
nand U42855 (N_42855,N_40283,N_40714);
nand U42856 (N_42856,N_40844,N_42279);
or U42857 (N_42857,N_42017,N_41481);
xnor U42858 (N_42858,N_42127,N_41740);
xnor U42859 (N_42859,N_40637,N_42194);
nand U42860 (N_42860,N_40136,N_41245);
nand U42861 (N_42861,N_40220,N_41624);
nor U42862 (N_42862,N_40268,N_42000);
nand U42863 (N_42863,N_40595,N_40808);
and U42864 (N_42864,N_40132,N_40299);
and U42865 (N_42865,N_40557,N_40185);
xor U42866 (N_42866,N_40739,N_42171);
nand U42867 (N_42867,N_41029,N_40424);
xor U42868 (N_42868,N_41398,N_40586);
and U42869 (N_42869,N_40093,N_41801);
or U42870 (N_42870,N_41136,N_40316);
nand U42871 (N_42871,N_41306,N_40341);
and U42872 (N_42872,N_41713,N_40113);
nand U42873 (N_42873,N_42108,N_40537);
and U42874 (N_42874,N_40958,N_41890);
or U42875 (N_42875,N_40727,N_42072);
nand U42876 (N_42876,N_41884,N_40335);
xor U42877 (N_42877,N_41057,N_41371);
nand U42878 (N_42878,N_41941,N_41812);
and U42879 (N_42879,N_41907,N_40786);
and U42880 (N_42880,N_41591,N_40622);
xnor U42881 (N_42881,N_40689,N_40187);
nor U42882 (N_42882,N_40835,N_41814);
or U42883 (N_42883,N_40915,N_41797);
or U42884 (N_42884,N_42269,N_41061);
nor U42885 (N_42885,N_42258,N_42190);
xnor U42886 (N_42886,N_42436,N_40484);
xnor U42887 (N_42887,N_40017,N_40199);
nor U42888 (N_42888,N_40640,N_40619);
nand U42889 (N_42889,N_42277,N_40374);
nand U42890 (N_42890,N_40793,N_40939);
and U42891 (N_42891,N_41131,N_41399);
and U42892 (N_42892,N_40709,N_40968);
xnor U42893 (N_42893,N_41163,N_41359);
or U42894 (N_42894,N_40688,N_41733);
or U42895 (N_42895,N_40162,N_42363);
xor U42896 (N_42896,N_40814,N_42461);
nand U42897 (N_42897,N_42119,N_41534);
nand U42898 (N_42898,N_41104,N_40292);
or U42899 (N_42899,N_40978,N_40859);
or U42900 (N_42900,N_41793,N_40411);
xor U42901 (N_42901,N_42444,N_42002);
nor U42902 (N_42902,N_40090,N_41231);
or U42903 (N_42903,N_40131,N_42381);
or U42904 (N_42904,N_42347,N_40554);
and U42905 (N_42905,N_41748,N_40165);
and U42906 (N_42906,N_41843,N_40137);
nor U42907 (N_42907,N_40485,N_40460);
nand U42908 (N_42908,N_40171,N_40038);
or U42909 (N_42909,N_42069,N_40012);
nor U42910 (N_42910,N_41046,N_40346);
and U42911 (N_42911,N_41601,N_41274);
and U42912 (N_42912,N_41707,N_41269);
xor U42913 (N_42913,N_41939,N_41970);
nor U42914 (N_42914,N_40997,N_40830);
xnor U42915 (N_42915,N_41983,N_40471);
nor U42916 (N_42916,N_41881,N_40079);
nor U42917 (N_42917,N_40785,N_40839);
or U42918 (N_42918,N_41049,N_42449);
or U42919 (N_42919,N_40473,N_40852);
and U42920 (N_42920,N_41391,N_41420);
and U42921 (N_42921,N_41153,N_41460);
nand U42922 (N_42922,N_41199,N_42096);
or U42923 (N_42923,N_40723,N_42137);
and U42924 (N_42924,N_40726,N_41554);
and U42925 (N_42925,N_42146,N_41434);
nand U42926 (N_42926,N_42302,N_40704);
nor U42927 (N_42927,N_40716,N_40061);
xnor U42928 (N_42928,N_40692,N_41634);
nor U42929 (N_42929,N_40487,N_41240);
nand U42930 (N_42930,N_42182,N_42073);
nor U42931 (N_42931,N_41525,N_41546);
nor U42932 (N_42932,N_41711,N_40691);
xnor U42933 (N_42933,N_42405,N_42342);
xor U42934 (N_42934,N_41986,N_41068);
xor U42935 (N_42935,N_41853,N_40752);
and U42936 (N_42936,N_41900,N_41766);
or U42937 (N_42937,N_41326,N_40349);
nor U42938 (N_42938,N_41493,N_40965);
xor U42939 (N_42939,N_41443,N_40274);
and U42940 (N_42940,N_40523,N_42079);
and U42941 (N_42941,N_40156,N_40453);
nand U42942 (N_42942,N_42420,N_41816);
xor U42943 (N_42943,N_41056,N_40202);
xor U42944 (N_42944,N_40180,N_41094);
xor U42945 (N_42945,N_41628,N_40216);
or U42946 (N_42946,N_40245,N_42163);
or U42947 (N_42947,N_41775,N_42118);
and U42948 (N_42948,N_42396,N_41677);
or U42949 (N_42949,N_42404,N_41609);
and U42950 (N_42950,N_40476,N_40872);
nor U42951 (N_42951,N_40538,N_41280);
nand U42952 (N_42952,N_40539,N_42210);
or U42953 (N_42953,N_40235,N_40681);
nor U42954 (N_42954,N_40161,N_40099);
and U42955 (N_42955,N_40300,N_42064);
and U42956 (N_42956,N_40294,N_41197);
and U42957 (N_42957,N_41765,N_41619);
or U42958 (N_42958,N_41790,N_41379);
nand U42959 (N_42959,N_40750,N_42407);
xnor U42960 (N_42960,N_42100,N_40222);
xor U42961 (N_42961,N_42047,N_41212);
nand U42962 (N_42962,N_40660,N_42296);
or U42963 (N_42963,N_41253,N_42317);
nand U42964 (N_42964,N_41366,N_40212);
and U42965 (N_42965,N_40412,N_41828);
nor U42966 (N_42966,N_40331,N_41173);
xor U42967 (N_42967,N_40976,N_40610);
nand U42968 (N_42968,N_42380,N_42454);
xor U42969 (N_42969,N_40898,N_40183);
xnor U42970 (N_42970,N_41625,N_40781);
nor U42971 (N_42971,N_41590,N_40383);
nand U42972 (N_42972,N_40837,N_40927);
and U42973 (N_42973,N_41209,N_41224);
or U42974 (N_42974,N_41058,N_40884);
nand U42975 (N_42975,N_42099,N_40040);
nand U42976 (N_42976,N_40819,N_42134);
or U42977 (N_42977,N_42259,N_40507);
nor U42978 (N_42978,N_41179,N_41835);
nand U42979 (N_42979,N_42349,N_40552);
nand U42980 (N_42980,N_40258,N_40102);
xor U42981 (N_42981,N_41806,N_42463);
or U42982 (N_42982,N_41115,N_41340);
nand U42983 (N_42983,N_42343,N_40112);
or U42984 (N_42984,N_40265,N_41234);
and U42985 (N_42985,N_41350,N_42432);
or U42986 (N_42986,N_40360,N_40478);
or U42987 (N_42987,N_42464,N_41098);
nor U42988 (N_42988,N_41335,N_42326);
nand U42989 (N_42989,N_41702,N_40654);
nand U42990 (N_42990,N_40492,N_41297);
or U42991 (N_42991,N_41117,N_40188);
nand U42992 (N_42992,N_41425,N_40596);
nor U42993 (N_42993,N_40944,N_42244);
xnor U42994 (N_42994,N_41175,N_41220);
nand U42995 (N_42995,N_41032,N_40564);
nand U42996 (N_42996,N_41466,N_40115);
nand U42997 (N_42997,N_41874,N_41502);
xor U42998 (N_42998,N_42305,N_40582);
or U42999 (N_42999,N_40362,N_40378);
or U43000 (N_43000,N_42459,N_40083);
or U43001 (N_43001,N_41851,N_42188);
and U43002 (N_43002,N_41517,N_42485);
nand U43003 (N_43003,N_40145,N_42387);
and U43004 (N_43004,N_42068,N_40877);
nand U43005 (N_43005,N_41718,N_40016);
nor U43006 (N_43006,N_42413,N_41839);
xnor U43007 (N_43007,N_40970,N_40123);
xor U43008 (N_43008,N_40301,N_40879);
or U43009 (N_43009,N_40543,N_41547);
nor U43010 (N_43010,N_40605,N_41918);
nand U43011 (N_43011,N_42048,N_40198);
nor U43012 (N_43012,N_40806,N_42267);
nand U43013 (N_43013,N_40592,N_42488);
nand U43014 (N_43014,N_41669,N_41164);
and U43015 (N_43015,N_42266,N_40071);
or U43016 (N_43016,N_40836,N_40098);
nand U43017 (N_43017,N_41247,N_42121);
xor U43018 (N_43018,N_41300,N_42324);
nand U43019 (N_43019,N_41603,N_42026);
nor U43020 (N_43020,N_41617,N_41382);
nor U43021 (N_43021,N_40231,N_40729);
nor U43022 (N_43022,N_41449,N_41250);
nor U43023 (N_43023,N_41864,N_41681);
nor U43024 (N_43024,N_41469,N_41523);
xnor U43025 (N_43025,N_41780,N_42036);
nand U43026 (N_43026,N_40159,N_42475);
or U43027 (N_43027,N_40434,N_42094);
and U43028 (N_43028,N_41915,N_40636);
nor U43029 (N_43029,N_41010,N_42434);
or U43030 (N_43030,N_42337,N_41973);
nand U43031 (N_43031,N_40887,N_41582);
or U43032 (N_43032,N_40657,N_42391);
nor U43033 (N_43033,N_40567,N_41189);
and U43034 (N_43034,N_41615,N_40444);
and U43035 (N_43035,N_40203,N_41962);
or U43036 (N_43036,N_40643,N_40324);
xnor U43037 (N_43037,N_41465,N_40842);
xnor U43038 (N_43038,N_40556,N_40620);
nor U43039 (N_43039,N_40455,N_42477);
xor U43040 (N_43040,N_40838,N_41762);
or U43041 (N_43041,N_40588,N_41886);
xnor U43042 (N_43042,N_41951,N_40311);
and U43043 (N_43043,N_41844,N_40291);
nand U43044 (N_43044,N_40295,N_40059);
nor U43045 (N_43045,N_41364,N_41279);
nand U43046 (N_43046,N_40014,N_40850);
or U43047 (N_43047,N_41885,N_41697);
and U43048 (N_43048,N_42247,N_42339);
nor U43049 (N_43049,N_40361,N_40687);
and U43050 (N_43050,N_41914,N_42209);
or U43051 (N_43051,N_41823,N_42254);
xor U43052 (N_43052,N_42144,N_40568);
xor U43053 (N_43053,N_41910,N_41298);
xor U43054 (N_43054,N_41361,N_42336);
xor U43055 (N_43055,N_40693,N_41265);
and U43056 (N_43056,N_40591,N_41008);
xnor U43057 (N_43057,N_40900,N_42278);
nor U43058 (N_43058,N_42123,N_42030);
nand U43059 (N_43059,N_41678,N_42409);
xor U43060 (N_43060,N_41530,N_41454);
xor U43061 (N_43061,N_40443,N_41998);
nand U43062 (N_43062,N_40594,N_40699);
or U43063 (N_43063,N_40664,N_41725);
xor U43064 (N_43064,N_41035,N_42243);
nand U43065 (N_43065,N_41602,N_41051);
xnor U43066 (N_43066,N_40638,N_41597);
nand U43067 (N_43067,N_42335,N_40181);
nor U43068 (N_43068,N_40544,N_41255);
xor U43069 (N_43069,N_41516,N_41887);
and U43070 (N_43070,N_41447,N_40841);
nor U43071 (N_43071,N_40420,N_40155);
xnor U43072 (N_43072,N_40573,N_40777);
nand U43073 (N_43073,N_40057,N_41820);
xor U43074 (N_43074,N_42494,N_41433);
xor U43075 (N_43075,N_40880,N_40649);
nor U43076 (N_43076,N_41728,N_42490);
nand U43077 (N_43077,N_41899,N_40550);
and U43078 (N_43078,N_42018,N_40152);
nand U43079 (N_43079,N_41670,N_41825);
xor U43080 (N_43080,N_41262,N_42226);
nor U43081 (N_43081,N_40070,N_42316);
and U43082 (N_43082,N_40160,N_41694);
xnor U43083 (N_43083,N_42276,N_40647);
and U43084 (N_43084,N_42275,N_42400);
nor U43085 (N_43085,N_40214,N_42264);
xor U43086 (N_43086,N_40069,N_42351);
nor U43087 (N_43087,N_41596,N_42470);
xnor U43088 (N_43088,N_41206,N_40816);
or U43089 (N_43089,N_40789,N_42345);
nand U43090 (N_43090,N_41572,N_41440);
xor U43091 (N_43091,N_40652,N_40332);
or U43092 (N_43092,N_41223,N_40563);
xor U43093 (N_43093,N_42439,N_40430);
nand U43094 (N_43094,N_40779,N_42054);
nor U43095 (N_43095,N_40821,N_41324);
nand U43096 (N_43096,N_41099,N_41985);
or U43097 (N_43097,N_41019,N_40250);
xnor U43098 (N_43098,N_40317,N_40771);
and U43099 (N_43099,N_42481,N_41958);
xor U43100 (N_43100,N_40021,N_41487);
nor U43101 (N_43101,N_40598,N_41266);
nor U43102 (N_43102,N_40095,N_42433);
and U43103 (N_43103,N_41698,N_42034);
or U43104 (N_43104,N_41264,N_40627);
nand U43105 (N_43105,N_41673,N_40339);
nor U43106 (N_43106,N_40576,N_41873);
nor U43107 (N_43107,N_41041,N_40462);
nand U43108 (N_43108,N_42450,N_40060);
and U43109 (N_43109,N_40290,N_41183);
and U43110 (N_43110,N_40045,N_41897);
xnor U43111 (N_43111,N_41288,N_41118);
xor U43112 (N_43112,N_41706,N_41289);
xor U43113 (N_43113,N_40046,N_40190);
xor U43114 (N_43114,N_42187,N_41868);
nor U43115 (N_43115,N_42390,N_40672);
xor U43116 (N_43116,N_41577,N_40002);
and U43117 (N_43117,N_41358,N_42340);
or U43118 (N_43118,N_42148,N_41407);
nor U43119 (N_43119,N_40407,N_40072);
nor U43120 (N_43120,N_41137,N_40562);
xnor U43121 (N_43121,N_40006,N_41645);
nand U43122 (N_43122,N_40431,N_40414);
nor U43123 (N_43123,N_41037,N_42128);
or U43124 (N_43124,N_40179,N_40846);
or U43125 (N_43125,N_41096,N_41815);
nor U43126 (N_43126,N_40353,N_41557);
nor U43127 (N_43127,N_40629,N_42120);
xor U43128 (N_43128,N_41181,N_40862);
nor U43129 (N_43129,N_41979,N_40600);
and U43130 (N_43130,N_41822,N_41688);
or U43131 (N_43131,N_40607,N_40108);
xnor U43132 (N_43132,N_40763,N_42471);
or U43133 (N_43133,N_40003,N_41919);
xnor U43134 (N_43134,N_41672,N_40858);
and U43135 (N_43135,N_42019,N_42327);
xnor U43136 (N_43136,N_40684,N_40712);
xor U43137 (N_43137,N_41296,N_40802);
nand U43138 (N_43138,N_41484,N_41258);
and U43139 (N_43139,N_40140,N_41452);
nor U43140 (N_43140,N_41720,N_40746);
and U43141 (N_43141,N_40400,N_40166);
nand U43142 (N_43142,N_42074,N_40368);
and U43143 (N_43143,N_41696,N_40047);
and U43144 (N_43144,N_40546,N_41435);
nor U43145 (N_43145,N_42446,N_40232);
or U43146 (N_43146,N_40784,N_40195);
or U43147 (N_43147,N_40310,N_41294);
xor U43148 (N_43148,N_41369,N_41185);
or U43149 (N_43149,N_41705,N_40987);
and U43150 (N_43150,N_42273,N_41263);
nand U43151 (N_43151,N_41894,N_40073);
xnor U43152 (N_43152,N_42116,N_40574);
and U43153 (N_43153,N_40685,N_41964);
xnor U43154 (N_43154,N_41385,N_41411);
xor U43155 (N_43155,N_42107,N_42282);
or U43156 (N_43156,N_42255,N_41556);
xor U43157 (N_43157,N_41054,N_40408);
nand U43158 (N_43158,N_40422,N_42300);
and U43159 (N_43159,N_40725,N_41965);
and U43160 (N_43160,N_41497,N_41834);
and U43161 (N_43161,N_42362,N_41769);
nand U43162 (N_43162,N_40772,N_41002);
xnor U43163 (N_43163,N_40505,N_42020);
or U43164 (N_43164,N_41858,N_41580);
or U43165 (N_43165,N_41303,N_41103);
nand U43166 (N_43166,N_40730,N_42262);
and U43167 (N_43167,N_41836,N_41594);
and U43168 (N_43168,N_41752,N_40911);
or U43169 (N_43169,N_42291,N_40734);
xor U43170 (N_43170,N_42176,N_41531);
nor U43171 (N_43171,N_41737,N_42455);
nor U43172 (N_43172,N_40921,N_41722);
nor U43173 (N_43173,N_41410,N_41842);
or U43174 (N_43174,N_40670,N_40519);
xor U43175 (N_43175,N_40812,N_40845);
or U43176 (N_43176,N_42271,N_40025);
xor U43177 (N_43177,N_40395,N_40458);
and U43178 (N_43178,N_40912,N_42383);
and U43179 (N_43179,N_40418,N_40768);
nand U43180 (N_43180,N_40315,N_40501);
xor U43181 (N_43181,N_40874,N_42474);
xnor U43182 (N_43182,N_40350,N_41776);
nor U43183 (N_43183,N_40117,N_40356);
and U43184 (N_43184,N_42261,N_40221);
xnor U43185 (N_43185,N_41059,N_42288);
xor U43186 (N_43186,N_42088,N_42131);
nand U43187 (N_43187,N_40499,N_41322);
and U43188 (N_43188,N_40148,N_42289);
nor U43189 (N_43189,N_41587,N_40493);
or U43190 (N_43190,N_42056,N_41841);
nand U43191 (N_43191,N_40572,N_42124);
or U43192 (N_43192,N_41124,N_40988);
and U43193 (N_43193,N_40043,N_41949);
xor U43194 (N_43194,N_40474,N_42394);
nand U43195 (N_43195,N_40169,N_40951);
nand U43196 (N_43196,N_40096,N_40371);
or U43197 (N_43197,N_40528,N_42201);
or U43198 (N_43198,N_41162,N_41213);
and U43199 (N_43199,N_41510,N_41539);
nor U43200 (N_43200,N_41821,N_40551);
and U43201 (N_43201,N_40578,N_40925);
or U43202 (N_43202,N_40373,N_42332);
xnor U43203 (N_43203,N_41774,N_41657);
xor U43204 (N_43204,N_41975,N_41977);
or U43205 (N_43205,N_42166,N_41063);
xnor U43206 (N_43206,N_40336,N_41208);
nor U43207 (N_43207,N_41963,N_41370);
and U43208 (N_43208,N_42355,N_42313);
or U43209 (N_43209,N_42075,N_42493);
nor U43210 (N_43210,N_41888,N_41047);
xor U43211 (N_43211,N_40770,N_40717);
nor U43212 (N_43212,N_42314,N_40533);
and U43213 (N_43213,N_40885,N_41778);
xnor U43214 (N_43214,N_40744,N_40508);
nor U43215 (N_43215,N_40969,N_40200);
nor U43216 (N_43216,N_41023,N_40218);
nand U43217 (N_43217,N_41044,N_40321);
nor U43218 (N_43218,N_40700,N_41744);
or U43219 (N_43219,N_40051,N_40394);
xor U43220 (N_43220,N_41191,N_41480);
and U43221 (N_43221,N_40340,N_41421);
nand U43222 (N_43222,N_40773,N_41025);
and U43223 (N_43223,N_41583,N_41108);
and U43224 (N_43224,N_41719,N_41352);
nand U43225 (N_43225,N_40834,N_42499);
or U43226 (N_43226,N_41654,N_41651);
nand U43227 (N_43227,N_41532,N_41809);
nand U43228 (N_43228,N_40239,N_42035);
nand U43229 (N_43229,N_40227,N_41033);
nand U43230 (N_43230,N_40977,N_40296);
nand U43231 (N_43231,N_40518,N_40064);
nor U43232 (N_43232,N_42003,N_41437);
and U43233 (N_43233,N_40041,N_42411);
or U43234 (N_43234,N_40297,N_41966);
and U43235 (N_43235,N_42027,N_40966);
xnor U43236 (N_43236,N_41757,N_40653);
xor U43237 (N_43237,N_42435,N_42482);
and U43238 (N_43238,N_41446,N_41529);
nor U43239 (N_43239,N_41127,N_40456);
and U43240 (N_43240,N_41564,N_41926);
nor U43241 (N_43241,N_40751,N_41584);
and U43242 (N_43242,N_40153,N_42423);
xor U43243 (N_43243,N_41513,N_42031);
or U43244 (N_43244,N_40517,N_40614);
nand U43245 (N_43245,N_41938,N_41995);
and U43246 (N_43246,N_40888,N_40665);
and U43247 (N_43247,N_41749,N_42301);
nand U43248 (N_43248,N_42392,N_42105);
or U43249 (N_43249,N_40990,N_40388);
and U43250 (N_43250,N_41348,N_40853);
nand U43251 (N_43251,N_42097,N_42161);
xor U43252 (N_43252,N_40613,N_40246);
nand U43253 (N_43253,N_41916,N_41830);
nor U43254 (N_43254,N_41520,N_40889);
xnor U43255 (N_43255,N_40511,N_40449);
and U43256 (N_43256,N_41380,N_41723);
nand U43257 (N_43257,N_42011,N_40039);
nand U43258 (N_43258,N_40882,N_41503);
or U43259 (N_43259,N_40125,N_42115);
nand U43260 (N_43260,N_40495,N_42225);
xor U43261 (N_43261,N_41618,N_41895);
and U43262 (N_43262,N_40870,N_42229);
or U43263 (N_43263,N_40211,N_41717);
and U43264 (N_43264,N_41637,N_42221);
xor U43265 (N_43265,N_40741,N_41408);
or U43266 (N_43266,N_41904,N_41075);
or U43267 (N_43267,N_40952,N_40249);
or U43268 (N_43268,N_40930,N_42165);
nand U43269 (N_43269,N_41558,N_42479);
nand U43270 (N_43270,N_41376,N_40074);
or U43271 (N_43271,N_42066,N_40429);
or U43272 (N_43272,N_40445,N_40344);
nor U43273 (N_43273,N_42341,N_41396);
nor U43274 (N_43274,N_40217,N_41924);
or U43275 (N_43275,N_40536,N_40659);
nand U43276 (N_43276,N_41158,N_41431);
or U43277 (N_43277,N_41082,N_40547);
or U43278 (N_43278,N_40333,N_41457);
nor U43279 (N_43279,N_40500,N_41439);
and U43280 (N_43280,N_41000,N_40205);
or U43281 (N_43281,N_40163,N_41969);
nor U43282 (N_43282,N_40397,N_42281);
or U43283 (N_43283,N_42364,N_40650);
nand U43284 (N_43284,N_41427,N_41507);
nand U43285 (N_43285,N_40855,N_41661);
or U43286 (N_43286,N_41174,N_42052);
nor U43287 (N_43287,N_40438,N_40516);
and U43288 (N_43288,N_40248,N_40502);
or U43289 (N_43289,N_40886,N_40213);
or U43290 (N_43290,N_42053,N_42322);
and U43291 (N_43291,N_42231,N_41579);
and U43292 (N_43292,N_40804,N_41125);
xnor U43293 (N_43293,N_41328,N_40680);
or U43294 (N_43294,N_40058,N_42315);
and U43295 (N_43295,N_40757,N_40263);
nand U43296 (N_43296,N_41112,N_41638);
nor U43297 (N_43297,N_41377,N_40512);
or U43298 (N_43298,N_41084,N_40237);
nand U43299 (N_43299,N_40766,N_42234);
and U43300 (N_43300,N_41309,N_40087);
xor U43301 (N_43301,N_40139,N_41473);
nand U43302 (N_43302,N_41905,N_40111);
nand U43303 (N_43303,N_41676,N_40947);
or U43304 (N_43304,N_41632,N_42419);
or U43305 (N_43305,N_41937,N_41071);
nor U43306 (N_43306,N_41195,N_40026);
xnor U43307 (N_43307,N_41947,N_40621);
xnor U43308 (N_43308,N_41750,N_40022);
and U43309 (N_43309,N_40869,N_41107);
nand U43310 (N_43310,N_41307,N_41403);
and U43311 (N_43311,N_42200,N_41519);
xor U43312 (N_43312,N_41463,N_41081);
and U43313 (N_43313,N_40797,N_41971);
nor U43314 (N_43314,N_40052,N_40890);
or U43315 (N_43315,N_42492,N_40566);
and U43316 (N_43316,N_40082,N_41342);
or U43317 (N_43317,N_40585,N_40994);
and U43318 (N_43318,N_42169,N_41860);
nor U43319 (N_43319,N_41144,N_41180);
and U43320 (N_43320,N_40720,N_41360);
and U43321 (N_43321,N_41343,N_41592);
nor U43322 (N_43322,N_40377,N_41968);
xor U43323 (N_43323,N_42174,N_42424);
or U43324 (N_43324,N_41018,N_42346);
and U43325 (N_43325,N_42181,N_41134);
xor U43326 (N_43326,N_40755,N_42441);
and U43327 (N_43327,N_41656,N_40875);
or U43328 (N_43328,N_40417,N_42223);
xor U43329 (N_43329,N_40949,N_40540);
and U43330 (N_43330,N_41064,N_40285);
xor U43331 (N_43331,N_40436,N_41586);
and U43332 (N_43332,N_40695,N_40475);
nand U43333 (N_43333,N_40326,N_41444);
nand U43334 (N_43334,N_42122,N_42159);
and U43335 (N_43335,N_40491,N_41088);
xnor U43336 (N_43336,N_41392,N_41943);
nand U43337 (N_43337,N_41353,N_40081);
xnor U43338 (N_43338,N_40856,N_41325);
xnor U43339 (N_43339,N_40998,N_42426);
nor U43340 (N_43340,N_41595,N_40646);
and U43341 (N_43341,N_41384,N_41518);
nor U43342 (N_43342,N_40184,N_42005);
nor U43343 (N_43343,N_40327,N_40267);
and U43344 (N_43344,N_40172,N_40522);
or U43345 (N_43345,N_41902,N_40446);
nor U43346 (N_43346,N_40866,N_42126);
xnor U43347 (N_43347,N_40175,N_40272);
and U43348 (N_43348,N_41471,N_41363);
nand U43349 (N_43349,N_41132,N_40954);
and U43350 (N_43350,N_41034,N_42193);
and U43351 (N_43351,N_42063,N_42032);
nand U43352 (N_43352,N_40606,N_41277);
nor U43353 (N_43353,N_42013,N_42050);
and U43354 (N_43354,N_40932,N_41021);
nor U43355 (N_43355,N_40302,N_42151);
xor U43356 (N_43356,N_42129,N_41746);
nor U43357 (N_43357,N_42167,N_40078);
and U43358 (N_43358,N_42149,N_40124);
xor U43359 (N_43359,N_42082,N_41031);
xor U43360 (N_43360,N_40244,N_42334);
nand U43361 (N_43361,N_42457,N_41599);
nor U43362 (N_43362,N_41870,N_42004);
nor U43363 (N_43363,N_41249,N_40464);
nand U43364 (N_43364,N_41470,N_41709);
and U43365 (N_43365,N_40141,N_41292);
and U43366 (N_43366,N_40284,N_41222);
or U43367 (N_43367,N_41271,N_42331);
and U43368 (N_43368,N_40534,N_41276);
nor U43369 (N_43369,N_41652,N_40897);
and U43370 (N_43370,N_41078,N_40345);
xor U43371 (N_43371,N_41972,N_40167);
and U43372 (N_43372,N_41847,N_42111);
or U43373 (N_43373,N_40928,N_42251);
or U43374 (N_43374,N_41387,N_42399);
or U43375 (N_43375,N_40174,N_40116);
or U43376 (N_43376,N_40498,N_40907);
xnor U43377 (N_43377,N_41759,N_40189);
and U43378 (N_43378,N_42098,N_42306);
xnor U43379 (N_43379,N_40273,N_41804);
xor U43380 (N_43380,N_40387,N_40847);
nand U43381 (N_43381,N_40206,N_40457);
or U43382 (N_43382,N_41613,N_40743);
nand U43383 (N_43383,N_41092,N_41878);
and U43384 (N_43384,N_40833,N_41600);
xor U43385 (N_43385,N_40832,N_42357);
or U43386 (N_43386,N_41261,N_41664);
and U43387 (N_43387,N_41691,N_42162);
nor U43388 (N_43388,N_40655,N_40762);
nand U43389 (N_43389,N_40479,N_41178);
and U43390 (N_43390,N_41585,N_42173);
xnor U43391 (N_43391,N_41211,N_42242);
xor U43392 (N_43392,N_40780,N_40004);
nor U43393 (N_43393,N_42438,N_41960);
or U43394 (N_43394,N_41627,N_40355);
nand U43395 (N_43395,N_40201,N_41235);
and U43396 (N_43396,N_42431,N_41442);
nor U43397 (N_43397,N_41126,N_41606);
or U43398 (N_43398,N_40686,N_40597);
or U43399 (N_43399,N_40661,N_41917);
or U43400 (N_43400,N_42062,N_40318);
nor U43401 (N_43401,N_40347,N_42304);
nor U43402 (N_43402,N_41533,N_42319);
and U43403 (N_43403,N_41819,N_41909);
and U43404 (N_43404,N_41869,N_41196);
xnor U43405 (N_43405,N_42369,N_42393);
nand U43406 (N_43406,N_40662,N_41024);
nand U43407 (N_43407,N_41537,N_41732);
and U43408 (N_43408,N_41188,N_41321);
or U43409 (N_43409,N_40224,N_41311);
nor U43410 (N_43410,N_41316,N_40920);
and U43411 (N_43411,N_42093,N_41571);
nand U43412 (N_43412,N_40133,N_42451);
nand U43413 (N_43413,N_40173,N_40974);
and U43414 (N_43414,N_42001,N_42092);
and U43415 (N_43415,N_40007,N_41315);
or U43416 (N_43416,N_41003,N_41141);
nand U43417 (N_43417,N_41006,N_41553);
xnor U43418 (N_43418,N_42309,N_40000);
xor U43419 (N_43419,N_40257,N_41074);
nor U43420 (N_43420,N_40698,N_41607);
nand U43421 (N_43421,N_41933,N_41168);
and U43422 (N_43422,N_41550,N_40701);
or U43423 (N_43423,N_42185,N_41854);
or U43424 (N_43424,N_42294,N_42373);
and U43425 (N_43425,N_41506,N_41194);
and U43426 (N_43426,N_41285,N_40448);
and U43427 (N_43427,N_40971,N_41040);
xor U43428 (N_43428,N_40226,N_41135);
nand U43429 (N_43429,N_41541,N_42044);
nand U43430 (N_43430,N_40673,N_40402);
and U43431 (N_43431,N_41204,N_40891);
nand U43432 (N_43432,N_41148,N_42418);
nor U43433 (N_43433,N_40702,N_41097);
nor U43434 (N_43434,N_40950,N_42102);
or U43435 (N_43435,N_40642,N_41650);
and U43436 (N_43436,N_40736,N_40403);
nor U43437 (N_43437,N_41156,N_41980);
nand U43438 (N_43438,N_40963,N_41467);
nand U43439 (N_43439,N_42140,N_40228);
xnor U43440 (N_43440,N_41622,N_42448);
nor U43441 (N_43441,N_40076,N_41016);
or U43442 (N_43442,N_40398,N_41724);
nor U43443 (N_43443,N_41552,N_41486);
and U43444 (N_43444,N_40732,N_40943);
or U43445 (N_43445,N_42303,N_41218);
xor U43446 (N_43446,N_42250,N_41704);
xor U43447 (N_43447,N_42150,N_42370);
nor U43448 (N_43448,N_40293,N_40774);
nor U43449 (N_43449,N_41504,N_40892);
nand U43450 (N_43450,N_41013,N_42395);
and U43451 (N_43451,N_41139,N_41409);
xnor U43452 (N_43452,N_40972,N_42215);
nand U43453 (N_43453,N_40531,N_40138);
nand U43454 (N_43454,N_40196,N_41811);
xor U43455 (N_43455,N_41521,N_41742);
nor U43456 (N_43456,N_41840,N_40904);
xnor U43457 (N_43457,N_40824,N_40583);
or U43458 (N_43458,N_41862,N_42263);
nand U43459 (N_43459,N_41621,N_40535);
nand U43460 (N_43460,N_42472,N_42227);
nand U43461 (N_43461,N_42156,N_42361);
nand U43462 (N_43462,N_40018,N_41453);
nor U43463 (N_43463,N_41500,N_41120);
nor U43464 (N_43464,N_41182,N_41508);
xnor U43465 (N_43465,N_41055,N_42428);
nor U43466 (N_43466,N_41485,N_41921);
or U43467 (N_43467,N_40929,N_41620);
xnor U43468 (N_43468,N_41920,N_42272);
nand U43469 (N_43469,N_40463,N_42015);
xnor U43470 (N_43470,N_40796,N_40960);
and U43471 (N_43471,N_40826,N_40787);
or U43472 (N_43472,N_40168,N_41167);
xnor U43473 (N_43473,N_41237,N_42217);
nor U43474 (N_43474,N_41418,N_42253);
nor U43475 (N_43475,N_40230,N_40447);
nand U43476 (N_43476,N_42350,N_41320);
nand U43477 (N_43477,N_42293,N_41942);
nor U43478 (N_43478,N_40354,N_40801);
nor U43479 (N_43479,N_41871,N_40329);
xor U43480 (N_43480,N_41782,N_42218);
nand U43481 (N_43481,N_41436,N_41699);
xnor U43482 (N_43482,N_40277,N_41758);
nor U43483 (N_43483,N_41867,N_40822);
nor U43484 (N_43484,N_40322,N_40697);
xor U43485 (N_43485,N_40823,N_40873);
nor U43486 (N_43486,N_41165,N_42360);
xnor U43487 (N_43487,N_41879,N_41067);
nand U43488 (N_43488,N_40800,N_40513);
nand U43489 (N_43489,N_42478,N_40050);
or U43490 (N_43490,N_40690,N_41087);
and U43491 (N_43491,N_40146,N_41630);
nor U43492 (N_43492,N_40128,N_42091);
or U43493 (N_43493,N_41414,N_42043);
xnor U43494 (N_43494,N_42153,N_41027);
or U43495 (N_43495,N_40084,N_41217);
and U43496 (N_43496,N_40956,N_42365);
xnor U43497 (N_43497,N_40381,N_41642);
and U43498 (N_43498,N_42078,N_40042);
nand U43499 (N_43499,N_40100,N_41693);
nor U43500 (N_43500,N_41252,N_42323);
xor U43501 (N_43501,N_41646,N_42484);
nand U43502 (N_43502,N_40450,N_41993);
xor U43503 (N_43503,N_40909,N_42180);
nand U43504 (N_43504,N_41419,N_41301);
nor U43505 (N_43505,N_40343,N_42333);
xor U43506 (N_43506,N_40896,N_41855);
xnor U43507 (N_43507,N_41014,N_40756);
and U43508 (N_43508,N_40633,N_42136);
or U43509 (N_43509,N_41259,N_41337);
nor U43510 (N_43510,N_41479,N_40416);
or U43511 (N_43511,N_41389,N_40309);
nand U43512 (N_43512,N_41788,N_41281);
and U43513 (N_43513,N_40553,N_40924);
nor U43514 (N_43514,N_42285,N_40208);
and U43515 (N_43515,N_41616,N_42046);
nand U43516 (N_43516,N_41295,N_40393);
nor U43517 (N_43517,N_40056,N_41653);
and U43518 (N_43518,N_41687,N_40379);
nor U43519 (N_43519,N_42437,N_41560);
nand U43520 (N_43520,N_40027,N_42445);
or U43521 (N_43521,N_40731,N_40459);
nand U43522 (N_43522,N_41848,N_41604);
xor U43523 (N_43523,N_42377,N_41934);
and U43524 (N_43524,N_41747,N_42233);
nand U43525 (N_43525,N_40242,N_40234);
or U43526 (N_43526,N_41244,N_41171);
nand U43527 (N_43527,N_40106,N_41346);
nor U43528 (N_43528,N_41710,N_41679);
or U43529 (N_43529,N_41028,N_42040);
or U43530 (N_43530,N_40504,N_41393);
xnor U43531 (N_43531,N_42265,N_40413);
or U43532 (N_43532,N_41570,N_40565);
xor U43533 (N_43533,N_42220,N_41959);
nand U43534 (N_43534,N_40409,N_41205);
nand U43535 (N_43535,N_41565,N_41397);
nand U43536 (N_43536,N_41548,N_41982);
and U43537 (N_43537,N_41800,N_41113);
nor U43538 (N_43538,N_41406,N_41109);
or U43539 (N_43539,N_40470,N_40118);
nor U43540 (N_43540,N_41540,N_42382);
nor U43541 (N_43541,N_41347,N_41142);
xor U43542 (N_43542,N_40737,N_40490);
or U43543 (N_43543,N_41432,N_40465);
and U43544 (N_43544,N_41383,N_42311);
nand U43545 (N_43545,N_42427,N_41779);
or U43546 (N_43546,N_41610,N_42016);
nand U43547 (N_43547,N_41286,N_42195);
and U43548 (N_43548,N_41499,N_40871);
nor U43549 (N_43549,N_41423,N_41957);
nand U43550 (N_43550,N_40094,N_42287);
and U43551 (N_43551,N_41715,N_40068);
xor U43552 (N_43552,N_40964,N_41636);
and U43553 (N_43553,N_40396,N_40676);
nand U43554 (N_43554,N_40542,N_41402);
nor U43555 (N_43555,N_40197,N_40055);
xor U43556 (N_43556,N_41754,N_41817);
and U43557 (N_43557,N_42249,N_40530);
xor U43558 (N_43558,N_42376,N_42049);
and U43559 (N_43559,N_40306,N_40593);
and U43560 (N_43560,N_41837,N_42101);
nand U43561 (N_43561,N_41930,N_41459);
nor U43562 (N_43562,N_41101,N_40127);
xnor U43563 (N_43563,N_40917,N_41119);
or U43564 (N_43564,N_40177,N_41373);
nand U43565 (N_43565,N_41065,N_40724);
or U43566 (N_43566,N_40682,N_40895);
nor U43567 (N_43567,N_41130,N_41372);
xor U43568 (N_43568,N_40276,N_40030);
and U43569 (N_43569,N_40480,N_41898);
xnor U43570 (N_43570,N_40390,N_42057);
nand U43571 (N_43571,N_40764,N_40151);
and U43572 (N_43572,N_41429,N_41846);
nor U43573 (N_43573,N_40745,N_40668);
or U43574 (N_43574,N_41345,N_41633);
and U43575 (N_43575,N_42095,N_40010);
xor U43576 (N_43576,N_40157,N_41229);
nor U43577 (N_43577,N_40451,N_40667);
or U43578 (N_43578,N_41201,N_41789);
and U43579 (N_43579,N_41177,N_40432);
xnor U43580 (N_43580,N_40515,N_41712);
nand U43581 (N_43581,N_40973,N_40674);
or U43582 (N_43582,N_40626,N_41810);
nor U43583 (N_43583,N_40466,N_41219);
nand U43584 (N_43584,N_42177,N_41488);
xnor U43585 (N_43585,N_40019,N_41458);
nor U43586 (N_43586,N_41287,N_40054);
or U43587 (N_43587,N_40721,N_42143);
and U43588 (N_43588,N_40053,N_40992);
nor U43589 (N_43589,N_42060,N_42237);
nand U43590 (N_43590,N_40876,N_40142);
xnor U43591 (N_43591,N_40067,N_41438);
or U43592 (N_43592,N_42252,N_40147);
nand U43593 (N_43593,N_42280,N_42410);
xnor U43594 (N_43594,N_40435,N_42260);
or U43595 (N_43595,N_41659,N_40372);
nor U43596 (N_43596,N_40287,N_41129);
or U43597 (N_43597,N_41785,N_42145);
nand U43598 (N_43598,N_40604,N_40894);
or U43599 (N_43599,N_40477,N_42416);
and U43600 (N_43600,N_41726,N_40488);
nand U43601 (N_43601,N_40253,N_40941);
nor U43602 (N_43602,N_42033,N_40497);
xor U43603 (N_43603,N_42157,N_41832);
and U43604 (N_43604,N_40426,N_40577);
nand U43605 (N_43605,N_40609,N_42329);
xor U43606 (N_43606,N_41608,N_40192);
xor U43607 (N_43607,N_40126,N_41753);
nor U43608 (N_43608,N_40840,N_40312);
and U43609 (N_43609,N_40798,N_42024);
or U43610 (N_43610,N_40384,N_40210);
or U43611 (N_43611,N_40579,N_40658);
nor U43612 (N_43612,N_41561,N_41091);
nand U43613 (N_43613,N_40352,N_41666);
xnor U43614 (N_43614,N_40486,N_41931);
xnor U43615 (N_43615,N_40584,N_41767);
and U43616 (N_43616,N_40364,N_42328);
or U43617 (N_43617,N_40748,N_40828);
and U43618 (N_43618,N_40307,N_40385);
nand U43619 (N_43619,N_41150,N_40931);
xnor U43620 (N_43620,N_41474,N_40256);
nor U43621 (N_43621,N_42402,N_41498);
nor U43622 (N_43622,N_41241,N_41187);
or U43623 (N_43623,N_42117,N_40769);
nor U43624 (N_43624,N_41524,N_40494);
or U43625 (N_43625,N_41338,N_41967);
or U43626 (N_43626,N_41536,N_41308);
nand U43627 (N_43627,N_40005,N_41242);
or U43628 (N_43628,N_41095,N_42292);
and U43629 (N_43629,N_41365,N_41478);
or U43630 (N_43630,N_41080,N_41430);
nand U43631 (N_43631,N_41675,N_40467);
nand U43632 (N_43632,N_42480,N_40031);
nand U43633 (N_43633,N_42429,N_40708);
xor U43634 (N_43634,N_42130,N_41741);
nand U43635 (N_43635,N_41001,N_42456);
nor U43636 (N_43636,N_41773,N_40366);
nand U43637 (N_43637,N_40910,N_42191);
nand U43638 (N_43638,N_42283,N_41374);
and U43639 (N_43639,N_40639,N_41339);
xor U43640 (N_43640,N_41186,N_40182);
xor U43641 (N_43641,N_42170,N_41122);
and U43642 (N_43642,N_40170,N_41598);
or U43643 (N_43643,N_41655,N_40602);
nand U43644 (N_43644,N_41593,N_41401);
nand U43645 (N_43645,N_40013,N_40548);
or U43646 (N_43646,N_42465,N_41908);
nand U43647 (N_43647,N_41482,N_41954);
nor U43648 (N_43648,N_40104,N_41004);
xor U43649 (N_43649,N_41323,N_40935);
and U43650 (N_43650,N_40623,N_42486);
nand U43651 (N_43651,N_42496,N_41578);
nand U43652 (N_43652,N_41945,N_41925);
nor U43653 (N_43653,N_40269,N_40034);
and U43654 (N_43654,N_41105,N_40817);
xor U43655 (N_43655,N_41772,N_41987);
nor U43656 (N_43656,N_42330,N_42071);
and U43657 (N_43657,N_40754,N_40738);
xor U43658 (N_43658,N_41330,N_40902);
nor U43659 (N_43659,N_40114,N_40107);
nor U43660 (N_43660,N_40848,N_40995);
xor U43661 (N_43661,N_40980,N_40191);
and U43662 (N_43662,N_42344,N_41994);
nand U43663 (N_43663,N_42037,N_40759);
nor U43664 (N_43664,N_42430,N_40696);
or U43665 (N_43665,N_40742,N_42241);
and U43666 (N_43666,N_40271,N_41036);
and U43667 (N_43667,N_40760,N_41319);
nand U43668 (N_43668,N_40678,N_41588);
or U43669 (N_43669,N_40863,N_42356);
and U43670 (N_43670,N_40934,N_41424);
nand U43671 (N_43671,N_41455,N_41629);
nor U43672 (N_43672,N_41304,N_40357);
xnor U43673 (N_43673,N_40775,N_41997);
xor U43674 (N_43674,N_42125,N_41805);
or U43675 (N_43675,N_41988,N_40545);
xor U43676 (N_43676,N_40603,N_41913);
nor U43677 (N_43677,N_41626,N_40338);
nor U43678 (N_43678,N_40261,N_41426);
or U43679 (N_43679,N_42458,N_40319);
and U43680 (N_43680,N_42198,N_41684);
xnor U43681 (N_43681,N_42213,N_40008);
nor U43682 (N_43682,N_41761,N_41877);
nand U43683 (N_43683,N_41011,N_41215);
nand U43684 (N_43684,N_41690,N_40305);
nand U43685 (N_43685,N_40857,N_41416);
or U43686 (N_43686,N_41246,N_41495);
nor U43687 (N_43687,N_41827,N_40827);
or U43688 (N_43688,N_40666,N_41152);
nand U43689 (N_43689,N_40810,N_41680);
nand U43690 (N_43690,N_40644,N_42154);
or U43691 (N_43691,N_41989,N_41771);
or U43692 (N_43692,N_40525,N_42196);
xor U43693 (N_43693,N_40129,N_42135);
nand U43694 (N_43694,N_40282,N_40795);
or U43695 (N_43695,N_41685,N_41662);
or U43696 (N_43696,N_42007,N_42353);
nor U43697 (N_43697,N_42375,N_41738);
or U43698 (N_43698,N_42268,N_40433);
or U43699 (N_43699,N_42142,N_41708);
or U43700 (N_43700,N_40298,N_40066);
and U43701 (N_43701,N_42029,N_40761);
nand U43702 (N_43702,N_42214,N_40001);
or U43703 (N_43703,N_41984,N_41133);
nand U43704 (N_43704,N_41225,N_41170);
and U43705 (N_43705,N_41017,N_41228);
or U43706 (N_43706,N_41703,N_40088);
xnor U43707 (N_43707,N_42320,N_41102);
nand U43708 (N_43708,N_41932,N_41214);
nand U43709 (N_43709,N_41070,N_42083);
xnor U43710 (N_43710,N_41512,N_40380);
xnor U43711 (N_43711,N_41146,N_42202);
xnor U43712 (N_43712,N_40942,N_41149);
xor U43713 (N_43713,N_41796,N_41996);
nor U43714 (N_43714,N_40829,N_40558);
nor U43715 (N_43715,N_41838,N_41689);
nand U43716 (N_43716,N_40035,N_42147);
nand U43717 (N_43717,N_41551,N_41310);
xor U43718 (N_43718,N_41501,N_41770);
or U43719 (N_43719,N_41668,N_42421);
nor U43720 (N_43720,N_40425,N_42398);
nand U43721 (N_43721,N_40549,N_41236);
xor U43722 (N_43722,N_42286,N_40303);
nor U43723 (N_43723,N_40767,N_41043);
or U43724 (N_43724,N_40439,N_41428);
xor U43725 (N_43725,N_41042,N_42417);
and U43726 (N_43726,N_40571,N_42358);
nand U43727 (N_43727,N_41050,N_40740);
nor U43728 (N_43728,N_41395,N_42406);
xor U43729 (N_43729,N_42006,N_41166);
nand U43730 (N_43730,N_41714,N_41683);
nand U43731 (N_43731,N_40009,N_42014);
and U43732 (N_43732,N_42495,N_40032);
xor U43733 (N_43733,N_40325,N_40158);
nor U43734 (N_43734,N_42104,N_40916);
and U43735 (N_43735,N_40176,N_41927);
nor U43736 (N_43736,N_41349,N_41872);
and U43737 (N_43737,N_42086,N_41527);
nand U43738 (N_43738,N_40616,N_42192);
nor U43739 (N_43739,N_40461,N_41417);
and U43740 (N_43740,N_41559,N_40957);
and U43741 (N_43741,N_40452,N_41808);
or U43742 (N_43742,N_41412,N_40024);
nand U43743 (N_43743,N_42207,N_40215);
nand U43744 (N_43744,N_40037,N_40314);
nand U43745 (N_43745,N_40865,N_40711);
or U43746 (N_43746,N_42295,N_41483);
nor U43747 (N_43747,N_40348,N_40376);
nor U43748 (N_43748,N_42203,N_41172);
nor U43749 (N_43749,N_42204,N_41535);
or U43750 (N_43750,N_42246,N_42428);
nand U43751 (N_43751,N_42215,N_41392);
xnor U43752 (N_43752,N_40408,N_40806);
xnor U43753 (N_43753,N_41259,N_40435);
or U43754 (N_43754,N_41142,N_42141);
nand U43755 (N_43755,N_41908,N_40739);
nand U43756 (N_43756,N_42111,N_41851);
nand U43757 (N_43757,N_41041,N_42120);
nor U43758 (N_43758,N_42456,N_41537);
or U43759 (N_43759,N_40170,N_40808);
and U43760 (N_43760,N_42048,N_41827);
nor U43761 (N_43761,N_41666,N_41072);
xor U43762 (N_43762,N_40336,N_41616);
nor U43763 (N_43763,N_42270,N_41622);
or U43764 (N_43764,N_42344,N_42245);
and U43765 (N_43765,N_40235,N_41691);
xnor U43766 (N_43766,N_42078,N_40033);
nor U43767 (N_43767,N_42457,N_40463);
or U43768 (N_43768,N_41402,N_41719);
and U43769 (N_43769,N_42418,N_41953);
xor U43770 (N_43770,N_41794,N_42362);
nor U43771 (N_43771,N_40678,N_40339);
nand U43772 (N_43772,N_40026,N_40627);
and U43773 (N_43773,N_40534,N_42477);
nand U43774 (N_43774,N_41551,N_41288);
nor U43775 (N_43775,N_40738,N_41166);
nand U43776 (N_43776,N_42489,N_42373);
nand U43777 (N_43777,N_42375,N_42305);
nand U43778 (N_43778,N_40264,N_40384);
or U43779 (N_43779,N_42008,N_40908);
and U43780 (N_43780,N_40276,N_40654);
and U43781 (N_43781,N_40417,N_42218);
nand U43782 (N_43782,N_42378,N_41239);
nand U43783 (N_43783,N_40428,N_40549);
or U43784 (N_43784,N_41427,N_41270);
nand U43785 (N_43785,N_40738,N_42102);
or U43786 (N_43786,N_40303,N_40909);
nand U43787 (N_43787,N_41262,N_41632);
nor U43788 (N_43788,N_41152,N_42238);
xnor U43789 (N_43789,N_42193,N_41122);
or U43790 (N_43790,N_41233,N_42075);
nor U43791 (N_43791,N_40540,N_41307);
xor U43792 (N_43792,N_42269,N_41027);
or U43793 (N_43793,N_41306,N_41102);
nor U43794 (N_43794,N_42496,N_40295);
nand U43795 (N_43795,N_40027,N_42266);
nand U43796 (N_43796,N_41495,N_41536);
xor U43797 (N_43797,N_41250,N_41565);
and U43798 (N_43798,N_42146,N_41876);
nor U43799 (N_43799,N_42493,N_40258);
xnor U43800 (N_43800,N_40093,N_42486);
xor U43801 (N_43801,N_41806,N_41485);
nor U43802 (N_43802,N_41020,N_41756);
nand U43803 (N_43803,N_40440,N_41484);
and U43804 (N_43804,N_41176,N_40103);
and U43805 (N_43805,N_41742,N_42197);
nand U43806 (N_43806,N_40287,N_41028);
nor U43807 (N_43807,N_41608,N_40014);
nand U43808 (N_43808,N_40225,N_41432);
nor U43809 (N_43809,N_41936,N_42208);
or U43810 (N_43810,N_40049,N_42426);
nand U43811 (N_43811,N_41089,N_40402);
nor U43812 (N_43812,N_41936,N_40691);
xnor U43813 (N_43813,N_42425,N_41882);
or U43814 (N_43814,N_40532,N_41108);
nand U43815 (N_43815,N_42095,N_40434);
or U43816 (N_43816,N_41679,N_40867);
or U43817 (N_43817,N_40747,N_41571);
or U43818 (N_43818,N_42445,N_40407);
and U43819 (N_43819,N_41290,N_40473);
nor U43820 (N_43820,N_42273,N_41353);
xor U43821 (N_43821,N_41526,N_42003);
or U43822 (N_43822,N_40615,N_41052);
or U43823 (N_43823,N_42024,N_41836);
xnor U43824 (N_43824,N_40737,N_40114);
and U43825 (N_43825,N_42257,N_40748);
nand U43826 (N_43826,N_42447,N_40532);
xor U43827 (N_43827,N_41778,N_41207);
or U43828 (N_43828,N_41915,N_40784);
or U43829 (N_43829,N_40974,N_40105);
nor U43830 (N_43830,N_40615,N_41965);
or U43831 (N_43831,N_40848,N_41516);
nand U43832 (N_43832,N_40989,N_40607);
xnor U43833 (N_43833,N_42367,N_40482);
or U43834 (N_43834,N_40688,N_41163);
nor U43835 (N_43835,N_42273,N_41673);
xor U43836 (N_43836,N_40487,N_41225);
and U43837 (N_43837,N_40564,N_40444);
nor U43838 (N_43838,N_41127,N_41806);
nand U43839 (N_43839,N_41585,N_41446);
xor U43840 (N_43840,N_40139,N_40278);
nor U43841 (N_43841,N_41189,N_41292);
nor U43842 (N_43842,N_42346,N_40146);
nor U43843 (N_43843,N_40285,N_41914);
and U43844 (N_43844,N_40383,N_42323);
xnor U43845 (N_43845,N_40830,N_40457);
xor U43846 (N_43846,N_40580,N_40090);
nand U43847 (N_43847,N_40073,N_42262);
xor U43848 (N_43848,N_42387,N_40082);
nor U43849 (N_43849,N_40568,N_42227);
xnor U43850 (N_43850,N_42484,N_41745);
and U43851 (N_43851,N_41773,N_40786);
nand U43852 (N_43852,N_41423,N_42095);
xor U43853 (N_43853,N_41338,N_40393);
nor U43854 (N_43854,N_42132,N_41537);
or U43855 (N_43855,N_42092,N_41155);
nand U43856 (N_43856,N_41157,N_40945);
xnor U43857 (N_43857,N_40492,N_41568);
or U43858 (N_43858,N_40202,N_40863);
xor U43859 (N_43859,N_40092,N_40711);
nor U43860 (N_43860,N_41499,N_40980);
and U43861 (N_43861,N_41889,N_41741);
nand U43862 (N_43862,N_41318,N_41556);
xnor U43863 (N_43863,N_42490,N_40227);
or U43864 (N_43864,N_41452,N_40538);
or U43865 (N_43865,N_40182,N_42304);
nor U43866 (N_43866,N_42301,N_41661);
xor U43867 (N_43867,N_40181,N_40359);
nor U43868 (N_43868,N_40931,N_41183);
nand U43869 (N_43869,N_41029,N_40231);
xnor U43870 (N_43870,N_40312,N_41512);
nor U43871 (N_43871,N_40053,N_41698);
nor U43872 (N_43872,N_40851,N_40385);
and U43873 (N_43873,N_40415,N_40660);
or U43874 (N_43874,N_41922,N_40523);
or U43875 (N_43875,N_42184,N_40983);
nor U43876 (N_43876,N_41329,N_40906);
nand U43877 (N_43877,N_42475,N_42162);
or U43878 (N_43878,N_41920,N_42029);
nand U43879 (N_43879,N_40917,N_42333);
nand U43880 (N_43880,N_40596,N_41277);
nand U43881 (N_43881,N_41226,N_40175);
and U43882 (N_43882,N_40899,N_41657);
and U43883 (N_43883,N_41895,N_40602);
nand U43884 (N_43884,N_40172,N_41753);
nor U43885 (N_43885,N_40272,N_40120);
xnor U43886 (N_43886,N_40117,N_42082);
nand U43887 (N_43887,N_40966,N_40283);
nor U43888 (N_43888,N_40215,N_40619);
and U43889 (N_43889,N_40761,N_41082);
nor U43890 (N_43890,N_41366,N_41027);
or U43891 (N_43891,N_41145,N_41182);
or U43892 (N_43892,N_40736,N_41444);
or U43893 (N_43893,N_40248,N_41910);
and U43894 (N_43894,N_40651,N_41200);
and U43895 (N_43895,N_41336,N_41755);
nand U43896 (N_43896,N_40676,N_42280);
nand U43897 (N_43897,N_40119,N_40173);
or U43898 (N_43898,N_41637,N_41001);
and U43899 (N_43899,N_41178,N_41081);
xor U43900 (N_43900,N_41777,N_40204);
nand U43901 (N_43901,N_41317,N_40565);
nand U43902 (N_43902,N_42128,N_41378);
nand U43903 (N_43903,N_40770,N_40510);
nor U43904 (N_43904,N_40374,N_40250);
nor U43905 (N_43905,N_41356,N_40278);
or U43906 (N_43906,N_40626,N_40045);
nor U43907 (N_43907,N_40812,N_41888);
and U43908 (N_43908,N_41269,N_40016);
xnor U43909 (N_43909,N_42039,N_41746);
xor U43910 (N_43910,N_41943,N_41534);
xor U43911 (N_43911,N_42431,N_40534);
and U43912 (N_43912,N_42163,N_40522);
nor U43913 (N_43913,N_41560,N_42442);
and U43914 (N_43914,N_40488,N_41800);
or U43915 (N_43915,N_42473,N_41170);
and U43916 (N_43916,N_41328,N_41885);
nor U43917 (N_43917,N_40683,N_42185);
xor U43918 (N_43918,N_40768,N_40692);
xnor U43919 (N_43919,N_40175,N_40506);
nor U43920 (N_43920,N_41806,N_40093);
xor U43921 (N_43921,N_40076,N_41660);
or U43922 (N_43922,N_40469,N_41246);
nor U43923 (N_43923,N_40261,N_41594);
and U43924 (N_43924,N_40497,N_40000);
and U43925 (N_43925,N_40068,N_40829);
xnor U43926 (N_43926,N_40985,N_42486);
nor U43927 (N_43927,N_41350,N_41785);
nand U43928 (N_43928,N_42253,N_41818);
and U43929 (N_43929,N_40757,N_40255);
nand U43930 (N_43930,N_40020,N_41632);
or U43931 (N_43931,N_41492,N_40338);
xor U43932 (N_43932,N_40529,N_40321);
and U43933 (N_43933,N_42071,N_41701);
or U43934 (N_43934,N_40711,N_42056);
nand U43935 (N_43935,N_40977,N_40585);
and U43936 (N_43936,N_41832,N_40708);
nor U43937 (N_43937,N_40104,N_40312);
or U43938 (N_43938,N_42392,N_41870);
nand U43939 (N_43939,N_41648,N_41959);
nor U43940 (N_43940,N_40819,N_41460);
or U43941 (N_43941,N_40233,N_40212);
nor U43942 (N_43942,N_42493,N_40159);
nor U43943 (N_43943,N_41286,N_42293);
xnor U43944 (N_43944,N_42458,N_42354);
xor U43945 (N_43945,N_41995,N_40920);
xor U43946 (N_43946,N_41663,N_41947);
xor U43947 (N_43947,N_41499,N_40766);
and U43948 (N_43948,N_40147,N_40230);
nand U43949 (N_43949,N_42247,N_40867);
or U43950 (N_43950,N_41913,N_41546);
or U43951 (N_43951,N_41056,N_41778);
nand U43952 (N_43952,N_40534,N_41155);
and U43953 (N_43953,N_40906,N_41891);
nor U43954 (N_43954,N_40037,N_41185);
nor U43955 (N_43955,N_40741,N_40662);
and U43956 (N_43956,N_40281,N_41805);
xnor U43957 (N_43957,N_41280,N_40469);
or U43958 (N_43958,N_41315,N_40699);
and U43959 (N_43959,N_40729,N_41861);
nand U43960 (N_43960,N_42138,N_41969);
xnor U43961 (N_43961,N_40681,N_40395);
nand U43962 (N_43962,N_41293,N_42226);
nor U43963 (N_43963,N_42400,N_42232);
and U43964 (N_43964,N_40397,N_40423);
nor U43965 (N_43965,N_41794,N_41253);
or U43966 (N_43966,N_41967,N_41127);
and U43967 (N_43967,N_42334,N_40375);
or U43968 (N_43968,N_40708,N_41137);
or U43969 (N_43969,N_40834,N_40579);
and U43970 (N_43970,N_40618,N_40444);
or U43971 (N_43971,N_40786,N_40993);
xor U43972 (N_43972,N_40482,N_41438);
xnor U43973 (N_43973,N_42291,N_40542);
nor U43974 (N_43974,N_40399,N_40411);
xor U43975 (N_43975,N_40887,N_42322);
and U43976 (N_43976,N_42336,N_41501);
and U43977 (N_43977,N_40834,N_42337);
or U43978 (N_43978,N_41377,N_40752);
nor U43979 (N_43979,N_41750,N_40505);
xor U43980 (N_43980,N_40273,N_40450);
and U43981 (N_43981,N_41893,N_41059);
nor U43982 (N_43982,N_40856,N_42017);
nand U43983 (N_43983,N_41563,N_40169);
or U43984 (N_43984,N_41690,N_40680);
xor U43985 (N_43985,N_41231,N_41773);
nand U43986 (N_43986,N_41970,N_41315);
nor U43987 (N_43987,N_41323,N_41567);
and U43988 (N_43988,N_41116,N_40311);
xnor U43989 (N_43989,N_41687,N_42296);
xor U43990 (N_43990,N_40344,N_41913);
and U43991 (N_43991,N_40234,N_41207);
and U43992 (N_43992,N_40075,N_40503);
and U43993 (N_43993,N_40307,N_42410);
or U43994 (N_43994,N_40058,N_41358);
nand U43995 (N_43995,N_41118,N_41522);
nand U43996 (N_43996,N_41924,N_42083);
xor U43997 (N_43997,N_41170,N_42195);
and U43998 (N_43998,N_42274,N_41429);
nand U43999 (N_43999,N_41448,N_42206);
or U44000 (N_44000,N_40901,N_40293);
nand U44001 (N_44001,N_41543,N_42045);
xnor U44002 (N_44002,N_41075,N_41785);
nand U44003 (N_44003,N_40238,N_40435);
nand U44004 (N_44004,N_40830,N_40068);
nand U44005 (N_44005,N_41642,N_41240);
nor U44006 (N_44006,N_40870,N_41151);
and U44007 (N_44007,N_40805,N_40775);
nor U44008 (N_44008,N_42466,N_41804);
and U44009 (N_44009,N_41502,N_42039);
xnor U44010 (N_44010,N_42258,N_40739);
or U44011 (N_44011,N_40714,N_40322);
nand U44012 (N_44012,N_42027,N_41726);
and U44013 (N_44013,N_41979,N_41173);
nor U44014 (N_44014,N_40172,N_41768);
nand U44015 (N_44015,N_40410,N_40419);
or U44016 (N_44016,N_41551,N_41970);
nand U44017 (N_44017,N_40286,N_41031);
or U44018 (N_44018,N_40630,N_40215);
and U44019 (N_44019,N_40188,N_41869);
xnor U44020 (N_44020,N_41450,N_42152);
xnor U44021 (N_44021,N_40993,N_40476);
and U44022 (N_44022,N_41607,N_40593);
xor U44023 (N_44023,N_40823,N_40720);
nor U44024 (N_44024,N_41322,N_42209);
nand U44025 (N_44025,N_41862,N_41773);
and U44026 (N_44026,N_42037,N_40544);
or U44027 (N_44027,N_41275,N_41801);
or U44028 (N_44028,N_42498,N_40340);
nand U44029 (N_44029,N_42335,N_40844);
or U44030 (N_44030,N_40385,N_40765);
xnor U44031 (N_44031,N_41144,N_41077);
and U44032 (N_44032,N_40392,N_41774);
or U44033 (N_44033,N_40107,N_40004);
and U44034 (N_44034,N_40382,N_42118);
nor U44035 (N_44035,N_42029,N_42320);
and U44036 (N_44036,N_41458,N_41697);
xnor U44037 (N_44037,N_41898,N_40143);
and U44038 (N_44038,N_42448,N_41590);
or U44039 (N_44039,N_41059,N_40245);
or U44040 (N_44040,N_41317,N_40360);
xnor U44041 (N_44041,N_41485,N_41080);
or U44042 (N_44042,N_41234,N_41641);
or U44043 (N_44043,N_42007,N_41657);
nor U44044 (N_44044,N_40328,N_40059);
or U44045 (N_44045,N_41448,N_40806);
and U44046 (N_44046,N_40395,N_42310);
nor U44047 (N_44047,N_41859,N_41941);
xor U44048 (N_44048,N_42364,N_40976);
xor U44049 (N_44049,N_42191,N_41065);
and U44050 (N_44050,N_40405,N_42448);
or U44051 (N_44051,N_41399,N_41949);
xnor U44052 (N_44052,N_40209,N_40835);
nor U44053 (N_44053,N_40521,N_40748);
or U44054 (N_44054,N_40874,N_41899);
and U44055 (N_44055,N_41986,N_40053);
and U44056 (N_44056,N_41073,N_42273);
xor U44057 (N_44057,N_40210,N_40627);
xor U44058 (N_44058,N_41105,N_40698);
nor U44059 (N_44059,N_41649,N_41836);
and U44060 (N_44060,N_41434,N_41107);
nor U44061 (N_44061,N_41255,N_40816);
or U44062 (N_44062,N_40080,N_40306);
or U44063 (N_44063,N_40806,N_41530);
nand U44064 (N_44064,N_40841,N_41865);
nand U44065 (N_44065,N_40102,N_41830);
xnor U44066 (N_44066,N_40101,N_40406);
or U44067 (N_44067,N_41786,N_40998);
and U44068 (N_44068,N_40983,N_40264);
xnor U44069 (N_44069,N_41372,N_40541);
or U44070 (N_44070,N_41849,N_41503);
nand U44071 (N_44071,N_42488,N_41226);
nand U44072 (N_44072,N_40456,N_40925);
or U44073 (N_44073,N_42143,N_41286);
nor U44074 (N_44074,N_41125,N_41602);
nor U44075 (N_44075,N_40977,N_40096);
or U44076 (N_44076,N_40026,N_42076);
and U44077 (N_44077,N_41423,N_40732);
or U44078 (N_44078,N_40062,N_40834);
xnor U44079 (N_44079,N_41132,N_40741);
nor U44080 (N_44080,N_40620,N_41912);
nor U44081 (N_44081,N_41213,N_41090);
xnor U44082 (N_44082,N_40556,N_42358);
and U44083 (N_44083,N_41091,N_40510);
or U44084 (N_44084,N_40944,N_41430);
nand U44085 (N_44085,N_41354,N_42053);
xnor U44086 (N_44086,N_41058,N_42399);
nand U44087 (N_44087,N_40269,N_42353);
nand U44088 (N_44088,N_42445,N_42490);
or U44089 (N_44089,N_42150,N_41910);
and U44090 (N_44090,N_40247,N_40716);
nand U44091 (N_44091,N_41250,N_42156);
nand U44092 (N_44092,N_41568,N_40350);
nand U44093 (N_44093,N_40711,N_40302);
nand U44094 (N_44094,N_41175,N_41844);
and U44095 (N_44095,N_40394,N_40170);
nor U44096 (N_44096,N_41987,N_41950);
xor U44097 (N_44097,N_41200,N_41463);
or U44098 (N_44098,N_41669,N_40655);
xnor U44099 (N_44099,N_40735,N_41873);
nor U44100 (N_44100,N_40768,N_41850);
nor U44101 (N_44101,N_40589,N_41074);
and U44102 (N_44102,N_41109,N_41928);
xor U44103 (N_44103,N_40456,N_40671);
or U44104 (N_44104,N_40411,N_41931);
nor U44105 (N_44105,N_40008,N_41978);
and U44106 (N_44106,N_40521,N_42226);
and U44107 (N_44107,N_40128,N_41062);
or U44108 (N_44108,N_41744,N_41535);
and U44109 (N_44109,N_40047,N_40496);
xor U44110 (N_44110,N_41402,N_41302);
xnor U44111 (N_44111,N_40250,N_41722);
or U44112 (N_44112,N_41540,N_40065);
nand U44113 (N_44113,N_41109,N_40423);
or U44114 (N_44114,N_41803,N_40910);
or U44115 (N_44115,N_41570,N_41254);
xor U44116 (N_44116,N_41531,N_42375);
and U44117 (N_44117,N_40543,N_41758);
and U44118 (N_44118,N_41971,N_41276);
or U44119 (N_44119,N_41913,N_41261);
xnor U44120 (N_44120,N_40658,N_41670);
nor U44121 (N_44121,N_40612,N_41616);
or U44122 (N_44122,N_42407,N_40059);
nor U44123 (N_44123,N_42424,N_42134);
xnor U44124 (N_44124,N_41977,N_40592);
nor U44125 (N_44125,N_42358,N_41325);
xor U44126 (N_44126,N_40514,N_42016);
xnor U44127 (N_44127,N_40226,N_40670);
nor U44128 (N_44128,N_40314,N_41717);
xor U44129 (N_44129,N_41162,N_41038);
and U44130 (N_44130,N_42299,N_40463);
nand U44131 (N_44131,N_41177,N_40135);
or U44132 (N_44132,N_40222,N_40237);
xor U44133 (N_44133,N_40685,N_40623);
xor U44134 (N_44134,N_42068,N_40411);
nand U44135 (N_44135,N_40642,N_41951);
nand U44136 (N_44136,N_40948,N_41080);
nor U44137 (N_44137,N_42025,N_41999);
xnor U44138 (N_44138,N_40648,N_40979);
nor U44139 (N_44139,N_41072,N_41492);
nand U44140 (N_44140,N_40288,N_41551);
xor U44141 (N_44141,N_42416,N_41470);
or U44142 (N_44142,N_41289,N_40321);
nand U44143 (N_44143,N_40928,N_40503);
nor U44144 (N_44144,N_42057,N_42122);
nor U44145 (N_44145,N_42379,N_41005);
nand U44146 (N_44146,N_42387,N_41548);
or U44147 (N_44147,N_40947,N_42117);
xnor U44148 (N_44148,N_40752,N_40164);
nor U44149 (N_44149,N_42212,N_40051);
nor U44150 (N_44150,N_40491,N_42240);
nor U44151 (N_44151,N_41381,N_41826);
nand U44152 (N_44152,N_41286,N_41789);
nor U44153 (N_44153,N_41965,N_40944);
nand U44154 (N_44154,N_42042,N_41519);
and U44155 (N_44155,N_41802,N_40762);
and U44156 (N_44156,N_41703,N_40253);
and U44157 (N_44157,N_42012,N_40785);
nor U44158 (N_44158,N_40907,N_42006);
nand U44159 (N_44159,N_40609,N_42286);
nand U44160 (N_44160,N_41542,N_40136);
nor U44161 (N_44161,N_41213,N_41543);
nand U44162 (N_44162,N_42481,N_40624);
nor U44163 (N_44163,N_41980,N_40032);
nor U44164 (N_44164,N_41747,N_41099);
nor U44165 (N_44165,N_40864,N_40675);
or U44166 (N_44166,N_40985,N_41722);
or U44167 (N_44167,N_42142,N_40251);
xnor U44168 (N_44168,N_41327,N_40670);
nor U44169 (N_44169,N_41818,N_40430);
or U44170 (N_44170,N_41765,N_40302);
nand U44171 (N_44171,N_41067,N_40187);
nand U44172 (N_44172,N_40655,N_40329);
xor U44173 (N_44173,N_41550,N_41847);
nand U44174 (N_44174,N_40423,N_41267);
and U44175 (N_44175,N_40283,N_41766);
and U44176 (N_44176,N_41809,N_42134);
or U44177 (N_44177,N_41261,N_40366);
xnor U44178 (N_44178,N_41269,N_40113);
or U44179 (N_44179,N_41300,N_41519);
xnor U44180 (N_44180,N_40719,N_42499);
and U44181 (N_44181,N_41530,N_40470);
or U44182 (N_44182,N_41495,N_40272);
and U44183 (N_44183,N_40631,N_40863);
nor U44184 (N_44184,N_41435,N_42220);
and U44185 (N_44185,N_40121,N_42088);
and U44186 (N_44186,N_41456,N_40687);
nor U44187 (N_44187,N_40160,N_41813);
nand U44188 (N_44188,N_42134,N_40391);
xnor U44189 (N_44189,N_40356,N_42300);
nor U44190 (N_44190,N_40788,N_42063);
nor U44191 (N_44191,N_40457,N_41396);
or U44192 (N_44192,N_40923,N_40157);
xor U44193 (N_44193,N_40340,N_40366);
nand U44194 (N_44194,N_40299,N_42226);
nor U44195 (N_44195,N_41648,N_40300);
xnor U44196 (N_44196,N_41305,N_40627);
and U44197 (N_44197,N_41030,N_42491);
xnor U44198 (N_44198,N_40949,N_40307);
and U44199 (N_44199,N_40430,N_42023);
xor U44200 (N_44200,N_40528,N_40309);
nor U44201 (N_44201,N_40013,N_41255);
xor U44202 (N_44202,N_41472,N_41350);
and U44203 (N_44203,N_41067,N_40546);
and U44204 (N_44204,N_40617,N_42098);
xor U44205 (N_44205,N_40887,N_40378);
nand U44206 (N_44206,N_41246,N_41979);
nor U44207 (N_44207,N_42161,N_40083);
xor U44208 (N_44208,N_42212,N_42462);
xor U44209 (N_44209,N_42126,N_41747);
or U44210 (N_44210,N_40502,N_40241);
xor U44211 (N_44211,N_40640,N_40856);
nand U44212 (N_44212,N_42163,N_40979);
and U44213 (N_44213,N_40647,N_40543);
nor U44214 (N_44214,N_41529,N_41408);
nand U44215 (N_44215,N_40092,N_42079);
xnor U44216 (N_44216,N_42197,N_41081);
nand U44217 (N_44217,N_42464,N_40417);
nor U44218 (N_44218,N_41009,N_40205);
xor U44219 (N_44219,N_42252,N_41317);
xnor U44220 (N_44220,N_42193,N_41896);
nand U44221 (N_44221,N_41221,N_40691);
nand U44222 (N_44222,N_41396,N_41778);
or U44223 (N_44223,N_42037,N_40541);
or U44224 (N_44224,N_41628,N_40195);
nand U44225 (N_44225,N_41742,N_40643);
nand U44226 (N_44226,N_42413,N_40618);
or U44227 (N_44227,N_40980,N_40461);
nor U44228 (N_44228,N_41485,N_40887);
xnor U44229 (N_44229,N_40600,N_41896);
nor U44230 (N_44230,N_40357,N_40569);
or U44231 (N_44231,N_40552,N_41256);
or U44232 (N_44232,N_42371,N_40480);
nor U44233 (N_44233,N_41913,N_41460);
nor U44234 (N_44234,N_41252,N_41052);
xnor U44235 (N_44235,N_40040,N_40516);
nor U44236 (N_44236,N_41913,N_41383);
xor U44237 (N_44237,N_40336,N_42067);
nand U44238 (N_44238,N_40350,N_40516);
and U44239 (N_44239,N_41167,N_40436);
and U44240 (N_44240,N_40880,N_40989);
nor U44241 (N_44241,N_41422,N_41233);
and U44242 (N_44242,N_42073,N_42119);
and U44243 (N_44243,N_41563,N_41792);
nand U44244 (N_44244,N_40451,N_41920);
nor U44245 (N_44245,N_41048,N_41927);
nand U44246 (N_44246,N_41069,N_42465);
nand U44247 (N_44247,N_40921,N_41267);
xor U44248 (N_44248,N_40299,N_41639);
nand U44249 (N_44249,N_40993,N_40805);
or U44250 (N_44250,N_41018,N_41102);
or U44251 (N_44251,N_40506,N_40314);
nor U44252 (N_44252,N_40425,N_41917);
xor U44253 (N_44253,N_42222,N_42385);
xnor U44254 (N_44254,N_40204,N_41546);
or U44255 (N_44255,N_41113,N_41863);
or U44256 (N_44256,N_40728,N_41283);
or U44257 (N_44257,N_41955,N_41527);
nand U44258 (N_44258,N_41789,N_41171);
and U44259 (N_44259,N_41409,N_40083);
xnor U44260 (N_44260,N_41971,N_40991);
xnor U44261 (N_44261,N_41765,N_41453);
or U44262 (N_44262,N_41677,N_41239);
xnor U44263 (N_44263,N_41269,N_42448);
and U44264 (N_44264,N_41773,N_42049);
and U44265 (N_44265,N_40705,N_42409);
or U44266 (N_44266,N_40547,N_41308);
and U44267 (N_44267,N_41118,N_41178);
or U44268 (N_44268,N_41225,N_40325);
xor U44269 (N_44269,N_40413,N_40195);
and U44270 (N_44270,N_41514,N_41348);
nand U44271 (N_44271,N_41067,N_40290);
xor U44272 (N_44272,N_40837,N_42230);
or U44273 (N_44273,N_40366,N_41323);
nand U44274 (N_44274,N_40640,N_41449);
or U44275 (N_44275,N_40261,N_40358);
xnor U44276 (N_44276,N_41985,N_41878);
or U44277 (N_44277,N_40920,N_41153);
nand U44278 (N_44278,N_42161,N_41502);
or U44279 (N_44279,N_40068,N_40414);
and U44280 (N_44280,N_41748,N_41306);
nand U44281 (N_44281,N_41464,N_41868);
or U44282 (N_44282,N_41652,N_40537);
and U44283 (N_44283,N_41958,N_41061);
or U44284 (N_44284,N_41311,N_41673);
nor U44285 (N_44285,N_40106,N_41813);
nand U44286 (N_44286,N_41568,N_40363);
or U44287 (N_44287,N_41000,N_40994);
or U44288 (N_44288,N_40126,N_41452);
and U44289 (N_44289,N_40256,N_41249);
xnor U44290 (N_44290,N_41972,N_40113);
nand U44291 (N_44291,N_40168,N_41165);
nand U44292 (N_44292,N_42164,N_41355);
xor U44293 (N_44293,N_40129,N_41649);
and U44294 (N_44294,N_41312,N_41226);
and U44295 (N_44295,N_41087,N_41239);
nand U44296 (N_44296,N_40663,N_41933);
nand U44297 (N_44297,N_41578,N_41078);
or U44298 (N_44298,N_41735,N_40130);
nand U44299 (N_44299,N_40956,N_42404);
xor U44300 (N_44300,N_41079,N_41713);
xnor U44301 (N_44301,N_40934,N_41075);
nand U44302 (N_44302,N_42173,N_40007);
xnor U44303 (N_44303,N_40481,N_41987);
nor U44304 (N_44304,N_40005,N_41021);
nor U44305 (N_44305,N_41396,N_41434);
and U44306 (N_44306,N_40251,N_40384);
nand U44307 (N_44307,N_40257,N_41058);
nand U44308 (N_44308,N_40388,N_41022);
xor U44309 (N_44309,N_41950,N_40731);
and U44310 (N_44310,N_40728,N_40462);
nand U44311 (N_44311,N_41679,N_41388);
nor U44312 (N_44312,N_41109,N_41447);
and U44313 (N_44313,N_40703,N_40719);
xor U44314 (N_44314,N_41255,N_40197);
xor U44315 (N_44315,N_40865,N_41335);
or U44316 (N_44316,N_40846,N_41822);
or U44317 (N_44317,N_41982,N_41738);
nor U44318 (N_44318,N_40976,N_42200);
nor U44319 (N_44319,N_40625,N_40042);
xor U44320 (N_44320,N_41316,N_41620);
nor U44321 (N_44321,N_41191,N_41067);
and U44322 (N_44322,N_41208,N_40778);
nor U44323 (N_44323,N_41036,N_41948);
xor U44324 (N_44324,N_41139,N_40163);
nor U44325 (N_44325,N_41623,N_40696);
xor U44326 (N_44326,N_41124,N_42053);
nor U44327 (N_44327,N_42341,N_40975);
and U44328 (N_44328,N_42408,N_40085);
nor U44329 (N_44329,N_41787,N_41468);
nand U44330 (N_44330,N_41374,N_42324);
nor U44331 (N_44331,N_41151,N_40281);
nand U44332 (N_44332,N_42353,N_41666);
nor U44333 (N_44333,N_41619,N_41992);
xor U44334 (N_44334,N_40672,N_42379);
or U44335 (N_44335,N_40437,N_42375);
or U44336 (N_44336,N_40472,N_40871);
nor U44337 (N_44337,N_40624,N_41143);
nor U44338 (N_44338,N_40153,N_40472);
and U44339 (N_44339,N_40513,N_41882);
or U44340 (N_44340,N_41117,N_41848);
nand U44341 (N_44341,N_41483,N_42452);
or U44342 (N_44342,N_41595,N_40495);
nor U44343 (N_44343,N_40718,N_42187);
and U44344 (N_44344,N_41163,N_40454);
xnor U44345 (N_44345,N_40958,N_42284);
xor U44346 (N_44346,N_41226,N_41013);
xor U44347 (N_44347,N_41588,N_41541);
xor U44348 (N_44348,N_40224,N_40519);
nand U44349 (N_44349,N_41682,N_41735);
nor U44350 (N_44350,N_41119,N_41261);
nand U44351 (N_44351,N_42260,N_42198);
nor U44352 (N_44352,N_40401,N_41996);
or U44353 (N_44353,N_42372,N_41741);
nor U44354 (N_44354,N_40040,N_41372);
nand U44355 (N_44355,N_41604,N_41978);
nor U44356 (N_44356,N_41380,N_41255);
nor U44357 (N_44357,N_40102,N_40703);
and U44358 (N_44358,N_40894,N_41429);
nand U44359 (N_44359,N_41075,N_41453);
xnor U44360 (N_44360,N_41944,N_40124);
or U44361 (N_44361,N_40194,N_41247);
or U44362 (N_44362,N_40528,N_40409);
nand U44363 (N_44363,N_41201,N_42068);
nor U44364 (N_44364,N_41569,N_40336);
or U44365 (N_44365,N_40080,N_41827);
and U44366 (N_44366,N_40063,N_40818);
nand U44367 (N_44367,N_42366,N_40994);
or U44368 (N_44368,N_41869,N_41990);
xnor U44369 (N_44369,N_40830,N_42193);
and U44370 (N_44370,N_40286,N_41868);
xnor U44371 (N_44371,N_40112,N_40002);
nand U44372 (N_44372,N_41476,N_40247);
or U44373 (N_44373,N_40231,N_41641);
or U44374 (N_44374,N_42284,N_42409);
nor U44375 (N_44375,N_42272,N_40789);
xnor U44376 (N_44376,N_41310,N_40865);
or U44377 (N_44377,N_40655,N_40857);
xor U44378 (N_44378,N_40388,N_40304);
nor U44379 (N_44379,N_40753,N_40910);
nor U44380 (N_44380,N_42280,N_40950);
or U44381 (N_44381,N_41202,N_40430);
and U44382 (N_44382,N_42354,N_41690);
and U44383 (N_44383,N_40103,N_42168);
xnor U44384 (N_44384,N_41319,N_40717);
xor U44385 (N_44385,N_40435,N_40442);
xor U44386 (N_44386,N_40023,N_40403);
xnor U44387 (N_44387,N_40542,N_40603);
and U44388 (N_44388,N_42222,N_41993);
nand U44389 (N_44389,N_41689,N_40604);
xnor U44390 (N_44390,N_42081,N_42476);
nand U44391 (N_44391,N_41043,N_41892);
or U44392 (N_44392,N_40772,N_40993);
xor U44393 (N_44393,N_41294,N_40420);
nand U44394 (N_44394,N_40722,N_40456);
and U44395 (N_44395,N_41937,N_41987);
nand U44396 (N_44396,N_40620,N_42194);
xnor U44397 (N_44397,N_40271,N_41285);
and U44398 (N_44398,N_42362,N_41818);
and U44399 (N_44399,N_40057,N_40411);
nand U44400 (N_44400,N_40045,N_41222);
nor U44401 (N_44401,N_41743,N_40159);
nand U44402 (N_44402,N_42029,N_42200);
nor U44403 (N_44403,N_40198,N_42006);
or U44404 (N_44404,N_40960,N_40387);
nand U44405 (N_44405,N_41110,N_42193);
xnor U44406 (N_44406,N_41272,N_40797);
or U44407 (N_44407,N_42135,N_40480);
and U44408 (N_44408,N_40390,N_41264);
nor U44409 (N_44409,N_40342,N_42355);
xnor U44410 (N_44410,N_41356,N_40719);
nor U44411 (N_44411,N_40515,N_41105);
nor U44412 (N_44412,N_40056,N_41364);
or U44413 (N_44413,N_42460,N_41734);
nand U44414 (N_44414,N_40738,N_41556);
and U44415 (N_44415,N_40737,N_41066);
nand U44416 (N_44416,N_41171,N_40212);
and U44417 (N_44417,N_41423,N_41704);
nand U44418 (N_44418,N_40829,N_41766);
nand U44419 (N_44419,N_41371,N_41459);
or U44420 (N_44420,N_42202,N_40873);
nand U44421 (N_44421,N_41768,N_40910);
nor U44422 (N_44422,N_40223,N_41710);
nor U44423 (N_44423,N_41902,N_40560);
nand U44424 (N_44424,N_42269,N_40773);
xnor U44425 (N_44425,N_40916,N_40069);
xor U44426 (N_44426,N_40720,N_41569);
nand U44427 (N_44427,N_40128,N_41147);
nor U44428 (N_44428,N_41195,N_40709);
and U44429 (N_44429,N_40688,N_41041);
nor U44430 (N_44430,N_42308,N_42092);
and U44431 (N_44431,N_40548,N_40761);
nor U44432 (N_44432,N_40776,N_40132);
xnor U44433 (N_44433,N_40012,N_41991);
xnor U44434 (N_44434,N_42229,N_41144);
nor U44435 (N_44435,N_41301,N_40648);
nor U44436 (N_44436,N_41866,N_41927);
nor U44437 (N_44437,N_41079,N_42439);
and U44438 (N_44438,N_40421,N_40834);
and U44439 (N_44439,N_42370,N_42126);
xor U44440 (N_44440,N_42323,N_41970);
xor U44441 (N_44441,N_42348,N_40669);
nor U44442 (N_44442,N_40574,N_40229);
nand U44443 (N_44443,N_41342,N_41773);
xor U44444 (N_44444,N_42021,N_40136);
or U44445 (N_44445,N_41675,N_42417);
or U44446 (N_44446,N_41373,N_40720);
or U44447 (N_44447,N_42422,N_40374);
nand U44448 (N_44448,N_41942,N_40797);
xor U44449 (N_44449,N_42192,N_42400);
nand U44450 (N_44450,N_41720,N_40683);
and U44451 (N_44451,N_42044,N_42473);
and U44452 (N_44452,N_41842,N_42378);
nand U44453 (N_44453,N_41194,N_41375);
nand U44454 (N_44454,N_41236,N_40140);
nand U44455 (N_44455,N_41748,N_42434);
or U44456 (N_44456,N_42015,N_41245);
nand U44457 (N_44457,N_42374,N_41241);
and U44458 (N_44458,N_40467,N_41546);
nand U44459 (N_44459,N_41063,N_40931);
and U44460 (N_44460,N_42323,N_40642);
nand U44461 (N_44461,N_40479,N_40138);
and U44462 (N_44462,N_42300,N_40157);
or U44463 (N_44463,N_41513,N_42200);
nor U44464 (N_44464,N_42399,N_41960);
xnor U44465 (N_44465,N_40412,N_41911);
or U44466 (N_44466,N_40190,N_41446);
nor U44467 (N_44467,N_41453,N_40273);
nor U44468 (N_44468,N_41328,N_41318);
xor U44469 (N_44469,N_41517,N_41800);
or U44470 (N_44470,N_41257,N_41938);
and U44471 (N_44471,N_41485,N_40829);
and U44472 (N_44472,N_40462,N_41073);
or U44473 (N_44473,N_42350,N_41741);
xor U44474 (N_44474,N_40798,N_41170);
and U44475 (N_44475,N_40693,N_41623);
nor U44476 (N_44476,N_40386,N_41272);
nand U44477 (N_44477,N_40358,N_41449);
nor U44478 (N_44478,N_41776,N_41754);
and U44479 (N_44479,N_41881,N_41645);
nand U44480 (N_44480,N_41380,N_41218);
or U44481 (N_44481,N_40938,N_40607);
and U44482 (N_44482,N_40735,N_42365);
and U44483 (N_44483,N_42440,N_42209);
and U44484 (N_44484,N_40509,N_41096);
xnor U44485 (N_44485,N_41226,N_40774);
xnor U44486 (N_44486,N_40702,N_41710);
nor U44487 (N_44487,N_41326,N_40343);
or U44488 (N_44488,N_42476,N_40523);
xnor U44489 (N_44489,N_40314,N_40387);
and U44490 (N_44490,N_40709,N_40143);
nand U44491 (N_44491,N_40229,N_40134);
nor U44492 (N_44492,N_41844,N_41779);
xnor U44493 (N_44493,N_41069,N_40659);
nand U44494 (N_44494,N_42051,N_41330);
or U44495 (N_44495,N_40205,N_41962);
nand U44496 (N_44496,N_41359,N_42494);
nor U44497 (N_44497,N_41769,N_42479);
or U44498 (N_44498,N_40972,N_40386);
nor U44499 (N_44499,N_41981,N_41717);
and U44500 (N_44500,N_42197,N_42192);
and U44501 (N_44501,N_40234,N_40883);
xor U44502 (N_44502,N_41582,N_41689);
xor U44503 (N_44503,N_42464,N_41831);
xor U44504 (N_44504,N_40447,N_42005);
nand U44505 (N_44505,N_40140,N_42421);
and U44506 (N_44506,N_40898,N_41223);
xor U44507 (N_44507,N_42024,N_41661);
or U44508 (N_44508,N_40944,N_41959);
nor U44509 (N_44509,N_40559,N_41231);
or U44510 (N_44510,N_40226,N_40234);
nand U44511 (N_44511,N_41428,N_42345);
nor U44512 (N_44512,N_41026,N_42337);
or U44513 (N_44513,N_41110,N_41912);
and U44514 (N_44514,N_41005,N_41857);
nand U44515 (N_44515,N_41455,N_41247);
xnor U44516 (N_44516,N_42394,N_41354);
nor U44517 (N_44517,N_42485,N_40588);
nor U44518 (N_44518,N_41050,N_42007);
or U44519 (N_44519,N_42418,N_42478);
and U44520 (N_44520,N_40267,N_41194);
nand U44521 (N_44521,N_41439,N_40302);
nand U44522 (N_44522,N_41519,N_41753);
and U44523 (N_44523,N_41532,N_41216);
and U44524 (N_44524,N_41423,N_41161);
and U44525 (N_44525,N_41824,N_41543);
and U44526 (N_44526,N_41763,N_42431);
nand U44527 (N_44527,N_40933,N_41847);
xnor U44528 (N_44528,N_41676,N_40208);
and U44529 (N_44529,N_41814,N_40420);
xnor U44530 (N_44530,N_42333,N_41560);
and U44531 (N_44531,N_40397,N_40577);
or U44532 (N_44532,N_41547,N_41124);
and U44533 (N_44533,N_41069,N_40114);
xor U44534 (N_44534,N_41892,N_40205);
nor U44535 (N_44535,N_40214,N_40740);
and U44536 (N_44536,N_40920,N_41305);
or U44537 (N_44537,N_40355,N_40432);
nand U44538 (N_44538,N_41882,N_42483);
nor U44539 (N_44539,N_40969,N_40099);
and U44540 (N_44540,N_41323,N_41695);
nand U44541 (N_44541,N_41540,N_41236);
nor U44542 (N_44542,N_41529,N_42244);
xnor U44543 (N_44543,N_40796,N_40874);
nor U44544 (N_44544,N_40911,N_41296);
xor U44545 (N_44545,N_41648,N_42085);
nor U44546 (N_44546,N_40329,N_40817);
nand U44547 (N_44547,N_42375,N_40225);
and U44548 (N_44548,N_41790,N_42263);
nor U44549 (N_44549,N_40861,N_41505);
or U44550 (N_44550,N_41828,N_40934);
xor U44551 (N_44551,N_41428,N_41736);
nor U44552 (N_44552,N_40520,N_41593);
nand U44553 (N_44553,N_41469,N_40668);
and U44554 (N_44554,N_40635,N_41677);
xor U44555 (N_44555,N_41940,N_41725);
and U44556 (N_44556,N_41417,N_40309);
nand U44557 (N_44557,N_41269,N_41235);
or U44558 (N_44558,N_42262,N_42485);
xor U44559 (N_44559,N_40454,N_41476);
and U44560 (N_44560,N_41233,N_42394);
or U44561 (N_44561,N_40764,N_42360);
or U44562 (N_44562,N_41248,N_40199);
and U44563 (N_44563,N_40415,N_40300);
and U44564 (N_44564,N_42048,N_41240);
nor U44565 (N_44565,N_42372,N_40229);
and U44566 (N_44566,N_42162,N_40537);
and U44567 (N_44567,N_40451,N_41037);
xnor U44568 (N_44568,N_40046,N_40841);
or U44569 (N_44569,N_40188,N_40816);
and U44570 (N_44570,N_41112,N_40081);
and U44571 (N_44571,N_41928,N_40168);
nor U44572 (N_44572,N_41590,N_41647);
nor U44573 (N_44573,N_41532,N_41766);
and U44574 (N_44574,N_40421,N_40983);
and U44575 (N_44575,N_40797,N_40275);
and U44576 (N_44576,N_41540,N_40822);
nor U44577 (N_44577,N_40819,N_41727);
nand U44578 (N_44578,N_41882,N_40305);
or U44579 (N_44579,N_40260,N_41330);
nor U44580 (N_44580,N_40835,N_41256);
and U44581 (N_44581,N_40728,N_41870);
nor U44582 (N_44582,N_41304,N_41384);
nor U44583 (N_44583,N_40385,N_42325);
xor U44584 (N_44584,N_41402,N_41045);
xnor U44585 (N_44585,N_41155,N_41903);
xor U44586 (N_44586,N_41124,N_41264);
nand U44587 (N_44587,N_41118,N_41719);
or U44588 (N_44588,N_40221,N_41197);
or U44589 (N_44589,N_41754,N_40111);
and U44590 (N_44590,N_40322,N_40623);
xor U44591 (N_44591,N_41752,N_40320);
nor U44592 (N_44592,N_40195,N_41037);
and U44593 (N_44593,N_40121,N_40570);
or U44594 (N_44594,N_41915,N_41257);
nand U44595 (N_44595,N_42033,N_41662);
and U44596 (N_44596,N_42043,N_42341);
nor U44597 (N_44597,N_40612,N_41505);
nor U44598 (N_44598,N_42269,N_40565);
or U44599 (N_44599,N_40764,N_41286);
nand U44600 (N_44600,N_41968,N_40056);
nand U44601 (N_44601,N_42465,N_41271);
nor U44602 (N_44602,N_40890,N_40465);
xor U44603 (N_44603,N_40430,N_41244);
and U44604 (N_44604,N_41608,N_40554);
nor U44605 (N_44605,N_42233,N_40490);
nand U44606 (N_44606,N_40912,N_41917);
or U44607 (N_44607,N_41996,N_42133);
or U44608 (N_44608,N_40763,N_40668);
nand U44609 (N_44609,N_42231,N_40672);
xnor U44610 (N_44610,N_41554,N_40883);
nor U44611 (N_44611,N_41114,N_41131);
nor U44612 (N_44612,N_41223,N_42043);
xnor U44613 (N_44613,N_41603,N_41833);
nand U44614 (N_44614,N_40004,N_42484);
nand U44615 (N_44615,N_40928,N_40834);
nor U44616 (N_44616,N_41265,N_40317);
nand U44617 (N_44617,N_42015,N_41839);
and U44618 (N_44618,N_42471,N_40385);
or U44619 (N_44619,N_42426,N_40983);
nand U44620 (N_44620,N_40336,N_41699);
nand U44621 (N_44621,N_42395,N_40510);
nor U44622 (N_44622,N_41143,N_42143);
nor U44623 (N_44623,N_41793,N_42470);
and U44624 (N_44624,N_41700,N_41562);
or U44625 (N_44625,N_40670,N_41272);
and U44626 (N_44626,N_42296,N_41929);
and U44627 (N_44627,N_40732,N_41723);
or U44628 (N_44628,N_40105,N_41459);
xor U44629 (N_44629,N_40369,N_40688);
nand U44630 (N_44630,N_40735,N_42028);
nand U44631 (N_44631,N_40397,N_40568);
nor U44632 (N_44632,N_41072,N_40822);
or U44633 (N_44633,N_40834,N_41475);
nor U44634 (N_44634,N_40121,N_41555);
nand U44635 (N_44635,N_40311,N_41222);
or U44636 (N_44636,N_41756,N_40472);
xor U44637 (N_44637,N_40552,N_40515);
nand U44638 (N_44638,N_41226,N_41868);
and U44639 (N_44639,N_40985,N_41503);
or U44640 (N_44640,N_41930,N_42420);
and U44641 (N_44641,N_40093,N_41613);
nor U44642 (N_44642,N_40138,N_41725);
and U44643 (N_44643,N_40749,N_40825);
and U44644 (N_44644,N_40252,N_42430);
xnor U44645 (N_44645,N_40657,N_41942);
and U44646 (N_44646,N_41708,N_41243);
or U44647 (N_44647,N_42042,N_42142);
xor U44648 (N_44648,N_41955,N_40928);
and U44649 (N_44649,N_41671,N_41991);
and U44650 (N_44650,N_40785,N_41222);
or U44651 (N_44651,N_41457,N_40546);
or U44652 (N_44652,N_40743,N_40438);
nor U44653 (N_44653,N_41588,N_42156);
nor U44654 (N_44654,N_40222,N_41144);
or U44655 (N_44655,N_40193,N_42434);
xor U44656 (N_44656,N_41412,N_41649);
xnor U44657 (N_44657,N_40792,N_42487);
nor U44658 (N_44658,N_40503,N_40378);
or U44659 (N_44659,N_42090,N_40198);
or U44660 (N_44660,N_41833,N_40709);
nand U44661 (N_44661,N_40309,N_40628);
and U44662 (N_44662,N_41165,N_41333);
nand U44663 (N_44663,N_42120,N_42305);
nor U44664 (N_44664,N_41243,N_40503);
and U44665 (N_44665,N_41471,N_40550);
xnor U44666 (N_44666,N_42027,N_41017);
xnor U44667 (N_44667,N_41097,N_41275);
or U44668 (N_44668,N_41930,N_40569);
nor U44669 (N_44669,N_40651,N_41001);
nor U44670 (N_44670,N_42406,N_40008);
nand U44671 (N_44671,N_40742,N_40161);
or U44672 (N_44672,N_42016,N_42154);
nor U44673 (N_44673,N_41994,N_41733);
nand U44674 (N_44674,N_41871,N_42014);
or U44675 (N_44675,N_40654,N_42313);
or U44676 (N_44676,N_42210,N_41137);
or U44677 (N_44677,N_40955,N_41148);
or U44678 (N_44678,N_40206,N_41032);
or U44679 (N_44679,N_41580,N_41430);
nand U44680 (N_44680,N_40731,N_42021);
or U44681 (N_44681,N_42154,N_40557);
xor U44682 (N_44682,N_41049,N_42463);
xnor U44683 (N_44683,N_41660,N_40791);
nand U44684 (N_44684,N_42361,N_40463);
and U44685 (N_44685,N_40671,N_41821);
xnor U44686 (N_44686,N_41628,N_41476);
and U44687 (N_44687,N_40467,N_42494);
and U44688 (N_44688,N_41371,N_42292);
nor U44689 (N_44689,N_40329,N_41271);
and U44690 (N_44690,N_41265,N_40407);
or U44691 (N_44691,N_42216,N_40019);
nand U44692 (N_44692,N_41804,N_41701);
nand U44693 (N_44693,N_41934,N_40080);
nor U44694 (N_44694,N_41415,N_41483);
and U44695 (N_44695,N_40740,N_41366);
nand U44696 (N_44696,N_40884,N_41882);
and U44697 (N_44697,N_41617,N_42479);
xor U44698 (N_44698,N_40108,N_42268);
and U44699 (N_44699,N_40256,N_40759);
nand U44700 (N_44700,N_40762,N_40553);
and U44701 (N_44701,N_40667,N_41465);
nand U44702 (N_44702,N_42342,N_42223);
xnor U44703 (N_44703,N_40779,N_41247);
or U44704 (N_44704,N_42173,N_42127);
nand U44705 (N_44705,N_40883,N_41684);
nand U44706 (N_44706,N_41583,N_41279);
nand U44707 (N_44707,N_42128,N_40250);
or U44708 (N_44708,N_40451,N_40422);
nor U44709 (N_44709,N_42275,N_40331);
nor U44710 (N_44710,N_40814,N_41779);
xnor U44711 (N_44711,N_40180,N_41722);
nor U44712 (N_44712,N_41991,N_42143);
or U44713 (N_44713,N_40485,N_41142);
or U44714 (N_44714,N_41461,N_41328);
nor U44715 (N_44715,N_40551,N_42289);
xnor U44716 (N_44716,N_41191,N_41216);
and U44717 (N_44717,N_42023,N_42175);
and U44718 (N_44718,N_40099,N_40308);
and U44719 (N_44719,N_40101,N_40770);
and U44720 (N_44720,N_42051,N_42113);
nor U44721 (N_44721,N_42466,N_40798);
nor U44722 (N_44722,N_41515,N_40927);
and U44723 (N_44723,N_40818,N_41603);
or U44724 (N_44724,N_41111,N_40948);
and U44725 (N_44725,N_40377,N_41551);
and U44726 (N_44726,N_42226,N_40799);
nor U44727 (N_44727,N_41990,N_41083);
xor U44728 (N_44728,N_40341,N_40938);
nand U44729 (N_44729,N_40865,N_40463);
nor U44730 (N_44730,N_40598,N_41455);
nor U44731 (N_44731,N_41707,N_41502);
and U44732 (N_44732,N_42140,N_41231);
and U44733 (N_44733,N_40909,N_41815);
or U44734 (N_44734,N_40103,N_41144);
nor U44735 (N_44735,N_41272,N_40926);
or U44736 (N_44736,N_41215,N_40557);
or U44737 (N_44737,N_42266,N_40425);
and U44738 (N_44738,N_41866,N_41635);
or U44739 (N_44739,N_40013,N_40462);
or U44740 (N_44740,N_42142,N_40105);
nor U44741 (N_44741,N_40665,N_41272);
nand U44742 (N_44742,N_40406,N_40305);
nand U44743 (N_44743,N_40399,N_41444);
or U44744 (N_44744,N_41860,N_40339);
nand U44745 (N_44745,N_40221,N_41843);
xnor U44746 (N_44746,N_41434,N_41088);
nor U44747 (N_44747,N_41374,N_40217);
xor U44748 (N_44748,N_42139,N_41792);
xor U44749 (N_44749,N_42329,N_41426);
xor U44750 (N_44750,N_40520,N_42350);
and U44751 (N_44751,N_41404,N_41424);
nand U44752 (N_44752,N_41722,N_40078);
xor U44753 (N_44753,N_41535,N_40653);
nand U44754 (N_44754,N_40786,N_40732);
nor U44755 (N_44755,N_41331,N_40567);
nand U44756 (N_44756,N_42010,N_40302);
nor U44757 (N_44757,N_40843,N_41321);
nor U44758 (N_44758,N_40559,N_40506);
nor U44759 (N_44759,N_41848,N_41923);
or U44760 (N_44760,N_40947,N_42098);
and U44761 (N_44761,N_40709,N_42229);
nor U44762 (N_44762,N_41552,N_40967);
xor U44763 (N_44763,N_41364,N_40452);
or U44764 (N_44764,N_42413,N_40049);
and U44765 (N_44765,N_40996,N_41487);
nand U44766 (N_44766,N_41193,N_41088);
nor U44767 (N_44767,N_40268,N_41549);
nor U44768 (N_44768,N_41367,N_42457);
nor U44769 (N_44769,N_40695,N_42219);
nor U44770 (N_44770,N_41159,N_41608);
or U44771 (N_44771,N_40639,N_41047);
nor U44772 (N_44772,N_41560,N_41889);
and U44773 (N_44773,N_42231,N_41828);
nand U44774 (N_44774,N_41272,N_42395);
and U44775 (N_44775,N_40531,N_41077);
and U44776 (N_44776,N_42445,N_41624);
or U44777 (N_44777,N_41456,N_41780);
or U44778 (N_44778,N_40550,N_42050);
and U44779 (N_44779,N_40896,N_41293);
nand U44780 (N_44780,N_40814,N_41477);
nor U44781 (N_44781,N_42371,N_41148);
xnor U44782 (N_44782,N_40057,N_42158);
xor U44783 (N_44783,N_40485,N_40122);
or U44784 (N_44784,N_40770,N_41725);
and U44785 (N_44785,N_41003,N_41520);
xor U44786 (N_44786,N_41522,N_41195);
and U44787 (N_44787,N_41385,N_42486);
and U44788 (N_44788,N_41569,N_40475);
or U44789 (N_44789,N_41036,N_40127);
xnor U44790 (N_44790,N_41661,N_40325);
nor U44791 (N_44791,N_42371,N_40211);
and U44792 (N_44792,N_41718,N_40519);
nand U44793 (N_44793,N_42496,N_41221);
nand U44794 (N_44794,N_40784,N_40893);
nand U44795 (N_44795,N_41605,N_41421);
nor U44796 (N_44796,N_40614,N_40347);
or U44797 (N_44797,N_41644,N_40658);
nor U44798 (N_44798,N_40017,N_40831);
and U44799 (N_44799,N_41052,N_42364);
and U44800 (N_44800,N_42441,N_41751);
xnor U44801 (N_44801,N_40610,N_41896);
xnor U44802 (N_44802,N_40284,N_42020);
and U44803 (N_44803,N_40525,N_42178);
nand U44804 (N_44804,N_42328,N_42055);
or U44805 (N_44805,N_41192,N_41912);
nand U44806 (N_44806,N_40210,N_41795);
and U44807 (N_44807,N_41145,N_40149);
nor U44808 (N_44808,N_40715,N_41591);
nor U44809 (N_44809,N_41012,N_42354);
nor U44810 (N_44810,N_40319,N_42038);
nand U44811 (N_44811,N_40355,N_40559);
xnor U44812 (N_44812,N_42283,N_41460);
or U44813 (N_44813,N_41718,N_42336);
xor U44814 (N_44814,N_42305,N_41628);
nand U44815 (N_44815,N_41928,N_40131);
or U44816 (N_44816,N_41162,N_40327);
nand U44817 (N_44817,N_41306,N_41307);
or U44818 (N_44818,N_40282,N_40220);
and U44819 (N_44819,N_42498,N_40654);
and U44820 (N_44820,N_40636,N_40469);
nand U44821 (N_44821,N_42470,N_41592);
nand U44822 (N_44822,N_42127,N_42001);
xnor U44823 (N_44823,N_41941,N_40649);
nor U44824 (N_44824,N_40010,N_40844);
nand U44825 (N_44825,N_41210,N_41602);
and U44826 (N_44826,N_40774,N_42484);
xnor U44827 (N_44827,N_40783,N_40513);
nand U44828 (N_44828,N_41507,N_41444);
nand U44829 (N_44829,N_40415,N_42111);
xor U44830 (N_44830,N_40909,N_41374);
nor U44831 (N_44831,N_41084,N_41155);
or U44832 (N_44832,N_40698,N_40106);
and U44833 (N_44833,N_42014,N_40416);
nand U44834 (N_44834,N_42408,N_40808);
xor U44835 (N_44835,N_41648,N_41365);
nor U44836 (N_44836,N_40446,N_42492);
xor U44837 (N_44837,N_40640,N_42131);
and U44838 (N_44838,N_41943,N_41434);
nand U44839 (N_44839,N_41914,N_42366);
or U44840 (N_44840,N_40160,N_41174);
xnor U44841 (N_44841,N_41981,N_40495);
nand U44842 (N_44842,N_41404,N_41833);
xnor U44843 (N_44843,N_40405,N_41535);
or U44844 (N_44844,N_40461,N_41319);
or U44845 (N_44845,N_41015,N_40128);
nand U44846 (N_44846,N_42306,N_40585);
xor U44847 (N_44847,N_40205,N_41804);
xor U44848 (N_44848,N_41378,N_41385);
or U44849 (N_44849,N_41781,N_41041);
and U44850 (N_44850,N_40420,N_40107);
nor U44851 (N_44851,N_42106,N_40200);
xor U44852 (N_44852,N_40797,N_40890);
or U44853 (N_44853,N_41484,N_41549);
nor U44854 (N_44854,N_40348,N_40013);
and U44855 (N_44855,N_40274,N_41636);
nor U44856 (N_44856,N_41531,N_40197);
or U44857 (N_44857,N_40436,N_40032);
xnor U44858 (N_44858,N_42439,N_40272);
nor U44859 (N_44859,N_40371,N_41536);
nor U44860 (N_44860,N_40708,N_41080);
and U44861 (N_44861,N_41112,N_40941);
xnor U44862 (N_44862,N_42251,N_41345);
xor U44863 (N_44863,N_40412,N_41528);
nor U44864 (N_44864,N_40146,N_40278);
or U44865 (N_44865,N_41236,N_40680);
xnor U44866 (N_44866,N_41579,N_41909);
nand U44867 (N_44867,N_41500,N_40619);
nor U44868 (N_44868,N_41422,N_40223);
and U44869 (N_44869,N_41823,N_42021);
and U44870 (N_44870,N_41543,N_40307);
xnor U44871 (N_44871,N_41290,N_40033);
xor U44872 (N_44872,N_41037,N_41026);
or U44873 (N_44873,N_41050,N_40630);
or U44874 (N_44874,N_40020,N_40850);
and U44875 (N_44875,N_41813,N_41967);
nor U44876 (N_44876,N_40978,N_40806);
or U44877 (N_44877,N_41173,N_41983);
xor U44878 (N_44878,N_40454,N_41477);
or U44879 (N_44879,N_41504,N_40047);
and U44880 (N_44880,N_41972,N_41585);
or U44881 (N_44881,N_41362,N_42256);
nand U44882 (N_44882,N_41520,N_40070);
and U44883 (N_44883,N_41706,N_41966);
and U44884 (N_44884,N_40952,N_40054);
nand U44885 (N_44885,N_41877,N_42384);
nor U44886 (N_44886,N_42081,N_40763);
nor U44887 (N_44887,N_40600,N_41006);
or U44888 (N_44888,N_41334,N_41679);
nand U44889 (N_44889,N_41307,N_40953);
nor U44890 (N_44890,N_40409,N_40649);
or U44891 (N_44891,N_40304,N_42044);
and U44892 (N_44892,N_41889,N_41115);
and U44893 (N_44893,N_40070,N_41864);
nand U44894 (N_44894,N_41871,N_42193);
nand U44895 (N_44895,N_40396,N_41259);
nor U44896 (N_44896,N_41938,N_41170);
nand U44897 (N_44897,N_42098,N_41985);
or U44898 (N_44898,N_42461,N_40152);
nand U44899 (N_44899,N_41165,N_41172);
xor U44900 (N_44900,N_42170,N_40615);
or U44901 (N_44901,N_40446,N_40385);
xnor U44902 (N_44902,N_41695,N_40596);
nand U44903 (N_44903,N_41351,N_40944);
and U44904 (N_44904,N_40170,N_41619);
and U44905 (N_44905,N_40085,N_41155);
xnor U44906 (N_44906,N_41189,N_41098);
xnor U44907 (N_44907,N_40392,N_40739);
nand U44908 (N_44908,N_40334,N_42212);
or U44909 (N_44909,N_40575,N_42153);
nor U44910 (N_44910,N_40849,N_41176);
or U44911 (N_44911,N_41817,N_40540);
and U44912 (N_44912,N_41727,N_41555);
nor U44913 (N_44913,N_42117,N_41891);
xnor U44914 (N_44914,N_40254,N_42378);
or U44915 (N_44915,N_40961,N_41253);
nand U44916 (N_44916,N_41832,N_41373);
xnor U44917 (N_44917,N_42460,N_40975);
nand U44918 (N_44918,N_41591,N_41895);
or U44919 (N_44919,N_40121,N_40512);
nand U44920 (N_44920,N_41688,N_42256);
nand U44921 (N_44921,N_40557,N_42279);
and U44922 (N_44922,N_42026,N_42145);
and U44923 (N_44923,N_42311,N_41170);
and U44924 (N_44924,N_41803,N_40651);
nand U44925 (N_44925,N_42497,N_41448);
nor U44926 (N_44926,N_42326,N_40816);
or U44927 (N_44927,N_42127,N_41719);
xor U44928 (N_44928,N_41836,N_40299);
xor U44929 (N_44929,N_41984,N_40984);
and U44930 (N_44930,N_41892,N_41939);
or U44931 (N_44931,N_41457,N_41860);
and U44932 (N_44932,N_41027,N_40709);
xor U44933 (N_44933,N_41654,N_40016);
and U44934 (N_44934,N_40300,N_41162);
xnor U44935 (N_44935,N_40758,N_41927);
or U44936 (N_44936,N_41122,N_40937);
nor U44937 (N_44937,N_40686,N_40941);
nor U44938 (N_44938,N_42471,N_41565);
nor U44939 (N_44939,N_42258,N_40290);
xnor U44940 (N_44940,N_42418,N_42448);
and U44941 (N_44941,N_40953,N_42459);
xor U44942 (N_44942,N_41337,N_40359);
nor U44943 (N_44943,N_42486,N_42159);
nand U44944 (N_44944,N_40293,N_41835);
nor U44945 (N_44945,N_41652,N_42017);
nor U44946 (N_44946,N_41184,N_41108);
and U44947 (N_44947,N_41903,N_41241);
nand U44948 (N_44948,N_41480,N_40802);
and U44949 (N_44949,N_41631,N_41892);
nand U44950 (N_44950,N_42151,N_40145);
nand U44951 (N_44951,N_41906,N_41801);
xnor U44952 (N_44952,N_42009,N_42353);
xnor U44953 (N_44953,N_42457,N_41484);
nor U44954 (N_44954,N_41482,N_40575);
nand U44955 (N_44955,N_40602,N_41179);
and U44956 (N_44956,N_42143,N_40155);
nor U44957 (N_44957,N_41271,N_40296);
nor U44958 (N_44958,N_41794,N_41518);
or U44959 (N_44959,N_42114,N_40136);
nand U44960 (N_44960,N_41830,N_40176);
nand U44961 (N_44961,N_40911,N_40645);
nor U44962 (N_44962,N_40865,N_42231);
nor U44963 (N_44963,N_41306,N_41902);
and U44964 (N_44964,N_40175,N_41796);
nand U44965 (N_44965,N_42255,N_42414);
nor U44966 (N_44966,N_41726,N_42168);
or U44967 (N_44967,N_41767,N_40216);
and U44968 (N_44968,N_40937,N_40694);
nand U44969 (N_44969,N_42108,N_42073);
xor U44970 (N_44970,N_41379,N_42263);
and U44971 (N_44971,N_42019,N_42018);
or U44972 (N_44972,N_41806,N_40024);
or U44973 (N_44973,N_42291,N_41669);
or U44974 (N_44974,N_40835,N_42276);
nor U44975 (N_44975,N_41415,N_41761);
nor U44976 (N_44976,N_41330,N_41421);
xnor U44977 (N_44977,N_40442,N_41787);
and U44978 (N_44978,N_40384,N_41925);
nand U44979 (N_44979,N_40903,N_41887);
and U44980 (N_44980,N_41159,N_41817);
or U44981 (N_44981,N_41234,N_40592);
nand U44982 (N_44982,N_41111,N_41208);
or U44983 (N_44983,N_42167,N_41589);
nor U44984 (N_44984,N_40606,N_40022);
nand U44985 (N_44985,N_41885,N_41110);
and U44986 (N_44986,N_41183,N_42161);
nand U44987 (N_44987,N_41775,N_42436);
xor U44988 (N_44988,N_42475,N_40083);
or U44989 (N_44989,N_41506,N_41165);
or U44990 (N_44990,N_40480,N_42189);
or U44991 (N_44991,N_41203,N_42361);
nand U44992 (N_44992,N_41559,N_40474);
nand U44993 (N_44993,N_41515,N_42397);
or U44994 (N_44994,N_41869,N_42345);
nand U44995 (N_44995,N_41575,N_40389);
nand U44996 (N_44996,N_40765,N_42381);
or U44997 (N_44997,N_42035,N_40125);
nand U44998 (N_44998,N_40548,N_41142);
xor U44999 (N_44999,N_41042,N_41805);
or U45000 (N_45000,N_43721,N_43073);
and U45001 (N_45001,N_43404,N_44369);
or U45002 (N_45002,N_44842,N_44513);
nor U45003 (N_45003,N_43262,N_43441);
xor U45004 (N_45004,N_43586,N_43329);
xnor U45005 (N_45005,N_43770,N_44496);
nand U45006 (N_45006,N_43622,N_44273);
xnor U45007 (N_45007,N_43896,N_44361);
xor U45008 (N_45008,N_43728,N_43264);
or U45009 (N_45009,N_42911,N_43410);
xnor U45010 (N_45010,N_44218,N_42908);
or U45011 (N_45011,N_43347,N_43708);
xor U45012 (N_45012,N_44300,N_42581);
xor U45013 (N_45013,N_44096,N_43711);
nor U45014 (N_45014,N_43575,N_43689);
or U45015 (N_45015,N_42561,N_42902);
nand U45016 (N_45016,N_43204,N_43255);
nor U45017 (N_45017,N_43312,N_44154);
and U45018 (N_45018,N_44325,N_44788);
nor U45019 (N_45019,N_44698,N_43577);
and U45020 (N_45020,N_42934,N_43341);
nor U45021 (N_45021,N_44954,N_44946);
or U45022 (N_45022,N_44538,N_42513);
or U45023 (N_45023,N_44399,N_42876);
nor U45024 (N_45024,N_44964,N_43185);
or U45025 (N_45025,N_44802,N_43106);
nand U45026 (N_45026,N_42963,N_42767);
nor U45027 (N_45027,N_44173,N_44792);
nor U45028 (N_45028,N_44515,N_44180);
nand U45029 (N_45029,N_44874,N_42759);
xor U45030 (N_45030,N_43716,N_43457);
and U45031 (N_45031,N_44326,N_43256);
and U45032 (N_45032,N_43922,N_42724);
or U45033 (N_45033,N_44799,N_44794);
and U45034 (N_45034,N_43873,N_44229);
and U45035 (N_45035,N_43701,N_44329);
nand U45036 (N_45036,N_43828,N_43836);
nand U45037 (N_45037,N_42900,N_44161);
nand U45038 (N_45038,N_44042,N_43832);
xnor U45039 (N_45039,N_43623,N_42854);
and U45040 (N_45040,N_43435,N_43222);
nand U45041 (N_45041,N_44729,N_44781);
and U45042 (N_45042,N_42933,N_44331);
xor U45043 (N_45043,N_42804,N_42906);
or U45044 (N_45044,N_43205,N_44335);
or U45045 (N_45045,N_43128,N_43574);
or U45046 (N_45046,N_43459,N_42922);
nor U45047 (N_45047,N_44672,N_43317);
and U45048 (N_45048,N_44424,N_42889);
nand U45049 (N_45049,N_43121,N_43150);
xor U45050 (N_45050,N_43501,N_42962);
or U45051 (N_45051,N_43985,N_44212);
and U45052 (N_45052,N_43562,N_42572);
nand U45053 (N_45053,N_44140,N_43334);
nand U45054 (N_45054,N_44742,N_44385);
nand U45055 (N_45055,N_43916,N_43883);
or U45056 (N_45056,N_44434,N_42744);
nand U45057 (N_45057,N_44535,N_44084);
or U45058 (N_45058,N_44452,N_44083);
or U45059 (N_45059,N_44055,N_42692);
nand U45060 (N_45060,N_42520,N_43880);
nand U45061 (N_45061,N_44275,N_43059);
or U45062 (N_45062,N_44391,N_42660);
and U45063 (N_45063,N_43432,N_44689);
nand U45064 (N_45064,N_43652,N_44172);
or U45065 (N_45065,N_43236,N_44403);
xnor U45066 (N_45066,N_42868,N_43738);
xnor U45067 (N_45067,N_44056,N_43902);
and U45068 (N_45068,N_42815,N_42618);
nand U45069 (N_45069,N_42931,N_43010);
xor U45070 (N_45070,N_43780,N_43585);
or U45071 (N_45071,N_42993,N_44857);
nor U45072 (N_45072,N_44838,N_44474);
or U45073 (N_45073,N_43162,N_43642);
and U45074 (N_45074,N_42687,N_44157);
and U45075 (N_45075,N_43012,N_43604);
and U45076 (N_45076,N_43066,N_42604);
xor U45077 (N_45077,N_44195,N_42644);
nand U45078 (N_45078,N_44904,N_44599);
and U45079 (N_45079,N_43451,N_44415);
and U45080 (N_45080,N_43176,N_44253);
nand U45081 (N_45081,N_44345,N_44339);
nor U45082 (N_45082,N_44031,N_42536);
and U45083 (N_45083,N_43508,N_42585);
nand U45084 (N_45084,N_43164,N_42826);
nor U45085 (N_45085,N_42949,N_43583);
nand U45086 (N_45086,N_44736,N_44882);
or U45087 (N_45087,N_44120,N_43438);
xnor U45088 (N_45088,N_42714,N_44125);
and U45089 (N_45089,N_44845,N_43251);
nand U45090 (N_45090,N_44576,N_44541);
and U45091 (N_45091,N_43151,N_44092);
or U45092 (N_45092,N_44859,N_44081);
nor U45093 (N_45093,N_43077,N_44138);
and U45094 (N_45094,N_43299,N_44468);
xor U45095 (N_45095,N_44628,N_43439);
or U45096 (N_45096,N_43300,N_44054);
nor U45097 (N_45097,N_43355,N_43821);
and U45098 (N_45098,N_44205,N_43303);
nand U45099 (N_45099,N_43384,N_42700);
or U45100 (N_45100,N_43993,N_42816);
nor U45101 (N_45101,N_43213,N_43744);
nand U45102 (N_45102,N_44871,N_43815);
nand U45103 (N_45103,N_44320,N_44019);
xor U45104 (N_45104,N_42723,N_43506);
xor U45105 (N_45105,N_44677,N_44841);
nand U45106 (N_45106,N_43265,N_42917);
nor U45107 (N_45107,N_44077,N_43816);
or U45108 (N_45108,N_44804,N_44421);
xor U45109 (N_45109,N_43737,N_43153);
nor U45110 (N_45110,N_42718,N_44309);
or U45111 (N_45111,N_42632,N_43216);
xor U45112 (N_45112,N_43041,N_42684);
or U45113 (N_45113,N_44316,N_43084);
nand U45114 (N_45114,N_42576,N_43311);
xnor U45115 (N_45115,N_43131,N_42909);
and U45116 (N_45116,N_43470,N_43136);
nand U45117 (N_45117,N_43129,N_42651);
nand U45118 (N_45118,N_44649,N_43759);
nand U45119 (N_45119,N_44133,N_44990);
xnor U45120 (N_45120,N_43733,N_44569);
nand U45121 (N_45121,N_43378,N_44759);
and U45122 (N_45122,N_42741,N_44503);
or U45123 (N_45123,N_43989,N_43923);
nand U45124 (N_45124,N_42831,N_43731);
nor U45125 (N_45125,N_42810,N_44485);
nor U45126 (N_45126,N_43812,N_42626);
nor U45127 (N_45127,N_42874,N_43603);
and U45128 (N_45128,N_42600,N_42838);
or U45129 (N_45129,N_44635,N_43418);
xor U45130 (N_45130,N_44997,N_43058);
or U45131 (N_45131,N_44302,N_43539);
nand U45132 (N_45132,N_44591,N_42664);
and U45133 (N_45133,N_44948,N_44923);
nand U45134 (N_45134,N_44010,N_44365);
nand U45135 (N_45135,N_42702,N_43067);
nand U45136 (N_45136,N_44596,N_44098);
nor U45137 (N_45137,N_44900,N_43643);
and U45138 (N_45138,N_43540,N_42515);
nor U45139 (N_45139,N_42596,N_44147);
nand U45140 (N_45140,N_43627,N_44961);
and U45141 (N_45141,N_43653,N_43638);
or U45142 (N_45142,N_43934,N_43807);
xor U45143 (N_45143,N_43482,N_43487);
nor U45144 (N_45144,N_42638,N_43290);
nor U45145 (N_45145,N_43805,N_43661);
and U45146 (N_45146,N_43633,N_44594);
nand U45147 (N_45147,N_44240,N_42637);
xnor U45148 (N_45148,N_42758,N_42983);
or U45149 (N_45149,N_43776,N_44289);
or U45150 (N_45150,N_43935,N_44484);
xor U45151 (N_45151,N_44370,N_43109);
xnor U45152 (N_45152,N_44855,N_43184);
nor U45153 (N_45153,N_43739,N_44749);
or U45154 (N_45154,N_44200,N_42849);
nor U45155 (N_45155,N_43849,N_43085);
nand U45156 (N_45156,N_42595,N_44294);
xor U45157 (N_45157,N_42850,N_44851);
nor U45158 (N_45158,N_44069,N_44895);
or U45159 (N_45159,N_43270,N_43709);
xnor U45160 (N_45160,N_43007,N_43964);
nor U45161 (N_45161,N_42589,N_42803);
nand U45162 (N_45162,N_43940,N_44561);
and U45163 (N_45163,N_42624,N_43336);
nand U45164 (N_45164,N_44057,N_43434);
nand U45165 (N_45165,N_43137,N_42777);
or U45166 (N_45166,N_43596,N_42806);
and U45167 (N_45167,N_44786,N_43226);
xnor U45168 (N_45168,N_43949,N_44975);
xnor U45169 (N_45169,N_43785,N_44824);
xnor U45170 (N_45170,N_43281,N_44566);
xor U45171 (N_45171,N_42739,N_44864);
and U45172 (N_45172,N_44626,N_44080);
xnor U45173 (N_45173,N_43760,N_44629);
nor U45174 (N_45174,N_44683,N_44268);
and U45175 (N_45175,N_43984,N_44521);
nor U45176 (N_45176,N_43907,N_43887);
xor U45177 (N_45177,N_43001,N_43833);
xnor U45178 (N_45178,N_42640,N_43302);
nor U45179 (N_45179,N_43296,N_42516);
nand U45180 (N_45180,N_43587,N_44870);
nor U45181 (N_45181,N_44165,N_44317);
and U45182 (N_45182,N_44723,N_43177);
nand U45183 (N_45183,N_44464,N_43551);
and U45184 (N_45184,N_44708,N_42689);
nor U45185 (N_45185,N_44518,N_43790);
and U45186 (N_45186,N_43552,N_44592);
and U45187 (N_45187,N_43869,N_43192);
nand U45188 (N_45188,N_43011,N_44145);
xnor U45189 (N_45189,N_43602,N_44658);
and U45190 (N_45190,N_42812,N_42558);
nor U45191 (N_45191,N_43096,N_44358);
xor U45192 (N_45192,N_44122,N_44686);
xnor U45193 (N_45193,N_43282,N_43283);
or U45194 (N_45194,N_44426,N_43474);
nor U45195 (N_45195,N_43069,N_43544);
nand U45196 (N_45196,N_44116,N_43771);
nand U45197 (N_45197,N_43367,N_42545);
or U45198 (N_45198,N_43693,N_44453);
xor U45199 (N_45199,N_44696,N_43820);
or U45200 (N_45200,N_44374,N_43690);
and U45201 (N_45201,N_43286,N_42981);
xnor U45202 (N_45202,N_44016,N_43895);
nand U45203 (N_45203,N_42552,N_43091);
or U45204 (N_45204,N_44706,N_43695);
nand U45205 (N_45205,N_43855,N_43301);
nor U45206 (N_45206,N_43114,N_44507);
nand U45207 (N_45207,N_44447,N_43169);
nor U45208 (N_45208,N_42623,N_42607);
xor U45209 (N_45209,N_43379,N_43996);
xnor U45210 (N_45210,N_43528,N_43571);
nor U45211 (N_45211,N_44030,N_43764);
nand U45212 (N_45212,N_44489,N_43829);
nor U45213 (N_45213,N_43972,N_43694);
nand U45214 (N_45214,N_43796,N_44292);
nor U45215 (N_45215,N_43092,N_43406);
nor U45216 (N_45216,N_43392,N_42913);
nand U45217 (N_45217,N_43699,N_43515);
nand U45218 (N_45218,N_43810,N_42837);
and U45219 (N_45219,N_44709,N_42857);
nor U45220 (N_45220,N_43080,N_44366);
nand U45221 (N_45221,N_43813,N_42650);
xor U45222 (N_45222,N_42997,N_43189);
and U45223 (N_45223,N_43068,N_43789);
xnor U45224 (N_45224,N_44201,N_44796);
and U45225 (N_45225,N_43182,N_42925);
xnor U45226 (N_45226,N_44045,N_43385);
or U45227 (N_45227,N_43013,N_44735);
nor U45228 (N_45228,N_44136,N_43635);
or U45229 (N_45229,N_43969,N_43202);
and U45230 (N_45230,N_43060,N_44048);
and U45231 (N_45231,N_42707,N_44621);
or U45232 (N_45232,N_44863,N_43391);
nand U45233 (N_45233,N_44891,N_43992);
nand U45234 (N_45234,N_44088,N_44390);
xnor U45235 (N_45235,N_44657,N_43580);
or U45236 (N_45236,N_43997,N_42659);
nand U45237 (N_45237,N_43518,N_44674);
xnor U45238 (N_45238,N_42742,N_42961);
xor U45239 (N_45239,N_43514,N_42609);
xnor U45240 (N_45240,N_44360,N_42706);
or U45241 (N_45241,N_43665,N_44356);
xor U45242 (N_45242,N_44440,N_44108);
nand U45243 (N_45243,N_42932,N_44710);
and U45244 (N_45244,N_42645,N_42508);
or U45245 (N_45245,N_42616,N_43030);
nand U45246 (N_45246,N_42699,N_43977);
and U45247 (N_45247,N_44494,N_43982);
nand U45248 (N_45248,N_44005,N_42543);
nor U45249 (N_45249,N_44527,N_44156);
nor U45250 (N_45250,N_43372,N_43473);
nor U45251 (N_45251,N_42952,N_44446);
nor U45252 (N_45252,N_42630,N_44359);
and U45253 (N_45253,N_44226,N_44101);
or U45254 (N_45254,N_43364,N_44957);
and U45255 (N_45255,N_43707,N_42903);
xnor U45256 (N_45256,N_43382,N_44504);
nand U45257 (N_45257,N_43932,N_42860);
nor U45258 (N_45258,N_43168,N_44304);
nand U45259 (N_45259,N_44064,N_43053);
nor U45260 (N_45260,N_43125,N_44328);
xor U45261 (N_45261,N_44892,N_44746);
or U45262 (N_45262,N_44579,N_42597);
or U45263 (N_45263,N_43970,N_42950);
and U45264 (N_45264,N_43083,N_44725);
and U45265 (N_45265,N_42780,N_43822);
nand U45266 (N_45266,N_43777,N_44624);
nand U45267 (N_45267,N_42918,N_43995);
xnor U45268 (N_45268,N_44004,N_44124);
nor U45269 (N_45269,N_44803,N_44000);
nor U45270 (N_45270,N_42720,N_44822);
nand U45271 (N_45271,N_44393,N_44667);
nor U45272 (N_45272,N_44071,N_43976);
nor U45273 (N_45273,N_44918,N_43803);
nor U45274 (N_45274,N_44298,N_43036);
xnor U45275 (N_45275,N_44694,N_43081);
and U45276 (N_45276,N_43043,N_43052);
nor U45277 (N_45277,N_44319,N_44992);
and U45278 (N_45278,N_44881,N_43858);
nor U45279 (N_45279,N_42652,N_43353);
and U45280 (N_45280,N_43107,N_43998);
and U45281 (N_45281,N_43843,N_44899);
and U45282 (N_45282,N_42987,N_43087);
nand U45283 (N_45283,N_44619,N_43867);
and U45284 (N_45284,N_44811,N_42795);
or U45285 (N_45285,N_44241,N_44903);
nor U45286 (N_45286,N_42984,N_43217);
nor U45287 (N_45287,N_44480,N_42691);
nand U45288 (N_45288,N_44297,N_43930);
and U45289 (N_45289,N_42786,N_43070);
xnor U45290 (N_45290,N_42677,N_44678);
nor U45291 (N_45291,N_44557,N_43878);
and U45292 (N_45292,N_44754,N_42731);
nand U45293 (N_45293,N_43297,N_44721);
xnor U45294 (N_45294,N_42639,N_44471);
nor U45295 (N_45295,N_42544,N_44753);
or U45296 (N_45296,N_43553,N_42512);
or U45297 (N_45297,N_42910,N_43090);
xnor U45298 (N_45298,N_44321,N_43399);
and U45299 (N_45299,N_44087,N_43720);
nor U45300 (N_45300,N_44565,N_42540);
or U45301 (N_45301,N_44828,N_44930);
nand U45302 (N_45302,N_43729,N_44431);
xor U45303 (N_45303,N_44276,N_43956);
and U45304 (N_45304,N_42856,N_42500);
xor U45305 (N_45305,N_43826,N_43187);
and U45306 (N_45306,N_44944,N_43675);
and U45307 (N_45307,N_44969,N_43327);
nor U45308 (N_45308,N_44301,N_43590);
xor U45309 (N_45309,N_44143,N_44648);
or U45310 (N_45310,N_42631,N_44763);
nor U45311 (N_45311,N_42915,N_44551);
nor U45312 (N_45312,N_44597,N_43304);
nand U45313 (N_45313,N_44656,N_44135);
xor U45314 (N_45314,N_43320,N_43914);
xor U45315 (N_45315,N_42822,N_42662);
nand U45316 (N_45316,N_44502,N_44916);
or U45317 (N_45317,N_43680,N_43337);
xnor U45318 (N_45318,N_44885,N_44931);
xnor U45319 (N_45319,N_44953,N_44430);
xnor U45320 (N_45320,N_42790,N_44266);
and U45321 (N_45321,N_43333,N_44442);
or U45322 (N_45322,N_44112,N_42878);
and U45323 (N_45323,N_44761,N_44979);
or U45324 (N_45324,N_43845,N_44872);
nor U45325 (N_45325,N_42887,N_43409);
nand U45326 (N_45326,N_44645,N_43240);
and U45327 (N_45327,N_44236,N_44843);
xnor U45328 (N_45328,N_44449,N_43948);
and U45329 (N_45329,N_43747,N_43783);
nand U45330 (N_45330,N_43498,N_44181);
or U45331 (N_45331,N_43545,N_42764);
and U45332 (N_45332,N_44014,N_44868);
nor U45333 (N_45333,N_43140,N_43274);
and U45334 (N_45334,N_43718,N_42892);
xor U45335 (N_45335,N_43062,N_42808);
xnor U45336 (N_45336,N_43028,N_44582);
or U45337 (N_45337,N_43079,N_43933);
and U45338 (N_45338,N_42970,N_43659);
or U45339 (N_45339,N_43157,N_44396);
and U45340 (N_45340,N_44704,N_43298);
nand U45341 (N_45341,N_42518,N_44663);
nor U45342 (N_45342,N_44281,N_42890);
and U45343 (N_45343,N_42549,N_43014);
nand U45344 (N_45344,N_43133,N_44549);
or U45345 (N_45345,N_44420,N_44978);
or U45346 (N_45346,N_43247,N_43322);
and U45347 (N_45347,N_44685,N_42912);
xor U45348 (N_45348,N_43448,N_44475);
or U45349 (N_45349,N_44970,N_44972);
and U45350 (N_45350,N_44270,N_44225);
or U45351 (N_45351,N_44085,N_42919);
nand U45352 (N_45352,N_44114,N_43521);
nand U45353 (N_45353,N_43316,N_44676);
xnor U45354 (N_45354,N_44210,N_44026);
xor U45355 (N_45355,N_44983,N_44196);
xnor U45356 (N_45356,N_44158,N_44137);
nor U45357 (N_45357,N_44738,N_44015);
or U45358 (N_45358,N_44939,N_42756);
xnor U45359 (N_45359,N_44230,N_43427);
or U45360 (N_45360,N_43231,N_44805);
nor U45361 (N_45361,N_42798,N_44717);
and U45362 (N_45362,N_43368,N_42665);
xnor U45363 (N_45363,N_43359,N_43033);
nor U45364 (N_45364,N_44833,N_43314);
xor U45365 (N_45365,N_44520,N_43152);
and U45366 (N_45366,N_42841,N_44884);
and U45367 (N_45367,N_42990,N_43775);
and U45368 (N_45368,N_43741,N_43403);
xor U45369 (N_45369,N_44966,N_43667);
nor U45370 (N_45370,N_43560,N_44126);
or U45371 (N_45371,N_44283,N_43363);
or U45372 (N_45372,N_43619,N_43126);
or U45373 (N_45373,N_43476,N_43509);
xor U45374 (N_45374,N_42907,N_42884);
xor U45375 (N_45375,N_43488,N_44634);
xnor U45376 (N_45376,N_44705,N_44911);
xor U45377 (N_45377,N_44510,N_42785);
nand U45378 (N_45378,N_42772,N_42783);
nand U45379 (N_45379,N_42958,N_43422);
nor U45380 (N_45380,N_43567,N_43851);
nor U45381 (N_45381,N_43749,N_43788);
xnor U45382 (N_45382,N_44595,N_43120);
xnor U45383 (N_45383,N_42740,N_43158);
or U45384 (N_45384,N_43513,N_44675);
nand U45385 (N_45385,N_44713,N_42567);
or U45386 (N_45386,N_42554,N_43962);
nand U45387 (N_45387,N_43987,N_44668);
and U45388 (N_45388,N_44888,N_44839);
and U45389 (N_45389,N_44233,N_44461);
nand U45390 (N_45390,N_43097,N_44740);
xor U45391 (N_45391,N_44901,N_42534);
xor U45392 (N_45392,N_43541,N_44347);
xnor U45393 (N_45393,N_44323,N_44248);
nor U45394 (N_45394,N_43980,N_42847);
or U45395 (N_45395,N_43955,N_43160);
and U45396 (N_45396,N_42619,N_43734);
or U45397 (N_45397,N_43724,N_44878);
nand U45398 (N_45398,N_43736,N_42974);
or U45399 (N_45399,N_42773,N_44915);
or U45400 (N_45400,N_44287,N_43559);
or U45401 (N_45401,N_44211,N_43674);
nor U45402 (N_45402,N_42673,N_44586);
and U45403 (N_45403,N_44183,N_42683);
and U45404 (N_45404,N_42846,N_42929);
xor U45405 (N_45405,N_42598,N_43573);
or U45406 (N_45406,N_44950,N_42730);
xor U45407 (N_45407,N_44247,N_44655);
nor U45408 (N_45408,N_42827,N_43357);
or U45409 (N_45409,N_43038,N_44422);
or U45410 (N_45410,N_43397,N_44076);
xnor U45411 (N_45411,N_43862,N_43871);
and U45412 (N_45412,N_42805,N_44741);
xnor U45413 (N_45413,N_43293,N_44581);
and U45414 (N_45414,N_44936,N_44039);
and U45415 (N_45415,N_44227,N_43257);
or U45416 (N_45416,N_44898,N_43877);
and U45417 (N_45417,N_44920,N_43852);
or U45418 (N_45418,N_43630,N_43782);
nor U45419 (N_45419,N_44777,N_43229);
and U45420 (N_45420,N_43913,N_43468);
nor U45421 (N_45421,N_42557,N_44558);
nand U45422 (N_45422,N_43755,N_44590);
nor U45423 (N_45423,N_43872,N_43318);
and U45424 (N_45424,N_43276,N_42694);
or U45425 (N_45425,N_42748,N_43496);
nand U45426 (N_45426,N_44144,N_43906);
xor U45427 (N_45427,N_42555,N_44271);
xor U45428 (N_45428,N_44651,N_44769);
xnor U45429 (N_45429,N_44531,N_44118);
xor U45430 (N_45430,N_44070,N_43389);
and U45431 (N_45431,N_43569,N_44783);
and U45432 (N_45432,N_44486,N_43212);
nand U45433 (N_45433,N_44318,N_42574);
and U45434 (N_45434,N_42882,N_44615);
or U45435 (N_45435,N_44179,N_44208);
and U45436 (N_45436,N_43889,N_43309);
and U45437 (N_45437,N_44261,N_42625);
and U45438 (N_45438,N_42590,N_42573);
and U45439 (N_45439,N_44330,N_43103);
nand U45440 (N_45440,N_43884,N_43032);
xor U45441 (N_45441,N_44718,N_44046);
nand U45442 (N_45442,N_44673,N_42503);
nor U45443 (N_45443,N_43328,N_43793);
xor U45444 (N_45444,N_43986,N_44896);
nor U45445 (N_45445,N_43864,N_43319);
or U45446 (N_45446,N_42845,N_43617);
nor U45447 (N_45447,N_42768,N_44379);
or U45448 (N_45448,N_44382,N_43668);
nor U45449 (N_45449,N_43047,N_43526);
or U45450 (N_45450,N_44130,N_43751);
and U45451 (N_45451,N_43792,N_43905);
xnor U45452 (N_45452,N_43655,N_44416);
nor U45453 (N_45453,N_44697,N_44780);
or U45454 (N_45454,N_43074,N_44109);
xnor U45455 (N_45455,N_43387,N_44355);
or U45456 (N_45456,N_42789,N_43108);
xnor U45457 (N_45457,N_42871,N_44166);
xor U45458 (N_45458,N_43095,N_44467);
nor U45459 (N_45459,N_43165,N_43965);
and U45460 (N_45460,N_43063,N_43576);
xnor U45461 (N_45461,N_43809,N_44061);
nand U45462 (N_45462,N_43154,N_43003);
and U45463 (N_45463,N_44745,N_44767);
or U45464 (N_45464,N_42797,N_44666);
nor U45465 (N_45465,N_44387,N_44222);
or U45466 (N_45466,N_44381,N_44831);
or U45467 (N_45467,N_44947,N_42843);
nor U45468 (N_45468,N_42899,N_42599);
nor U45469 (N_45469,N_43598,N_44282);
and U45470 (N_45470,N_43522,N_43542);
or U45471 (N_45471,N_43436,N_42979);
nor U45472 (N_45472,N_44540,N_44193);
and U45473 (N_45473,N_44938,N_42710);
nand U45474 (N_45474,N_43774,N_42943);
or U45475 (N_45475,N_44025,N_43188);
xor U45476 (N_45476,N_44216,N_44349);
nand U45477 (N_45477,N_43344,N_44907);
and U45478 (N_45478,N_44530,N_43658);
xor U45479 (N_45479,N_44100,N_44768);
and U45480 (N_45480,N_43072,N_44034);
or U45481 (N_45481,N_44257,N_44231);
and U45482 (N_45482,N_43988,N_44752);
xnor U45483 (N_45483,N_43768,N_42666);
nor U45484 (N_45484,N_44073,N_44217);
or U45485 (N_45485,N_44996,N_44963);
and U45486 (N_45486,N_42914,N_42788);
and U45487 (N_45487,N_44198,N_44760);
or U45488 (N_45488,N_43897,N_42769);
xnor U45489 (N_45489,N_44989,N_44880);
xnor U45490 (N_45490,N_43929,N_42794);
nand U45491 (N_45491,N_44984,N_43315);
or U45492 (N_45492,N_43719,N_43786);
xnor U45493 (N_45493,N_43424,N_43161);
and U45494 (N_45494,N_44052,N_43237);
nor U45495 (N_45495,N_42813,N_42828);
xnor U45496 (N_45496,N_42733,N_44798);
or U45497 (N_45497,N_43742,N_42824);
nand U45498 (N_45498,N_44607,N_43191);
xnor U45499 (N_45499,N_44568,N_44693);
xnor U45500 (N_45500,N_43022,N_44601);
nor U45501 (N_45501,N_42541,N_44127);
and U45502 (N_45502,N_42553,N_43629);
nand U45503 (N_45503,N_44889,N_44679);
nand U45504 (N_45504,N_43863,N_44498);
or U45505 (N_45505,N_42746,N_43477);
xor U45506 (N_45506,N_43479,N_44778);
xnor U45507 (N_45507,N_43859,N_42861);
xor U45508 (N_45508,N_43149,N_43974);
nor U45509 (N_45509,N_43287,N_44800);
and U45510 (N_45510,N_43263,N_43447);
or U45511 (N_45511,N_43691,N_42667);
xor U45512 (N_45512,N_44357,N_42947);
and U45513 (N_45513,N_44460,N_43565);
nor U45514 (N_45514,N_42655,N_43846);
xor U45515 (N_45515,N_44747,N_44436);
or U45516 (N_45516,N_42762,N_44040);
and U45517 (N_45517,N_43279,N_43795);
or U45518 (N_45518,N_44351,N_43208);
nor U45519 (N_45519,N_42749,N_44701);
nor U45520 (N_45520,N_44921,N_43093);
and U45521 (N_45521,N_42605,N_43163);
xnor U45522 (N_45522,N_44620,N_44750);
and U45523 (N_45523,N_44734,N_44336);
or U45524 (N_45524,N_42593,N_42923);
or U45525 (N_45525,N_44327,N_42757);
nor U45526 (N_45526,N_43750,N_44574);
and U45527 (N_45527,N_43346,N_43454);
nand U45528 (N_45528,N_44219,N_44184);
nand U45529 (N_45529,N_44263,N_43275);
and U45530 (N_45530,N_42940,N_43049);
nand U45531 (N_45531,N_42770,N_43469);
or U45532 (N_45532,N_42701,N_42737);
nor U45533 (N_45533,N_44945,N_43610);
or U45534 (N_45534,N_42760,N_43866);
nor U45535 (N_45535,N_44876,N_44623);
nand U45536 (N_45536,N_44239,N_43706);
or U45537 (N_45537,N_42743,N_44714);
xnor U45538 (N_45538,N_43171,N_43609);
nor U45539 (N_45539,N_44646,N_43115);
and U45540 (N_45540,N_43278,N_44067);
xor U45541 (N_45541,N_44252,N_43102);
nand U45542 (N_45542,N_43650,N_44692);
nor U45543 (N_45543,N_43860,N_44913);
xnor U45544 (N_45544,N_42862,N_43402);
nor U45545 (N_45545,N_44570,N_43383);
nor U45546 (N_45546,N_42867,N_44417);
or U45547 (N_45547,N_43549,N_44762);
nor U45548 (N_45548,N_43321,N_42643);
or U45549 (N_45549,N_42591,N_42620);
nor U45550 (N_45550,N_42728,N_44008);
and U45551 (N_45551,N_43040,N_44131);
nand U45552 (N_45552,N_42654,N_42627);
and U45553 (N_45553,N_44825,N_43966);
nand U45554 (N_45554,N_43183,N_43599);
and U45555 (N_45555,N_43766,N_44307);
and U45556 (N_45556,N_43443,N_43681);
xnor U45557 (N_45557,N_44631,N_42784);
or U45558 (N_45558,N_42975,N_44886);
and U45559 (N_45559,N_44063,N_43639);
and U45560 (N_45560,N_43957,N_43745);
nand U45561 (N_45561,N_42679,N_44603);
xor U45562 (N_45562,N_44524,N_43692);
nand U45563 (N_45563,N_44012,N_44378);
and U45564 (N_45564,N_44593,N_44203);
nand U45565 (N_45565,N_44238,N_44097);
nor U45566 (N_45566,N_42953,N_44512);
nand U45567 (N_45567,N_43330,N_43124);
xor U45568 (N_45568,N_43017,N_43611);
or U45569 (N_45569,N_44680,N_44371);
and U45570 (N_45570,N_43112,N_44829);
or U45571 (N_45571,N_43398,N_43006);
or U45572 (N_45572,N_42656,N_43767);
nand U45573 (N_45573,N_42719,N_44353);
xor U45574 (N_45574,N_42825,N_42542);
and U45575 (N_45575,N_44625,N_43370);
and U45576 (N_45576,N_44338,N_43641);
nor U45577 (N_45577,N_44785,N_44142);
nor U45578 (N_45578,N_43348,N_44712);
nor U45579 (N_45579,N_44977,N_44837);
nand U45580 (N_45580,N_44633,N_44472);
and U45581 (N_45581,N_44299,N_44149);
nor U45582 (N_45582,N_43462,N_43752);
or U45583 (N_45583,N_44584,N_42603);
nor U45584 (N_45584,N_43313,N_44974);
and U45585 (N_45585,N_42752,N_44772);
xor U45586 (N_45586,N_43220,N_43142);
xor U45587 (N_45587,N_43503,N_43221);
nand U45588 (N_45588,N_43563,N_43682);
or U45589 (N_45589,N_44727,N_44826);
xor U45590 (N_45590,N_43952,N_43145);
or U45591 (N_45591,N_44234,N_42525);
xor U45592 (N_45592,N_43730,N_42550);
and U45593 (N_45593,N_44079,N_42509);
nand U45594 (N_45594,N_43890,N_44563);
nand U45595 (N_45595,N_42930,N_44443);
and U45596 (N_45596,N_42880,N_43360);
nand U45597 (N_45597,N_42649,N_44389);
and U45598 (N_45598,N_43825,N_43620);
and U45599 (N_45599,N_43472,N_44169);
and U45600 (N_45600,N_44505,N_44894);
nor U45601 (N_45601,N_42898,N_42965);
nor U45602 (N_45602,N_42592,N_42866);
or U45603 (N_45603,N_43122,N_43156);
and U45604 (N_45604,N_43582,N_44103);
nor U45605 (N_45605,N_43277,N_44779);
xor U45606 (N_45606,N_43307,N_43248);
nand U45607 (N_45607,N_42885,N_43938);
xnor U45608 (N_45608,N_42865,N_42506);
or U45609 (N_45609,N_43511,N_42935);
nand U45610 (N_45610,N_42575,N_44258);
xor U45611 (N_45611,N_44707,N_44265);
and U45612 (N_45612,N_44532,N_43148);
nor U45613 (N_45613,N_42661,N_44782);
nor U45614 (N_45614,N_44908,N_43533);
and U45615 (N_45615,N_43478,N_43198);
nand U45616 (N_45616,N_43483,N_43394);
xnor U45617 (N_45617,N_42792,N_43735);
and U45618 (N_45618,N_44095,N_42583);
and U45619 (N_45619,N_44820,N_44139);
and U45620 (N_45620,N_42569,N_44267);
or U45621 (N_45621,N_44167,N_44830);
xnor U45622 (N_45622,N_44795,N_43717);
xor U45623 (N_45623,N_44852,N_43566);
and U45624 (N_45624,N_42968,N_42897);
nand U45625 (N_45625,N_43361,N_43524);
xor U45626 (N_45626,N_43688,N_44414);
xor U45627 (N_45627,N_43193,N_43663);
and U45628 (N_45628,N_43570,N_43159);
nand U45629 (N_45629,N_42502,N_43271);
and U45630 (N_45630,N_44600,N_43016);
nor U45631 (N_45631,N_43376,N_43525);
and U45632 (N_45632,N_42991,N_43676);
or U45633 (N_45633,N_43640,N_44246);
xor U45634 (N_45634,N_43250,N_43910);
and U45635 (N_45635,N_44435,N_44341);
xor U45636 (N_45636,N_42566,N_42998);
nor U45637 (N_45637,N_42778,N_42729);
nor U45638 (N_45638,N_42941,N_44726);
xor U45639 (N_45639,N_43794,N_44699);
and U45640 (N_45640,N_44428,N_43686);
nor U45641 (N_45641,N_43267,N_44419);
and U45642 (N_45642,N_43892,N_44832);
nand U45643 (N_45643,N_43207,N_44410);
or U45644 (N_45644,N_43076,N_43417);
xnor U45645 (N_45645,N_42966,N_43197);
xor U45646 (N_45646,N_44571,N_42834);
and U45647 (N_45647,N_43677,N_43272);
and U45648 (N_45648,N_43211,N_44639);
xnor U45649 (N_45649,N_43349,N_43340);
nand U45650 (N_45650,N_44438,N_43517);
nor U45651 (N_45651,N_44711,N_44243);
xor U45652 (N_45652,N_44223,N_43536);
and U45653 (N_45653,N_43891,N_43754);
nor U45654 (N_45654,N_43614,N_43345);
and U45655 (N_45655,N_42524,N_43179);
or U45656 (N_45656,N_43261,N_44511);
xor U45657 (N_45657,N_43224,N_44481);
and U45658 (N_45658,N_43113,N_43885);
or U45659 (N_45659,N_43761,N_43463);
and U45660 (N_45660,N_44716,N_42571);
and U45661 (N_45661,N_44809,N_44577);
and U45662 (N_45662,N_43882,N_44703);
nand U45663 (N_45663,N_44854,N_42675);
and U45664 (N_45664,N_43039,N_44956);
or U45665 (N_45665,N_43763,N_44691);
xnor U45666 (N_45666,N_43480,N_42685);
nor U45667 (N_45667,N_44191,N_42836);
nand U45668 (N_45668,N_42705,N_43444);
and U45669 (N_45669,N_43983,N_44102);
nand U45670 (N_45670,N_44013,N_44962);
nand U45671 (N_45671,N_43830,N_43351);
nand U45672 (N_45672,N_43134,N_43823);
nand U45673 (N_45673,N_42951,N_43294);
xnor U45674 (N_45674,N_42537,N_44395);
nand U45675 (N_45675,N_44821,N_44117);
and U45676 (N_45676,N_44072,N_43141);
and U45677 (N_45677,N_43139,N_44342);
and U45678 (N_45678,N_43243,N_42988);
or U45679 (N_45679,N_44279,N_43797);
xor U45680 (N_45680,N_44652,N_43900);
nor U45681 (N_45681,N_43078,N_44988);
nand U45682 (N_45682,N_43118,N_44305);
nand U45683 (N_45683,N_44731,N_44090);
and U45684 (N_45684,N_43791,N_43502);
or U45685 (N_45685,N_43266,N_43854);
xnor U45686 (N_45686,N_44847,N_43031);
and U45687 (N_45687,N_44910,N_44002);
or U45688 (N_45688,N_43835,N_44372);
xnor U45689 (N_45689,N_43657,N_42528);
nor U45690 (N_45690,N_42672,N_44555);
nor U45691 (N_45691,N_43558,N_44280);
and U45692 (N_45692,N_42864,N_43684);
and U45693 (N_45693,N_43492,N_42657);
and U45694 (N_45694,N_44024,N_44380);
or U45695 (N_45695,N_43415,N_44836);
xnor U45696 (N_45696,N_44458,N_44980);
nor U45697 (N_45697,N_44751,N_43086);
and U45698 (N_45698,N_43252,N_43029);
nand U45699 (N_45699,N_43507,N_44099);
nand U45700 (N_45700,N_44286,N_44400);
nand U45701 (N_45701,N_44580,N_44290);
or U45702 (N_45702,N_44991,N_43362);
nand U45703 (N_45703,N_43273,N_43740);
or U45704 (N_45704,N_43756,N_43595);
xnor U45705 (N_45705,N_43917,N_43801);
and U45706 (N_45706,N_42617,N_44020);
nor U45707 (N_45707,N_44288,N_42634);
nand U45708 (N_45708,N_43101,N_43722);
nand U45709 (N_45709,N_44695,N_42578);
nor U45710 (N_45710,N_42964,N_43071);
and U45711 (N_45711,N_44748,N_44844);
nand U45712 (N_45712,N_44251,N_44495);
or U45713 (N_45713,N_44413,N_43591);
and U45714 (N_45714,N_43704,N_44094);
nand U45715 (N_45715,N_43426,N_44044);
xor U45716 (N_45716,N_44255,N_43561);
nor U45717 (N_45717,N_43146,N_43456);
xor U45718 (N_45718,N_44423,N_42835);
or U45719 (N_45719,N_44533,N_42873);
and U45720 (N_45720,N_43234,N_42716);
xor U45721 (N_45721,N_42776,N_43094);
or U45722 (N_45722,N_43230,N_42944);
nand U45723 (N_45723,N_43490,N_42959);
xor U45724 (N_45724,N_44875,N_43110);
or U45725 (N_45725,N_43116,N_43325);
and U45726 (N_45726,N_43753,N_42895);
or U45727 (N_45727,N_43429,N_44638);
or U45728 (N_45728,N_44641,N_44627);
nand U45729 (N_45729,N_43475,N_43214);
or U45730 (N_45730,N_42697,N_42879);
and U45731 (N_45731,N_43850,N_44810);
and U45732 (N_45732,N_44959,N_43493);
or U45733 (N_45733,N_43909,N_42960);
xor U45734 (N_45734,N_44773,N_44982);
xnor U45735 (N_45735,N_44425,N_42976);
or U45736 (N_45736,N_44684,N_43848);
and U45737 (N_45737,N_43632,N_43589);
nor U45738 (N_45738,N_44121,N_43645);
and U45739 (N_45739,N_43608,N_43894);
nor U45740 (N_45740,N_43626,N_44311);
nor U45741 (N_45741,N_43433,N_44148);
nor U45742 (N_45742,N_44765,N_44150);
nand U45743 (N_45743,N_43365,N_42829);
and U45744 (N_45744,N_43235,N_43381);
xnor U45745 (N_45745,N_44564,N_42717);
xnor U45746 (N_45746,N_42559,N_44700);
xor U45747 (N_45747,N_44324,N_44877);
nor U45748 (N_45748,N_42791,N_44032);
xor U45749 (N_45749,N_43950,N_43990);
or U45750 (N_45750,N_44801,N_43666);
nor U45751 (N_45751,N_43099,N_43564);
xor U45752 (N_45752,N_43893,N_42755);
nand U45753 (N_45753,N_44214,N_44572);
or U45754 (N_45754,N_43697,N_43554);
xnor U45755 (N_45755,N_44346,N_43664);
nor U45756 (N_45756,N_42920,N_42504);
nand U45757 (N_45757,N_43242,N_44187);
or U45758 (N_45758,N_44632,N_43180);
nor U45759 (N_45759,N_44616,N_44364);
or U45760 (N_45760,N_44278,N_44537);
nand U45761 (N_45761,N_44993,N_43841);
xor U45762 (N_45762,N_43037,N_42830);
or U45763 (N_45763,N_43971,N_43034);
or U45764 (N_45764,N_42766,N_44291);
xnor U45765 (N_45765,N_44614,N_43486);
nand U45766 (N_45766,N_43332,N_44797);
or U45767 (N_45767,N_44254,N_44522);
and U45768 (N_45768,N_44134,N_43831);
or U45769 (N_45769,N_44861,N_44587);
xor U45770 (N_45770,N_43065,N_44106);
or U45771 (N_45771,N_44146,N_43819);
nand U45772 (N_45772,N_43407,N_44732);
nor U45773 (N_45773,N_44968,N_44334);
xnor U45774 (N_45774,N_42811,N_44194);
and U45775 (N_45775,N_44604,N_44958);
or U45776 (N_45776,N_44650,N_44644);
xnor U45777 (N_45777,N_43015,N_42611);
nand U45778 (N_45778,N_44482,N_42969);
nor U45779 (N_45779,N_44017,N_43411);
xor U45780 (N_45780,N_42703,N_44766);
and U45781 (N_45781,N_43901,N_42648);
xor U45782 (N_45782,N_44322,N_44995);
and U45783 (N_45783,N_43147,N_42989);
xor U45784 (N_45784,N_44905,N_44373);
nand U45785 (N_45785,N_42765,N_44444);
and U45786 (N_45786,N_44035,N_43117);
nand U45787 (N_45787,N_43414,N_43280);
xor U45788 (N_45788,N_43994,N_43834);
and U45789 (N_45789,N_44893,N_44866);
or U45790 (N_45790,N_44499,N_43292);
or U45791 (N_45791,N_42852,N_44919);
or U45792 (N_45792,N_44089,N_44622);
nand U45793 (N_45793,N_44929,N_44162);
and U45794 (N_45794,N_44439,N_44476);
xor U45795 (N_45795,N_43827,N_44284);
xnor U45796 (N_45796,N_42642,N_43408);
or U45797 (N_45797,N_44029,N_44562);
or U45798 (N_45798,N_44999,N_42926);
nand U45799 (N_45799,N_42529,N_43921);
or U45800 (N_45800,N_44724,N_44559);
nand U45801 (N_45801,N_44433,N_42738);
nor U45802 (N_45802,N_42818,N_44509);
nor U45803 (N_45803,N_42533,N_43857);
or U45804 (N_45804,N_44743,N_43172);
or U45805 (N_45805,N_44544,N_43504);
nor U45806 (N_45806,N_42647,N_44160);
nor U45807 (N_45807,N_43430,N_44059);
xnor U45808 (N_45808,N_44189,N_43817);
nor U45809 (N_45809,N_44491,N_44459);
or U45810 (N_45810,N_42551,N_44058);
or U45811 (N_45811,N_44237,N_43285);
nor U45812 (N_45812,N_42995,N_42948);
nor U45813 (N_45813,N_44155,N_44483);
or U45814 (N_45814,N_44909,N_44661);
or U45815 (N_45815,N_44865,N_43918);
or U45816 (N_45816,N_43616,N_42711);
and U45817 (N_45817,N_44981,N_44477);
nand U45818 (N_45818,N_42779,N_44548);
or U45819 (N_45819,N_44647,N_44618);
nand U45820 (N_45820,N_42967,N_44492);
and U45821 (N_45821,N_42510,N_43814);
and U45822 (N_45822,N_43757,N_43042);
xnor U45823 (N_45823,N_44432,N_43915);
nand U45824 (N_45824,N_44343,N_42587);
nor U45825 (N_45825,N_44119,N_44470);
nor U45826 (N_45826,N_44879,N_43532);
xor U45827 (N_45827,N_44517,N_44985);
nand U45828 (N_45828,N_43200,N_43847);
xor U45829 (N_45829,N_42565,N_42690);
xnor U45830 (N_45830,N_44250,N_43875);
or U45831 (N_45831,N_44812,N_44277);
and U45832 (N_45832,N_43098,N_43865);
and U45833 (N_45833,N_42851,N_43529);
and U45834 (N_45834,N_44466,N_44308);
nand U45835 (N_45835,N_42735,N_42531);
xnor U45836 (N_45836,N_43350,N_43898);
xor U45837 (N_45837,N_42601,N_43698);
nand U45838 (N_45838,N_43019,N_43607);
nand U45839 (N_45839,N_44409,N_44259);
and U45840 (N_45840,N_43778,N_44550);
xor U45841 (N_45841,N_43100,N_44091);
nand U45842 (N_45842,N_44897,N_43572);
or U45843 (N_45843,N_44197,N_44406);
nand U45844 (N_45844,N_43371,N_44965);
xnor U45845 (N_45845,N_43519,N_44937);
nand U45846 (N_45846,N_44164,N_44914);
or U45847 (N_45847,N_44552,N_44869);
nor U45848 (N_45848,N_42924,N_44368);
nor U45849 (N_45849,N_44719,N_44141);
and U45850 (N_45850,N_43636,N_44412);
or U45851 (N_45851,N_43352,N_42713);
xor U45852 (N_45852,N_42688,N_42921);
xor U45853 (N_45853,N_43465,N_44313);
nand U45854 (N_45854,N_44405,N_43055);
nand U45855 (N_45855,N_43725,N_42817);
or U45856 (N_45856,N_42863,N_43555);
nand U45857 (N_45857,N_44285,N_44152);
or U45858 (N_45858,N_43765,N_43615);
nand U45859 (N_45859,N_44429,N_43339);
nor U45860 (N_45860,N_42870,N_44455);
xnor U45861 (N_45861,N_44352,N_43497);
nand U45862 (N_45862,N_43625,N_42821);
xor U45863 (N_45863,N_44500,N_43175);
nand U45864 (N_45864,N_43186,N_44793);
or U45865 (N_45865,N_43442,N_43354);
nand U45866 (N_45866,N_43061,N_43453);
or U45867 (N_45867,N_42658,N_43144);
and U45868 (N_45868,N_44404,N_43802);
xor U45869 (N_45869,N_43646,N_44589);
nand U45870 (N_45870,N_44850,N_43556);
and U45871 (N_45871,N_43516,N_43132);
or U45872 (N_45872,N_43947,N_43968);
xnor U45873 (N_45873,N_42646,N_44556);
or U45874 (N_45874,N_42937,N_43908);
xnor U45875 (N_45875,N_44037,N_43057);
or U45876 (N_45876,N_44204,N_44344);
xnor U45877 (N_45877,N_43600,N_43936);
nor U45878 (N_45878,N_44041,N_44151);
and U45879 (N_45879,N_44525,N_44078);
xnor U45880 (N_45880,N_43258,N_44720);
or U45881 (N_45881,N_44224,N_44060);
xnor U45882 (N_45882,N_42793,N_44022);
nand U45883 (N_45883,N_42547,N_43375);
nor U45884 (N_45884,N_43170,N_44840);
nor U45885 (N_45885,N_44526,N_43838);
xnor U45886 (N_45886,N_43678,N_43326);
nor U45887 (N_45887,N_43648,N_43206);
xor U45888 (N_45888,N_43051,N_44175);
or U45889 (N_45889,N_44488,N_44835);
nor U45890 (N_45890,N_44506,N_44295);
or U45891 (N_45891,N_43215,N_43225);
xor U45892 (N_45892,N_43440,N_43238);
or U45893 (N_45893,N_44737,N_44862);
or U45894 (N_45894,N_43662,N_42807);
xor U45895 (N_45895,N_43000,N_43395);
xor U45896 (N_45896,N_44573,N_43904);
nand U45897 (N_45897,N_42568,N_44926);
and U45898 (N_45898,N_43550,N_42514);
xnor U45899 (N_45899,N_44671,N_43592);
nor U45900 (N_45900,N_43975,N_43715);
nor U45901 (N_45901,N_42844,N_44228);
xnor U45902 (N_45902,N_43806,N_43405);
or U45903 (N_45903,N_43961,N_42840);
xor U45904 (N_45904,N_43374,N_42501);
or U45905 (N_45905,N_43811,N_43369);
nor U45906 (N_45906,N_43416,N_42992);
and U45907 (N_45907,N_42745,N_43924);
or U45908 (N_45908,N_44508,N_43605);
and U45909 (N_45909,N_44971,N_44848);
and U45910 (N_45910,N_43269,N_43644);
nor U45911 (N_45911,N_44928,N_44036);
xnor U45912 (N_45912,N_42548,N_44976);
and U45913 (N_45913,N_44445,N_43510);
xor U45914 (N_45914,N_43723,N_44994);
or U45915 (N_45915,N_44182,N_42736);
nor U45916 (N_45916,N_44171,N_44111);
or U45917 (N_45917,N_42883,N_42750);
nand U45918 (N_45918,N_42888,N_44817);
nand U45919 (N_45919,N_44264,N_43194);
nor U45920 (N_45920,N_44375,N_42505);
nand U45921 (N_45921,N_43631,N_42698);
nor U45922 (N_45922,N_42872,N_42751);
xnor U45923 (N_45923,N_44662,N_44986);
nor U45924 (N_45924,N_43773,N_44543);
nor U45925 (N_45925,N_43714,N_43244);
nor U45926 (N_45926,N_42734,N_44943);
xor U45927 (N_45927,N_43581,N_44722);
nand U45928 (N_45928,N_43941,N_44546);
nand U45929 (N_45929,N_43960,N_43702);
nor U45930 (N_45930,N_43669,N_44462);
and U45931 (N_45931,N_43259,N_42610);
or U45932 (N_45932,N_42858,N_43911);
and U45933 (N_45933,N_43289,N_44033);
nor U45934 (N_45934,N_44849,N_43762);
and U45935 (N_45935,N_44049,N_44858);
nor U45936 (N_45936,N_44516,N_42833);
and U45937 (N_45937,N_43104,N_43366);
nor U45938 (N_45938,N_42796,N_42753);
xnor U45939 (N_45939,N_43288,N_44110);
xnor U45940 (N_45940,N_42653,N_44728);
xor U45941 (N_45941,N_43951,N_43173);
or U45942 (N_45942,N_44038,N_43306);
and U45943 (N_45943,N_43166,N_42763);
and U45944 (N_45944,N_43135,N_42996);
xnor U45945 (N_45945,N_43388,N_44867);
nor U45946 (N_45946,N_44186,N_42628);
xor U45947 (N_45947,N_44602,N_43461);
nand U45948 (N_45948,N_44942,N_44935);
or U45949 (N_45949,N_43840,N_44873);
and U45950 (N_45950,N_44654,N_43612);
and U45951 (N_45951,N_44190,N_43579);
and U45952 (N_45952,N_42535,N_43223);
nand U45953 (N_45953,N_44397,N_44383);
nor U45954 (N_45954,N_44170,N_42721);
nand U45955 (N_45955,N_43925,N_43649);
and U45956 (N_45956,N_43945,N_43928);
nor U45957 (N_45957,N_42955,N_43881);
and U45958 (N_45958,N_42564,N_44272);
nor U45959 (N_45959,N_42839,N_42938);
or U45960 (N_45960,N_43531,N_44664);
and U45961 (N_45961,N_44808,N_42781);
nor U45962 (N_45962,N_44856,N_43937);
xnor U45963 (N_45963,N_44104,N_43035);
or U45964 (N_45964,N_43568,N_43853);
xnor U45965 (N_45965,N_42761,N_43241);
nor U45966 (N_45966,N_43481,N_44846);
nor U45967 (N_45967,N_42978,N_43421);
xnor U45968 (N_45968,N_43547,N_42820);
nor U45969 (N_45969,N_43377,N_43870);
and U45970 (N_45970,N_43048,N_44643);
or U45971 (N_45971,N_42875,N_44715);
or U45972 (N_45972,N_44764,N_43588);
or U45973 (N_45973,N_44260,N_43861);
or U45974 (N_45974,N_42855,N_44807);
or U45975 (N_45975,N_43253,N_44973);
and U45976 (N_45976,N_44199,N_42704);
nand U45977 (N_45977,N_43494,N_44027);
or U45978 (N_45978,N_43199,N_44617);
or U45979 (N_45979,N_43005,N_44598);
and U45980 (N_45980,N_43449,N_44043);
nor U45981 (N_45981,N_42517,N_44469);
nor U45982 (N_45982,N_44553,N_44367);
nand U45983 (N_45983,N_44613,N_43452);
and U45984 (N_45984,N_43523,N_44771);
or U45985 (N_45985,N_44086,N_43445);
or U45986 (N_45986,N_42681,N_44128);
and U45987 (N_45987,N_44758,N_44384);
nand U45988 (N_45988,N_43393,N_43842);
nor U45989 (N_45989,N_42546,N_43958);
and U45990 (N_45990,N_42663,N_44456);
and U45991 (N_45991,N_43331,N_42869);
or U45992 (N_45992,N_44448,N_44739);
nor U45993 (N_45993,N_42708,N_44068);
and U45994 (N_45994,N_43050,N_43467);
nor U45995 (N_45995,N_44790,N_43868);
xor U45996 (N_45996,N_43044,N_44611);
and U45997 (N_45997,N_43500,N_44757);
or U45998 (N_45998,N_43088,N_42775);
and U45999 (N_45999,N_42511,N_42747);
nor U46000 (N_46000,N_43021,N_42842);
or U46001 (N_46001,N_44610,N_44787);
or U46002 (N_46002,N_43358,N_44823);
nor U46003 (N_46003,N_43613,N_44376);
xnor U46004 (N_46004,N_43155,N_44411);
nor U46005 (N_46005,N_42612,N_42693);
xor U46006 (N_46006,N_44153,N_43784);
and U46007 (N_46007,N_44534,N_43373);
nand U46008 (N_46008,N_43748,N_43683);
nor U46009 (N_46009,N_43800,N_43685);
xor U46010 (N_46010,N_44348,N_44791);
nand U46011 (N_46011,N_42771,N_42999);
xor U46012 (N_46012,N_44784,N_43946);
or U46013 (N_46013,N_43594,N_42994);
nand U46014 (N_46014,N_43338,N_42972);
and U46015 (N_46015,N_44262,N_43660);
nor U46016 (N_46016,N_43726,N_44437);
nand U46017 (N_46017,N_43484,N_43167);
or U46018 (N_46018,N_44123,N_44925);
xnor U46019 (N_46019,N_42819,N_43026);
or U46020 (N_46020,N_43233,N_44932);
nor U46021 (N_46021,N_44774,N_44296);
nand U46022 (N_46022,N_42939,N_43705);
nor U46023 (N_46023,N_42891,N_44021);
or U46024 (N_46024,N_43978,N_44232);
or U46025 (N_46025,N_44244,N_43386);
xor U46026 (N_46026,N_43174,N_44215);
xnor U46027 (N_46027,N_44006,N_42715);
or U46028 (N_46028,N_44354,N_43130);
and U46029 (N_46029,N_43249,N_44637);
and U46030 (N_46030,N_42727,N_43291);
or U46031 (N_46031,N_44479,N_43027);
xnor U46032 (N_46032,N_44107,N_42539);
nor U46033 (N_46033,N_44402,N_44770);
nand U46034 (N_46034,N_42636,N_44221);
xnor U46035 (N_46035,N_42622,N_42521);
or U46036 (N_46036,N_43431,N_43546);
or U46037 (N_46037,N_42800,N_43245);
nand U46038 (N_46038,N_42722,N_44642);
or U46039 (N_46039,N_42674,N_44755);
xnor U46040 (N_46040,N_43578,N_42881);
nor U46041 (N_46041,N_44733,N_44609);
or U46042 (N_46042,N_44386,N_43412);
nand U46043 (N_46043,N_44934,N_44202);
and U46044 (N_46044,N_44902,N_42712);
or U46045 (N_46045,N_42823,N_44912);
or U46046 (N_46046,N_43203,N_43505);
nor U46047 (N_46047,N_43284,N_42614);
nand U46048 (N_46048,N_44585,N_43618);
xnor U46049 (N_46049,N_43593,N_44818);
and U46050 (N_46050,N_42602,N_43127);
and U46051 (N_46051,N_43926,N_44545);
nand U46052 (N_46052,N_43876,N_42832);
or U46053 (N_46053,N_43844,N_44514);
nor U46054 (N_46054,N_44363,N_43953);
nand U46055 (N_46055,N_42936,N_44407);
nand U46056 (N_46056,N_44163,N_43557);
or U46057 (N_46057,N_43499,N_43981);
nand U46058 (N_46058,N_44575,N_42582);
or U46059 (N_46059,N_43824,N_44310);
nand U46060 (N_46060,N_43628,N_43295);
xnor U46061 (N_46061,N_43342,N_43323);
and U46062 (N_46062,N_43425,N_44998);
nand U46063 (N_46063,N_43839,N_44941);
or U46064 (N_46064,N_43743,N_44185);
and U46065 (N_46065,N_43919,N_44529);
nand U46066 (N_46066,N_42973,N_44220);
xnor U46067 (N_46067,N_43209,N_44209);
or U46068 (N_46068,N_43672,N_42980);
nand U46069 (N_46069,N_43419,N_42530);
xnor U46070 (N_46070,N_43420,N_43712);
or U46071 (N_46071,N_42696,N_43651);
and U46072 (N_46072,N_42893,N_44952);
or U46073 (N_46073,N_43075,N_43584);
and U46074 (N_46074,N_44256,N_44340);
and U46075 (N_46075,N_43009,N_42527);
nor U46076 (N_46076,N_44567,N_42945);
or U46077 (N_46077,N_43888,N_43046);
and U46078 (N_46078,N_44523,N_43210);
or U46079 (N_46079,N_44132,N_43025);
and U46080 (N_46080,N_43228,N_43181);
and U46081 (N_46081,N_43727,N_42956);
nor U46082 (N_46082,N_43056,N_42613);
and U46083 (N_46083,N_43700,N_43232);
or U46084 (N_46084,N_43943,N_43512);
or U46085 (N_46085,N_42621,N_43746);
nand U46086 (N_46086,N_43973,N_44776);
or U46087 (N_46087,N_44192,N_43798);
and U46088 (N_46088,N_43856,N_43713);
nand U46089 (N_46089,N_44539,N_42577);
xnor U46090 (N_46090,N_44547,N_44853);
or U46091 (N_46091,N_44605,N_42927);
nand U46092 (N_46092,N_43624,N_44274);
nand U46093 (N_46093,N_43396,N_43004);
nand U46094 (N_46094,N_43942,N_42507);
or U46095 (N_46095,N_44377,N_42668);
nand U46096 (N_46096,N_44519,N_44050);
nand U46097 (N_46097,N_43491,N_44473);
xor U46098 (N_46098,N_44249,N_44408);
xnor U46099 (N_46099,N_44113,N_44806);
xnor U46100 (N_46100,N_42523,N_42519);
xnor U46101 (N_46101,N_43268,N_44065);
or U46102 (N_46102,N_43455,N_42556);
and U46103 (N_46103,N_43190,N_43089);
or U46104 (N_46104,N_43310,N_42848);
xnor U46105 (N_46105,N_42916,N_42801);
nand U46106 (N_46106,N_43818,N_43787);
xnor U46107 (N_46107,N_42669,N_43710);
and U46108 (N_46108,N_44659,N_44501);
xnor U46109 (N_46109,N_42799,N_44815);
xor U46110 (N_46110,N_42633,N_42686);
or U46111 (N_46111,N_43979,N_43495);
or U46112 (N_46112,N_42905,N_44924);
and U46113 (N_46113,N_43606,N_42680);
or U46114 (N_46114,N_44670,N_43196);
or U46115 (N_46115,N_44213,N_42682);
nand U46116 (N_46116,N_43437,N_43201);
nor U46117 (N_46117,N_42971,N_43024);
xor U46118 (N_46118,N_44536,N_43837);
xnor U46119 (N_46119,N_42584,N_43959);
nor U46120 (N_46120,N_44206,N_44465);
xnor U46121 (N_46121,N_43654,N_43530);
xnor U46122 (N_46122,N_43527,N_44636);
and U46123 (N_46123,N_43808,N_43601);
nor U46124 (N_46124,N_42986,N_43045);
xnor U46125 (N_46125,N_44242,N_44009);
and U46126 (N_46126,N_43671,N_43769);
or U46127 (N_46127,N_43413,N_42579);
nand U46128 (N_46128,N_44949,N_42946);
xnor U46129 (N_46129,N_44814,N_44159);
or U46130 (N_46130,N_44332,N_43305);
nand U46131 (N_46131,N_44960,N_43471);
nor U46132 (N_46132,N_43920,N_44682);
or U46133 (N_46133,N_42522,N_43178);
nand U46134 (N_46134,N_43246,N_44681);
nor U46135 (N_46135,N_44554,N_43912);
xnor U46136 (N_46136,N_43647,N_44168);
and U46137 (N_46137,N_43018,N_42608);
nor U46138 (N_46138,N_42560,N_43380);
xor U46139 (N_46139,N_44337,N_44207);
xnor U46140 (N_46140,N_44312,N_43903);
or U46141 (N_46141,N_43963,N_42580);
and U46142 (N_46142,N_42586,N_44478);
or U46143 (N_46143,N_43020,N_44490);
and U46144 (N_46144,N_44398,N_42802);
and U46145 (N_46145,N_44235,N_43335);
nor U46146 (N_46146,N_44450,N_44028);
and U46147 (N_46147,N_43944,N_44394);
and U46148 (N_46148,N_43064,N_44454);
nor U46149 (N_46149,N_44463,N_43489);
or U46150 (N_46150,N_42814,N_43991);
and U46151 (N_46151,N_43637,N_42957);
nor U46152 (N_46152,N_44018,N_43670);
nor U46153 (N_46153,N_44688,N_44074);
or U46154 (N_46154,N_44578,N_42896);
or U46155 (N_46155,N_44441,N_42670);
nand U46156 (N_46156,N_44987,N_42526);
or U46157 (N_46157,N_44188,N_42886);
nand U46158 (N_46158,N_44303,N_44306);
and U46159 (N_46159,N_44047,N_43260);
or U46160 (N_46160,N_43123,N_43779);
xor U46161 (N_46161,N_42678,N_43537);
nand U46162 (N_46162,N_43899,N_44813);
and U46163 (N_46163,N_43543,N_44744);
and U46164 (N_46164,N_43143,N_42985);
nand U46165 (N_46165,N_44560,N_42809);
or U46166 (N_46166,N_44333,N_43781);
and U46167 (N_46167,N_43227,N_43967);
nand U46168 (N_46168,N_42853,N_44011);
nor U46169 (N_46169,N_44653,N_43219);
nand U46170 (N_46170,N_43886,N_44612);
nand U46171 (N_46171,N_44115,N_44883);
or U46172 (N_46172,N_43656,N_44427);
nor U46173 (N_46173,N_44927,N_43772);
nand U46174 (N_46174,N_44906,N_42859);
or U46175 (N_46175,N_43008,N_42709);
and U46176 (N_46176,N_44608,N_43254);
nor U46177 (N_46177,N_43999,N_43634);
xor U46178 (N_46178,N_43239,N_43390);
xnor U46179 (N_46179,N_42532,N_44775);
and U46180 (N_46180,N_43023,N_43927);
xor U46181 (N_46181,N_44690,N_44967);
nand U46182 (N_46182,N_43466,N_43450);
and U46183 (N_46183,N_44314,N_42606);
and U46184 (N_46184,N_44401,N_43082);
nand U46185 (N_46185,N_43520,N_44588);
or U46186 (N_46186,N_44542,N_44293);
nor U46187 (N_46187,N_42695,N_43105);
and U46188 (N_46188,N_44388,N_44392);
nor U46189 (N_46189,N_44177,N_43119);
or U46190 (N_46190,N_44819,N_44789);
xor U46191 (N_46191,N_44756,N_44129);
or U46192 (N_46192,N_44487,N_44933);
xnor U46193 (N_46193,N_44315,N_43874);
or U46194 (N_46194,N_43538,N_44493);
nor U46195 (N_46195,N_44497,N_43548);
nand U46196 (N_46196,N_42615,N_43401);
nand U46197 (N_46197,N_43111,N_44702);
and U46198 (N_46198,N_43621,N_42562);
nand U46199 (N_46199,N_43799,N_44003);
or U46200 (N_46200,N_42754,N_44827);
and U46201 (N_46201,N_44860,N_44082);
or U46202 (N_46202,N_44660,N_43485);
or U46203 (N_46203,N_44105,N_43687);
nand U46204 (N_46204,N_42635,N_44816);
and U46205 (N_46205,N_43879,N_42588);
nand U46206 (N_46206,N_43931,N_44093);
nor U46207 (N_46207,N_42725,N_44606);
nor U46208 (N_46208,N_44955,N_44665);
and U46209 (N_46209,N_42726,N_43597);
or U46210 (N_46210,N_42954,N_44583);
or U46211 (N_46211,N_44528,N_44001);
xnor U46212 (N_46212,N_44457,N_43324);
and U46213 (N_46213,N_42732,N_43308);
nand U46214 (N_46214,N_44350,N_42894);
xnor U46215 (N_46215,N_44640,N_43954);
xor U46216 (N_46216,N_42942,N_44730);
or U46217 (N_46217,N_42877,N_43535);
nand U46218 (N_46218,N_44178,N_42538);
nand U46219 (N_46219,N_42787,N_44687);
or U46220 (N_46220,N_43534,N_42570);
nor U46221 (N_46221,N_44062,N_44245);
xnor U46222 (N_46222,N_42982,N_43458);
nand U46223 (N_46223,N_43696,N_44951);
and U46224 (N_46224,N_43460,N_44362);
xnor U46225 (N_46225,N_43002,N_44176);
nand U46226 (N_46226,N_43343,N_42671);
nand U46227 (N_46227,N_42977,N_43218);
or U46228 (N_46228,N_44630,N_43400);
nand U46229 (N_46229,N_42676,N_44075);
nor U46230 (N_46230,N_44917,N_44834);
nand U46231 (N_46231,N_43138,N_42782);
and U46232 (N_46232,N_44418,N_43356);
nand U46233 (N_46233,N_44451,N_43804);
xor U46234 (N_46234,N_43758,N_43464);
or U46235 (N_46235,N_44269,N_42641);
and U46236 (N_46236,N_42901,N_44051);
and U46237 (N_46237,N_44922,N_43673);
and U46238 (N_46238,N_44066,N_42594);
nor U46239 (N_46239,N_42629,N_44890);
nand U46240 (N_46240,N_43446,N_43428);
nand U46241 (N_46241,N_43423,N_42928);
or U46242 (N_46242,N_43679,N_44053);
or U46243 (N_46243,N_44023,N_44887);
nand U46244 (N_46244,N_43195,N_44669);
and U46245 (N_46245,N_43939,N_42904);
xor U46246 (N_46246,N_43703,N_42563);
xnor U46247 (N_46247,N_42774,N_44007);
and U46248 (N_46248,N_44940,N_44174);
or U46249 (N_46249,N_43054,N_43732);
or U46250 (N_46250,N_43997,N_44115);
or U46251 (N_46251,N_43543,N_44789);
or U46252 (N_46252,N_42801,N_44170);
and U46253 (N_46253,N_43887,N_44387);
nand U46254 (N_46254,N_43209,N_42975);
nand U46255 (N_46255,N_44676,N_42540);
xor U46256 (N_46256,N_43772,N_42861);
xnor U46257 (N_46257,N_44532,N_43807);
nor U46258 (N_46258,N_44568,N_43613);
or U46259 (N_46259,N_42862,N_44230);
nor U46260 (N_46260,N_44705,N_43938);
nand U46261 (N_46261,N_44155,N_44653);
nand U46262 (N_46262,N_42747,N_44814);
and U46263 (N_46263,N_43291,N_44707);
and U46264 (N_46264,N_42633,N_43012);
and U46265 (N_46265,N_44063,N_44375);
nand U46266 (N_46266,N_43778,N_43003);
or U46267 (N_46267,N_43201,N_44227);
or U46268 (N_46268,N_44351,N_43436);
nand U46269 (N_46269,N_43834,N_44471);
and U46270 (N_46270,N_43980,N_43979);
nand U46271 (N_46271,N_44996,N_44469);
xnor U46272 (N_46272,N_44507,N_43847);
xor U46273 (N_46273,N_44484,N_43068);
and U46274 (N_46274,N_42972,N_43329);
and U46275 (N_46275,N_43663,N_44217);
or U46276 (N_46276,N_43053,N_44584);
and U46277 (N_46277,N_43308,N_44027);
and U46278 (N_46278,N_44652,N_44866);
and U46279 (N_46279,N_44526,N_43881);
and U46280 (N_46280,N_42687,N_42660);
and U46281 (N_46281,N_44463,N_43866);
nand U46282 (N_46282,N_44548,N_44690);
and U46283 (N_46283,N_42530,N_42561);
xnor U46284 (N_46284,N_43099,N_44568);
or U46285 (N_46285,N_44511,N_43605);
and U46286 (N_46286,N_44686,N_44169);
and U46287 (N_46287,N_44042,N_42840);
or U46288 (N_46288,N_44212,N_44187);
nor U46289 (N_46289,N_44436,N_42953);
nand U46290 (N_46290,N_43790,N_44865);
or U46291 (N_46291,N_44030,N_44183);
nand U46292 (N_46292,N_44693,N_44116);
or U46293 (N_46293,N_42810,N_42990);
nand U46294 (N_46294,N_43873,N_43341);
nor U46295 (N_46295,N_42886,N_43816);
or U46296 (N_46296,N_43223,N_43781);
and U46297 (N_46297,N_44680,N_44085);
xnor U46298 (N_46298,N_43063,N_43700);
or U46299 (N_46299,N_44537,N_44263);
nand U46300 (N_46300,N_44031,N_44823);
and U46301 (N_46301,N_43838,N_44218);
nor U46302 (N_46302,N_42904,N_43430);
nor U46303 (N_46303,N_44500,N_44248);
or U46304 (N_46304,N_43896,N_44639);
nor U46305 (N_46305,N_42566,N_44659);
xor U46306 (N_46306,N_44696,N_44225);
and U46307 (N_46307,N_43632,N_42930);
nand U46308 (N_46308,N_42901,N_42533);
or U46309 (N_46309,N_43669,N_44495);
or U46310 (N_46310,N_43407,N_42503);
xnor U46311 (N_46311,N_44621,N_43390);
or U46312 (N_46312,N_43814,N_42743);
nor U46313 (N_46313,N_43294,N_44715);
or U46314 (N_46314,N_43095,N_43484);
and U46315 (N_46315,N_44984,N_42531);
or U46316 (N_46316,N_44706,N_42874);
and U46317 (N_46317,N_44445,N_43181);
nor U46318 (N_46318,N_44518,N_42876);
nor U46319 (N_46319,N_42917,N_43544);
and U46320 (N_46320,N_42959,N_44645);
and U46321 (N_46321,N_43333,N_44137);
nor U46322 (N_46322,N_44528,N_42989);
xnor U46323 (N_46323,N_42954,N_43967);
or U46324 (N_46324,N_43141,N_43004);
or U46325 (N_46325,N_44655,N_44728);
or U46326 (N_46326,N_43284,N_42818);
or U46327 (N_46327,N_42665,N_44949);
or U46328 (N_46328,N_43426,N_42534);
or U46329 (N_46329,N_43956,N_43793);
xnor U46330 (N_46330,N_44852,N_43481);
nand U46331 (N_46331,N_43330,N_44384);
xnor U46332 (N_46332,N_44381,N_42951);
xor U46333 (N_46333,N_44327,N_42998);
or U46334 (N_46334,N_42759,N_44957);
nor U46335 (N_46335,N_43955,N_43299);
nand U46336 (N_46336,N_43902,N_44331);
or U46337 (N_46337,N_44635,N_42760);
and U46338 (N_46338,N_44509,N_43321);
nand U46339 (N_46339,N_44009,N_43748);
nand U46340 (N_46340,N_42966,N_44828);
and U46341 (N_46341,N_44838,N_43912);
nor U46342 (N_46342,N_42501,N_43636);
or U46343 (N_46343,N_43606,N_44511);
or U46344 (N_46344,N_44771,N_44417);
nor U46345 (N_46345,N_43995,N_44986);
nor U46346 (N_46346,N_43095,N_43279);
or U46347 (N_46347,N_43984,N_42578);
or U46348 (N_46348,N_44501,N_44318);
nand U46349 (N_46349,N_44189,N_42932);
nand U46350 (N_46350,N_42728,N_44159);
nand U46351 (N_46351,N_42772,N_43849);
and U46352 (N_46352,N_43920,N_42649);
nand U46353 (N_46353,N_43717,N_42820);
and U46354 (N_46354,N_44074,N_43229);
nand U46355 (N_46355,N_42603,N_43085);
xor U46356 (N_46356,N_43300,N_44906);
nand U46357 (N_46357,N_43190,N_42937);
nor U46358 (N_46358,N_44343,N_43304);
nor U46359 (N_46359,N_44422,N_43282);
nor U46360 (N_46360,N_42638,N_42726);
nor U46361 (N_46361,N_44382,N_43661);
nor U46362 (N_46362,N_43150,N_42730);
or U46363 (N_46363,N_43776,N_43057);
nor U46364 (N_46364,N_44226,N_44631);
xor U46365 (N_46365,N_44379,N_44214);
nand U46366 (N_46366,N_44899,N_44503);
or U46367 (N_46367,N_44343,N_44565);
or U46368 (N_46368,N_44260,N_44951);
or U46369 (N_46369,N_43871,N_44330);
nand U46370 (N_46370,N_44864,N_44306);
or U46371 (N_46371,N_43154,N_44834);
or U46372 (N_46372,N_43514,N_42975);
xnor U46373 (N_46373,N_43695,N_42500);
nor U46374 (N_46374,N_43599,N_44774);
nor U46375 (N_46375,N_42942,N_42632);
nor U46376 (N_46376,N_44599,N_44738);
nand U46377 (N_46377,N_43223,N_44529);
and U46378 (N_46378,N_43113,N_44847);
nand U46379 (N_46379,N_44460,N_44642);
or U46380 (N_46380,N_43109,N_42655);
and U46381 (N_46381,N_44755,N_44141);
nand U46382 (N_46382,N_42857,N_43209);
xor U46383 (N_46383,N_42574,N_43526);
or U46384 (N_46384,N_43062,N_42685);
nor U46385 (N_46385,N_44545,N_44267);
and U46386 (N_46386,N_43634,N_42869);
and U46387 (N_46387,N_44086,N_42732);
and U46388 (N_46388,N_44769,N_44838);
and U46389 (N_46389,N_43422,N_44968);
or U46390 (N_46390,N_43227,N_43097);
or U46391 (N_46391,N_44400,N_43681);
xnor U46392 (N_46392,N_43391,N_44741);
or U46393 (N_46393,N_44282,N_43752);
and U46394 (N_46394,N_44646,N_43349);
nand U46395 (N_46395,N_42815,N_43627);
nor U46396 (N_46396,N_43637,N_43827);
or U46397 (N_46397,N_44489,N_43238);
nand U46398 (N_46398,N_44236,N_43586);
xnor U46399 (N_46399,N_43042,N_44236);
and U46400 (N_46400,N_42501,N_44790);
nor U46401 (N_46401,N_43212,N_43798);
or U46402 (N_46402,N_42936,N_44342);
and U46403 (N_46403,N_44600,N_44774);
and U46404 (N_46404,N_43936,N_44018);
or U46405 (N_46405,N_43828,N_44649);
or U46406 (N_46406,N_42577,N_42976);
nor U46407 (N_46407,N_43813,N_44464);
and U46408 (N_46408,N_42677,N_42886);
or U46409 (N_46409,N_42558,N_43939);
nor U46410 (N_46410,N_43472,N_43746);
nor U46411 (N_46411,N_43798,N_44011);
nand U46412 (N_46412,N_44990,N_43520);
and U46413 (N_46413,N_43951,N_43403);
nand U46414 (N_46414,N_44277,N_44829);
nor U46415 (N_46415,N_44256,N_44891);
nand U46416 (N_46416,N_44798,N_43734);
nand U46417 (N_46417,N_44076,N_42516);
nand U46418 (N_46418,N_43770,N_43147);
nor U46419 (N_46419,N_44659,N_44918);
and U46420 (N_46420,N_44530,N_42983);
or U46421 (N_46421,N_44323,N_44783);
xnor U46422 (N_46422,N_44126,N_44823);
and U46423 (N_46423,N_44316,N_44654);
xor U46424 (N_46424,N_44777,N_42635);
xor U46425 (N_46425,N_43280,N_44752);
or U46426 (N_46426,N_42868,N_42747);
xnor U46427 (N_46427,N_43578,N_44083);
nor U46428 (N_46428,N_43414,N_44944);
xnor U46429 (N_46429,N_43705,N_44890);
and U46430 (N_46430,N_44228,N_44234);
nor U46431 (N_46431,N_42955,N_44881);
xor U46432 (N_46432,N_43120,N_44273);
nor U46433 (N_46433,N_43561,N_42609);
nand U46434 (N_46434,N_43979,N_43744);
and U46435 (N_46435,N_43557,N_43775);
xnor U46436 (N_46436,N_43099,N_43084);
or U46437 (N_46437,N_43529,N_43826);
nand U46438 (N_46438,N_43814,N_43722);
and U46439 (N_46439,N_42638,N_44894);
and U46440 (N_46440,N_43940,N_42750);
nand U46441 (N_46441,N_43172,N_42644);
nor U46442 (N_46442,N_43697,N_44741);
nand U46443 (N_46443,N_44732,N_44751);
nor U46444 (N_46444,N_42570,N_44095);
xnor U46445 (N_46445,N_43171,N_44532);
nand U46446 (N_46446,N_44847,N_44403);
xnor U46447 (N_46447,N_43502,N_44087);
or U46448 (N_46448,N_44909,N_44063);
nor U46449 (N_46449,N_44741,N_43124);
nand U46450 (N_46450,N_43692,N_44911);
xnor U46451 (N_46451,N_44872,N_43856);
or U46452 (N_46452,N_44646,N_42829);
nor U46453 (N_46453,N_44917,N_43561);
xor U46454 (N_46454,N_44503,N_43516);
nor U46455 (N_46455,N_43510,N_44265);
xor U46456 (N_46456,N_44960,N_43457);
or U46457 (N_46457,N_42835,N_43238);
and U46458 (N_46458,N_43188,N_42737);
xor U46459 (N_46459,N_44852,N_42756);
nor U46460 (N_46460,N_43306,N_44275);
and U46461 (N_46461,N_44906,N_43917);
or U46462 (N_46462,N_44526,N_43366);
nor U46463 (N_46463,N_42620,N_43132);
or U46464 (N_46464,N_44988,N_44312);
nor U46465 (N_46465,N_43775,N_44435);
nor U46466 (N_46466,N_42819,N_42909);
and U46467 (N_46467,N_44040,N_43038);
or U46468 (N_46468,N_43834,N_43620);
xnor U46469 (N_46469,N_42909,N_44272);
and U46470 (N_46470,N_43469,N_43821);
nor U46471 (N_46471,N_44716,N_43269);
nor U46472 (N_46472,N_42831,N_44353);
nand U46473 (N_46473,N_44505,N_43204);
nand U46474 (N_46474,N_44757,N_43696);
xnor U46475 (N_46475,N_44701,N_43015);
xor U46476 (N_46476,N_43948,N_44796);
and U46477 (N_46477,N_43843,N_43966);
xnor U46478 (N_46478,N_43592,N_44297);
or U46479 (N_46479,N_43065,N_43381);
nand U46480 (N_46480,N_43317,N_42680);
nand U46481 (N_46481,N_44799,N_44583);
or U46482 (N_46482,N_44203,N_44836);
and U46483 (N_46483,N_44502,N_44148);
or U46484 (N_46484,N_43145,N_44556);
xor U46485 (N_46485,N_43037,N_42627);
nor U46486 (N_46486,N_43383,N_44033);
xnor U46487 (N_46487,N_44588,N_43857);
nor U46488 (N_46488,N_42599,N_43709);
xor U46489 (N_46489,N_43830,N_42766);
xnor U46490 (N_46490,N_44923,N_43493);
nor U46491 (N_46491,N_43246,N_42985);
nor U46492 (N_46492,N_42795,N_44088);
nor U46493 (N_46493,N_43078,N_44408);
nand U46494 (N_46494,N_43921,N_42634);
and U46495 (N_46495,N_44826,N_44646);
or U46496 (N_46496,N_43573,N_44844);
and U46497 (N_46497,N_44906,N_43834);
and U46498 (N_46498,N_44213,N_43623);
nor U46499 (N_46499,N_43053,N_44872);
xor U46500 (N_46500,N_42692,N_44148);
nor U46501 (N_46501,N_44487,N_44535);
nor U46502 (N_46502,N_44591,N_43033);
xnor U46503 (N_46503,N_43453,N_44207);
and U46504 (N_46504,N_42696,N_43991);
and U46505 (N_46505,N_43235,N_43225);
or U46506 (N_46506,N_44501,N_44200);
xnor U46507 (N_46507,N_43153,N_44879);
and U46508 (N_46508,N_42822,N_43544);
and U46509 (N_46509,N_43763,N_44939);
nand U46510 (N_46510,N_43402,N_43331);
or U46511 (N_46511,N_44271,N_44978);
nor U46512 (N_46512,N_43627,N_43179);
nor U46513 (N_46513,N_44377,N_43142);
or U46514 (N_46514,N_43164,N_42991);
nor U46515 (N_46515,N_43488,N_44288);
nor U46516 (N_46516,N_42627,N_44569);
or U46517 (N_46517,N_43779,N_44582);
nand U46518 (N_46518,N_43850,N_43192);
nand U46519 (N_46519,N_42538,N_43714);
and U46520 (N_46520,N_44898,N_44185);
nor U46521 (N_46521,N_44843,N_44368);
nand U46522 (N_46522,N_44636,N_44183);
nor U46523 (N_46523,N_44710,N_42738);
and U46524 (N_46524,N_44298,N_42533);
or U46525 (N_46525,N_42791,N_44246);
and U46526 (N_46526,N_44438,N_43784);
nor U46527 (N_46527,N_43053,N_43456);
xnor U46528 (N_46528,N_43331,N_44690);
nand U46529 (N_46529,N_44730,N_43655);
nor U46530 (N_46530,N_43855,N_44478);
and U46531 (N_46531,N_44221,N_43602);
or U46532 (N_46532,N_43047,N_43638);
nand U46533 (N_46533,N_44253,N_44440);
xor U46534 (N_46534,N_43305,N_44488);
nor U46535 (N_46535,N_42612,N_44001);
nand U46536 (N_46536,N_44267,N_44676);
and U46537 (N_46537,N_43697,N_42763);
or U46538 (N_46538,N_43043,N_44075);
xor U46539 (N_46539,N_43112,N_43767);
and U46540 (N_46540,N_42888,N_43906);
or U46541 (N_46541,N_43291,N_43412);
xor U46542 (N_46542,N_43181,N_44343);
or U46543 (N_46543,N_42944,N_44987);
and U46544 (N_46544,N_43132,N_43642);
xor U46545 (N_46545,N_42838,N_44897);
and U46546 (N_46546,N_44616,N_44803);
xor U46547 (N_46547,N_44423,N_44657);
xnor U46548 (N_46548,N_44441,N_42695);
xor U46549 (N_46549,N_43471,N_44267);
nor U46550 (N_46550,N_42549,N_44811);
nand U46551 (N_46551,N_42728,N_42786);
nand U46552 (N_46552,N_44849,N_44746);
and U46553 (N_46553,N_43190,N_44218);
nand U46554 (N_46554,N_44500,N_44950);
xnor U46555 (N_46555,N_44172,N_42908);
and U46556 (N_46556,N_43755,N_43561);
nand U46557 (N_46557,N_43194,N_43012);
or U46558 (N_46558,N_44303,N_42775);
nor U46559 (N_46559,N_43192,N_43799);
nor U46560 (N_46560,N_44598,N_43463);
nor U46561 (N_46561,N_44129,N_42944);
and U46562 (N_46562,N_42536,N_43571);
nor U46563 (N_46563,N_42721,N_43466);
and U46564 (N_46564,N_43126,N_44624);
xnor U46565 (N_46565,N_42742,N_44229);
or U46566 (N_46566,N_43615,N_44373);
nand U46567 (N_46567,N_43199,N_43511);
and U46568 (N_46568,N_42953,N_44005);
or U46569 (N_46569,N_42617,N_44166);
nor U46570 (N_46570,N_44029,N_43380);
nor U46571 (N_46571,N_43551,N_43831);
nor U46572 (N_46572,N_44060,N_44320);
nor U46573 (N_46573,N_44273,N_43696);
or U46574 (N_46574,N_43568,N_43474);
or U46575 (N_46575,N_44511,N_43947);
or U46576 (N_46576,N_43959,N_44864);
and U46577 (N_46577,N_42959,N_42566);
nor U46578 (N_46578,N_44203,N_44131);
nor U46579 (N_46579,N_44340,N_44130);
nand U46580 (N_46580,N_43657,N_44320);
and U46581 (N_46581,N_43456,N_43617);
nand U46582 (N_46582,N_42788,N_44591);
or U46583 (N_46583,N_43063,N_43391);
or U46584 (N_46584,N_43765,N_43062);
and U46585 (N_46585,N_43604,N_43035);
xor U46586 (N_46586,N_43691,N_43700);
nor U46587 (N_46587,N_43937,N_42877);
nor U46588 (N_46588,N_42599,N_44629);
and U46589 (N_46589,N_44210,N_43981);
nor U46590 (N_46590,N_42874,N_42597);
nand U46591 (N_46591,N_42934,N_43696);
nand U46592 (N_46592,N_44853,N_44724);
nor U46593 (N_46593,N_42680,N_44830);
nand U46594 (N_46594,N_43178,N_44213);
or U46595 (N_46595,N_43846,N_44990);
nand U46596 (N_46596,N_42981,N_43221);
xor U46597 (N_46597,N_43473,N_42889);
or U46598 (N_46598,N_44810,N_44228);
nand U46599 (N_46599,N_43418,N_44763);
nand U46600 (N_46600,N_43775,N_42618);
or U46601 (N_46601,N_44562,N_44309);
nor U46602 (N_46602,N_44685,N_42884);
or U46603 (N_46603,N_44845,N_43116);
nand U46604 (N_46604,N_43645,N_43250);
or U46605 (N_46605,N_44686,N_42924);
xor U46606 (N_46606,N_43943,N_43665);
nor U46607 (N_46607,N_43091,N_43241);
xor U46608 (N_46608,N_43696,N_42592);
and U46609 (N_46609,N_44698,N_42625);
or U46610 (N_46610,N_43462,N_44073);
nor U46611 (N_46611,N_44412,N_44902);
or U46612 (N_46612,N_44269,N_43399);
nor U46613 (N_46613,N_42616,N_43521);
xor U46614 (N_46614,N_44688,N_44166);
nor U46615 (N_46615,N_44396,N_44981);
nor U46616 (N_46616,N_44114,N_43368);
nand U46617 (N_46617,N_44650,N_43395);
or U46618 (N_46618,N_42692,N_42914);
xor U46619 (N_46619,N_43878,N_43121);
or U46620 (N_46620,N_44617,N_43205);
xor U46621 (N_46621,N_43351,N_43500);
and U46622 (N_46622,N_44780,N_43349);
xnor U46623 (N_46623,N_43966,N_44761);
nor U46624 (N_46624,N_43406,N_44587);
or U46625 (N_46625,N_44122,N_44058);
xnor U46626 (N_46626,N_43217,N_43378);
nand U46627 (N_46627,N_43902,N_44350);
nor U46628 (N_46628,N_43061,N_43330);
nand U46629 (N_46629,N_44886,N_43439);
and U46630 (N_46630,N_43767,N_43244);
or U46631 (N_46631,N_44350,N_44284);
or U46632 (N_46632,N_43840,N_44539);
or U46633 (N_46633,N_43800,N_43053);
or U46634 (N_46634,N_44380,N_44334);
nand U46635 (N_46635,N_43239,N_44683);
xor U46636 (N_46636,N_43719,N_43977);
xnor U46637 (N_46637,N_43873,N_44572);
or U46638 (N_46638,N_43466,N_44612);
nor U46639 (N_46639,N_44683,N_42682);
xor U46640 (N_46640,N_42927,N_43938);
nor U46641 (N_46641,N_44038,N_44783);
nand U46642 (N_46642,N_43501,N_44200);
xnor U46643 (N_46643,N_43302,N_44938);
or U46644 (N_46644,N_44676,N_44055);
xor U46645 (N_46645,N_42691,N_43849);
xnor U46646 (N_46646,N_44090,N_42570);
or U46647 (N_46647,N_43224,N_43128);
nand U46648 (N_46648,N_42913,N_43770);
nor U46649 (N_46649,N_44559,N_44426);
or U46650 (N_46650,N_43965,N_44377);
and U46651 (N_46651,N_42649,N_42946);
or U46652 (N_46652,N_42843,N_43859);
nand U46653 (N_46653,N_43938,N_42998);
nor U46654 (N_46654,N_43894,N_44349);
and U46655 (N_46655,N_43044,N_44180);
or U46656 (N_46656,N_43206,N_44451);
nor U46657 (N_46657,N_43878,N_44082);
xor U46658 (N_46658,N_43309,N_43026);
nor U46659 (N_46659,N_43086,N_44843);
nand U46660 (N_46660,N_44111,N_44671);
nor U46661 (N_46661,N_42976,N_43097);
or U46662 (N_46662,N_42973,N_43690);
nand U46663 (N_46663,N_44316,N_43172);
nand U46664 (N_46664,N_42691,N_43919);
or U46665 (N_46665,N_43568,N_42732);
and U46666 (N_46666,N_43028,N_43230);
or U46667 (N_46667,N_44496,N_44298);
or U46668 (N_46668,N_44756,N_44493);
nand U46669 (N_46669,N_44531,N_44440);
xor U46670 (N_46670,N_44704,N_44371);
and U46671 (N_46671,N_44198,N_43491);
nor U46672 (N_46672,N_44177,N_44838);
nor U46673 (N_46673,N_44644,N_42949);
nand U46674 (N_46674,N_42596,N_44955);
nand U46675 (N_46675,N_43519,N_44568);
and U46676 (N_46676,N_42909,N_42559);
or U46677 (N_46677,N_44138,N_43855);
or U46678 (N_46678,N_42733,N_44652);
and U46679 (N_46679,N_43382,N_44268);
xnor U46680 (N_46680,N_44610,N_43414);
xor U46681 (N_46681,N_42932,N_44786);
nand U46682 (N_46682,N_44909,N_42803);
xnor U46683 (N_46683,N_43872,N_42787);
or U46684 (N_46684,N_43565,N_43521);
nand U46685 (N_46685,N_43656,N_43902);
or U46686 (N_46686,N_43604,N_43121);
nor U46687 (N_46687,N_43481,N_43958);
nand U46688 (N_46688,N_42505,N_44013);
nor U46689 (N_46689,N_43804,N_44201);
and U46690 (N_46690,N_42583,N_44781);
nor U46691 (N_46691,N_44287,N_43979);
nor U46692 (N_46692,N_42669,N_44437);
xnor U46693 (N_46693,N_44310,N_43176);
xor U46694 (N_46694,N_44268,N_44732);
nand U46695 (N_46695,N_44533,N_43856);
or U46696 (N_46696,N_44910,N_42742);
nor U46697 (N_46697,N_42956,N_42796);
nand U46698 (N_46698,N_43982,N_43858);
nor U46699 (N_46699,N_43161,N_44683);
and U46700 (N_46700,N_44407,N_44795);
nand U46701 (N_46701,N_44292,N_43683);
xnor U46702 (N_46702,N_43979,N_44307);
and U46703 (N_46703,N_42922,N_42911);
nor U46704 (N_46704,N_43119,N_43029);
xnor U46705 (N_46705,N_42876,N_43492);
or U46706 (N_46706,N_44604,N_44335);
or U46707 (N_46707,N_44675,N_44169);
nand U46708 (N_46708,N_44053,N_44842);
nand U46709 (N_46709,N_44570,N_43388);
xnor U46710 (N_46710,N_44665,N_43634);
or U46711 (N_46711,N_43666,N_44418);
nand U46712 (N_46712,N_42525,N_43177);
xnor U46713 (N_46713,N_44942,N_44864);
and U46714 (N_46714,N_43292,N_42567);
nor U46715 (N_46715,N_42978,N_43812);
and U46716 (N_46716,N_43876,N_43665);
and U46717 (N_46717,N_43942,N_43921);
nor U46718 (N_46718,N_43705,N_42723);
and U46719 (N_46719,N_44035,N_43290);
nand U46720 (N_46720,N_44551,N_44196);
or U46721 (N_46721,N_43156,N_43123);
nor U46722 (N_46722,N_44616,N_43153);
or U46723 (N_46723,N_42713,N_44646);
nand U46724 (N_46724,N_43575,N_42676);
or U46725 (N_46725,N_43993,N_42857);
nand U46726 (N_46726,N_43364,N_43687);
xor U46727 (N_46727,N_43060,N_44960);
or U46728 (N_46728,N_43892,N_42613);
xor U46729 (N_46729,N_43316,N_44755);
nand U46730 (N_46730,N_44325,N_44986);
nor U46731 (N_46731,N_43785,N_43388);
xnor U46732 (N_46732,N_42872,N_42752);
or U46733 (N_46733,N_43353,N_42847);
nor U46734 (N_46734,N_44204,N_44176);
and U46735 (N_46735,N_43993,N_43525);
nor U46736 (N_46736,N_42729,N_43491);
or U46737 (N_46737,N_43348,N_44361);
nor U46738 (N_46738,N_44892,N_42819);
and U46739 (N_46739,N_44793,N_44145);
nand U46740 (N_46740,N_44842,N_43560);
nand U46741 (N_46741,N_44877,N_44876);
nor U46742 (N_46742,N_44531,N_44039);
or U46743 (N_46743,N_42556,N_44321);
nor U46744 (N_46744,N_43768,N_42612);
nand U46745 (N_46745,N_43686,N_44875);
xnor U46746 (N_46746,N_43707,N_42854);
or U46747 (N_46747,N_44817,N_42813);
nand U46748 (N_46748,N_43318,N_43626);
nor U46749 (N_46749,N_44308,N_43553);
and U46750 (N_46750,N_44039,N_44212);
nor U46751 (N_46751,N_43927,N_43412);
nor U46752 (N_46752,N_43351,N_43221);
nand U46753 (N_46753,N_44967,N_44466);
xor U46754 (N_46754,N_43513,N_43844);
xnor U46755 (N_46755,N_44401,N_42938);
nand U46756 (N_46756,N_43439,N_44421);
nand U46757 (N_46757,N_43715,N_42817);
nand U46758 (N_46758,N_44587,N_43215);
xnor U46759 (N_46759,N_43437,N_42695);
nor U46760 (N_46760,N_43402,N_43240);
xor U46761 (N_46761,N_44606,N_43375);
nor U46762 (N_46762,N_44979,N_43694);
or U46763 (N_46763,N_44372,N_44933);
and U46764 (N_46764,N_44645,N_44839);
and U46765 (N_46765,N_44965,N_42733);
or U46766 (N_46766,N_44192,N_42510);
nor U46767 (N_46767,N_43336,N_44934);
nor U46768 (N_46768,N_44484,N_44327);
xor U46769 (N_46769,N_44616,N_43302);
nand U46770 (N_46770,N_44961,N_43413);
nor U46771 (N_46771,N_42771,N_43357);
nor U46772 (N_46772,N_44446,N_43249);
or U46773 (N_46773,N_44561,N_44565);
xnor U46774 (N_46774,N_42968,N_42871);
and U46775 (N_46775,N_43500,N_43225);
xnor U46776 (N_46776,N_44152,N_43582);
nand U46777 (N_46777,N_42642,N_43579);
xnor U46778 (N_46778,N_42540,N_44120);
and U46779 (N_46779,N_44499,N_44400);
nand U46780 (N_46780,N_44992,N_44395);
or U46781 (N_46781,N_44340,N_44966);
nand U46782 (N_46782,N_44412,N_44278);
nor U46783 (N_46783,N_44704,N_44664);
nor U46784 (N_46784,N_43721,N_43248);
xnor U46785 (N_46785,N_44260,N_44877);
nand U46786 (N_46786,N_43997,N_44341);
or U46787 (N_46787,N_44900,N_42947);
and U46788 (N_46788,N_44339,N_43368);
xnor U46789 (N_46789,N_44424,N_44477);
nand U46790 (N_46790,N_44432,N_44945);
xor U46791 (N_46791,N_44224,N_43977);
xor U46792 (N_46792,N_44935,N_44305);
xnor U46793 (N_46793,N_44285,N_42914);
xor U46794 (N_46794,N_43181,N_43880);
xor U46795 (N_46795,N_43284,N_44837);
xor U46796 (N_46796,N_44427,N_43854);
or U46797 (N_46797,N_43669,N_43968);
nor U46798 (N_46798,N_44812,N_44620);
nand U46799 (N_46799,N_44610,N_44597);
xor U46800 (N_46800,N_43449,N_43890);
and U46801 (N_46801,N_44054,N_43043);
and U46802 (N_46802,N_43261,N_44114);
nand U46803 (N_46803,N_42580,N_44704);
xor U46804 (N_46804,N_44094,N_43041);
or U46805 (N_46805,N_42842,N_43258);
nand U46806 (N_46806,N_44262,N_44952);
and U46807 (N_46807,N_44874,N_43790);
nor U46808 (N_46808,N_42970,N_44757);
nand U46809 (N_46809,N_42820,N_43097);
nor U46810 (N_46810,N_43292,N_43965);
nor U46811 (N_46811,N_44460,N_43881);
nor U46812 (N_46812,N_44503,N_44977);
nor U46813 (N_46813,N_44166,N_44771);
nand U46814 (N_46814,N_42691,N_43041);
xor U46815 (N_46815,N_44849,N_42867);
and U46816 (N_46816,N_43065,N_42625);
and U46817 (N_46817,N_42557,N_42918);
or U46818 (N_46818,N_43187,N_43227);
nand U46819 (N_46819,N_43495,N_44620);
or U46820 (N_46820,N_43269,N_44259);
and U46821 (N_46821,N_44817,N_44806);
nand U46822 (N_46822,N_44629,N_43627);
nand U46823 (N_46823,N_44405,N_43237);
nor U46824 (N_46824,N_43960,N_43551);
and U46825 (N_46825,N_42968,N_44988);
or U46826 (N_46826,N_43384,N_43996);
nand U46827 (N_46827,N_42968,N_43818);
or U46828 (N_46828,N_42529,N_44484);
or U46829 (N_46829,N_44411,N_43910);
or U46830 (N_46830,N_44221,N_42755);
and U46831 (N_46831,N_44253,N_44946);
xnor U46832 (N_46832,N_43463,N_43932);
nand U46833 (N_46833,N_44528,N_43878);
xor U46834 (N_46834,N_44732,N_44801);
or U46835 (N_46835,N_44144,N_44380);
or U46836 (N_46836,N_44936,N_42550);
or U46837 (N_46837,N_44044,N_42549);
xor U46838 (N_46838,N_44911,N_44029);
nor U46839 (N_46839,N_42588,N_43590);
or U46840 (N_46840,N_44810,N_44571);
and U46841 (N_46841,N_42762,N_44714);
nand U46842 (N_46842,N_43251,N_42829);
nor U46843 (N_46843,N_42730,N_43483);
or U46844 (N_46844,N_44359,N_42985);
nand U46845 (N_46845,N_44484,N_43091);
and U46846 (N_46846,N_43958,N_43581);
xnor U46847 (N_46847,N_42695,N_44042);
xor U46848 (N_46848,N_43170,N_43982);
nor U46849 (N_46849,N_44519,N_44696);
xnor U46850 (N_46850,N_43626,N_43185);
nand U46851 (N_46851,N_43633,N_44602);
xor U46852 (N_46852,N_43090,N_43285);
and U46853 (N_46853,N_42974,N_44247);
nor U46854 (N_46854,N_43124,N_43376);
or U46855 (N_46855,N_42641,N_44126);
or U46856 (N_46856,N_44836,N_43239);
and U46857 (N_46857,N_44294,N_42719);
nand U46858 (N_46858,N_43298,N_43000);
xor U46859 (N_46859,N_42970,N_43024);
and U46860 (N_46860,N_43630,N_44142);
nor U46861 (N_46861,N_44509,N_43419);
and U46862 (N_46862,N_44713,N_44144);
nor U46863 (N_46863,N_42543,N_43205);
and U46864 (N_46864,N_44572,N_44031);
or U46865 (N_46865,N_44667,N_42914);
nor U46866 (N_46866,N_42717,N_44800);
nand U46867 (N_46867,N_44905,N_44704);
nand U46868 (N_46868,N_44624,N_44117);
nor U46869 (N_46869,N_42986,N_44961);
or U46870 (N_46870,N_43544,N_43208);
nor U46871 (N_46871,N_44467,N_43250);
nand U46872 (N_46872,N_42943,N_43018);
or U46873 (N_46873,N_43415,N_44777);
nand U46874 (N_46874,N_44198,N_44781);
nand U46875 (N_46875,N_42693,N_43424);
xnor U46876 (N_46876,N_43693,N_43526);
xor U46877 (N_46877,N_43059,N_43226);
and U46878 (N_46878,N_43880,N_43037);
nor U46879 (N_46879,N_43554,N_42767);
and U46880 (N_46880,N_44315,N_43160);
and U46881 (N_46881,N_44841,N_43851);
or U46882 (N_46882,N_44163,N_43387);
nand U46883 (N_46883,N_43842,N_43782);
nor U46884 (N_46884,N_44049,N_43140);
or U46885 (N_46885,N_43024,N_42903);
or U46886 (N_46886,N_42797,N_43742);
or U46887 (N_46887,N_43762,N_44908);
and U46888 (N_46888,N_44887,N_44501);
or U46889 (N_46889,N_42580,N_42612);
and U46890 (N_46890,N_43589,N_44375);
nor U46891 (N_46891,N_43354,N_43382);
nand U46892 (N_46892,N_44498,N_43242);
xor U46893 (N_46893,N_43116,N_44013);
nor U46894 (N_46894,N_44872,N_42768);
nand U46895 (N_46895,N_44252,N_44497);
or U46896 (N_46896,N_43035,N_43570);
nor U46897 (N_46897,N_43913,N_44602);
nand U46898 (N_46898,N_44106,N_43516);
and U46899 (N_46899,N_44298,N_42708);
nand U46900 (N_46900,N_43724,N_44729);
and U46901 (N_46901,N_44467,N_44361);
or U46902 (N_46902,N_43856,N_43262);
or U46903 (N_46903,N_42937,N_43812);
nor U46904 (N_46904,N_42667,N_43799);
nor U46905 (N_46905,N_43962,N_42786);
nand U46906 (N_46906,N_44735,N_42907);
or U46907 (N_46907,N_42585,N_43179);
xnor U46908 (N_46908,N_42841,N_44245);
and U46909 (N_46909,N_42602,N_43228);
nand U46910 (N_46910,N_44091,N_44478);
nand U46911 (N_46911,N_44877,N_44032);
or U46912 (N_46912,N_43558,N_43094);
or U46913 (N_46913,N_43130,N_43889);
xor U46914 (N_46914,N_42506,N_42961);
nor U46915 (N_46915,N_43104,N_44919);
nand U46916 (N_46916,N_42723,N_44384);
xnor U46917 (N_46917,N_43814,N_43877);
or U46918 (N_46918,N_43604,N_43957);
and U46919 (N_46919,N_44607,N_44902);
and U46920 (N_46920,N_43803,N_43502);
nor U46921 (N_46921,N_44371,N_44630);
nand U46922 (N_46922,N_43973,N_44305);
nand U46923 (N_46923,N_44590,N_43936);
xor U46924 (N_46924,N_44245,N_43624);
or U46925 (N_46925,N_43969,N_43872);
nor U46926 (N_46926,N_44591,N_44784);
nor U46927 (N_46927,N_44403,N_43253);
nor U46928 (N_46928,N_42873,N_42564);
nor U46929 (N_46929,N_44100,N_43259);
nor U46930 (N_46930,N_44033,N_44508);
xnor U46931 (N_46931,N_44931,N_43210);
xnor U46932 (N_46932,N_43660,N_43954);
nand U46933 (N_46933,N_44185,N_43848);
xor U46934 (N_46934,N_44057,N_44263);
nand U46935 (N_46935,N_43095,N_42746);
or U46936 (N_46936,N_43649,N_44909);
and U46937 (N_46937,N_44884,N_44002);
or U46938 (N_46938,N_44757,N_43907);
xnor U46939 (N_46939,N_44621,N_44265);
nand U46940 (N_46940,N_43921,N_44475);
xnor U46941 (N_46941,N_44546,N_44029);
or U46942 (N_46942,N_44977,N_44020);
xnor U46943 (N_46943,N_42510,N_44878);
or U46944 (N_46944,N_43431,N_43446);
xor U46945 (N_46945,N_43327,N_44986);
nor U46946 (N_46946,N_44760,N_44707);
and U46947 (N_46947,N_43010,N_42538);
or U46948 (N_46948,N_44290,N_43814);
or U46949 (N_46949,N_43709,N_44225);
xnor U46950 (N_46950,N_43834,N_44736);
nand U46951 (N_46951,N_43259,N_43306);
xnor U46952 (N_46952,N_44817,N_42996);
or U46953 (N_46953,N_44719,N_44548);
or U46954 (N_46954,N_43531,N_42827);
nor U46955 (N_46955,N_44530,N_44757);
nand U46956 (N_46956,N_44276,N_42861);
nor U46957 (N_46957,N_44255,N_44454);
nand U46958 (N_46958,N_44581,N_42618);
nor U46959 (N_46959,N_43452,N_44315);
or U46960 (N_46960,N_43806,N_43915);
nand U46961 (N_46961,N_44489,N_44487);
xnor U46962 (N_46962,N_44214,N_42973);
nor U46963 (N_46963,N_43624,N_44532);
xnor U46964 (N_46964,N_43923,N_43327);
and U46965 (N_46965,N_44209,N_44036);
nor U46966 (N_46966,N_42742,N_43874);
nor U46967 (N_46967,N_43502,N_44875);
and U46968 (N_46968,N_44033,N_42503);
and U46969 (N_46969,N_43768,N_43179);
nand U46970 (N_46970,N_43749,N_42870);
or U46971 (N_46971,N_43451,N_43755);
or U46972 (N_46972,N_44493,N_43371);
nand U46973 (N_46973,N_43835,N_43880);
xnor U46974 (N_46974,N_44131,N_44274);
and U46975 (N_46975,N_44671,N_44270);
nand U46976 (N_46976,N_44609,N_44020);
nand U46977 (N_46977,N_43487,N_44529);
nand U46978 (N_46978,N_44527,N_43865);
and U46979 (N_46979,N_43366,N_43037);
nor U46980 (N_46980,N_43460,N_43741);
or U46981 (N_46981,N_43995,N_44322);
xor U46982 (N_46982,N_43884,N_42916);
xor U46983 (N_46983,N_44388,N_43105);
xor U46984 (N_46984,N_44092,N_43731);
nor U46985 (N_46985,N_42979,N_44337);
nor U46986 (N_46986,N_44767,N_44502);
xor U46987 (N_46987,N_44911,N_44884);
and U46988 (N_46988,N_42791,N_43927);
or U46989 (N_46989,N_43872,N_42858);
and U46990 (N_46990,N_44410,N_42792);
xnor U46991 (N_46991,N_43076,N_42504);
xnor U46992 (N_46992,N_42733,N_43884);
nand U46993 (N_46993,N_44643,N_44218);
nand U46994 (N_46994,N_44551,N_44741);
nand U46995 (N_46995,N_42535,N_44017);
nand U46996 (N_46996,N_42680,N_43360);
or U46997 (N_46997,N_43499,N_43562);
nand U46998 (N_46998,N_44589,N_43688);
nand U46999 (N_46999,N_44845,N_44443);
xnor U47000 (N_47000,N_44151,N_42812);
xor U47001 (N_47001,N_44175,N_43879);
nand U47002 (N_47002,N_42897,N_44014);
and U47003 (N_47003,N_44578,N_44954);
xor U47004 (N_47004,N_44409,N_44470);
xor U47005 (N_47005,N_43408,N_42765);
or U47006 (N_47006,N_44732,N_42657);
and U47007 (N_47007,N_42717,N_44414);
xor U47008 (N_47008,N_44549,N_44412);
nor U47009 (N_47009,N_44710,N_44040);
or U47010 (N_47010,N_44936,N_42597);
xor U47011 (N_47011,N_43442,N_43874);
nor U47012 (N_47012,N_44276,N_44823);
or U47013 (N_47013,N_42834,N_43096);
or U47014 (N_47014,N_42653,N_43289);
xnor U47015 (N_47015,N_43060,N_42983);
nor U47016 (N_47016,N_44456,N_43205);
or U47017 (N_47017,N_43488,N_44441);
nand U47018 (N_47018,N_44820,N_42691);
or U47019 (N_47019,N_44663,N_42903);
xor U47020 (N_47020,N_43332,N_42986);
xnor U47021 (N_47021,N_43212,N_42688);
and U47022 (N_47022,N_44392,N_43030);
xnor U47023 (N_47023,N_44704,N_44296);
nand U47024 (N_47024,N_43538,N_44474);
xnor U47025 (N_47025,N_44158,N_43312);
nand U47026 (N_47026,N_42718,N_44926);
nor U47027 (N_47027,N_44198,N_42819);
nand U47028 (N_47028,N_42991,N_43982);
nor U47029 (N_47029,N_43476,N_44107);
or U47030 (N_47030,N_43826,N_43662);
nand U47031 (N_47031,N_43568,N_44143);
nor U47032 (N_47032,N_43900,N_43637);
nor U47033 (N_47033,N_42531,N_42587);
xnor U47034 (N_47034,N_43485,N_43696);
nor U47035 (N_47035,N_42570,N_42959);
nor U47036 (N_47036,N_42595,N_43068);
nor U47037 (N_47037,N_43513,N_43516);
nor U47038 (N_47038,N_44761,N_44468);
xnor U47039 (N_47039,N_42719,N_42617);
nand U47040 (N_47040,N_42957,N_43017);
xor U47041 (N_47041,N_42998,N_43831);
xor U47042 (N_47042,N_43821,N_42976);
xnor U47043 (N_47043,N_43533,N_43365);
nor U47044 (N_47044,N_42998,N_44394);
or U47045 (N_47045,N_43999,N_43090);
nor U47046 (N_47046,N_43011,N_42879);
and U47047 (N_47047,N_43679,N_44898);
nor U47048 (N_47048,N_42997,N_42879);
xor U47049 (N_47049,N_43298,N_44687);
xor U47050 (N_47050,N_44757,N_42538);
nor U47051 (N_47051,N_43790,N_44941);
and U47052 (N_47052,N_42593,N_43756);
nor U47053 (N_47053,N_44063,N_44736);
nand U47054 (N_47054,N_42962,N_44018);
and U47055 (N_47055,N_43846,N_43785);
or U47056 (N_47056,N_43937,N_44346);
nor U47057 (N_47057,N_42551,N_42597);
xnor U47058 (N_47058,N_43751,N_44843);
or U47059 (N_47059,N_42935,N_43225);
or U47060 (N_47060,N_44026,N_43101);
and U47061 (N_47061,N_43821,N_44545);
and U47062 (N_47062,N_43394,N_42630);
xnor U47063 (N_47063,N_43673,N_44067);
xnor U47064 (N_47064,N_44960,N_44646);
nor U47065 (N_47065,N_43820,N_43114);
or U47066 (N_47066,N_44137,N_44386);
xor U47067 (N_47067,N_44797,N_43918);
xor U47068 (N_47068,N_43479,N_42715);
xor U47069 (N_47069,N_43120,N_44641);
xnor U47070 (N_47070,N_44841,N_44977);
nor U47071 (N_47071,N_44708,N_42943);
xor U47072 (N_47072,N_42784,N_44862);
and U47073 (N_47073,N_43777,N_44667);
xnor U47074 (N_47074,N_42949,N_44129);
xor U47075 (N_47075,N_44272,N_44373);
nor U47076 (N_47076,N_44720,N_42873);
and U47077 (N_47077,N_42879,N_42573);
or U47078 (N_47078,N_43074,N_43344);
xnor U47079 (N_47079,N_43646,N_43768);
xor U47080 (N_47080,N_43091,N_43621);
nand U47081 (N_47081,N_44022,N_44606);
or U47082 (N_47082,N_43863,N_43619);
and U47083 (N_47083,N_42898,N_44817);
nor U47084 (N_47084,N_44496,N_42564);
xor U47085 (N_47085,N_43266,N_44305);
and U47086 (N_47086,N_43415,N_44763);
xnor U47087 (N_47087,N_44954,N_44369);
nand U47088 (N_47088,N_44610,N_42684);
or U47089 (N_47089,N_42645,N_43807);
xnor U47090 (N_47090,N_44612,N_44275);
xnor U47091 (N_47091,N_44637,N_42658);
nor U47092 (N_47092,N_42792,N_43529);
and U47093 (N_47093,N_44243,N_43667);
nor U47094 (N_47094,N_43142,N_43778);
nor U47095 (N_47095,N_43864,N_43262);
xnor U47096 (N_47096,N_42990,N_43762);
xor U47097 (N_47097,N_43849,N_44043);
nor U47098 (N_47098,N_43280,N_42737);
nand U47099 (N_47099,N_43948,N_44658);
or U47100 (N_47100,N_43834,N_42708);
nor U47101 (N_47101,N_43937,N_43582);
nor U47102 (N_47102,N_44881,N_44924);
or U47103 (N_47103,N_43652,N_42867);
nand U47104 (N_47104,N_43975,N_42704);
xor U47105 (N_47105,N_44731,N_43862);
or U47106 (N_47106,N_43042,N_42795);
and U47107 (N_47107,N_43249,N_43959);
and U47108 (N_47108,N_44698,N_44737);
xnor U47109 (N_47109,N_43894,N_44187);
and U47110 (N_47110,N_43537,N_44207);
xor U47111 (N_47111,N_43429,N_43116);
nand U47112 (N_47112,N_43111,N_42890);
and U47113 (N_47113,N_42657,N_44698);
nor U47114 (N_47114,N_43616,N_44923);
or U47115 (N_47115,N_43889,N_43929);
nand U47116 (N_47116,N_43852,N_44055);
or U47117 (N_47117,N_43003,N_44552);
and U47118 (N_47118,N_44180,N_44537);
nand U47119 (N_47119,N_43809,N_43346);
and U47120 (N_47120,N_42969,N_43515);
and U47121 (N_47121,N_44758,N_42836);
nand U47122 (N_47122,N_44555,N_44020);
nand U47123 (N_47123,N_44769,N_43349);
nand U47124 (N_47124,N_44494,N_42806);
nor U47125 (N_47125,N_43597,N_43913);
or U47126 (N_47126,N_44446,N_43217);
xnor U47127 (N_47127,N_44863,N_44091);
and U47128 (N_47128,N_44377,N_44770);
xnor U47129 (N_47129,N_42772,N_44919);
and U47130 (N_47130,N_43477,N_43155);
and U47131 (N_47131,N_42891,N_43983);
and U47132 (N_47132,N_44169,N_44203);
xor U47133 (N_47133,N_44111,N_44502);
nor U47134 (N_47134,N_43045,N_42643);
nor U47135 (N_47135,N_44143,N_44535);
or U47136 (N_47136,N_44423,N_44745);
or U47137 (N_47137,N_43597,N_44480);
and U47138 (N_47138,N_43097,N_42771);
nor U47139 (N_47139,N_44611,N_44312);
nand U47140 (N_47140,N_43617,N_44343);
nor U47141 (N_47141,N_44145,N_43033);
nand U47142 (N_47142,N_43673,N_43892);
nor U47143 (N_47143,N_43175,N_42841);
nand U47144 (N_47144,N_44463,N_44582);
or U47145 (N_47145,N_44665,N_42867);
xnor U47146 (N_47146,N_43987,N_43770);
or U47147 (N_47147,N_44758,N_44147);
and U47148 (N_47148,N_44748,N_44921);
and U47149 (N_47149,N_44789,N_42939);
xor U47150 (N_47150,N_44789,N_43685);
nor U47151 (N_47151,N_43836,N_44206);
nand U47152 (N_47152,N_44681,N_44050);
or U47153 (N_47153,N_44170,N_43521);
or U47154 (N_47154,N_43020,N_43300);
and U47155 (N_47155,N_42670,N_44671);
or U47156 (N_47156,N_43826,N_43111);
and U47157 (N_47157,N_44409,N_43689);
and U47158 (N_47158,N_44068,N_44284);
nand U47159 (N_47159,N_43848,N_44242);
nor U47160 (N_47160,N_44505,N_42584);
nand U47161 (N_47161,N_43537,N_44073);
or U47162 (N_47162,N_43252,N_42880);
nand U47163 (N_47163,N_42938,N_43142);
and U47164 (N_47164,N_43302,N_42613);
and U47165 (N_47165,N_44163,N_43427);
nor U47166 (N_47166,N_42964,N_43142);
and U47167 (N_47167,N_43434,N_43996);
xor U47168 (N_47168,N_43027,N_43468);
xor U47169 (N_47169,N_43146,N_43587);
nand U47170 (N_47170,N_43656,N_44591);
or U47171 (N_47171,N_44359,N_42984);
nor U47172 (N_47172,N_43973,N_42754);
nand U47173 (N_47173,N_44553,N_43705);
or U47174 (N_47174,N_44640,N_42781);
or U47175 (N_47175,N_43512,N_42704);
or U47176 (N_47176,N_44334,N_44177);
nor U47177 (N_47177,N_42864,N_43561);
nand U47178 (N_47178,N_42696,N_42862);
nand U47179 (N_47179,N_43449,N_43066);
nand U47180 (N_47180,N_43578,N_42958);
nor U47181 (N_47181,N_43186,N_44191);
xor U47182 (N_47182,N_43938,N_44765);
nor U47183 (N_47183,N_43720,N_42529);
nor U47184 (N_47184,N_42894,N_44846);
xnor U47185 (N_47185,N_43420,N_43728);
and U47186 (N_47186,N_43984,N_43693);
and U47187 (N_47187,N_43294,N_43761);
nor U47188 (N_47188,N_43979,N_43304);
nor U47189 (N_47189,N_42989,N_43241);
xor U47190 (N_47190,N_44893,N_43710);
nand U47191 (N_47191,N_44956,N_43937);
xor U47192 (N_47192,N_43411,N_44136);
nor U47193 (N_47193,N_44256,N_42849);
nor U47194 (N_47194,N_43881,N_43382);
nand U47195 (N_47195,N_44900,N_44366);
nand U47196 (N_47196,N_44431,N_43442);
nor U47197 (N_47197,N_44104,N_44755);
and U47198 (N_47198,N_43553,N_43403);
and U47199 (N_47199,N_43874,N_42623);
and U47200 (N_47200,N_42562,N_43285);
nor U47201 (N_47201,N_43316,N_44310);
nand U47202 (N_47202,N_44596,N_43712);
xor U47203 (N_47203,N_44233,N_43244);
xor U47204 (N_47204,N_42807,N_42564);
and U47205 (N_47205,N_42512,N_43481);
xor U47206 (N_47206,N_43573,N_44893);
and U47207 (N_47207,N_43057,N_44254);
or U47208 (N_47208,N_44079,N_44015);
xor U47209 (N_47209,N_42645,N_43467);
nand U47210 (N_47210,N_42776,N_43476);
and U47211 (N_47211,N_43048,N_43236);
or U47212 (N_47212,N_44090,N_43298);
or U47213 (N_47213,N_44191,N_43830);
nor U47214 (N_47214,N_43824,N_44837);
or U47215 (N_47215,N_42881,N_42567);
or U47216 (N_47216,N_43214,N_43096);
nand U47217 (N_47217,N_42869,N_44947);
and U47218 (N_47218,N_44257,N_43302);
xor U47219 (N_47219,N_43782,N_43137);
nor U47220 (N_47220,N_43625,N_43104);
xnor U47221 (N_47221,N_44608,N_44571);
xnor U47222 (N_47222,N_42661,N_42563);
xor U47223 (N_47223,N_43795,N_44266);
xor U47224 (N_47224,N_42779,N_43470);
and U47225 (N_47225,N_42927,N_43959);
nand U47226 (N_47226,N_44833,N_44398);
nand U47227 (N_47227,N_44974,N_43828);
nor U47228 (N_47228,N_43814,N_44412);
and U47229 (N_47229,N_43225,N_44343);
nor U47230 (N_47230,N_43442,N_42781);
or U47231 (N_47231,N_43577,N_44851);
nand U47232 (N_47232,N_44818,N_42825);
xnor U47233 (N_47233,N_44250,N_44752);
nor U47234 (N_47234,N_42923,N_42515);
and U47235 (N_47235,N_43298,N_43441);
or U47236 (N_47236,N_43966,N_43453);
nand U47237 (N_47237,N_44954,N_42552);
nand U47238 (N_47238,N_43462,N_43125);
xnor U47239 (N_47239,N_43383,N_44413);
or U47240 (N_47240,N_44491,N_43554);
or U47241 (N_47241,N_43248,N_43983);
nand U47242 (N_47242,N_44569,N_44121);
nor U47243 (N_47243,N_43414,N_44816);
nor U47244 (N_47244,N_43118,N_42897);
or U47245 (N_47245,N_44545,N_44390);
nor U47246 (N_47246,N_43266,N_44030);
nand U47247 (N_47247,N_43790,N_44848);
nand U47248 (N_47248,N_43410,N_43571);
nand U47249 (N_47249,N_42614,N_43057);
nand U47250 (N_47250,N_44020,N_43250);
and U47251 (N_47251,N_43791,N_43289);
xor U47252 (N_47252,N_44924,N_43461);
nor U47253 (N_47253,N_44758,N_43337);
nor U47254 (N_47254,N_43323,N_44708);
or U47255 (N_47255,N_44636,N_43213);
or U47256 (N_47256,N_44179,N_42843);
or U47257 (N_47257,N_42956,N_43751);
nand U47258 (N_47258,N_43260,N_44156);
and U47259 (N_47259,N_43196,N_43304);
nand U47260 (N_47260,N_44922,N_42995);
or U47261 (N_47261,N_44876,N_44088);
and U47262 (N_47262,N_43559,N_43171);
xor U47263 (N_47263,N_44507,N_44406);
nand U47264 (N_47264,N_43635,N_44928);
xnor U47265 (N_47265,N_43089,N_43918);
or U47266 (N_47266,N_43505,N_42942);
xnor U47267 (N_47267,N_44904,N_42615);
or U47268 (N_47268,N_43272,N_44476);
xnor U47269 (N_47269,N_43211,N_44088);
nand U47270 (N_47270,N_42628,N_42979);
nor U47271 (N_47271,N_43367,N_43362);
xor U47272 (N_47272,N_44137,N_43908);
xor U47273 (N_47273,N_43812,N_43928);
nand U47274 (N_47274,N_44757,N_42514);
or U47275 (N_47275,N_43143,N_43731);
or U47276 (N_47276,N_43163,N_44382);
and U47277 (N_47277,N_42514,N_43819);
nand U47278 (N_47278,N_44126,N_42834);
and U47279 (N_47279,N_43919,N_44585);
xor U47280 (N_47280,N_44939,N_43606);
and U47281 (N_47281,N_42684,N_43061);
nor U47282 (N_47282,N_42612,N_44486);
nor U47283 (N_47283,N_43505,N_44656);
or U47284 (N_47284,N_43101,N_44936);
xor U47285 (N_47285,N_43115,N_43343);
nand U47286 (N_47286,N_43860,N_44089);
or U47287 (N_47287,N_42819,N_43953);
nor U47288 (N_47288,N_43754,N_44334);
nand U47289 (N_47289,N_44865,N_42958);
and U47290 (N_47290,N_43560,N_42527);
and U47291 (N_47291,N_43305,N_42952);
and U47292 (N_47292,N_42949,N_42737);
and U47293 (N_47293,N_43472,N_44103);
xnor U47294 (N_47294,N_44722,N_43019);
nor U47295 (N_47295,N_44768,N_42580);
or U47296 (N_47296,N_44831,N_44062);
or U47297 (N_47297,N_42906,N_44931);
and U47298 (N_47298,N_44745,N_43294);
nor U47299 (N_47299,N_43056,N_43330);
xor U47300 (N_47300,N_43407,N_43860);
and U47301 (N_47301,N_44930,N_43628);
xnor U47302 (N_47302,N_43259,N_42845);
nor U47303 (N_47303,N_44593,N_44881);
or U47304 (N_47304,N_42622,N_44841);
nor U47305 (N_47305,N_44177,N_43746);
xor U47306 (N_47306,N_43135,N_44342);
xor U47307 (N_47307,N_43403,N_42694);
or U47308 (N_47308,N_44211,N_44600);
and U47309 (N_47309,N_43677,N_43012);
xor U47310 (N_47310,N_44512,N_44744);
nand U47311 (N_47311,N_43672,N_44175);
xor U47312 (N_47312,N_44356,N_44679);
nand U47313 (N_47313,N_44165,N_43995);
xnor U47314 (N_47314,N_43237,N_44025);
and U47315 (N_47315,N_43992,N_43645);
or U47316 (N_47316,N_44987,N_43195);
xnor U47317 (N_47317,N_43248,N_44668);
and U47318 (N_47318,N_43031,N_43989);
or U47319 (N_47319,N_42961,N_43133);
and U47320 (N_47320,N_43964,N_44827);
or U47321 (N_47321,N_43265,N_43712);
or U47322 (N_47322,N_43711,N_43281);
xnor U47323 (N_47323,N_44344,N_43601);
and U47324 (N_47324,N_43818,N_43067);
and U47325 (N_47325,N_43889,N_43181);
xor U47326 (N_47326,N_44257,N_43387);
or U47327 (N_47327,N_43912,N_42696);
nor U47328 (N_47328,N_43972,N_43615);
xor U47329 (N_47329,N_43185,N_43246);
xor U47330 (N_47330,N_44690,N_44123);
nor U47331 (N_47331,N_43572,N_44053);
or U47332 (N_47332,N_44013,N_44980);
and U47333 (N_47333,N_44368,N_43311);
xnor U47334 (N_47334,N_43678,N_43795);
and U47335 (N_47335,N_44750,N_44825);
and U47336 (N_47336,N_42591,N_44029);
xnor U47337 (N_47337,N_44213,N_44835);
and U47338 (N_47338,N_44584,N_44960);
nand U47339 (N_47339,N_43938,N_44076);
xnor U47340 (N_47340,N_43619,N_43874);
nor U47341 (N_47341,N_43378,N_44422);
and U47342 (N_47342,N_44967,N_42999);
xnor U47343 (N_47343,N_44279,N_42773);
nor U47344 (N_47344,N_42622,N_43364);
xor U47345 (N_47345,N_43909,N_43090);
nand U47346 (N_47346,N_44441,N_44462);
xor U47347 (N_47347,N_44158,N_44673);
nor U47348 (N_47348,N_42763,N_43533);
nor U47349 (N_47349,N_44569,N_42757);
or U47350 (N_47350,N_44116,N_43536);
and U47351 (N_47351,N_44685,N_44187);
nand U47352 (N_47352,N_43301,N_42548);
nand U47353 (N_47353,N_44102,N_43734);
and U47354 (N_47354,N_44786,N_43906);
xor U47355 (N_47355,N_42540,N_44396);
xnor U47356 (N_47356,N_42779,N_43730);
and U47357 (N_47357,N_43724,N_44799);
xnor U47358 (N_47358,N_44234,N_44106);
xnor U47359 (N_47359,N_43402,N_43203);
nand U47360 (N_47360,N_43522,N_43198);
nand U47361 (N_47361,N_43423,N_43743);
nand U47362 (N_47362,N_43663,N_44003);
nor U47363 (N_47363,N_42854,N_43565);
and U47364 (N_47364,N_44461,N_43080);
and U47365 (N_47365,N_44506,N_43756);
xnor U47366 (N_47366,N_42541,N_43226);
nor U47367 (N_47367,N_44088,N_44310);
and U47368 (N_47368,N_43153,N_44768);
or U47369 (N_47369,N_44589,N_43930);
xnor U47370 (N_47370,N_44321,N_42982);
nor U47371 (N_47371,N_44917,N_44251);
and U47372 (N_47372,N_44347,N_44022);
or U47373 (N_47373,N_44680,N_42604);
or U47374 (N_47374,N_43808,N_44259);
nand U47375 (N_47375,N_44529,N_42896);
or U47376 (N_47376,N_44845,N_43884);
or U47377 (N_47377,N_42642,N_44478);
xor U47378 (N_47378,N_43023,N_43709);
or U47379 (N_47379,N_44831,N_44326);
and U47380 (N_47380,N_44349,N_43070);
nor U47381 (N_47381,N_44230,N_43428);
and U47382 (N_47382,N_43738,N_43421);
nor U47383 (N_47383,N_43404,N_43072);
nor U47384 (N_47384,N_44540,N_44575);
and U47385 (N_47385,N_44239,N_44604);
and U47386 (N_47386,N_44808,N_43288);
nor U47387 (N_47387,N_44867,N_44435);
nor U47388 (N_47388,N_44678,N_42899);
nand U47389 (N_47389,N_44492,N_43035);
xor U47390 (N_47390,N_43187,N_43426);
xnor U47391 (N_47391,N_42682,N_44896);
xnor U47392 (N_47392,N_43621,N_44263);
or U47393 (N_47393,N_43798,N_42688);
nor U47394 (N_47394,N_43212,N_42597);
nor U47395 (N_47395,N_43472,N_43604);
or U47396 (N_47396,N_43932,N_44033);
nor U47397 (N_47397,N_42966,N_43475);
nor U47398 (N_47398,N_42865,N_44872);
and U47399 (N_47399,N_44231,N_44934);
and U47400 (N_47400,N_42907,N_44161);
nor U47401 (N_47401,N_42886,N_43138);
or U47402 (N_47402,N_42686,N_44809);
nor U47403 (N_47403,N_43864,N_43643);
nor U47404 (N_47404,N_42880,N_43903);
nand U47405 (N_47405,N_43898,N_43724);
nor U47406 (N_47406,N_44573,N_42672);
or U47407 (N_47407,N_43850,N_42513);
or U47408 (N_47408,N_43455,N_43274);
nor U47409 (N_47409,N_43832,N_44842);
or U47410 (N_47410,N_43940,N_44529);
nor U47411 (N_47411,N_44612,N_44122);
nand U47412 (N_47412,N_42822,N_43139);
and U47413 (N_47413,N_43966,N_42986);
or U47414 (N_47414,N_42945,N_44139);
or U47415 (N_47415,N_44862,N_44777);
xor U47416 (N_47416,N_43604,N_44421);
or U47417 (N_47417,N_44869,N_42920);
nor U47418 (N_47418,N_42829,N_44169);
and U47419 (N_47419,N_44021,N_44433);
xor U47420 (N_47420,N_43898,N_43485);
nand U47421 (N_47421,N_44226,N_44187);
and U47422 (N_47422,N_43896,N_43630);
and U47423 (N_47423,N_44611,N_43613);
nand U47424 (N_47424,N_43284,N_42786);
or U47425 (N_47425,N_43109,N_44924);
nor U47426 (N_47426,N_42694,N_43348);
nor U47427 (N_47427,N_42670,N_43709);
and U47428 (N_47428,N_43639,N_42975);
or U47429 (N_47429,N_42772,N_43844);
and U47430 (N_47430,N_44641,N_44289);
xor U47431 (N_47431,N_44962,N_43050);
xnor U47432 (N_47432,N_43251,N_43441);
or U47433 (N_47433,N_44128,N_42798);
nor U47434 (N_47434,N_43813,N_44163);
and U47435 (N_47435,N_43402,N_43650);
nand U47436 (N_47436,N_43905,N_43809);
or U47437 (N_47437,N_42942,N_44831);
and U47438 (N_47438,N_42688,N_44136);
and U47439 (N_47439,N_44326,N_42687);
nor U47440 (N_47440,N_43033,N_42869);
and U47441 (N_47441,N_43227,N_42808);
nor U47442 (N_47442,N_43221,N_44980);
and U47443 (N_47443,N_43164,N_43469);
nor U47444 (N_47444,N_42516,N_44607);
and U47445 (N_47445,N_43391,N_43866);
xor U47446 (N_47446,N_42636,N_43031);
nand U47447 (N_47447,N_43201,N_42968);
nand U47448 (N_47448,N_44329,N_44640);
and U47449 (N_47449,N_44484,N_44820);
xnor U47450 (N_47450,N_43655,N_43224);
or U47451 (N_47451,N_44616,N_44695);
xor U47452 (N_47452,N_43909,N_43575);
nand U47453 (N_47453,N_43957,N_44670);
nand U47454 (N_47454,N_43104,N_44872);
xor U47455 (N_47455,N_44185,N_42610);
nor U47456 (N_47456,N_44104,N_44306);
nor U47457 (N_47457,N_44992,N_44464);
and U47458 (N_47458,N_44519,N_42928);
nand U47459 (N_47459,N_42959,N_43861);
xnor U47460 (N_47460,N_43523,N_44432);
or U47461 (N_47461,N_44973,N_44615);
nand U47462 (N_47462,N_43416,N_44610);
nand U47463 (N_47463,N_42762,N_42801);
or U47464 (N_47464,N_44836,N_44296);
or U47465 (N_47465,N_44384,N_43789);
nor U47466 (N_47466,N_43096,N_44483);
nor U47467 (N_47467,N_44287,N_43222);
and U47468 (N_47468,N_44336,N_42565);
xor U47469 (N_47469,N_44051,N_43618);
nand U47470 (N_47470,N_43738,N_43896);
and U47471 (N_47471,N_44652,N_44368);
nand U47472 (N_47472,N_42827,N_43937);
nand U47473 (N_47473,N_44225,N_43562);
nor U47474 (N_47474,N_44903,N_44667);
or U47475 (N_47475,N_43009,N_44939);
xor U47476 (N_47476,N_44982,N_44354);
and U47477 (N_47477,N_44351,N_42709);
xnor U47478 (N_47478,N_42506,N_44085);
or U47479 (N_47479,N_43880,N_43058);
xnor U47480 (N_47480,N_43090,N_43415);
or U47481 (N_47481,N_42885,N_43775);
nor U47482 (N_47482,N_43298,N_44544);
and U47483 (N_47483,N_42586,N_43944);
and U47484 (N_47484,N_43624,N_42683);
xor U47485 (N_47485,N_44297,N_44063);
nor U47486 (N_47486,N_44982,N_42592);
nor U47487 (N_47487,N_44742,N_44186);
nand U47488 (N_47488,N_44560,N_43661);
nor U47489 (N_47489,N_44323,N_44898);
and U47490 (N_47490,N_43217,N_42608);
nor U47491 (N_47491,N_44613,N_43758);
or U47492 (N_47492,N_42951,N_43394);
nand U47493 (N_47493,N_43065,N_44841);
nand U47494 (N_47494,N_42816,N_44783);
nand U47495 (N_47495,N_43756,N_42921);
xnor U47496 (N_47496,N_44882,N_43846);
nor U47497 (N_47497,N_44468,N_44662);
or U47498 (N_47498,N_42673,N_43564);
nand U47499 (N_47499,N_44816,N_42607);
and U47500 (N_47500,N_46722,N_45836);
and U47501 (N_47501,N_46417,N_46712);
nor U47502 (N_47502,N_45480,N_45007);
nor U47503 (N_47503,N_45419,N_46308);
and U47504 (N_47504,N_46669,N_46327);
nand U47505 (N_47505,N_47195,N_46470);
nand U47506 (N_47506,N_46189,N_46320);
or U47507 (N_47507,N_45244,N_46093);
nand U47508 (N_47508,N_45665,N_46268);
or U47509 (N_47509,N_45631,N_45871);
nor U47510 (N_47510,N_45863,N_47261);
and U47511 (N_47511,N_47116,N_45979);
xnor U47512 (N_47512,N_45864,N_45664);
xor U47513 (N_47513,N_45336,N_47349);
nand U47514 (N_47514,N_45744,N_45512);
xnor U47515 (N_47515,N_45596,N_46517);
nor U47516 (N_47516,N_47136,N_45049);
nor U47517 (N_47517,N_46210,N_45261);
nor U47518 (N_47518,N_46905,N_45453);
xor U47519 (N_47519,N_45893,N_45442);
nand U47520 (N_47520,N_45354,N_47313);
xor U47521 (N_47521,N_46205,N_46435);
or U47522 (N_47522,N_46059,N_47166);
and U47523 (N_47523,N_46812,N_47318);
or U47524 (N_47524,N_45643,N_45425);
and U47525 (N_47525,N_47455,N_45878);
nor U47526 (N_47526,N_47023,N_46472);
nor U47527 (N_47527,N_46975,N_47452);
nand U47528 (N_47528,N_45868,N_47167);
nor U47529 (N_47529,N_45200,N_47079);
nand U47530 (N_47530,N_45750,N_45048);
nand U47531 (N_47531,N_46816,N_45950);
or U47532 (N_47532,N_45167,N_45745);
nand U47533 (N_47533,N_46265,N_45296);
nor U47534 (N_47534,N_46491,N_47286);
and U47535 (N_47535,N_46895,N_46989);
and U47536 (N_47536,N_46706,N_45806);
nand U47537 (N_47537,N_46565,N_45133);
or U47538 (N_47538,N_46777,N_47225);
nand U47539 (N_47539,N_46430,N_46645);
nor U47540 (N_47540,N_46578,N_45498);
nand U47541 (N_47541,N_46527,N_46376);
nand U47542 (N_47542,N_46525,N_45972);
nor U47543 (N_47543,N_47105,N_47255);
and U47544 (N_47544,N_47087,N_46882);
nand U47545 (N_47545,N_46735,N_46571);
and U47546 (N_47546,N_45809,N_45628);
xor U47547 (N_47547,N_46555,N_45513);
or U47548 (N_47548,N_46022,N_47338);
and U47549 (N_47549,N_46450,N_45392);
nand U47550 (N_47550,N_46971,N_46233);
xnor U47551 (N_47551,N_46631,N_46587);
nor U47552 (N_47552,N_45753,N_46613);
nand U47553 (N_47553,N_45931,N_47353);
nand U47554 (N_47554,N_45873,N_45627);
xor U47555 (N_47555,N_46532,N_45340);
and U47556 (N_47556,N_45918,N_45349);
xor U47557 (N_47557,N_46946,N_46674);
and U47558 (N_47558,N_45091,N_45082);
xnor U47559 (N_47559,N_45090,N_46064);
nor U47560 (N_47560,N_46090,N_45071);
and U47561 (N_47561,N_45074,N_47182);
xnor U47562 (N_47562,N_46909,N_46838);
nand U47563 (N_47563,N_45062,N_46299);
nor U47564 (N_47564,N_46862,N_46158);
or U47565 (N_47565,N_45834,N_45667);
and U47566 (N_47566,N_46643,N_45487);
nand U47567 (N_47567,N_45663,N_46634);
nor U47568 (N_47568,N_45684,N_45781);
or U47569 (N_47569,N_46419,N_47153);
nor U47570 (N_47570,N_45333,N_45535);
and U47571 (N_47571,N_46237,N_45678);
nand U47572 (N_47572,N_45112,N_45951);
xor U47573 (N_47573,N_46983,N_46902);
nor U47574 (N_47574,N_45479,N_45465);
nor U47575 (N_47575,N_45367,N_46732);
or U47576 (N_47576,N_47330,N_46904);
nor U47577 (N_47577,N_47265,N_46951);
xor U47578 (N_47578,N_45694,N_47326);
nand U47579 (N_47579,N_46958,N_45636);
nor U47580 (N_47580,N_45120,N_46918);
xnor U47581 (N_47581,N_46508,N_47333);
nand U47582 (N_47582,N_45433,N_46745);
xnor U47583 (N_47583,N_45175,N_47275);
nor U47584 (N_47584,N_45242,N_45432);
or U47585 (N_47585,N_45788,N_46938);
nor U47586 (N_47586,N_46206,N_45124);
nand U47587 (N_47587,N_45289,N_45592);
nor U47588 (N_47588,N_46744,N_45517);
xor U47589 (N_47589,N_45867,N_46025);
nand U47590 (N_47590,N_46992,N_46252);
nor U47591 (N_47591,N_46843,N_45552);
xor U47592 (N_47592,N_47289,N_46341);
nor U47593 (N_47593,N_45227,N_45073);
nor U47594 (N_47594,N_46139,N_45875);
nand U47595 (N_47595,N_46344,N_47483);
and U47596 (N_47596,N_46941,N_46316);
and U47597 (N_47597,N_47430,N_46700);
nor U47598 (N_47598,N_45219,N_46468);
nand U47599 (N_47599,N_47253,N_46833);
nand U47600 (N_47600,N_46442,N_45445);
xor U47601 (N_47601,N_45356,N_47207);
nor U47602 (N_47602,N_47017,N_46134);
xor U47603 (N_47603,N_47325,N_45718);
nand U47604 (N_47604,N_45658,N_46209);
nor U47605 (N_47605,N_45965,N_46774);
xor U47606 (N_47606,N_46784,N_46600);
nor U47607 (N_47607,N_45539,N_45096);
nand U47608 (N_47608,N_47071,N_45383);
nand U47609 (N_47609,N_46590,N_46378);
nand U47610 (N_47610,N_46962,N_47061);
and U47611 (N_47611,N_46692,N_45942);
or U47612 (N_47612,N_46225,N_46171);
or U47613 (N_47613,N_46231,N_45571);
nor U47614 (N_47614,N_46754,N_46760);
or U47615 (N_47615,N_45524,N_47106);
xnor U47616 (N_47616,N_45766,N_46884);
nand U47617 (N_47617,N_45110,N_47141);
nand U47618 (N_47618,N_45825,N_45856);
nor U47619 (N_47619,N_47357,N_46543);
nand U47620 (N_47620,N_46329,N_45474);
xor U47621 (N_47621,N_46602,N_45443);
and U47622 (N_47622,N_46597,N_46293);
or U47623 (N_47623,N_46827,N_45786);
and U47624 (N_47624,N_47189,N_46428);
nor U47625 (N_47625,N_46787,N_46886);
and U47626 (N_47626,N_45258,N_46803);
and U47627 (N_47627,N_45176,N_46390);
nor U47628 (N_47628,N_46551,N_46738);
nand U47629 (N_47629,N_45095,N_46421);
nand U47630 (N_47630,N_46924,N_45174);
or U47631 (N_47631,N_47216,N_46709);
and U47632 (N_47632,N_47276,N_46452);
or U47633 (N_47633,N_46808,N_47047);
xor U47634 (N_47634,N_45463,N_47347);
nor U47635 (N_47635,N_46516,N_45970);
and U47636 (N_47636,N_46057,N_46739);
nor U47637 (N_47637,N_47468,N_45317);
and U47638 (N_47638,N_47285,N_45015);
nand U47639 (N_47639,N_47191,N_46708);
nand U47640 (N_47640,N_46748,N_46496);
or U47641 (N_47641,N_46557,N_45136);
xnor U47642 (N_47642,N_45936,N_46098);
nand U47643 (N_47643,N_47142,N_45906);
xnor U47644 (N_47644,N_46074,N_46141);
or U47645 (N_47645,N_45382,N_45470);
nor U47646 (N_47646,N_45689,N_45464);
xor U47647 (N_47647,N_45923,N_45917);
nand U47648 (N_47648,N_45012,N_46050);
nand U47649 (N_47649,N_45758,N_45948);
xnor U47650 (N_47650,N_46072,N_45471);
nor U47651 (N_47651,N_46668,N_46312);
nor U47652 (N_47652,N_47193,N_45975);
and U47653 (N_47653,N_47200,N_46250);
xor U47654 (N_47654,N_46153,N_47376);
xnor U47655 (N_47655,N_46832,N_47158);
or U47656 (N_47656,N_46475,N_46907);
or U47657 (N_47657,N_46004,N_46878);
xnor U47658 (N_47658,N_47161,N_45288);
or U47659 (N_47659,N_46531,N_45222);
xnor U47660 (N_47660,N_45169,N_45104);
xnor U47661 (N_47661,N_47054,N_45985);
nor U47662 (N_47662,N_45191,N_45661);
nand U47663 (N_47663,N_45251,N_46718);
nand U47664 (N_47664,N_45248,N_47089);
xnor U47665 (N_47665,N_46815,N_46092);
or U47666 (N_47666,N_45599,N_45990);
nand U47667 (N_47667,N_47108,N_46552);
nand U47668 (N_47668,N_47438,N_45347);
and U47669 (N_47669,N_45605,N_45737);
or U47670 (N_47670,N_46337,N_46349);
nor U47671 (N_47671,N_46103,N_46805);
or U47672 (N_47672,N_45780,N_46730);
or U47673 (N_47673,N_46725,N_45114);
and U47674 (N_47674,N_46868,N_46023);
nor U47675 (N_47675,N_46829,N_46936);
and U47676 (N_47676,N_46279,N_46498);
nor U47677 (N_47677,N_45804,N_45092);
nor U47678 (N_47678,N_46288,N_46129);
nor U47679 (N_47679,N_45041,N_46016);
or U47680 (N_47680,N_45139,N_46203);
xnor U47681 (N_47681,N_46703,N_45327);
and U47682 (N_47682,N_46467,N_47145);
xor U47683 (N_47683,N_45763,N_46284);
nor U47684 (N_47684,N_47323,N_45037);
nor U47685 (N_47685,N_47282,N_47043);
or U47686 (N_47686,N_45971,N_45277);
xor U47687 (N_47687,N_46729,N_46121);
and U47688 (N_47688,N_45156,N_46786);
and U47689 (N_47689,N_47209,N_46304);
nor U47690 (N_47690,N_45282,N_46647);
xnor U47691 (N_47691,N_45003,N_45161);
xor U47692 (N_47692,N_46236,N_46949);
xnor U47693 (N_47693,N_45707,N_45125);
or U47694 (N_47694,N_45103,N_46133);
or U47695 (N_47695,N_46441,N_45185);
and U47696 (N_47696,N_45920,N_45500);
xnor U47697 (N_47697,N_45572,N_45439);
or U47698 (N_47698,N_47477,N_45325);
xor U47699 (N_47699,N_45947,N_45118);
nand U47700 (N_47700,N_47097,N_45397);
nand U47701 (N_47701,N_47025,N_46996);
nor U47702 (N_47702,N_46906,N_45388);
xor U47703 (N_47703,N_46202,N_45884);
and U47704 (N_47704,N_46056,N_46926);
and U47705 (N_47705,N_45771,N_46144);
nand U47706 (N_47706,N_46124,N_46753);
nor U47707 (N_47707,N_45673,N_46953);
nor U47708 (N_47708,N_46523,N_46569);
xor U47709 (N_47709,N_45712,N_45623);
xor U47710 (N_47710,N_45431,N_47311);
xor U47711 (N_47711,N_46545,N_45329);
and U47712 (N_47712,N_46086,N_47434);
nand U47713 (N_47713,N_46686,N_45818);
xnor U47714 (N_47714,N_45391,N_45536);
xor U47715 (N_47715,N_45608,N_45014);
and U47716 (N_47716,N_46876,N_47082);
nor U47717 (N_47717,N_45020,N_45373);
or U47718 (N_47718,N_46285,N_45900);
nand U47719 (N_47719,N_47143,N_46095);
nand U47720 (N_47720,N_47059,N_45057);
or U47721 (N_47721,N_46822,N_45768);
nor U47722 (N_47722,N_46873,N_47171);
nand U47723 (N_47723,N_46084,N_45241);
xor U47724 (N_47724,N_46656,N_46561);
nor U47725 (N_47725,N_47174,N_45348);
or U47726 (N_47726,N_45466,N_45494);
or U47727 (N_47727,N_46264,N_46995);
xor U47728 (N_47728,N_46781,N_46967);
and U47729 (N_47729,N_46179,N_47331);
nand U47730 (N_47730,N_46658,N_45764);
nor U47731 (N_47731,N_46679,N_45220);
nand U47732 (N_47732,N_45098,N_46782);
nand U47733 (N_47733,N_46954,N_46834);
xnor U47734 (N_47734,N_47493,N_45430);
and U47735 (N_47735,N_45591,N_45675);
and U47736 (N_47736,N_46038,N_46506);
xnor U47737 (N_47737,N_46529,N_46020);
or U47738 (N_47738,N_47044,N_46934);
or U47739 (N_47739,N_46639,N_46006);
or U47740 (N_47740,N_47274,N_47283);
nand U47741 (N_47741,N_47442,N_45668);
and U47742 (N_47742,N_47203,N_46877);
nor U47743 (N_47743,N_45701,N_46355);
or U47744 (N_47744,N_47354,N_45314);
nor U47745 (N_47745,N_47155,N_47366);
xor U47746 (N_47746,N_45696,N_47443);
nor U47747 (N_47747,N_46969,N_45145);
and U47748 (N_47748,N_45190,N_46903);
nand U47749 (N_47749,N_46823,N_46794);
or U47750 (N_47750,N_47410,N_46388);
and U47751 (N_47751,N_46535,N_46610);
nor U47752 (N_47752,N_45759,N_46033);
nor U47753 (N_47753,N_46977,N_45787);
xor U47754 (N_47754,N_47169,N_46885);
xnor U47755 (N_47755,N_47341,N_45569);
and U47756 (N_47756,N_46193,N_46190);
nand U47757 (N_47757,N_46112,N_45642);
or U47758 (N_47758,N_46150,N_46110);
xnor U47759 (N_47759,N_46397,N_45243);
xnor U47760 (N_47760,N_46125,N_46979);
nor U47761 (N_47761,N_46240,N_45400);
nor U47762 (N_47762,N_45761,N_45656);
and U47763 (N_47763,N_47399,N_47495);
or U47764 (N_47764,N_46858,N_45278);
nand U47765 (N_47765,N_46069,N_46401);
or U47766 (N_47766,N_45000,N_46861);
nor U47767 (N_47767,N_47221,N_45719);
or U47768 (N_47768,N_45529,N_47026);
and U47769 (N_47769,N_47473,N_45021);
nor U47770 (N_47770,N_46117,N_47369);
and U47771 (N_47771,N_47236,N_45089);
or U47772 (N_47772,N_46440,N_46165);
nor U47773 (N_47773,N_46721,N_46292);
and U47774 (N_47774,N_46598,N_45024);
and U47775 (N_47775,N_45973,N_46601);
and U47776 (N_47776,N_46260,N_46661);
and U47777 (N_47777,N_45937,N_45410);
and U47778 (N_47778,N_47303,N_46772);
nand U47779 (N_47779,N_46177,N_46502);
and U47780 (N_47780,N_45616,N_46961);
xor U47781 (N_47781,N_47428,N_45308);
nand U47782 (N_47782,N_45724,N_45823);
or U47783 (N_47783,N_45032,N_45259);
or U47784 (N_47784,N_46461,N_46769);
nand U47785 (N_47785,N_46290,N_45618);
nor U47786 (N_47786,N_45651,N_46447);
nand U47787 (N_47787,N_45757,N_47383);
xnor U47788 (N_47788,N_47472,N_45217);
or U47789 (N_47789,N_47295,N_45444);
and U47790 (N_47790,N_45484,N_47280);
xor U47791 (N_47791,N_46194,N_46364);
nand U47792 (N_47792,N_47441,N_46889);
nor U47793 (N_47793,N_46495,N_46955);
xnor U47794 (N_47794,N_45551,N_45413);
nor U47795 (N_47795,N_45793,N_45612);
xor U47796 (N_47796,N_47407,N_45921);
nand U47797 (N_47797,N_46615,N_46762);
nand U47798 (N_47798,N_45727,N_46159);
xnor U47799 (N_47799,N_47304,N_45914);
and U47800 (N_47800,N_46462,N_45546);
and U47801 (N_47801,N_45803,N_45141);
xor U47802 (N_47802,N_46415,N_45047);
or U47803 (N_47803,N_45025,N_46314);
or U47804 (N_47804,N_46514,N_45137);
nor U47805 (N_47805,N_46881,N_45202);
and U47806 (N_47806,N_47034,N_47154);
nor U47807 (N_47807,N_46148,N_45322);
and U47808 (N_47808,N_45235,N_45832);
nand U47809 (N_47809,N_45997,N_47462);
or U47810 (N_47810,N_45518,N_45849);
or U47811 (N_47811,N_46581,N_45850);
nand U47812 (N_47812,N_46296,N_46383);
or U47813 (N_47813,N_45581,N_46638);
or U47814 (N_47814,N_46576,N_46997);
xor U47815 (N_47815,N_45194,N_45983);
nor U47816 (N_47816,N_45426,N_46046);
and U47817 (N_47817,N_45009,N_46717);
xor U47818 (N_47818,N_47273,N_45609);
and U47819 (N_47819,N_45648,N_45215);
xnor U47820 (N_47820,N_46431,N_46008);
xnor U47821 (N_47821,N_46132,N_47078);
nand U47822 (N_47822,N_45507,N_45550);
nor U47823 (N_47823,N_47422,N_45943);
or U47824 (N_47824,N_47279,N_47228);
nor U47825 (N_47825,N_47086,N_47481);
nor U47826 (N_47826,N_47467,N_46653);
or U47827 (N_47827,N_46908,N_46809);
and U47828 (N_47828,N_45967,N_45102);
xnor U47829 (N_47829,N_45326,N_47309);
and U47830 (N_47830,N_45735,N_45252);
nand U47831 (N_47831,N_46437,N_46648);
or U47832 (N_47832,N_45741,N_45495);
nor U47833 (N_47833,N_45239,N_47450);
or U47834 (N_47834,N_45929,N_47117);
xnor U47835 (N_47835,N_45690,N_46389);
and U47836 (N_47836,N_47316,N_46524);
and U47837 (N_47837,N_45221,N_46277);
or U47838 (N_47838,N_46584,N_46677);
nand U47839 (N_47839,N_45515,N_46088);
nor U47840 (N_47840,N_45894,N_45820);
nand U47841 (N_47841,N_46330,N_45127);
and U47842 (N_47842,N_45740,N_45401);
nand U47843 (N_47843,N_47464,N_46328);
xnor U47844 (N_47844,N_45926,N_45122);
nor U47845 (N_47845,N_47220,N_45455);
and U47846 (N_47846,N_45417,N_45105);
and U47847 (N_47847,N_45010,N_45903);
nor U47848 (N_47848,N_46505,N_47440);
and U47849 (N_47849,N_45398,N_46019);
nand U47850 (N_47850,N_47498,N_45891);
and U47851 (N_47851,N_45418,N_47489);
nor U47852 (N_47852,N_45146,N_45055);
and U47853 (N_47853,N_46374,N_45414);
or U47854 (N_47854,N_46494,N_46040);
xor U47855 (N_47855,N_47270,N_47342);
nand U47856 (N_47856,N_47425,N_46254);
and U47857 (N_47857,N_45813,N_45980);
or U47858 (N_47858,N_46985,N_46258);
nand U47859 (N_47859,N_46164,N_46411);
nor U47860 (N_47860,N_45944,N_46119);
or U47861 (N_47861,N_45595,N_45113);
or U47862 (N_47862,N_45538,N_47198);
xor U47863 (N_47863,N_46840,N_45530);
nand U47864 (N_47864,N_46800,N_46935);
xnor U47865 (N_47865,N_46499,N_45094);
nor U47866 (N_47866,N_45794,N_47242);
nor U47867 (N_47867,N_45059,N_47256);
xnor U47868 (N_47868,N_46222,N_46306);
nand U47869 (N_47869,N_45304,N_46097);
and U47870 (N_47870,N_45162,N_47126);
nand U47871 (N_47871,N_46649,N_47094);
nor U47872 (N_47872,N_45170,N_46066);
and U47873 (N_47873,N_46562,N_45692);
and U47874 (N_47874,N_47192,N_45924);
or U47875 (N_47875,N_47496,N_45674);
nor U47876 (N_47876,N_47490,N_47360);
nor U47877 (N_47877,N_45478,N_46990);
or U47878 (N_47878,N_45669,N_45065);
nor U47879 (N_47879,N_46965,N_45229);
nor U47880 (N_47880,N_45755,N_46939);
and U47881 (N_47881,N_45160,N_45896);
xnor U47882 (N_47882,N_46298,N_45468);
nand U47883 (N_47883,N_47214,N_45188);
and U47884 (N_47884,N_46695,N_45607);
nand U47885 (N_47885,N_46670,N_45353);
nor U47886 (N_47886,N_45149,N_46262);
or U47887 (N_47887,N_46127,N_47343);
xnor U47888 (N_47888,N_47235,N_45423);
nor U47889 (N_47889,N_45729,N_45840);
xor U47890 (N_47890,N_45361,N_45912);
and U47891 (N_47891,N_46187,N_46465);
nor U47892 (N_47892,N_46080,N_46436);
nor U47893 (N_47893,N_46195,N_47476);
nor U47894 (N_47894,N_47057,N_47243);
or U47895 (N_47895,N_45441,N_46434);
nor U47896 (N_47896,N_46636,N_46872);
nand U47897 (N_47897,N_45109,N_46563);
nand U47898 (N_47898,N_46333,N_46911);
and U47899 (N_47899,N_45998,N_45152);
nand U47900 (N_47900,N_46247,N_45790);
nand U47901 (N_47901,N_46303,N_47437);
and U47902 (N_47902,N_46269,N_46849);
xor U47903 (N_47903,N_47446,N_45670);
nor U47904 (N_47904,N_45231,N_46572);
and U47905 (N_47905,N_47085,N_46487);
xor U47906 (N_47906,N_45331,N_45715);
nor U47907 (N_47907,N_46566,N_46497);
nand U47908 (N_47908,N_46783,N_47172);
xor U47909 (N_47909,N_45532,N_46375);
or U47910 (N_47910,N_47239,N_45387);
xnor U47911 (N_47911,N_46931,N_46807);
xor U47912 (N_47912,N_46507,N_45654);
xnor U47913 (N_47913,N_46035,N_46414);
or U47914 (N_47914,N_46361,N_46830);
nor U47915 (N_47915,N_45533,N_45201);
nand U47916 (N_47916,N_46342,N_46313);
and U47917 (N_47917,N_45240,N_45974);
nor U47918 (N_47918,N_45290,N_47277);
nand U47919 (N_47919,N_45386,N_46272);
nand U47920 (N_47920,N_45380,N_45862);
and U47921 (N_47921,N_45534,N_45352);
or U47922 (N_47922,N_46646,N_45403);
xor U47923 (N_47923,N_45454,N_45343);
and U47924 (N_47924,N_45427,N_47188);
or U47925 (N_47925,N_45482,N_46409);
or U47926 (N_47926,N_45063,N_45449);
xnor U47927 (N_47927,N_45457,N_45580);
or U47928 (N_47928,N_45377,N_45779);
xor U47929 (N_47929,N_47077,N_45205);
xor U47930 (N_47930,N_46232,N_46002);
nand U47931 (N_47931,N_45826,N_45540);
nor U47932 (N_47932,N_46973,N_47164);
and U47933 (N_47933,N_46256,N_45143);
xnor U47934 (N_47934,N_45323,N_47014);
nor U47935 (N_47935,N_46652,N_46404);
nand U47936 (N_47936,N_47305,N_45379);
xnor U47937 (N_47937,N_47069,N_45526);
or U47938 (N_47938,N_46131,N_46261);
or U47939 (N_47939,N_46458,N_45519);
or U47940 (N_47940,N_45742,N_47453);
xor U47941 (N_47941,N_47372,N_46896);
nor U47942 (N_47942,N_47393,N_46140);
or U47943 (N_47943,N_46180,N_46920);
nor U47944 (N_47944,N_45281,N_46609);
or U47945 (N_47945,N_45368,N_46888);
nor U47946 (N_47946,N_45301,N_46867);
xnor U47947 (N_47947,N_47226,N_45123);
nand U47948 (N_47948,N_46053,N_46844);
nand U47949 (N_47949,N_46287,N_45691);
and U47950 (N_47950,N_45560,N_46077);
nor U47951 (N_47951,N_46152,N_46795);
nand U47952 (N_47952,N_46947,N_45385);
nor U47953 (N_47953,N_46591,N_46244);
and U47954 (N_47954,N_46412,N_47262);
nor U47955 (N_47955,N_47395,N_46693);
xor U47956 (N_47956,N_45469,N_45237);
and U47957 (N_47957,N_47184,N_45004);
or U47958 (N_47958,N_47412,N_47392);
nor U47959 (N_47959,N_47118,N_47063);
nand U47960 (N_47960,N_47083,N_46410);
xor U47961 (N_47961,N_46914,N_45869);
and U47962 (N_47962,N_46104,N_47321);
nand U47963 (N_47963,N_45837,N_46301);
xor U47964 (N_47964,N_45203,N_46013);
xor U47965 (N_47965,N_47478,N_45275);
and U47966 (N_47966,N_46900,N_46549);
xnor U47967 (N_47967,N_45134,N_46338);
nand U47968 (N_47968,N_47474,N_45624);
and U47969 (N_47969,N_47456,N_45283);
nor U47970 (N_47970,N_47370,N_46922);
nand U47971 (N_47971,N_45859,N_45611);
and U47972 (N_47972,N_47170,N_46921);
or U47973 (N_47973,N_46765,N_46100);
or U47974 (N_47974,N_46325,N_45585);
and U47975 (N_47975,N_45216,N_45316);
and U47976 (N_47976,N_45357,N_47486);
and U47977 (N_47977,N_47045,N_46460);
or U47978 (N_47978,N_45877,N_45557);
and U47979 (N_47979,N_45785,N_46605);
and U47980 (N_47980,N_45119,N_45762);
xnor U47981 (N_47981,N_46398,N_47218);
and U47982 (N_47982,N_45026,N_45197);
or U47983 (N_47983,N_46477,N_46763);
nand U47984 (N_47984,N_45365,N_45841);
and U47985 (N_47985,N_46220,N_46974);
or U47986 (N_47986,N_45969,N_46281);
and U47987 (N_47987,N_45559,N_45196);
xnor U47988 (N_47988,N_45360,N_46122);
or U47989 (N_47989,N_45590,N_45001);
xor U47990 (N_47990,N_45922,N_46276);
or U47991 (N_47991,N_46758,N_45842);
xnor U47992 (N_47992,N_45472,N_46094);
and U47993 (N_47993,N_45698,N_47092);
xnor U47994 (N_47994,N_47140,N_46752);
nand U47995 (N_47995,N_47436,N_46522);
nor U47996 (N_47996,N_46928,N_45051);
nand U47997 (N_47997,N_45284,N_45263);
or U47998 (N_47998,N_46170,N_46887);
and U47999 (N_47999,N_45582,N_45371);
nand U48000 (N_48000,N_46893,N_45456);
or U48001 (N_48001,N_46459,N_45638);
and U48002 (N_48002,N_45435,N_47367);
nor U48003 (N_48003,N_46620,N_46484);
nor U48004 (N_48004,N_45030,N_45556);
nand U48005 (N_48005,N_46317,N_46537);
nor U48006 (N_48006,N_45218,N_47396);
and U48007 (N_48007,N_45086,N_46335);
nand U48008 (N_48008,N_46676,N_46925);
nand U48009 (N_48009,N_45135,N_46446);
nand U48010 (N_48010,N_47127,N_46628);
nand U48011 (N_48011,N_45491,N_45565);
nand U48012 (N_48012,N_47049,N_46396);
nand U48013 (N_48013,N_45399,N_45271);
or U48014 (N_48014,N_46612,N_45600);
nand U48015 (N_48015,N_47006,N_45866);
and U48016 (N_48016,N_47028,N_45262);
nand U48017 (N_48017,N_45671,N_46845);
xor U48018 (N_48018,N_47130,N_47397);
and U48019 (N_48019,N_46149,N_47038);
nand U48020 (N_48020,N_46257,N_45537);
nor U48021 (N_48021,N_45475,N_47009);
and U48022 (N_48022,N_46988,N_46115);
nand U48023 (N_48023,N_47156,N_47135);
nand U48024 (N_48024,N_46423,N_47109);
nor U48025 (N_48025,N_45374,N_46055);
or U48026 (N_48026,N_45492,N_46749);
or U48027 (N_48027,N_46542,N_47074);
or U48028 (N_48028,N_45111,N_46061);
or U48029 (N_48029,N_45531,N_46444);
nand U48030 (N_48030,N_46854,N_46981);
nand U48031 (N_48031,N_46466,N_46607);
xnor U48032 (N_48032,N_46229,N_45952);
xnor U48033 (N_48033,N_45601,N_45774);
xnor U48034 (N_48034,N_46818,N_46780);
or U48035 (N_48035,N_45976,N_47314);
nand U48036 (N_48036,N_46650,N_47091);
or U48037 (N_48037,N_46245,N_46366);
nor U48038 (N_48038,N_46720,N_46003);
nand U48039 (N_48039,N_45816,N_46583);
xor U48040 (N_48040,N_45760,N_46624);
nand U48041 (N_48041,N_47252,N_47013);
nand U48042 (N_48042,N_45097,N_46336);
nand U48043 (N_48043,N_45428,N_47004);
or U48044 (N_48044,N_47281,N_45140);
or U48045 (N_48045,N_47124,N_46633);
nor U48046 (N_48046,N_47335,N_45064);
xor U48047 (N_48047,N_47202,N_47211);
and U48048 (N_48048,N_47199,N_46091);
nor U48049 (N_48049,N_47012,N_46511);
nor U48050 (N_48050,N_46196,N_45044);
nor U48051 (N_48051,N_46326,N_46021);
and U48052 (N_48052,N_45730,N_45812);
or U48053 (N_48053,N_45264,N_46356);
and U48054 (N_48054,N_47042,N_46406);
and U48055 (N_48055,N_46369,N_46041);
nand U48056 (N_48056,N_47249,N_46479);
or U48057 (N_48057,N_45299,N_47458);
nor U48058 (N_48058,N_46207,N_45452);
nor U48059 (N_48059,N_46663,N_46391);
or U48060 (N_48060,N_46146,N_47445);
xor U48061 (N_48061,N_45851,N_46901);
nor U48062 (N_48062,N_47463,N_46533);
nor U48063 (N_48063,N_46595,N_46048);
or U48064 (N_48064,N_46109,N_45748);
xnor U48065 (N_48065,N_47128,N_45228);
and U48066 (N_48066,N_45725,N_45083);
xnor U48067 (N_48067,N_47010,N_46968);
or U48068 (N_48068,N_45652,N_47329);
or U48069 (N_48069,N_46184,N_45687);
or U48070 (N_48070,N_47151,N_47173);
or U48071 (N_48071,N_45933,N_45293);
nor U48072 (N_48072,N_45236,N_46482);
nor U48073 (N_48073,N_46539,N_46185);
nand U48074 (N_48074,N_47352,N_47241);
xnor U48075 (N_48075,N_45320,N_46315);
nand U48076 (N_48076,N_47100,N_45378);
xnor U48077 (N_48077,N_46300,N_46667);
xor U48078 (N_48078,N_45233,N_45728);
or U48079 (N_48079,N_45568,N_46474);
nor U48080 (N_48080,N_47324,N_47389);
nand U48081 (N_48081,N_46183,N_46167);
nand U48082 (N_48082,N_47138,N_45946);
nand U48083 (N_48083,N_45459,N_45751);
nor U48084 (N_48084,N_45662,N_45959);
or U48085 (N_48085,N_45265,N_46821);
and U48086 (N_48086,N_45831,N_46802);
nand U48087 (N_48087,N_45366,N_46420);
and U48088 (N_48088,N_45558,N_45625);
nor U48089 (N_48089,N_45968,N_45722);
nand U48090 (N_48090,N_45930,N_45076);
and U48091 (N_48091,N_45306,N_46156);
nor U48092 (N_48092,N_45364,N_45958);
xor U48093 (N_48093,N_45328,N_45710);
and U48094 (N_48094,N_45807,N_46513);
nor U48095 (N_48095,N_47254,N_46987);
nand U48096 (N_48096,N_45060,N_47248);
nor U48097 (N_48097,N_45503,N_46181);
or U48098 (N_48098,N_46501,N_45649);
xor U48099 (N_48099,N_45409,N_45892);
nand U48100 (N_48100,N_45376,N_45525);
nand U48101 (N_48101,N_47084,N_46520);
and U48102 (N_48102,N_46831,N_46696);
nor U48103 (N_48103,N_45610,N_46847);
or U48104 (N_48104,N_46480,N_47264);
and U48105 (N_48105,N_46012,N_46972);
or U48106 (N_48106,N_45126,N_46427);
or U48107 (N_48107,N_45198,N_45870);
nand U48108 (N_48108,N_46182,N_46123);
nand U48109 (N_48109,N_46814,N_45838);
nor U48110 (N_48110,N_46734,N_47417);
xor U48111 (N_48111,N_46826,N_46898);
xor U48112 (N_48112,N_45158,N_46626);
xnor U48113 (N_48113,N_45286,N_46850);
xnor U48114 (N_48114,N_46702,N_45372);
and U48115 (N_48115,N_45440,N_45801);
or U48116 (N_48116,N_45700,N_47148);
nor U48117 (N_48117,N_45270,N_46295);
or U48118 (N_48118,N_47426,N_46916);
or U48119 (N_48119,N_45230,N_46963);
nor U48120 (N_48120,N_46548,N_47177);
nor U48121 (N_48121,N_45319,N_46943);
xnor U48122 (N_48122,N_46200,N_46451);
xnor U48123 (N_48123,N_45783,N_45986);
xor U48124 (N_48124,N_47390,N_46560);
and U48125 (N_48125,N_47051,N_45370);
xor U48126 (N_48126,N_46836,N_45462);
nand U48127 (N_48127,N_45318,N_46354);
xnor U48128 (N_48128,N_46864,N_47245);
xnor U48129 (N_48129,N_45412,N_45645);
or U48130 (N_48130,N_46363,N_46596);
xor U48131 (N_48131,N_46169,N_47457);
nand U48132 (N_48132,N_45053,N_45274);
nand U48133 (N_48133,N_46332,N_46614);
xor U48134 (N_48134,N_45738,N_46286);
or U48135 (N_48135,N_47373,N_46034);
xor U48136 (N_48136,N_45876,N_45106);
xor U48137 (N_48137,N_45705,N_46318);
nand U48138 (N_48138,N_46622,N_47433);
or U48139 (N_48139,N_47288,N_47301);
nand U48140 (N_48140,N_46028,N_47224);
nand U48141 (N_48141,N_46768,N_46155);
and U48142 (N_48142,N_46280,N_45938);
nand U48143 (N_48143,N_47336,N_45827);
xor U48144 (N_48144,N_45042,N_45593);
xnor U48145 (N_48145,N_45527,N_46689);
nor U48146 (N_48146,N_47423,N_46007);
or U48147 (N_48147,N_45437,N_47284);
or U48148 (N_48148,N_47419,N_47293);
xor U48149 (N_48149,N_46359,N_46603);
nor U48150 (N_48150,N_47053,N_47133);
xor U48151 (N_48151,N_46932,N_45522);
nor U48152 (N_48152,N_47016,N_45576);
xnor U48153 (N_48153,N_46945,N_45545);
nor U48154 (N_48154,N_45548,N_45819);
xnor U48155 (N_48155,N_47206,N_46348);
nor U48156 (N_48156,N_46485,N_45606);
or U48157 (N_48157,N_46087,N_46456);
xor U48158 (N_48158,N_46740,N_46340);
and U48159 (N_48159,N_45155,N_46585);
nor U48160 (N_48160,N_45544,N_45285);
xnor U48161 (N_48161,N_45257,N_45346);
or U48162 (N_48162,N_46799,N_46789);
and U48163 (N_48163,N_45736,N_46687);
nand U48164 (N_48164,N_45359,N_46915);
nor U48165 (N_48165,N_46559,N_45509);
xnor U48166 (N_48166,N_46682,N_47027);
xor U48167 (N_48167,N_46851,N_45038);
nand U48168 (N_48168,N_46510,N_45117);
xor U48169 (N_48169,N_46933,N_45486);
xor U48170 (N_48170,N_45775,N_45206);
nand U48171 (N_48171,N_45415,N_45888);
or U48172 (N_48172,N_45254,N_45630);
xnor U48173 (N_48173,N_46071,N_45626);
or U48174 (N_48174,N_46278,N_45050);
or U48175 (N_48175,N_45996,N_45991);
nand U48176 (N_48176,N_46422,N_45273);
nand U48177 (N_48177,N_46089,N_47230);
and U48178 (N_48178,N_45685,N_46589);
xor U48179 (N_48179,N_45436,N_45798);
nand U48180 (N_48180,N_45199,N_46067);
nor U48181 (N_48181,N_47292,N_47011);
xnor U48182 (N_48182,N_45511,N_46345);
or U48183 (N_48183,N_46358,N_46418);
nor U48184 (N_48184,N_47185,N_45256);
xor U48185 (N_48185,N_45178,N_45496);
xnor U48186 (N_48186,N_46493,N_45054);
nor U48187 (N_48187,N_46757,N_46011);
or U48188 (N_48188,N_45901,N_45887);
nand U48189 (N_48189,N_47150,N_46913);
nand U48190 (N_48190,N_46635,N_46099);
xnor U48191 (N_48191,N_47110,N_46357);
or U48192 (N_48192,N_47015,N_45767);
nor U48193 (N_48193,N_47339,N_47232);
or U48194 (N_48194,N_45072,N_46813);
nor U48195 (N_48195,N_45928,N_46393);
or U48196 (N_48196,N_45132,N_46065);
or U48197 (N_48197,N_47056,N_46764);
nand U48198 (N_48198,N_45573,N_46641);
or U48199 (N_48199,N_47146,N_46727);
and U48200 (N_48200,N_46439,N_46713);
nand U48201 (N_48201,N_45776,N_45695);
xnor U48202 (N_48202,N_46360,N_46828);
and U48203 (N_48203,N_47421,N_47413);
xor U48204 (N_48204,N_46917,N_46394);
nand U48205 (N_48205,N_47411,N_46793);
and U48206 (N_48206,N_46554,N_47394);
nor U48207 (N_48207,N_45702,N_45192);
and U48208 (N_48208,N_46956,N_46168);
or U48209 (N_48209,N_47040,N_47068);
xor U48210 (N_48210,N_47424,N_46592);
xor U48211 (N_48211,N_46515,N_45902);
nand U48212 (N_48212,N_46835,N_45619);
nor U48213 (N_48213,N_46970,N_45287);
and U48214 (N_48214,N_45660,N_46899);
xor U48215 (N_48215,N_45267,N_45028);
nand U48216 (N_48216,N_47008,N_47222);
nand U48217 (N_48217,N_46509,N_47340);
nand U48218 (N_48218,N_45334,N_45238);
and U48219 (N_48219,N_46761,N_46416);
or U48220 (N_48220,N_47119,N_45335);
nand U48221 (N_48221,N_47296,N_46604);
and U48222 (N_48222,N_47359,N_47361);
and U48223 (N_48223,N_47186,N_45956);
nor U48224 (N_48224,N_45617,N_46213);
xor U48225 (N_48225,N_45210,N_45731);
nor U48226 (N_48226,N_45756,N_47487);
nand U48227 (N_48227,N_45303,N_45822);
and U48228 (N_48228,N_46798,N_45232);
or U48229 (N_48229,N_45846,N_47227);
or U48230 (N_48230,N_46319,N_46352);
xor U48231 (N_48231,N_45321,N_46688);
nor U48232 (N_48232,N_47033,N_45337);
xnor U48233 (N_48233,N_45088,N_45080);
and U48234 (N_48234,N_47259,N_45772);
or U48235 (N_48235,N_45148,N_45406);
nand U48236 (N_48236,N_45844,N_46483);
and U48237 (N_48237,N_45659,N_45186);
or U48238 (N_48238,N_46302,N_45182);
nor U48239 (N_48239,N_46930,N_47307);
nor U48240 (N_48240,N_46683,N_45693);
and U48241 (N_48241,N_46944,N_46950);
nor U48242 (N_48242,N_46534,N_45784);
nor U48243 (N_48243,N_45204,N_47479);
and U48244 (N_48244,N_45005,N_46120);
or U48245 (N_48245,N_46385,N_47266);
nand U48246 (N_48246,N_47121,N_46910);
xor U48247 (N_48247,N_45575,N_46756);
and U48248 (N_48248,N_47197,N_46825);
or U48249 (N_48249,N_47196,N_45085);
nand U48250 (N_48250,N_45598,N_47090);
nand U48251 (N_48251,N_46018,N_46731);
nand U48252 (N_48252,N_45898,N_46403);
xor U48253 (N_48253,N_46714,N_45481);
xnor U48254 (N_48254,N_46108,N_47050);
and U48255 (N_48255,N_46438,N_47064);
xnor U48256 (N_48256,N_45603,N_46755);
xnor U48257 (N_48257,N_45193,N_47234);
nor U48258 (N_48258,N_46579,N_47448);
nand U48259 (N_48259,N_45294,N_45554);
and U48260 (N_48260,N_45882,N_47175);
nor U48261 (N_48261,N_45602,N_47002);
and U48262 (N_48262,N_47260,N_45108);
xor U48263 (N_48263,N_47246,N_47469);
and U48264 (N_48264,N_45429,N_45514);
xnor U48265 (N_48265,N_45138,N_46518);
nand U48266 (N_48266,N_45075,N_46891);
nand U48267 (N_48267,N_46062,N_46387);
xnor U48268 (N_48268,N_45650,N_45966);
and U48269 (N_48269,N_46157,N_45338);
or U48270 (N_48270,N_46266,N_46346);
nand U48271 (N_48271,N_46392,N_47065);
xnor U48272 (N_48272,N_47388,N_46982);
xnor U48273 (N_48273,N_47374,N_46937);
xor U48274 (N_48274,N_46307,N_47067);
xnor U48275 (N_48275,N_46424,N_45396);
and U48276 (N_48276,N_45613,N_46178);
or U48277 (N_48277,N_45987,N_45164);
and U48278 (N_48278,N_45907,N_45963);
xor U48279 (N_48279,N_46792,N_45635);
and U48280 (N_48280,N_46172,N_46044);
or U48281 (N_48281,N_45808,N_46224);
nand U48282 (N_48282,N_46841,N_46984);
or U48283 (N_48283,N_46678,N_46143);
and U48284 (N_48284,N_46043,N_46353);
xnor U48285 (N_48285,N_46655,N_45578);
or U48286 (N_48286,N_46837,N_45008);
xnor U48287 (N_48287,N_45982,N_45504);
xnor U48288 (N_48288,N_46052,N_46894);
nand U48289 (N_48289,N_45384,N_46544);
and U48290 (N_48290,N_47201,N_46619);
or U48291 (N_48291,N_45587,N_45172);
nor U48292 (N_48292,N_45795,N_45395);
nand U48293 (N_48293,N_46453,N_46215);
xnor U48294 (N_48294,N_46608,N_47075);
nor U48295 (N_48295,N_46351,N_47297);
or U48296 (N_48296,N_45260,N_45422);
nand U48297 (N_48297,N_46801,N_46082);
and U48298 (N_48298,N_45330,N_46386);
xnor U48299 (N_48299,N_46657,N_47400);
nor U48300 (N_48300,N_47107,N_46275);
or U48301 (N_48301,N_45168,N_46690);
or U48302 (N_48302,N_46724,N_46640);
nor U48303 (N_48303,N_46005,N_46654);
or U48304 (N_48304,N_45734,N_47217);
nand U48305 (N_48305,N_46788,N_47088);
nor U48306 (N_48306,N_45011,N_45508);
xnor U48307 (N_48307,N_45066,N_45056);
and U48308 (N_48308,N_45978,N_45821);
xnor U48309 (N_48309,N_47346,N_45477);
and U48310 (N_48310,N_45817,N_47312);
and U48311 (N_48311,N_46454,N_46241);
nor U48312 (N_48312,N_47408,N_45390);
nor U48313 (N_48313,N_46379,N_45189);
or U48314 (N_48314,N_45954,N_46289);
nand U48315 (N_48315,N_47378,N_46443);
nand U48316 (N_48316,N_46031,N_46230);
nand U48317 (N_48317,N_45789,N_47365);
xnor U48318 (N_48318,N_47021,N_46239);
or U48319 (N_48319,N_45144,N_45183);
or U48320 (N_48320,N_45208,N_47037);
and U48321 (N_48321,N_46723,N_47299);
nor U48322 (N_48322,N_47157,N_45639);
and U48323 (N_48323,N_45543,N_46611);
xor U48324 (N_48324,N_45067,N_46381);
and U48325 (N_48325,N_45679,N_47240);
nand U48326 (N_48326,N_46347,N_45101);
xnor U48327 (N_48327,N_47247,N_46489);
nor U48328 (N_48328,N_45013,N_45358);
and U48329 (N_48329,N_46892,N_46234);
nand U48330 (N_48330,N_45115,N_46672);
xor U48331 (N_48331,N_45309,N_46478);
nand U48332 (N_48332,N_45029,N_46796);
or U48333 (N_48333,N_46166,N_46161);
or U48334 (N_48334,N_45280,N_45579);
nand U48335 (N_48335,N_45023,N_45586);
nor U48336 (N_48336,N_46101,N_47039);
xnor U48337 (N_48337,N_46856,N_47095);
nand U48338 (N_48338,N_46001,N_47076);
nand U48339 (N_48339,N_45681,N_46546);
nand U48340 (N_48340,N_45225,N_47454);
or U48341 (N_48341,N_46309,N_45224);
nand U48342 (N_48342,N_45493,N_47380);
or U48343 (N_48343,N_46321,N_46570);
nor U48344 (N_48344,N_45860,N_45516);
nand U48345 (N_48345,N_47497,N_47345);
or U48346 (N_48346,N_47272,N_46147);
or U48347 (N_48347,N_46685,N_45653);
or U48348 (N_48348,N_46449,N_45940);
or U48349 (N_48349,N_46282,N_46399);
and U48350 (N_48350,N_45362,N_46114);
and U48351 (N_48351,N_46865,N_47459);
nand U48352 (N_48352,N_45899,N_46201);
and U48353 (N_48353,N_45855,N_47451);
or U48354 (N_48354,N_45084,N_47144);
nor U48355 (N_48355,N_45988,N_46130);
nor U48356 (N_48356,N_45989,N_45814);
xor U48357 (N_48357,N_45721,N_45570);
nand U48358 (N_48358,N_47058,N_46526);
and U48359 (N_48359,N_46577,N_47268);
or U48360 (N_48360,N_47070,N_47005);
nand U48361 (N_48361,N_45476,N_45555);
nand U48362 (N_48362,N_46223,N_46883);
nor U48363 (N_48363,N_45709,N_45226);
xor U48364 (N_48364,N_46469,N_45297);
and U48365 (N_48365,N_45880,N_47355);
and U48366 (N_48366,N_46929,N_45389);
nand U48367 (N_48367,N_45935,N_46448);
nor U48368 (N_48368,N_45087,N_46273);
or U48369 (N_48369,N_47048,N_46547);
xnor U48370 (N_48370,N_46558,N_46659);
nor U48371 (N_48371,N_46580,N_45852);
xor U48372 (N_48372,N_45939,N_46037);
nor U48373 (N_48373,N_45523,N_46297);
nor U48374 (N_48374,N_45393,N_45791);
xnor U48375 (N_48375,N_46015,N_46574);
nor U48376 (N_48376,N_45036,N_47465);
nand U48377 (N_48377,N_45394,N_45615);
and U48378 (N_48378,N_46890,N_45909);
or U48379 (N_48379,N_46957,N_46274);
or U48380 (N_48380,N_46105,N_47250);
nand U48381 (N_48381,N_46463,N_46039);
and U48382 (N_48382,N_45839,N_47060);
nor U48383 (N_48383,N_47190,N_46785);
and U48384 (N_48384,N_46075,N_46488);
or U48385 (N_48385,N_46637,N_45448);
nor U48386 (N_48386,N_45485,N_46283);
or U48387 (N_48387,N_46618,N_45717);
nand U48388 (N_48388,N_47139,N_46707);
nand U48389 (N_48389,N_47123,N_45874);
and U48390 (N_48390,N_46644,N_45577);
and U48391 (N_48391,N_46912,N_45885);
and U48392 (N_48392,N_46235,N_46630);
nor U48393 (N_48393,N_47332,N_45212);
nand U48394 (N_48394,N_46863,N_45276);
and U48395 (N_48395,N_45910,N_46750);
nor U48396 (N_48396,N_45058,N_45061);
and U48397 (N_48397,N_46671,N_46311);
and U48398 (N_48398,N_47229,N_45574);
xnor U48399 (N_48399,N_46599,N_46528);
nand U48400 (N_48400,N_47215,N_47168);
or U48401 (N_48401,N_45810,N_46625);
or U48402 (N_48402,N_46500,N_47480);
xnor U48403 (N_48403,N_45655,N_47178);
nor U48404 (N_48404,N_45310,N_45154);
and U48405 (N_48405,N_46214,N_47238);
nor U48406 (N_48406,N_45157,N_45131);
xor U48407 (N_48407,N_45018,N_45369);
or U48408 (N_48408,N_46076,N_45686);
nand U48409 (N_48409,N_45777,N_45295);
or U48410 (N_48410,N_46594,N_47187);
nor U48411 (N_48411,N_45905,N_46408);
nand U48412 (N_48412,N_46948,N_47036);
xor U48413 (N_48413,N_45778,N_45640);
xnor U48414 (N_48414,N_46384,N_45677);
nand U48415 (N_48415,N_45733,N_45253);
xnor U48416 (N_48416,N_46804,N_46976);
and U48417 (N_48417,N_45614,N_47194);
nor U48418 (N_48418,N_46163,N_45890);
or U48419 (N_48419,N_46042,N_46192);
xor U48420 (N_48420,N_47449,N_46617);
and U48421 (N_48421,N_45833,N_46365);
xor U48422 (N_48422,N_46853,N_45883);
nor U48423 (N_48423,N_45726,N_46759);
nor U48424 (N_48424,N_45853,N_46490);
nor U48425 (N_48425,N_46136,N_47485);
nand U48426 (N_48426,N_45187,N_45068);
or U48427 (N_48427,N_45932,N_45647);
nor U48428 (N_48428,N_45043,N_46719);
nor U48429 (N_48429,N_45797,N_45099);
and U48430 (N_48430,N_45960,N_45069);
nor U48431 (N_48431,N_45408,N_46073);
or U48432 (N_48432,N_46897,N_45147);
nor U48433 (N_48433,N_46047,N_47431);
xnor U48434 (N_48434,N_45311,N_46536);
nand U48435 (N_48435,N_45246,N_45830);
xor U48436 (N_48436,N_47460,N_46839);
xor U48437 (N_48437,N_46063,N_46162);
nand U48438 (N_48438,N_47470,N_45255);
nor U48439 (N_48439,N_46664,N_46540);
xnor U48440 (N_48440,N_45720,N_45027);
xor U48441 (N_48441,N_45159,N_47384);
nor U48442 (N_48442,N_47018,N_45703);
and U48443 (N_48443,N_47233,N_47080);
and U48444 (N_48444,N_46107,N_45467);
nand U48445 (N_48445,N_45739,N_46871);
nor U48446 (N_48446,N_46869,N_45324);
xor U48447 (N_48447,N_45528,N_45171);
nor U48448 (N_48448,N_47205,N_46323);
nor U48449 (N_48449,N_45116,N_45886);
xor U48450 (N_48450,N_46964,N_46198);
or U48451 (N_48451,N_45796,N_45897);
nand U48452 (N_48452,N_46952,N_46026);
and U48453 (N_48453,N_47387,N_46567);
xnor U48454 (N_48454,N_45107,N_47403);
and U48455 (N_48455,N_45824,N_46530);
xnor U48456 (N_48456,N_46029,N_47237);
or U48457 (N_48457,N_45447,N_47163);
nor U48458 (N_48458,N_47073,N_46267);
nand U48459 (N_48459,N_47294,N_47319);
nor U48460 (N_48460,N_46219,N_45799);
nor U48461 (N_48461,N_46228,N_47405);
and U48462 (N_48462,N_45451,N_45446);
nand U48463 (N_48463,N_47371,N_45142);
nand U48464 (N_48464,N_46698,N_45723);
xor U48465 (N_48465,N_46564,N_47291);
nor U48466 (N_48466,N_47492,N_47398);
or U48467 (N_48467,N_47055,N_46138);
nand U48468 (N_48468,N_46036,N_45405);
or U48469 (N_48469,N_47415,N_46691);
xnor U48470 (N_48470,N_46259,N_46221);
nor U48471 (N_48471,N_46660,N_47102);
or U48472 (N_48472,N_45402,N_45033);
xnor U48473 (N_48473,N_45927,N_45584);
nand U48474 (N_48474,N_47104,N_46694);
xor U48475 (N_48475,N_46588,N_47271);
nand U48476 (N_48476,N_45889,N_46154);
or U48477 (N_48477,N_45501,N_45207);
nand U48478 (N_48478,N_46980,N_46746);
nor U48479 (N_48479,N_47062,N_45502);
and U48480 (N_48480,N_47204,N_46305);
xnor U48481 (N_48481,N_46824,N_46629);
nor U48482 (N_48482,N_47484,N_47499);
or U48483 (N_48483,N_46820,N_46705);
or U48484 (N_48484,N_47114,N_46217);
xnor U48485 (N_48485,N_45594,N_46778);
nor U48486 (N_48486,N_47099,N_46736);
nor U48487 (N_48487,N_45747,N_47429);
nand U48488 (N_48488,N_47404,N_46870);
and U48489 (N_48489,N_45247,N_47244);
and U48490 (N_48490,N_45473,N_45881);
and U48491 (N_48491,N_46771,N_47401);
and U48492 (N_48492,N_47447,N_46227);
nor U48493 (N_48493,N_46846,N_46492);
nor U48494 (N_48494,N_45828,N_45506);
or U48495 (N_48495,N_45743,N_47317);
nand U48496 (N_48496,N_45434,N_45800);
nor U48497 (N_48497,N_45341,N_45017);
nand U48498 (N_48498,N_45714,N_45292);
and U48499 (N_48499,N_46726,N_45567);
xor U48500 (N_48500,N_47420,N_46078);
nor U48501 (N_48501,N_47134,N_46111);
xnor U48502 (N_48502,N_47181,N_45315);
or U48503 (N_48503,N_45424,N_45350);
and U48504 (N_48504,N_46070,N_45597);
nor U48505 (N_48505,N_46249,N_46322);
nor U48506 (N_48506,N_45450,N_45184);
xnor U48507 (N_48507,N_45765,N_45351);
nor U48508 (N_48508,N_45195,N_45621);
and U48509 (N_48509,N_46923,N_47129);
nor U48510 (N_48510,N_47491,N_45070);
xnor U48511 (N_48511,N_45749,N_45815);
and U48512 (N_48512,N_46817,N_46457);
xor U48513 (N_48513,N_47427,N_46135);
and U48514 (N_48514,N_47251,N_46733);
and U48515 (N_48515,N_46860,N_45919);
or U48516 (N_48516,N_45438,N_45847);
and U48517 (N_48517,N_45130,N_45994);
and U48518 (N_48518,N_45505,N_46550);
and U48519 (N_48519,N_47180,N_46791);
or U48520 (N_48520,N_46191,N_47111);
nor U48521 (N_48521,N_46176,N_47375);
nand U48522 (N_48522,N_45019,N_45993);
or U48523 (N_48523,N_46697,N_46334);
or U48524 (N_48524,N_46142,N_45541);
nor U48525 (N_48525,N_47031,N_45040);
nor U48526 (N_48526,N_47302,N_47308);
nor U48527 (N_48527,N_45302,N_45835);
and U48528 (N_48528,N_45564,N_45355);
and U48529 (N_48529,N_47125,N_45266);
and U48530 (N_48530,N_47219,N_45250);
and U48531 (N_48531,N_46174,N_45984);
nor U48532 (N_48532,N_47269,N_45497);
nand U48533 (N_48533,N_46362,N_45272);
xnor U48534 (N_48534,N_46742,N_47231);
nand U48535 (N_48535,N_47391,N_45079);
nor U48536 (N_48536,N_46464,N_46248);
xor U48537 (N_48537,N_46582,N_47032);
xor U48538 (N_48538,N_45925,N_47041);
or U48539 (N_48539,N_45179,N_46291);
nand U48540 (N_48540,N_46331,N_46204);
and U48541 (N_48541,N_46102,N_45699);
and U48542 (N_48542,N_45081,N_47385);
nor U48543 (N_48543,N_45547,N_46538);
nor U48544 (N_48544,N_45632,N_47212);
or U48545 (N_48545,N_46238,N_46819);
nor U48546 (N_48546,N_47379,N_46218);
or U48547 (N_48547,N_46024,N_46875);
or U48548 (N_48548,N_46991,N_47103);
xor U48549 (N_48549,N_45666,N_47377);
nand U48550 (N_48550,N_46400,N_46049);
nor U48551 (N_48551,N_45173,N_47344);
nand U48552 (N_48552,N_45682,N_46113);
and U48553 (N_48553,N_45957,N_45553);
and U48554 (N_48554,N_46553,N_45421);
nand U48555 (N_48555,N_47165,N_47081);
nor U48556 (N_48556,N_47439,N_47382);
nor U48557 (N_48557,N_47471,N_47113);
nor U48558 (N_48558,N_45381,N_47267);
xnor U48559 (N_48559,N_45934,N_45052);
nand U48560 (N_48560,N_45046,N_46779);
or U48561 (N_48561,N_45313,N_47183);
nor U48562 (N_48562,N_47052,N_45214);
and U48563 (N_48563,N_45634,N_45039);
and U48564 (N_48564,N_45520,N_47176);
and U48565 (N_48565,N_47159,N_45848);
and U48566 (N_48566,N_45077,N_47147);
nor U48567 (N_48567,N_47152,N_45407);
xor U48568 (N_48568,N_46993,N_45857);
or U48569 (N_48569,N_47416,N_46010);
or U48570 (N_48570,N_45035,N_47315);
or U48571 (N_48571,N_45209,N_46797);
and U48572 (N_48572,N_45561,N_45298);
xor U48573 (N_48573,N_45811,N_47322);
xor U48574 (N_48574,N_47263,N_46711);
xnor U48575 (N_48575,N_45629,N_46246);
xnor U48576 (N_48576,N_46699,N_46211);
nand U48577 (N_48577,N_46014,N_47351);
nand U48578 (N_48578,N_45908,N_47093);
and U48579 (N_48579,N_46096,N_46481);
nor U48580 (N_48580,N_46271,N_45704);
or U48581 (N_48581,N_46848,N_45915);
nor U48582 (N_48582,N_45488,N_46642);
and U48583 (N_48583,N_46106,N_47482);
xnor U48584 (N_48584,N_45510,N_47290);
or U48585 (N_48585,N_45961,N_47098);
nor U48586 (N_48586,N_46126,N_46575);
xor U48587 (N_48587,N_45093,N_47368);
xor U48588 (N_48588,N_47358,N_46085);
nand U48589 (N_48589,N_47101,N_45583);
xor U48590 (N_48590,N_46519,N_45641);
or U48591 (N_48591,N_46767,N_45644);
and U48592 (N_48592,N_46978,N_45461);
nand U48593 (N_48593,N_46741,N_46175);
nand U48594 (N_48594,N_46445,N_45746);
or U48595 (N_48595,N_45633,N_47402);
nor U48596 (N_48596,N_45688,N_47364);
and U48597 (N_48597,N_46137,N_47475);
nand U48598 (N_48598,N_47320,N_46433);
xor U48599 (N_48599,N_47003,N_45411);
nand U48600 (N_48600,N_46919,N_46866);
and U48601 (N_48601,N_47461,N_47179);
and U48602 (N_48602,N_45305,N_45911);
and U48603 (N_48603,N_47210,N_46242);
or U48604 (N_48604,N_46251,N_46471);
nand U48605 (N_48605,N_45163,N_45344);
or U48606 (N_48606,N_46058,N_46402);
or U48607 (N_48607,N_46373,N_47386);
or U48608 (N_48608,N_47414,N_46504);
xnor U48609 (N_48609,N_46627,N_46060);
and U48610 (N_48610,N_45249,N_47072);
xor U48611 (N_48611,N_46343,N_45805);
xnor U48612 (N_48612,N_46068,N_47112);
nor U48613 (N_48613,N_46350,N_47306);
nand U48614 (N_48614,N_46770,N_45363);
xnor U48615 (N_48615,N_45672,N_46568);
nand U48616 (N_48616,N_47258,N_46429);
nand U48617 (N_48617,N_47162,N_46651);
nor U48618 (N_48618,N_46368,N_45589);
and U48619 (N_48619,N_46473,N_46743);
nor U48620 (N_48620,N_46160,N_46998);
xnor U48621 (N_48621,N_46382,N_47362);
xnor U48622 (N_48622,N_45150,N_46673);
nand U48623 (N_48623,N_45916,N_47035);
xor U48624 (N_48624,N_45620,N_45680);
xnor U48625 (N_48625,N_46879,N_47337);
xnor U48626 (N_48626,N_47160,N_45460);
xor U48627 (N_48627,N_45307,N_47020);
or U48628 (N_48628,N_45121,N_45490);
or U48629 (N_48629,N_45782,N_45002);
or U48630 (N_48630,N_47122,N_46081);
nand U48631 (N_48631,N_45683,N_46675);
and U48632 (N_48632,N_46051,N_47131);
and U48633 (N_48633,N_46371,N_46212);
xor U48634 (N_48634,N_45770,N_45792);
nor U48635 (N_48635,N_45181,N_45291);
and U48636 (N_48636,N_45773,N_46573);
or U48637 (N_48637,N_45312,N_47149);
or U48638 (N_48638,N_45697,N_45879);
nand U48639 (N_48639,N_46666,N_47418);
nand U48640 (N_48640,N_46766,N_45375);
or U48641 (N_48641,N_45416,N_46367);
nand U48642 (N_48642,N_45872,N_47381);
nand U48643 (N_48643,N_47001,N_45031);
nor U48644 (N_48644,N_45151,N_47029);
nand U48645 (N_48645,N_45854,N_46216);
or U48646 (N_48646,N_46186,N_46811);
nor U48647 (N_48647,N_46425,N_47000);
xnor U48648 (N_48648,N_45802,N_47208);
xnor U48649 (N_48649,N_47406,N_46662);
or U48650 (N_48650,N_45016,N_46045);
and U48651 (N_48651,N_45342,N_46665);
nor U48652 (N_48652,N_46857,N_47310);
nor U48653 (N_48653,N_45006,N_46000);
or U48654 (N_48654,N_45962,N_45499);
xor U48655 (N_48655,N_45964,N_45676);
or U48656 (N_48656,N_45657,N_46521);
and U48657 (N_48657,N_46370,N_47046);
nand U48658 (N_48658,N_45022,N_47298);
and U48659 (N_48659,N_45100,N_46199);
or U48660 (N_48660,N_45420,N_46197);
or U48661 (N_48661,N_45861,N_45129);
and U48662 (N_48662,N_47115,N_45332);
xor U48663 (N_48663,N_47300,N_47287);
xnor U48664 (N_48664,N_46874,N_47137);
nor U48665 (N_48665,N_46118,N_45166);
or U48666 (N_48666,N_46455,N_47356);
xor U48667 (N_48667,N_46017,N_46486);
and U48668 (N_48668,N_45521,N_46079);
xor U48669 (N_48669,N_46054,N_45769);
nand U48670 (N_48670,N_46255,N_47494);
xnor U48671 (N_48671,N_46593,N_46188);
and U48672 (N_48672,N_45034,N_46927);
or U48673 (N_48673,N_45752,N_45706);
nor U48674 (N_48674,N_46959,N_46775);
nand U48675 (N_48675,N_46173,N_46395);
nand U48676 (N_48676,N_46806,N_45829);
xnor U48677 (N_48677,N_46715,N_46413);
or U48678 (N_48678,N_45646,N_46226);
or U48679 (N_48679,N_46027,N_45549);
nand U48680 (N_48680,N_47278,N_46632);
nor U48681 (N_48681,N_45945,N_46556);
nor U48682 (N_48682,N_47120,N_45895);
nor U48683 (N_48683,N_46586,N_46855);
or U48684 (N_48684,N_46681,N_45234);
nand U48685 (N_48685,N_45339,N_47328);
nand U48686 (N_48686,N_46751,N_46324);
nand U48687 (N_48687,N_46116,N_47132);
and U48688 (N_48688,N_46747,N_45268);
or U48689 (N_48689,N_46940,N_46339);
nor U48690 (N_48690,N_46616,N_45180);
nor U48691 (N_48691,N_45845,N_46503);
and U48692 (N_48692,N_46432,N_45953);
nor U48693 (N_48693,N_45732,N_46710);
and U48694 (N_48694,N_46684,N_45588);
or U48695 (N_48695,N_47466,N_46966);
and U48696 (N_48696,N_45345,N_46810);
or U48697 (N_48697,N_46737,N_46728);
and U48698 (N_48698,N_46380,N_46030);
nand U48699 (N_48699,N_47223,N_46704);
nand U48700 (N_48700,N_45279,N_45604);
nor U48701 (N_48701,N_45865,N_45904);
nand U48702 (N_48702,N_46623,N_46032);
nand U48703 (N_48703,N_46270,N_46680);
nor U48704 (N_48704,N_46407,N_46942);
xor U48705 (N_48705,N_47019,N_47350);
and U48706 (N_48706,N_46151,N_46842);
and U48707 (N_48707,N_46960,N_46128);
and U48708 (N_48708,N_47334,N_47257);
nor U48709 (N_48709,N_47435,N_45843);
xor U48710 (N_48710,N_45563,N_45622);
nor U48711 (N_48711,N_46701,N_46512);
xnor U48712 (N_48712,N_46606,N_46377);
xor U48713 (N_48713,N_45754,N_45992);
and U48714 (N_48714,N_46880,N_45177);
xnor U48715 (N_48715,N_45713,N_45458);
and U48716 (N_48716,N_46986,N_45955);
nor U48717 (N_48717,N_46541,N_45999);
and U48718 (N_48718,N_47432,N_45716);
or U48719 (N_48719,N_46208,N_46405);
and U48720 (N_48720,N_46426,N_47348);
nor U48721 (N_48721,N_45542,N_45078);
xnor U48722 (N_48722,N_47444,N_46294);
nor U48723 (N_48723,N_46476,N_45483);
and U48724 (N_48724,N_45949,N_47327);
xor U48725 (N_48725,N_45300,N_46790);
or U48726 (N_48726,N_46776,N_45223);
and U48727 (N_48727,N_45995,N_47022);
nor U48728 (N_48728,N_46372,N_45708);
nor U48729 (N_48729,N_45165,N_47024);
or U48730 (N_48730,N_46621,N_46310);
and U48731 (N_48731,N_45128,N_46009);
xnor U48732 (N_48732,N_47066,N_46994);
nand U48733 (N_48733,N_45977,N_47488);
nor U48734 (N_48734,N_47363,N_45711);
nor U48735 (N_48735,N_46773,N_45637);
and U48736 (N_48736,N_46083,N_45489);
or U48737 (N_48737,N_45562,N_46253);
nor U48738 (N_48738,N_46145,N_47096);
or U48739 (N_48739,N_46263,N_47007);
and U48740 (N_48740,N_47213,N_45566);
nor U48741 (N_48741,N_45941,N_46999);
and U48742 (N_48742,N_47030,N_46852);
and U48743 (N_48743,N_45045,N_45404);
and U48744 (N_48744,N_45913,N_45153);
or U48745 (N_48745,N_47409,N_45211);
or U48746 (N_48746,N_45858,N_45981);
xor U48747 (N_48747,N_46859,N_46243);
nor U48748 (N_48748,N_45269,N_45213);
xnor U48749 (N_48749,N_45245,N_46716);
nand U48750 (N_48750,N_45630,N_46727);
or U48751 (N_48751,N_45352,N_46743);
xor U48752 (N_48752,N_45350,N_46044);
nand U48753 (N_48753,N_45922,N_46164);
or U48754 (N_48754,N_46596,N_45821);
nand U48755 (N_48755,N_45270,N_45106);
or U48756 (N_48756,N_45266,N_47473);
or U48757 (N_48757,N_46970,N_46762);
xnor U48758 (N_48758,N_47373,N_46658);
xor U48759 (N_48759,N_45964,N_45863);
nand U48760 (N_48760,N_45014,N_45737);
nand U48761 (N_48761,N_45571,N_45075);
xor U48762 (N_48762,N_45595,N_47011);
or U48763 (N_48763,N_45542,N_45275);
and U48764 (N_48764,N_46238,N_46458);
xnor U48765 (N_48765,N_45998,N_46080);
xnor U48766 (N_48766,N_45677,N_46569);
nor U48767 (N_48767,N_45324,N_46905);
and U48768 (N_48768,N_46527,N_46833);
nor U48769 (N_48769,N_46978,N_45629);
nand U48770 (N_48770,N_45941,N_45469);
and U48771 (N_48771,N_46472,N_45932);
and U48772 (N_48772,N_46481,N_45475);
nor U48773 (N_48773,N_45742,N_45675);
or U48774 (N_48774,N_45627,N_46912);
xor U48775 (N_48775,N_47207,N_45637);
nor U48776 (N_48776,N_46238,N_45435);
or U48777 (N_48777,N_47059,N_46241);
or U48778 (N_48778,N_45525,N_46443);
xnor U48779 (N_48779,N_45458,N_45452);
nand U48780 (N_48780,N_46135,N_46484);
nor U48781 (N_48781,N_47322,N_45563);
nand U48782 (N_48782,N_45345,N_46527);
nand U48783 (N_48783,N_46021,N_45307);
or U48784 (N_48784,N_45217,N_45009);
and U48785 (N_48785,N_47453,N_45154);
nand U48786 (N_48786,N_47258,N_45454);
and U48787 (N_48787,N_46754,N_45815);
nor U48788 (N_48788,N_46264,N_45506);
nor U48789 (N_48789,N_47095,N_45265);
nand U48790 (N_48790,N_45860,N_47256);
xor U48791 (N_48791,N_46603,N_45319);
nor U48792 (N_48792,N_46683,N_45768);
xor U48793 (N_48793,N_46255,N_47097);
or U48794 (N_48794,N_46657,N_45061);
xnor U48795 (N_48795,N_47397,N_45109);
nor U48796 (N_48796,N_47109,N_46445);
nand U48797 (N_48797,N_46025,N_45565);
xor U48798 (N_48798,N_45608,N_46954);
or U48799 (N_48799,N_45149,N_45674);
and U48800 (N_48800,N_45900,N_45807);
xnor U48801 (N_48801,N_46237,N_45469);
nor U48802 (N_48802,N_47328,N_47181);
nor U48803 (N_48803,N_45359,N_45713);
and U48804 (N_48804,N_46578,N_46481);
or U48805 (N_48805,N_45174,N_45518);
nand U48806 (N_48806,N_46781,N_46424);
or U48807 (N_48807,N_45677,N_47189);
nand U48808 (N_48808,N_45561,N_45825);
or U48809 (N_48809,N_46659,N_45867);
and U48810 (N_48810,N_45137,N_46142);
nand U48811 (N_48811,N_47304,N_47384);
xor U48812 (N_48812,N_45723,N_45417);
or U48813 (N_48813,N_46091,N_46421);
or U48814 (N_48814,N_45614,N_45023);
and U48815 (N_48815,N_46389,N_47255);
and U48816 (N_48816,N_47082,N_45928);
nand U48817 (N_48817,N_46943,N_47161);
and U48818 (N_48818,N_46511,N_45842);
or U48819 (N_48819,N_46491,N_45975);
xor U48820 (N_48820,N_45163,N_46211);
nor U48821 (N_48821,N_47361,N_46167);
xor U48822 (N_48822,N_45452,N_45528);
or U48823 (N_48823,N_47111,N_45401);
xor U48824 (N_48824,N_46436,N_47174);
nor U48825 (N_48825,N_46554,N_47138);
nand U48826 (N_48826,N_45737,N_46004);
xor U48827 (N_48827,N_45009,N_45934);
nor U48828 (N_48828,N_45879,N_46421);
nor U48829 (N_48829,N_47081,N_45368);
and U48830 (N_48830,N_46171,N_45795);
nor U48831 (N_48831,N_46279,N_46285);
nand U48832 (N_48832,N_45149,N_45379);
xnor U48833 (N_48833,N_47041,N_47119);
xor U48834 (N_48834,N_47091,N_46676);
nor U48835 (N_48835,N_47301,N_45144);
nand U48836 (N_48836,N_45794,N_45103);
xnor U48837 (N_48837,N_47210,N_46797);
and U48838 (N_48838,N_45987,N_45979);
or U48839 (N_48839,N_47349,N_45484);
or U48840 (N_48840,N_46865,N_46383);
nor U48841 (N_48841,N_46874,N_46737);
nor U48842 (N_48842,N_46379,N_46818);
and U48843 (N_48843,N_46281,N_46320);
and U48844 (N_48844,N_47366,N_47437);
or U48845 (N_48845,N_45868,N_46467);
or U48846 (N_48846,N_46229,N_45959);
nor U48847 (N_48847,N_45816,N_45460);
and U48848 (N_48848,N_46223,N_47444);
xnor U48849 (N_48849,N_47254,N_45488);
xnor U48850 (N_48850,N_46529,N_46051);
nand U48851 (N_48851,N_45647,N_45186);
nand U48852 (N_48852,N_45159,N_47354);
xor U48853 (N_48853,N_45499,N_46420);
or U48854 (N_48854,N_46547,N_46185);
nor U48855 (N_48855,N_46591,N_45158);
nor U48856 (N_48856,N_45180,N_46981);
and U48857 (N_48857,N_46375,N_46249);
or U48858 (N_48858,N_45628,N_47131);
nand U48859 (N_48859,N_45719,N_46282);
nor U48860 (N_48860,N_46111,N_45165);
xnor U48861 (N_48861,N_45709,N_46358);
nand U48862 (N_48862,N_46203,N_46052);
and U48863 (N_48863,N_47235,N_46995);
nand U48864 (N_48864,N_46488,N_46863);
or U48865 (N_48865,N_46431,N_45123);
nand U48866 (N_48866,N_45710,N_46242);
xnor U48867 (N_48867,N_46590,N_45648);
nand U48868 (N_48868,N_45317,N_47353);
nor U48869 (N_48869,N_47343,N_46612);
or U48870 (N_48870,N_47127,N_47063);
and U48871 (N_48871,N_47349,N_46434);
and U48872 (N_48872,N_46259,N_47024);
or U48873 (N_48873,N_46940,N_46412);
or U48874 (N_48874,N_46635,N_47412);
nor U48875 (N_48875,N_46321,N_45452);
and U48876 (N_48876,N_47257,N_46616);
nand U48877 (N_48877,N_46856,N_47011);
and U48878 (N_48878,N_46792,N_47124);
and U48879 (N_48879,N_45940,N_47273);
and U48880 (N_48880,N_46522,N_46515);
xnor U48881 (N_48881,N_45644,N_46425);
nand U48882 (N_48882,N_46303,N_45990);
or U48883 (N_48883,N_45953,N_46471);
nand U48884 (N_48884,N_46951,N_47294);
or U48885 (N_48885,N_45779,N_47453);
xor U48886 (N_48886,N_46440,N_46914);
or U48887 (N_48887,N_45037,N_45464);
nor U48888 (N_48888,N_46703,N_45363);
and U48889 (N_48889,N_45845,N_46012);
xnor U48890 (N_48890,N_46821,N_45963);
or U48891 (N_48891,N_46162,N_45403);
and U48892 (N_48892,N_46326,N_45563);
or U48893 (N_48893,N_46409,N_45887);
nor U48894 (N_48894,N_45360,N_47052);
nand U48895 (N_48895,N_45645,N_45737);
xnor U48896 (N_48896,N_47082,N_45201);
xnor U48897 (N_48897,N_47403,N_45673);
nor U48898 (N_48898,N_45468,N_45566);
xnor U48899 (N_48899,N_45099,N_46049);
and U48900 (N_48900,N_46793,N_45704);
or U48901 (N_48901,N_45404,N_45234);
nand U48902 (N_48902,N_45378,N_46732);
or U48903 (N_48903,N_46131,N_45327);
and U48904 (N_48904,N_46029,N_45440);
nor U48905 (N_48905,N_45196,N_46743);
or U48906 (N_48906,N_46153,N_45827);
or U48907 (N_48907,N_45522,N_45551);
and U48908 (N_48908,N_45594,N_45230);
xnor U48909 (N_48909,N_46068,N_45736);
and U48910 (N_48910,N_45804,N_46987);
and U48911 (N_48911,N_45767,N_45971);
or U48912 (N_48912,N_46179,N_46283);
nor U48913 (N_48913,N_46045,N_45971);
nand U48914 (N_48914,N_45776,N_46006);
or U48915 (N_48915,N_46720,N_46617);
nor U48916 (N_48916,N_45758,N_45848);
nand U48917 (N_48917,N_46151,N_46392);
and U48918 (N_48918,N_45939,N_46129);
or U48919 (N_48919,N_46275,N_47035);
nor U48920 (N_48920,N_46790,N_46098);
nor U48921 (N_48921,N_47040,N_45112);
and U48922 (N_48922,N_47481,N_45397);
xor U48923 (N_48923,N_46618,N_47271);
xnor U48924 (N_48924,N_45881,N_47385);
or U48925 (N_48925,N_46747,N_47222);
nor U48926 (N_48926,N_45662,N_45530);
and U48927 (N_48927,N_47201,N_46501);
nand U48928 (N_48928,N_46373,N_47299);
xor U48929 (N_48929,N_46952,N_46656);
nand U48930 (N_48930,N_47088,N_45607);
nand U48931 (N_48931,N_46272,N_45635);
nand U48932 (N_48932,N_47285,N_46141);
nand U48933 (N_48933,N_47328,N_46758);
and U48934 (N_48934,N_45244,N_46013);
xor U48935 (N_48935,N_45226,N_46990);
nor U48936 (N_48936,N_45406,N_47258);
nand U48937 (N_48937,N_47201,N_46265);
nand U48938 (N_48938,N_45870,N_45993);
nor U48939 (N_48939,N_45363,N_45922);
and U48940 (N_48940,N_47366,N_45689);
xnor U48941 (N_48941,N_47459,N_45581);
xor U48942 (N_48942,N_47214,N_45183);
nor U48943 (N_48943,N_46929,N_45740);
or U48944 (N_48944,N_45844,N_45157);
nand U48945 (N_48945,N_47332,N_47198);
and U48946 (N_48946,N_45890,N_45297);
nand U48947 (N_48947,N_47395,N_46331);
xnor U48948 (N_48948,N_47351,N_46170);
and U48949 (N_48949,N_45915,N_45220);
nand U48950 (N_48950,N_45274,N_47385);
nor U48951 (N_48951,N_46460,N_46944);
and U48952 (N_48952,N_45927,N_45492);
and U48953 (N_48953,N_45000,N_46945);
nor U48954 (N_48954,N_45132,N_46130);
xnor U48955 (N_48955,N_45276,N_45615);
and U48956 (N_48956,N_46860,N_46169);
or U48957 (N_48957,N_45439,N_46752);
nand U48958 (N_48958,N_46027,N_46936);
nor U48959 (N_48959,N_46131,N_45749);
nand U48960 (N_48960,N_46080,N_45343);
and U48961 (N_48961,N_46568,N_45294);
and U48962 (N_48962,N_46714,N_47354);
nand U48963 (N_48963,N_46358,N_47007);
or U48964 (N_48964,N_46648,N_45350);
nand U48965 (N_48965,N_47005,N_46725);
and U48966 (N_48966,N_46434,N_45054);
xnor U48967 (N_48967,N_47451,N_45300);
xor U48968 (N_48968,N_46533,N_46627);
nor U48969 (N_48969,N_45437,N_47091);
or U48970 (N_48970,N_46491,N_47155);
nand U48971 (N_48971,N_46188,N_45718);
xnor U48972 (N_48972,N_46857,N_45972);
and U48973 (N_48973,N_46780,N_46704);
nand U48974 (N_48974,N_46964,N_45496);
nand U48975 (N_48975,N_46816,N_46302);
or U48976 (N_48976,N_46032,N_47452);
xnor U48977 (N_48977,N_45179,N_47448);
and U48978 (N_48978,N_47179,N_47173);
nor U48979 (N_48979,N_46489,N_45898);
or U48980 (N_48980,N_46069,N_45206);
nand U48981 (N_48981,N_45925,N_45757);
nor U48982 (N_48982,N_46602,N_45536);
nor U48983 (N_48983,N_45907,N_47176);
nor U48984 (N_48984,N_45308,N_47040);
xnor U48985 (N_48985,N_46093,N_45376);
nand U48986 (N_48986,N_47191,N_46887);
or U48987 (N_48987,N_45317,N_46994);
nor U48988 (N_48988,N_47438,N_46457);
xor U48989 (N_48989,N_46328,N_47310);
and U48990 (N_48990,N_46461,N_45435);
and U48991 (N_48991,N_46793,N_46975);
or U48992 (N_48992,N_46551,N_45456);
xor U48993 (N_48993,N_46368,N_45258);
or U48994 (N_48994,N_45378,N_45995);
xor U48995 (N_48995,N_46473,N_45813);
nor U48996 (N_48996,N_45393,N_45268);
or U48997 (N_48997,N_47068,N_47466);
nor U48998 (N_48998,N_45001,N_45550);
xnor U48999 (N_48999,N_45870,N_46458);
nor U49000 (N_49000,N_45652,N_45968);
nand U49001 (N_49001,N_45051,N_46387);
nor U49002 (N_49002,N_45820,N_45299);
nand U49003 (N_49003,N_45311,N_45194);
nand U49004 (N_49004,N_46350,N_45222);
nand U49005 (N_49005,N_46877,N_46992);
nand U49006 (N_49006,N_45845,N_47383);
xor U49007 (N_49007,N_46911,N_45111);
or U49008 (N_49008,N_47181,N_45989);
xnor U49009 (N_49009,N_45010,N_47167);
or U49010 (N_49010,N_46689,N_47428);
nand U49011 (N_49011,N_46146,N_46740);
xnor U49012 (N_49012,N_46247,N_47427);
xor U49013 (N_49013,N_47392,N_45588);
or U49014 (N_49014,N_45445,N_45269);
and U49015 (N_49015,N_45817,N_47164);
nand U49016 (N_49016,N_45864,N_46432);
nor U49017 (N_49017,N_45856,N_46076);
and U49018 (N_49018,N_46753,N_46741);
or U49019 (N_49019,N_46917,N_45361);
or U49020 (N_49020,N_46810,N_45716);
nor U49021 (N_49021,N_46676,N_46847);
xnor U49022 (N_49022,N_47060,N_45815);
or U49023 (N_49023,N_47450,N_46120);
nor U49024 (N_49024,N_46499,N_46707);
or U49025 (N_49025,N_46283,N_45513);
xnor U49026 (N_49026,N_45565,N_47141);
or U49027 (N_49027,N_45886,N_47228);
and U49028 (N_49028,N_45340,N_45870);
nor U49029 (N_49029,N_45714,N_46495);
xor U49030 (N_49030,N_46125,N_45000);
xor U49031 (N_49031,N_47085,N_45342);
xnor U49032 (N_49032,N_46724,N_45068);
nand U49033 (N_49033,N_47364,N_46341);
xnor U49034 (N_49034,N_46735,N_46964);
nor U49035 (N_49035,N_47445,N_47278);
nand U49036 (N_49036,N_45442,N_46947);
xnor U49037 (N_49037,N_47486,N_47497);
xor U49038 (N_49038,N_47411,N_45071);
and U49039 (N_49039,N_47318,N_46774);
and U49040 (N_49040,N_47411,N_45673);
nor U49041 (N_49041,N_45137,N_46389);
nor U49042 (N_49042,N_45908,N_46031);
nor U49043 (N_49043,N_46136,N_45354);
nand U49044 (N_49044,N_45160,N_47246);
and U49045 (N_49045,N_46275,N_47125);
and U49046 (N_49046,N_46698,N_45111);
xor U49047 (N_49047,N_46792,N_46185);
nor U49048 (N_49048,N_45976,N_46786);
nand U49049 (N_49049,N_47192,N_45312);
nand U49050 (N_49050,N_46489,N_46125);
nor U49051 (N_49051,N_47498,N_46228);
and U49052 (N_49052,N_47441,N_46725);
xor U49053 (N_49053,N_45289,N_45405);
nand U49054 (N_49054,N_47088,N_46888);
or U49055 (N_49055,N_46869,N_46711);
nand U49056 (N_49056,N_45525,N_45137);
nand U49057 (N_49057,N_46153,N_46902);
nand U49058 (N_49058,N_45850,N_45222);
xnor U49059 (N_49059,N_46269,N_45071);
and U49060 (N_49060,N_45974,N_45970);
xnor U49061 (N_49061,N_46129,N_47346);
xor U49062 (N_49062,N_46976,N_45568);
or U49063 (N_49063,N_46555,N_45194);
nor U49064 (N_49064,N_46556,N_45732);
xnor U49065 (N_49065,N_46250,N_46934);
and U49066 (N_49066,N_45843,N_46263);
nand U49067 (N_49067,N_45532,N_47469);
and U49068 (N_49068,N_46705,N_45939);
and U49069 (N_49069,N_45672,N_46598);
nor U49070 (N_49070,N_46467,N_46724);
and U49071 (N_49071,N_45417,N_45231);
xor U49072 (N_49072,N_45700,N_46120);
xnor U49073 (N_49073,N_46359,N_47125);
nor U49074 (N_49074,N_45216,N_46137);
nand U49075 (N_49075,N_46906,N_45728);
and U49076 (N_49076,N_47125,N_47002);
xnor U49077 (N_49077,N_46288,N_45446);
and U49078 (N_49078,N_45190,N_45767);
nand U49079 (N_49079,N_45952,N_45903);
nor U49080 (N_49080,N_45852,N_47213);
nand U49081 (N_49081,N_46095,N_47482);
or U49082 (N_49082,N_46294,N_46886);
nand U49083 (N_49083,N_45290,N_46017);
and U49084 (N_49084,N_45515,N_45111);
xnor U49085 (N_49085,N_45701,N_47364);
or U49086 (N_49086,N_45677,N_45245);
and U49087 (N_49087,N_45499,N_45193);
nor U49088 (N_49088,N_46512,N_45090);
nand U49089 (N_49089,N_45406,N_47254);
nor U49090 (N_49090,N_47248,N_45124);
xnor U49091 (N_49091,N_47226,N_45365);
nand U49092 (N_49092,N_47160,N_45763);
nor U49093 (N_49093,N_46212,N_46388);
or U49094 (N_49094,N_46571,N_47184);
nor U49095 (N_49095,N_46058,N_45285);
and U49096 (N_49096,N_47185,N_46722);
nand U49097 (N_49097,N_46207,N_46206);
nand U49098 (N_49098,N_45032,N_46860);
xnor U49099 (N_49099,N_45990,N_45938);
nor U49100 (N_49100,N_46597,N_45764);
nor U49101 (N_49101,N_47147,N_45038);
or U49102 (N_49102,N_45771,N_45866);
xor U49103 (N_49103,N_47205,N_45555);
xnor U49104 (N_49104,N_46543,N_46222);
nor U49105 (N_49105,N_46079,N_46035);
nor U49106 (N_49106,N_46977,N_45373);
and U49107 (N_49107,N_46418,N_47052);
and U49108 (N_49108,N_47196,N_46023);
nor U49109 (N_49109,N_47131,N_47178);
or U49110 (N_49110,N_47431,N_45326);
xor U49111 (N_49111,N_46998,N_47165);
nor U49112 (N_49112,N_46174,N_45883);
nor U49113 (N_49113,N_46834,N_46428);
nor U49114 (N_49114,N_45565,N_45392);
xnor U49115 (N_49115,N_45081,N_46001);
nor U49116 (N_49116,N_46487,N_45592);
and U49117 (N_49117,N_47188,N_46978);
and U49118 (N_49118,N_46931,N_45659);
xor U49119 (N_49119,N_45240,N_45724);
nand U49120 (N_49120,N_45942,N_47220);
or U49121 (N_49121,N_45145,N_47228);
and U49122 (N_49122,N_46836,N_46339);
nor U49123 (N_49123,N_45173,N_45998);
or U49124 (N_49124,N_46653,N_47284);
and U49125 (N_49125,N_46501,N_47040);
nor U49126 (N_49126,N_46846,N_47049);
and U49127 (N_49127,N_45923,N_46727);
and U49128 (N_49128,N_45537,N_45696);
or U49129 (N_49129,N_47254,N_47473);
or U49130 (N_49130,N_45355,N_46974);
xor U49131 (N_49131,N_45029,N_46084);
xnor U49132 (N_49132,N_46991,N_46953);
or U49133 (N_49133,N_45714,N_45984);
or U49134 (N_49134,N_46907,N_46313);
nand U49135 (N_49135,N_46565,N_46960);
or U49136 (N_49136,N_46369,N_46720);
and U49137 (N_49137,N_46763,N_45229);
nand U49138 (N_49138,N_45438,N_47239);
or U49139 (N_49139,N_46027,N_46885);
xor U49140 (N_49140,N_46630,N_47002);
nor U49141 (N_49141,N_46343,N_47303);
and U49142 (N_49142,N_45341,N_46097);
xor U49143 (N_49143,N_46345,N_46552);
and U49144 (N_49144,N_47287,N_46867);
xnor U49145 (N_49145,N_45673,N_47016);
or U49146 (N_49146,N_45003,N_45369);
or U49147 (N_49147,N_47000,N_45971);
nand U49148 (N_49148,N_46625,N_45421);
or U49149 (N_49149,N_46013,N_45675);
xor U49150 (N_49150,N_45747,N_46965);
nor U49151 (N_49151,N_46108,N_46971);
xor U49152 (N_49152,N_46430,N_45784);
xnor U49153 (N_49153,N_46225,N_45516);
or U49154 (N_49154,N_45591,N_46064);
and U49155 (N_49155,N_46510,N_47008);
xor U49156 (N_49156,N_47033,N_46947);
xor U49157 (N_49157,N_46351,N_45625);
nand U49158 (N_49158,N_46194,N_45235);
nor U49159 (N_49159,N_46249,N_45639);
or U49160 (N_49160,N_45416,N_46873);
or U49161 (N_49161,N_46293,N_46678);
or U49162 (N_49162,N_47265,N_46651);
xnor U49163 (N_49163,N_46723,N_46797);
or U49164 (N_49164,N_45716,N_46805);
nor U49165 (N_49165,N_45488,N_45165);
and U49166 (N_49166,N_45549,N_46155);
nor U49167 (N_49167,N_47446,N_45273);
xor U49168 (N_49168,N_45916,N_45780);
or U49169 (N_49169,N_45808,N_45661);
nor U49170 (N_49170,N_46860,N_47406);
nor U49171 (N_49171,N_45619,N_46208);
and U49172 (N_49172,N_47137,N_47402);
or U49173 (N_49173,N_46169,N_46808);
nor U49174 (N_49174,N_47028,N_46640);
nand U49175 (N_49175,N_45022,N_47195);
or U49176 (N_49176,N_47226,N_46816);
xor U49177 (N_49177,N_45861,N_47483);
or U49178 (N_49178,N_45528,N_45664);
nor U49179 (N_49179,N_45435,N_45473);
nor U49180 (N_49180,N_47367,N_46451);
or U49181 (N_49181,N_46726,N_45688);
xnor U49182 (N_49182,N_45683,N_47245);
xnor U49183 (N_49183,N_46766,N_45963);
xnor U49184 (N_49184,N_45790,N_45040);
nor U49185 (N_49185,N_47114,N_45635);
xor U49186 (N_49186,N_46612,N_46020);
xnor U49187 (N_49187,N_46634,N_46415);
xnor U49188 (N_49188,N_46797,N_47457);
and U49189 (N_49189,N_45759,N_46658);
or U49190 (N_49190,N_45855,N_47290);
or U49191 (N_49191,N_46228,N_45490);
and U49192 (N_49192,N_45302,N_45780);
and U49193 (N_49193,N_46353,N_47388);
nor U49194 (N_49194,N_46714,N_47378);
nand U49195 (N_49195,N_46753,N_46401);
nand U49196 (N_49196,N_47260,N_46531);
nor U49197 (N_49197,N_46029,N_46581);
nor U49198 (N_49198,N_45019,N_45865);
xor U49199 (N_49199,N_45316,N_46285);
and U49200 (N_49200,N_45619,N_46964);
nand U49201 (N_49201,N_46121,N_45981);
or U49202 (N_49202,N_45610,N_45723);
or U49203 (N_49203,N_47005,N_47349);
or U49204 (N_49204,N_45432,N_45241);
nor U49205 (N_49205,N_45538,N_45542);
nor U49206 (N_49206,N_46711,N_45302);
nand U49207 (N_49207,N_47493,N_47175);
nand U49208 (N_49208,N_45367,N_45930);
nor U49209 (N_49209,N_46690,N_45722);
nand U49210 (N_49210,N_45132,N_47249);
nor U49211 (N_49211,N_47138,N_45545);
xnor U49212 (N_49212,N_45085,N_45916);
nand U49213 (N_49213,N_46684,N_47354);
xnor U49214 (N_49214,N_46267,N_45158);
or U49215 (N_49215,N_46901,N_46336);
or U49216 (N_49216,N_47479,N_45212);
nand U49217 (N_49217,N_46577,N_45123);
nand U49218 (N_49218,N_45913,N_45768);
nor U49219 (N_49219,N_45921,N_47217);
xor U49220 (N_49220,N_47485,N_46658);
nor U49221 (N_49221,N_46965,N_46494);
and U49222 (N_49222,N_45420,N_45439);
and U49223 (N_49223,N_46506,N_47133);
or U49224 (N_49224,N_47117,N_46454);
xnor U49225 (N_49225,N_46237,N_45329);
and U49226 (N_49226,N_47195,N_46767);
xnor U49227 (N_49227,N_45321,N_46296);
or U49228 (N_49228,N_46585,N_46402);
nand U49229 (N_49229,N_46221,N_47042);
nor U49230 (N_49230,N_45518,N_46494);
and U49231 (N_49231,N_45378,N_45259);
and U49232 (N_49232,N_46718,N_46706);
and U49233 (N_49233,N_45803,N_47395);
nor U49234 (N_49234,N_46374,N_45291);
xnor U49235 (N_49235,N_45377,N_47162);
nor U49236 (N_49236,N_46892,N_45968);
and U49237 (N_49237,N_47208,N_46936);
or U49238 (N_49238,N_45219,N_45195);
and U49239 (N_49239,N_46831,N_46100);
or U49240 (N_49240,N_47397,N_45191);
nand U49241 (N_49241,N_45479,N_46571);
nor U49242 (N_49242,N_47152,N_46352);
xnor U49243 (N_49243,N_45992,N_46937);
xnor U49244 (N_49244,N_46041,N_46345);
nor U49245 (N_49245,N_46791,N_45589);
and U49246 (N_49246,N_45158,N_46397);
xnor U49247 (N_49247,N_46808,N_46089);
nor U49248 (N_49248,N_46828,N_46816);
xnor U49249 (N_49249,N_45096,N_46776);
or U49250 (N_49250,N_45611,N_45534);
xnor U49251 (N_49251,N_45062,N_46886);
nand U49252 (N_49252,N_45017,N_47380);
xor U49253 (N_49253,N_47370,N_45581);
xnor U49254 (N_49254,N_46588,N_46067);
or U49255 (N_49255,N_46908,N_46993);
xor U49256 (N_49256,N_45785,N_46919);
nand U49257 (N_49257,N_46504,N_46567);
nand U49258 (N_49258,N_46321,N_45222);
xor U49259 (N_49259,N_46441,N_45862);
or U49260 (N_49260,N_47064,N_45652);
and U49261 (N_49261,N_45256,N_45584);
and U49262 (N_49262,N_46426,N_46672);
and U49263 (N_49263,N_45603,N_46667);
or U49264 (N_49264,N_46016,N_46051);
nand U49265 (N_49265,N_47395,N_45751);
nand U49266 (N_49266,N_46656,N_47006);
xor U49267 (N_49267,N_46657,N_45470);
nand U49268 (N_49268,N_46840,N_45939);
xnor U49269 (N_49269,N_46961,N_46998);
xor U49270 (N_49270,N_46354,N_47275);
xnor U49271 (N_49271,N_45941,N_46587);
and U49272 (N_49272,N_45836,N_47193);
xnor U49273 (N_49273,N_46400,N_46620);
and U49274 (N_49274,N_47141,N_45033);
or U49275 (N_49275,N_45362,N_46368);
nand U49276 (N_49276,N_47200,N_47196);
nand U49277 (N_49277,N_46781,N_46710);
and U49278 (N_49278,N_45788,N_47397);
or U49279 (N_49279,N_46784,N_45444);
nand U49280 (N_49280,N_46153,N_45459);
and U49281 (N_49281,N_45681,N_46287);
xor U49282 (N_49282,N_46993,N_46727);
xnor U49283 (N_49283,N_47166,N_45855);
xnor U49284 (N_49284,N_45586,N_46139);
and U49285 (N_49285,N_45490,N_45012);
and U49286 (N_49286,N_45786,N_46009);
nand U49287 (N_49287,N_47450,N_47461);
xnor U49288 (N_49288,N_45585,N_45666);
or U49289 (N_49289,N_45906,N_47014);
xnor U49290 (N_49290,N_46848,N_45321);
xor U49291 (N_49291,N_45446,N_46744);
nor U49292 (N_49292,N_46551,N_47435);
nand U49293 (N_49293,N_47301,N_47263);
and U49294 (N_49294,N_46986,N_46558);
xnor U49295 (N_49295,N_46208,N_46878);
and U49296 (N_49296,N_45601,N_46361);
and U49297 (N_49297,N_45149,N_46538);
or U49298 (N_49298,N_46046,N_45961);
nand U49299 (N_49299,N_45199,N_46890);
nor U49300 (N_49300,N_45059,N_45602);
or U49301 (N_49301,N_45425,N_45406);
and U49302 (N_49302,N_46024,N_46193);
nor U49303 (N_49303,N_45536,N_47115);
or U49304 (N_49304,N_45507,N_47427);
or U49305 (N_49305,N_45087,N_46772);
nand U49306 (N_49306,N_45595,N_45597);
xnor U49307 (N_49307,N_45169,N_47082);
and U49308 (N_49308,N_45626,N_47255);
nor U49309 (N_49309,N_46422,N_45210);
or U49310 (N_49310,N_45889,N_45738);
and U49311 (N_49311,N_45871,N_47150);
or U49312 (N_49312,N_47192,N_46423);
or U49313 (N_49313,N_45271,N_47011);
nor U49314 (N_49314,N_46637,N_46213);
or U49315 (N_49315,N_47415,N_46933);
xnor U49316 (N_49316,N_45297,N_45588);
and U49317 (N_49317,N_45575,N_46280);
xor U49318 (N_49318,N_45229,N_45685);
or U49319 (N_49319,N_45971,N_46481);
or U49320 (N_49320,N_46958,N_47489);
xnor U49321 (N_49321,N_47082,N_45657);
nand U49322 (N_49322,N_46398,N_47047);
and U49323 (N_49323,N_46516,N_47109);
or U49324 (N_49324,N_45095,N_46497);
nor U49325 (N_49325,N_47067,N_46854);
nor U49326 (N_49326,N_47039,N_47061);
nand U49327 (N_49327,N_46530,N_45545);
nor U49328 (N_49328,N_45016,N_45593);
nand U49329 (N_49329,N_46605,N_45148);
xnor U49330 (N_49330,N_45381,N_47419);
or U49331 (N_49331,N_46467,N_45170);
nor U49332 (N_49332,N_46129,N_46869);
or U49333 (N_49333,N_46587,N_46207);
and U49334 (N_49334,N_46450,N_45311);
xor U49335 (N_49335,N_45199,N_46474);
or U49336 (N_49336,N_47246,N_46264);
or U49337 (N_49337,N_45106,N_46492);
xor U49338 (N_49338,N_45039,N_45736);
nand U49339 (N_49339,N_45316,N_47326);
and U49340 (N_49340,N_47086,N_46664);
nor U49341 (N_49341,N_45855,N_47480);
nor U49342 (N_49342,N_46022,N_46203);
and U49343 (N_49343,N_46803,N_46233);
nor U49344 (N_49344,N_46480,N_45637);
xnor U49345 (N_49345,N_46332,N_46019);
or U49346 (N_49346,N_46014,N_46025);
or U49347 (N_49347,N_47118,N_46117);
xnor U49348 (N_49348,N_45644,N_46510);
nand U49349 (N_49349,N_46565,N_45859);
nand U49350 (N_49350,N_46272,N_47468);
xor U49351 (N_49351,N_45516,N_46028);
xor U49352 (N_49352,N_46974,N_46921);
xor U49353 (N_49353,N_45932,N_45314);
or U49354 (N_49354,N_46933,N_45805);
nor U49355 (N_49355,N_47084,N_46794);
nor U49356 (N_49356,N_45193,N_45304);
nand U49357 (N_49357,N_46693,N_46266);
and U49358 (N_49358,N_45679,N_46874);
and U49359 (N_49359,N_47063,N_46722);
or U49360 (N_49360,N_46791,N_45484);
and U49361 (N_49361,N_45767,N_45377);
and U49362 (N_49362,N_46760,N_47116);
nor U49363 (N_49363,N_47331,N_47386);
and U49364 (N_49364,N_47014,N_45379);
nand U49365 (N_49365,N_46130,N_46907);
and U49366 (N_49366,N_45288,N_47301);
and U49367 (N_49367,N_45771,N_47079);
or U49368 (N_49368,N_45103,N_45382);
or U49369 (N_49369,N_45915,N_46315);
xnor U49370 (N_49370,N_47263,N_46329);
or U49371 (N_49371,N_45726,N_47458);
and U49372 (N_49372,N_47368,N_46905);
or U49373 (N_49373,N_46312,N_45744);
and U49374 (N_49374,N_45904,N_46337);
xnor U49375 (N_49375,N_45675,N_46199);
and U49376 (N_49376,N_47422,N_45274);
nor U49377 (N_49377,N_47161,N_45564);
xnor U49378 (N_49378,N_46736,N_46795);
and U49379 (N_49379,N_45820,N_46993);
nor U49380 (N_49380,N_45513,N_46581);
xor U49381 (N_49381,N_46853,N_45508);
nand U49382 (N_49382,N_46203,N_46210);
nand U49383 (N_49383,N_46137,N_45539);
or U49384 (N_49384,N_45647,N_46842);
nand U49385 (N_49385,N_47135,N_46998);
nor U49386 (N_49386,N_46065,N_46661);
nor U49387 (N_49387,N_47219,N_45578);
xor U49388 (N_49388,N_47024,N_45642);
xor U49389 (N_49389,N_45085,N_46320);
and U49390 (N_49390,N_45892,N_45335);
nand U49391 (N_49391,N_45404,N_45140);
or U49392 (N_49392,N_46248,N_45036);
or U49393 (N_49393,N_45976,N_45657);
xor U49394 (N_49394,N_45993,N_45415);
or U49395 (N_49395,N_45386,N_45569);
nor U49396 (N_49396,N_45537,N_45151);
nand U49397 (N_49397,N_45400,N_45845);
nor U49398 (N_49398,N_46763,N_46268);
or U49399 (N_49399,N_45838,N_45246);
nand U49400 (N_49400,N_46685,N_45070);
xnor U49401 (N_49401,N_45247,N_45194);
and U49402 (N_49402,N_46162,N_45234);
xor U49403 (N_49403,N_47110,N_45554);
and U49404 (N_49404,N_45797,N_46944);
xnor U49405 (N_49405,N_46473,N_46874);
nor U49406 (N_49406,N_45190,N_46539);
nand U49407 (N_49407,N_47161,N_47277);
and U49408 (N_49408,N_46790,N_45291);
or U49409 (N_49409,N_46149,N_45629);
nand U49410 (N_49410,N_46730,N_45897);
nand U49411 (N_49411,N_47429,N_45374);
or U49412 (N_49412,N_47256,N_46753);
and U49413 (N_49413,N_45219,N_45053);
nand U49414 (N_49414,N_47355,N_47175);
nor U49415 (N_49415,N_45605,N_47243);
xor U49416 (N_49416,N_45775,N_45966);
nor U49417 (N_49417,N_46786,N_45831);
and U49418 (N_49418,N_47132,N_46369);
nand U49419 (N_49419,N_47402,N_46219);
xnor U49420 (N_49420,N_45034,N_45533);
nor U49421 (N_49421,N_45124,N_45030);
or U49422 (N_49422,N_45291,N_46070);
and U49423 (N_49423,N_46909,N_45719);
nand U49424 (N_49424,N_46832,N_45248);
or U49425 (N_49425,N_46701,N_45967);
xor U49426 (N_49426,N_46751,N_45939);
or U49427 (N_49427,N_47022,N_45354);
and U49428 (N_49428,N_46111,N_45886);
or U49429 (N_49429,N_46840,N_45193);
nand U49430 (N_49430,N_45786,N_46363);
nor U49431 (N_49431,N_45315,N_46151);
and U49432 (N_49432,N_45412,N_45768);
nand U49433 (N_49433,N_45736,N_46371);
and U49434 (N_49434,N_46886,N_46659);
and U49435 (N_49435,N_46944,N_45960);
xor U49436 (N_49436,N_45032,N_45741);
nor U49437 (N_49437,N_46054,N_46060);
nand U49438 (N_49438,N_46807,N_46149);
nand U49439 (N_49439,N_45461,N_45883);
nand U49440 (N_49440,N_47128,N_46021);
nor U49441 (N_49441,N_45699,N_46291);
and U49442 (N_49442,N_46570,N_47423);
xor U49443 (N_49443,N_45611,N_46503);
nand U49444 (N_49444,N_45831,N_46550);
nand U49445 (N_49445,N_45564,N_46390);
nor U49446 (N_49446,N_47386,N_45464);
nand U49447 (N_49447,N_46571,N_45376);
and U49448 (N_49448,N_46179,N_45606);
nand U49449 (N_49449,N_47174,N_47240);
and U49450 (N_49450,N_46746,N_45140);
and U49451 (N_49451,N_46913,N_45237);
and U49452 (N_49452,N_46182,N_46895);
nor U49453 (N_49453,N_46292,N_47306);
or U49454 (N_49454,N_45578,N_47055);
nor U49455 (N_49455,N_45074,N_46016);
and U49456 (N_49456,N_46560,N_45694);
or U49457 (N_49457,N_45836,N_46168);
nor U49458 (N_49458,N_45977,N_46372);
nand U49459 (N_49459,N_45568,N_46052);
and U49460 (N_49460,N_45435,N_47465);
or U49461 (N_49461,N_47159,N_45435);
xnor U49462 (N_49462,N_45277,N_47352);
nor U49463 (N_49463,N_45145,N_45065);
nor U49464 (N_49464,N_46447,N_47165);
or U49465 (N_49465,N_47482,N_45238);
nor U49466 (N_49466,N_46573,N_47160);
nand U49467 (N_49467,N_47437,N_45352);
or U49468 (N_49468,N_45457,N_46216);
and U49469 (N_49469,N_47224,N_46966);
or U49470 (N_49470,N_47075,N_45931);
xnor U49471 (N_49471,N_45459,N_46082);
nor U49472 (N_49472,N_45425,N_46856);
nor U49473 (N_49473,N_45620,N_46916);
and U49474 (N_49474,N_45460,N_45168);
or U49475 (N_49475,N_47301,N_45700);
or U49476 (N_49476,N_45710,N_45056);
nand U49477 (N_49477,N_45793,N_45384);
nor U49478 (N_49478,N_47477,N_47105);
or U49479 (N_49479,N_46268,N_46092);
xor U49480 (N_49480,N_45523,N_45731);
nand U49481 (N_49481,N_46800,N_45320);
nor U49482 (N_49482,N_45733,N_47227);
or U49483 (N_49483,N_47216,N_46359);
xnor U49484 (N_49484,N_45084,N_47021);
or U49485 (N_49485,N_46349,N_46743);
or U49486 (N_49486,N_46934,N_47281);
nand U49487 (N_49487,N_45614,N_46396);
nand U49488 (N_49488,N_46167,N_45824);
nand U49489 (N_49489,N_45010,N_45114);
xnor U49490 (N_49490,N_45563,N_46285);
nor U49491 (N_49491,N_46577,N_46615);
or U49492 (N_49492,N_45417,N_46604);
xor U49493 (N_49493,N_47411,N_45699);
nand U49494 (N_49494,N_47387,N_45113);
or U49495 (N_49495,N_46744,N_45532);
nor U49496 (N_49496,N_45014,N_46757);
or U49497 (N_49497,N_45613,N_45652);
or U49498 (N_49498,N_45075,N_47392);
or U49499 (N_49499,N_47205,N_46618);
xor U49500 (N_49500,N_45332,N_46236);
and U49501 (N_49501,N_45823,N_45054);
xnor U49502 (N_49502,N_46481,N_45521);
xnor U49503 (N_49503,N_46347,N_46721);
nand U49504 (N_49504,N_46747,N_45752);
nor U49505 (N_49505,N_46099,N_45208);
nand U49506 (N_49506,N_45657,N_45826);
xor U49507 (N_49507,N_46361,N_46749);
and U49508 (N_49508,N_45388,N_47367);
or U49509 (N_49509,N_45072,N_46899);
xor U49510 (N_49510,N_45513,N_45257);
and U49511 (N_49511,N_46887,N_45619);
or U49512 (N_49512,N_46168,N_45362);
or U49513 (N_49513,N_45144,N_45596);
nand U49514 (N_49514,N_45369,N_46301);
xnor U49515 (N_49515,N_46869,N_46045);
nor U49516 (N_49516,N_46868,N_45778);
nor U49517 (N_49517,N_46856,N_46566);
nand U49518 (N_49518,N_46436,N_45648);
nand U49519 (N_49519,N_46495,N_46334);
nor U49520 (N_49520,N_45947,N_46445);
or U49521 (N_49521,N_47364,N_47190);
nor U49522 (N_49522,N_47132,N_47008);
and U49523 (N_49523,N_45930,N_46204);
nand U49524 (N_49524,N_45769,N_45879);
nor U49525 (N_49525,N_46383,N_46133);
and U49526 (N_49526,N_46680,N_46305);
nand U49527 (N_49527,N_45364,N_45913);
nand U49528 (N_49528,N_47066,N_46361);
and U49529 (N_49529,N_46896,N_46499);
xnor U49530 (N_49530,N_47300,N_45061);
and U49531 (N_49531,N_45901,N_46131);
and U49532 (N_49532,N_45563,N_46558);
xnor U49533 (N_49533,N_45045,N_46642);
nor U49534 (N_49534,N_47161,N_47187);
nand U49535 (N_49535,N_45321,N_45372);
nand U49536 (N_49536,N_46956,N_46255);
nand U49537 (N_49537,N_47007,N_46617);
and U49538 (N_49538,N_46258,N_45866);
and U49539 (N_49539,N_47403,N_46110);
and U49540 (N_49540,N_45438,N_45152);
xor U49541 (N_49541,N_45778,N_46783);
nand U49542 (N_49542,N_46970,N_45969);
nand U49543 (N_49543,N_47286,N_46507);
or U49544 (N_49544,N_47465,N_47133);
xor U49545 (N_49545,N_46283,N_46756);
and U49546 (N_49546,N_46621,N_46036);
xnor U49547 (N_49547,N_47412,N_47405);
xnor U49548 (N_49548,N_46442,N_47448);
and U49549 (N_49549,N_46625,N_46134);
nand U49550 (N_49550,N_46382,N_46885);
nand U49551 (N_49551,N_45395,N_45819);
or U49552 (N_49552,N_46619,N_46728);
xor U49553 (N_49553,N_45307,N_45048);
nand U49554 (N_49554,N_47436,N_47416);
xor U49555 (N_49555,N_45707,N_45536);
or U49556 (N_49556,N_46077,N_45369);
xnor U49557 (N_49557,N_46730,N_47299);
xor U49558 (N_49558,N_47348,N_45739);
xnor U49559 (N_49559,N_45566,N_45726);
nand U49560 (N_49560,N_46560,N_46586);
nand U49561 (N_49561,N_45253,N_47212);
xor U49562 (N_49562,N_46919,N_45584);
or U49563 (N_49563,N_46796,N_47202);
or U49564 (N_49564,N_46318,N_46321);
nand U49565 (N_49565,N_46450,N_46886);
and U49566 (N_49566,N_47424,N_46480);
or U49567 (N_49567,N_47284,N_46133);
or U49568 (N_49568,N_45018,N_45325);
and U49569 (N_49569,N_45068,N_45985);
or U49570 (N_49570,N_47249,N_46613);
xor U49571 (N_49571,N_46366,N_45233);
nor U49572 (N_49572,N_47060,N_45153);
nor U49573 (N_49573,N_46471,N_46937);
and U49574 (N_49574,N_45099,N_46312);
or U49575 (N_49575,N_47314,N_46295);
or U49576 (N_49576,N_46298,N_46828);
nand U49577 (N_49577,N_45649,N_45986);
nand U49578 (N_49578,N_45643,N_45239);
xnor U49579 (N_49579,N_45915,N_45948);
or U49580 (N_49580,N_47192,N_45621);
nor U49581 (N_49581,N_46811,N_45297);
xor U49582 (N_49582,N_46436,N_47031);
xor U49583 (N_49583,N_46150,N_46613);
and U49584 (N_49584,N_46713,N_46141);
nor U49585 (N_49585,N_45582,N_46542);
nand U49586 (N_49586,N_47214,N_46079);
nand U49587 (N_49587,N_45426,N_47298);
or U49588 (N_49588,N_47139,N_45559);
nor U49589 (N_49589,N_46487,N_45085);
and U49590 (N_49590,N_45323,N_46944);
or U49591 (N_49591,N_45784,N_46836);
or U49592 (N_49592,N_46920,N_45354);
nor U49593 (N_49593,N_46243,N_46791);
xnor U49594 (N_49594,N_45199,N_46107);
nand U49595 (N_49595,N_46318,N_47441);
and U49596 (N_49596,N_47485,N_47328);
and U49597 (N_49597,N_47255,N_46196);
nor U49598 (N_49598,N_45226,N_45940);
or U49599 (N_49599,N_47499,N_45769);
xnor U49600 (N_49600,N_45958,N_47487);
xor U49601 (N_49601,N_46748,N_46423);
or U49602 (N_49602,N_46399,N_46198);
and U49603 (N_49603,N_46985,N_46064);
nor U49604 (N_49604,N_46780,N_45135);
or U49605 (N_49605,N_46838,N_45107);
and U49606 (N_49606,N_46032,N_46743);
and U49607 (N_49607,N_45054,N_46680);
and U49608 (N_49608,N_47008,N_45404);
nor U49609 (N_49609,N_45253,N_45783);
or U49610 (N_49610,N_45498,N_46047);
and U49611 (N_49611,N_45938,N_47387);
nor U49612 (N_49612,N_47164,N_46090);
and U49613 (N_49613,N_45952,N_46674);
and U49614 (N_49614,N_45616,N_47496);
and U49615 (N_49615,N_46487,N_46774);
and U49616 (N_49616,N_46450,N_47064);
nand U49617 (N_49617,N_46193,N_47364);
and U49618 (N_49618,N_46613,N_46408);
or U49619 (N_49619,N_46071,N_45903);
xnor U49620 (N_49620,N_47302,N_46436);
xor U49621 (N_49621,N_45052,N_47024);
nand U49622 (N_49622,N_47330,N_45732);
nor U49623 (N_49623,N_46824,N_46085);
xnor U49624 (N_49624,N_46688,N_46916);
nor U49625 (N_49625,N_46891,N_46097);
xor U49626 (N_49626,N_45505,N_47359);
nor U49627 (N_49627,N_46497,N_47430);
nor U49628 (N_49628,N_45702,N_46261);
nand U49629 (N_49629,N_46132,N_46297);
nand U49630 (N_49630,N_45215,N_45566);
and U49631 (N_49631,N_46203,N_45525);
nor U49632 (N_49632,N_47141,N_46898);
and U49633 (N_49633,N_46780,N_46647);
nand U49634 (N_49634,N_45379,N_45825);
or U49635 (N_49635,N_46949,N_46196);
nand U49636 (N_49636,N_46720,N_46124);
xor U49637 (N_49637,N_45351,N_45867);
or U49638 (N_49638,N_47260,N_46909);
or U49639 (N_49639,N_46150,N_45819);
and U49640 (N_49640,N_46834,N_45489);
nand U49641 (N_49641,N_46610,N_45228);
xnor U49642 (N_49642,N_45258,N_46982);
and U49643 (N_49643,N_46833,N_45487);
or U49644 (N_49644,N_45158,N_45406);
nand U49645 (N_49645,N_46151,N_47300);
or U49646 (N_49646,N_46179,N_46447);
or U49647 (N_49647,N_45355,N_45005);
nor U49648 (N_49648,N_45757,N_46567);
nand U49649 (N_49649,N_45636,N_46848);
nand U49650 (N_49650,N_45487,N_45386);
nor U49651 (N_49651,N_45607,N_47078);
and U49652 (N_49652,N_47477,N_45926);
nand U49653 (N_49653,N_46568,N_46291);
nor U49654 (N_49654,N_45420,N_46225);
and U49655 (N_49655,N_45612,N_46500);
xnor U49656 (N_49656,N_46948,N_46294);
and U49657 (N_49657,N_46826,N_45369);
xnor U49658 (N_49658,N_45361,N_46040);
nand U49659 (N_49659,N_47207,N_46893);
nand U49660 (N_49660,N_47355,N_45562);
nand U49661 (N_49661,N_45528,N_45203);
nor U49662 (N_49662,N_46332,N_45200);
xnor U49663 (N_49663,N_45447,N_45812);
nor U49664 (N_49664,N_46824,N_46630);
xor U49665 (N_49665,N_47222,N_46681);
nand U49666 (N_49666,N_46117,N_46567);
nand U49667 (N_49667,N_45407,N_46656);
and U49668 (N_49668,N_45046,N_47216);
or U49669 (N_49669,N_46482,N_46150);
and U49670 (N_49670,N_45212,N_45216);
or U49671 (N_49671,N_46510,N_46102);
xor U49672 (N_49672,N_46933,N_47362);
or U49673 (N_49673,N_46069,N_45223);
or U49674 (N_49674,N_45646,N_45336);
nor U49675 (N_49675,N_45818,N_47294);
xnor U49676 (N_49676,N_46761,N_46397);
or U49677 (N_49677,N_46194,N_47030);
or U49678 (N_49678,N_46041,N_46277);
and U49679 (N_49679,N_46490,N_46647);
nor U49680 (N_49680,N_45825,N_45035);
nor U49681 (N_49681,N_45442,N_45104);
nor U49682 (N_49682,N_47048,N_45526);
xor U49683 (N_49683,N_46062,N_45134);
and U49684 (N_49684,N_46720,N_46002);
xor U49685 (N_49685,N_46700,N_46445);
xnor U49686 (N_49686,N_47025,N_45820);
nor U49687 (N_49687,N_45452,N_46158);
nand U49688 (N_49688,N_46446,N_45791);
and U49689 (N_49689,N_47050,N_46996);
xor U49690 (N_49690,N_45481,N_46477);
and U49691 (N_49691,N_46529,N_46008);
nand U49692 (N_49692,N_46387,N_46405);
or U49693 (N_49693,N_45357,N_46444);
nor U49694 (N_49694,N_45849,N_47200);
and U49695 (N_49695,N_45646,N_46952);
nor U49696 (N_49696,N_47453,N_45463);
xor U49697 (N_49697,N_46362,N_45352);
or U49698 (N_49698,N_45162,N_47454);
or U49699 (N_49699,N_46262,N_46496);
or U49700 (N_49700,N_47350,N_46029);
and U49701 (N_49701,N_47038,N_45109);
nor U49702 (N_49702,N_45595,N_47456);
xnor U49703 (N_49703,N_47173,N_47482);
xor U49704 (N_49704,N_45387,N_45218);
xnor U49705 (N_49705,N_45446,N_45926);
and U49706 (N_49706,N_45673,N_47456);
xor U49707 (N_49707,N_45525,N_46345);
xnor U49708 (N_49708,N_45787,N_45778);
xnor U49709 (N_49709,N_46415,N_46631);
or U49710 (N_49710,N_45904,N_45070);
and U49711 (N_49711,N_45816,N_47024);
or U49712 (N_49712,N_46090,N_45111);
and U49713 (N_49713,N_46012,N_45883);
and U49714 (N_49714,N_47235,N_45157);
xor U49715 (N_49715,N_45206,N_47179);
nand U49716 (N_49716,N_45369,N_45244);
xnor U49717 (N_49717,N_46435,N_46706);
nand U49718 (N_49718,N_47145,N_47227);
nor U49719 (N_49719,N_47287,N_46412);
nand U49720 (N_49720,N_45445,N_46406);
and U49721 (N_49721,N_45261,N_46478);
nand U49722 (N_49722,N_46143,N_45189);
xor U49723 (N_49723,N_45517,N_45028);
and U49724 (N_49724,N_45597,N_45846);
or U49725 (N_49725,N_46535,N_46356);
nor U49726 (N_49726,N_47347,N_46173);
or U49727 (N_49727,N_46976,N_46767);
and U49728 (N_49728,N_47390,N_47210);
xnor U49729 (N_49729,N_47162,N_47025);
and U49730 (N_49730,N_45962,N_47325);
nand U49731 (N_49731,N_46721,N_46236);
and U49732 (N_49732,N_46590,N_46716);
or U49733 (N_49733,N_45386,N_45791);
and U49734 (N_49734,N_45186,N_46466);
xnor U49735 (N_49735,N_47036,N_46512);
or U49736 (N_49736,N_45458,N_46387);
xor U49737 (N_49737,N_45384,N_45721);
nor U49738 (N_49738,N_47229,N_45213);
and U49739 (N_49739,N_45296,N_46581);
and U49740 (N_49740,N_47290,N_47193);
nor U49741 (N_49741,N_46507,N_45765);
and U49742 (N_49742,N_45964,N_45949);
nor U49743 (N_49743,N_45201,N_45649);
nor U49744 (N_49744,N_45768,N_45281);
nor U49745 (N_49745,N_45293,N_45057);
and U49746 (N_49746,N_47016,N_45173);
nor U49747 (N_49747,N_46046,N_47172);
nor U49748 (N_49748,N_47245,N_46349);
xnor U49749 (N_49749,N_46858,N_45050);
xnor U49750 (N_49750,N_46003,N_45130);
nor U49751 (N_49751,N_46838,N_45968);
and U49752 (N_49752,N_45964,N_46926);
nand U49753 (N_49753,N_46417,N_45380);
and U49754 (N_49754,N_46539,N_47387);
or U49755 (N_49755,N_45307,N_46627);
xor U49756 (N_49756,N_45555,N_47169);
and U49757 (N_49757,N_46262,N_46521);
nand U49758 (N_49758,N_45367,N_45964);
nor U49759 (N_49759,N_46231,N_45714);
or U49760 (N_49760,N_45650,N_47353);
or U49761 (N_49761,N_45414,N_45850);
nand U49762 (N_49762,N_45960,N_46189);
xor U49763 (N_49763,N_45993,N_46888);
xnor U49764 (N_49764,N_45849,N_45549);
nand U49765 (N_49765,N_47038,N_46286);
nand U49766 (N_49766,N_45746,N_45995);
nand U49767 (N_49767,N_45277,N_45486);
nor U49768 (N_49768,N_46479,N_46758);
and U49769 (N_49769,N_46405,N_45751);
nand U49770 (N_49770,N_46837,N_46731);
xor U49771 (N_49771,N_45958,N_47203);
nor U49772 (N_49772,N_46792,N_45823);
nor U49773 (N_49773,N_45337,N_47339);
and U49774 (N_49774,N_46147,N_46104);
nor U49775 (N_49775,N_47119,N_47278);
xor U49776 (N_49776,N_45995,N_45450);
nor U49777 (N_49777,N_45645,N_45973);
xnor U49778 (N_49778,N_46097,N_45520);
nand U49779 (N_49779,N_46943,N_47251);
or U49780 (N_49780,N_46780,N_46360);
and U49781 (N_49781,N_45092,N_45294);
nand U49782 (N_49782,N_46350,N_47318);
nor U49783 (N_49783,N_46207,N_45167);
and U49784 (N_49784,N_46065,N_46582);
and U49785 (N_49785,N_45508,N_45040);
nand U49786 (N_49786,N_46304,N_46108);
nor U49787 (N_49787,N_46165,N_45229);
or U49788 (N_49788,N_46070,N_47356);
or U49789 (N_49789,N_45916,N_45139);
xnor U49790 (N_49790,N_47293,N_45904);
nor U49791 (N_49791,N_46611,N_46070);
xnor U49792 (N_49792,N_46488,N_46999);
or U49793 (N_49793,N_46262,N_46399);
xnor U49794 (N_49794,N_46968,N_47304);
xnor U49795 (N_49795,N_45128,N_45676);
or U49796 (N_49796,N_46285,N_46659);
nand U49797 (N_49797,N_45536,N_47105);
nor U49798 (N_49798,N_45185,N_46478);
and U49799 (N_49799,N_45093,N_46752);
and U49800 (N_49800,N_45706,N_46571);
or U49801 (N_49801,N_46641,N_46415);
and U49802 (N_49802,N_46147,N_45578);
and U49803 (N_49803,N_46607,N_46435);
and U49804 (N_49804,N_47470,N_46209);
nor U49805 (N_49805,N_45137,N_45671);
xor U49806 (N_49806,N_46736,N_45197);
or U49807 (N_49807,N_45630,N_47258);
or U49808 (N_49808,N_45561,N_45339);
nor U49809 (N_49809,N_46997,N_45444);
xnor U49810 (N_49810,N_47043,N_45404);
and U49811 (N_49811,N_46371,N_47035);
nand U49812 (N_49812,N_46424,N_47375);
or U49813 (N_49813,N_45613,N_45247);
or U49814 (N_49814,N_45940,N_46189);
xor U49815 (N_49815,N_46776,N_45469);
nor U49816 (N_49816,N_46801,N_46244);
xnor U49817 (N_49817,N_45093,N_45035);
xnor U49818 (N_49818,N_46950,N_47145);
or U49819 (N_49819,N_45479,N_46433);
or U49820 (N_49820,N_45402,N_45112);
nand U49821 (N_49821,N_46975,N_45786);
and U49822 (N_49822,N_47401,N_47002);
or U49823 (N_49823,N_47470,N_45841);
nor U49824 (N_49824,N_46922,N_47246);
and U49825 (N_49825,N_46676,N_45729);
or U49826 (N_49826,N_47099,N_46682);
nand U49827 (N_49827,N_47331,N_45715);
and U49828 (N_49828,N_46333,N_46459);
nand U49829 (N_49829,N_45574,N_46446);
xor U49830 (N_49830,N_47090,N_46452);
nor U49831 (N_49831,N_45766,N_45515);
or U49832 (N_49832,N_45811,N_46658);
and U49833 (N_49833,N_46890,N_45188);
nor U49834 (N_49834,N_45893,N_47303);
and U49835 (N_49835,N_45475,N_46356);
and U49836 (N_49836,N_45957,N_45469);
nor U49837 (N_49837,N_47470,N_45490);
nor U49838 (N_49838,N_45528,N_45279);
or U49839 (N_49839,N_45541,N_46885);
xor U49840 (N_49840,N_47199,N_46151);
nand U49841 (N_49841,N_47424,N_47310);
nor U49842 (N_49842,N_47236,N_47284);
and U49843 (N_49843,N_46944,N_46117);
or U49844 (N_49844,N_45741,N_46109);
or U49845 (N_49845,N_47252,N_45794);
and U49846 (N_49846,N_45701,N_45889);
nand U49847 (N_49847,N_46483,N_45435);
xor U49848 (N_49848,N_46576,N_45409);
or U49849 (N_49849,N_47121,N_47091);
xor U49850 (N_49850,N_46838,N_45131);
nor U49851 (N_49851,N_46814,N_46091);
nor U49852 (N_49852,N_45140,N_45474);
or U49853 (N_49853,N_45873,N_45233);
xor U49854 (N_49854,N_45940,N_45427);
nand U49855 (N_49855,N_47086,N_45633);
xor U49856 (N_49856,N_46904,N_45206);
nand U49857 (N_49857,N_46399,N_46618);
xor U49858 (N_49858,N_47026,N_45979);
nand U49859 (N_49859,N_46333,N_46932);
or U49860 (N_49860,N_45648,N_45360);
nand U49861 (N_49861,N_47084,N_45373);
and U49862 (N_49862,N_45654,N_46349);
xnor U49863 (N_49863,N_45835,N_45446);
nand U49864 (N_49864,N_46947,N_47444);
nand U49865 (N_49865,N_47427,N_46706);
xnor U49866 (N_49866,N_46248,N_46243);
nor U49867 (N_49867,N_46664,N_47061);
nand U49868 (N_49868,N_45187,N_47269);
nor U49869 (N_49869,N_45539,N_46843);
nand U49870 (N_49870,N_46666,N_46771);
xor U49871 (N_49871,N_47427,N_46317);
xnor U49872 (N_49872,N_46064,N_45769);
and U49873 (N_49873,N_45861,N_46483);
xnor U49874 (N_49874,N_46822,N_46146);
nand U49875 (N_49875,N_46818,N_46872);
nand U49876 (N_49876,N_45887,N_45135);
or U49877 (N_49877,N_46735,N_47083);
and U49878 (N_49878,N_46362,N_45740);
nor U49879 (N_49879,N_46660,N_45782);
and U49880 (N_49880,N_46544,N_47048);
xor U49881 (N_49881,N_46415,N_46422);
nor U49882 (N_49882,N_45181,N_46633);
or U49883 (N_49883,N_46839,N_46592);
xor U49884 (N_49884,N_45667,N_45840);
and U49885 (N_49885,N_46891,N_46547);
nand U49886 (N_49886,N_45313,N_45304);
and U49887 (N_49887,N_45887,N_46281);
or U49888 (N_49888,N_47408,N_45236);
or U49889 (N_49889,N_45788,N_45735);
nand U49890 (N_49890,N_45687,N_45493);
nand U49891 (N_49891,N_45040,N_46879);
and U49892 (N_49892,N_45868,N_47358);
nand U49893 (N_49893,N_45260,N_45295);
or U49894 (N_49894,N_45840,N_47252);
xnor U49895 (N_49895,N_45533,N_46574);
xnor U49896 (N_49896,N_46052,N_46810);
nor U49897 (N_49897,N_45670,N_45705);
nand U49898 (N_49898,N_46904,N_46105);
xor U49899 (N_49899,N_45563,N_45935);
or U49900 (N_49900,N_47015,N_45788);
nor U49901 (N_49901,N_46087,N_45818);
and U49902 (N_49902,N_46759,N_45035);
xor U49903 (N_49903,N_47092,N_45425);
nor U49904 (N_49904,N_47332,N_46987);
nand U49905 (N_49905,N_45621,N_46342);
xor U49906 (N_49906,N_46157,N_45375);
xor U49907 (N_49907,N_45550,N_47090);
and U49908 (N_49908,N_46313,N_45821);
and U49909 (N_49909,N_47471,N_46742);
xnor U49910 (N_49910,N_46024,N_45589);
nand U49911 (N_49911,N_47286,N_47338);
nor U49912 (N_49912,N_46042,N_45998);
nand U49913 (N_49913,N_46541,N_45602);
xor U49914 (N_49914,N_45012,N_45178);
and U49915 (N_49915,N_47486,N_46517);
and U49916 (N_49916,N_45259,N_45190);
nand U49917 (N_49917,N_45315,N_47333);
xor U49918 (N_49918,N_46059,N_45552);
nand U49919 (N_49919,N_47252,N_47366);
or U49920 (N_49920,N_45840,N_45355);
nor U49921 (N_49921,N_46285,N_47034);
nor U49922 (N_49922,N_46039,N_46898);
xnor U49923 (N_49923,N_46758,N_46459);
and U49924 (N_49924,N_47347,N_46867);
nand U49925 (N_49925,N_46305,N_47350);
nand U49926 (N_49926,N_46204,N_46275);
xnor U49927 (N_49927,N_46278,N_45486);
nor U49928 (N_49928,N_46756,N_45420);
nand U49929 (N_49929,N_45514,N_45545);
nand U49930 (N_49930,N_46748,N_45481);
nor U49931 (N_49931,N_46025,N_45053);
and U49932 (N_49932,N_45694,N_45460);
nor U49933 (N_49933,N_45409,N_46989);
xor U49934 (N_49934,N_46413,N_45202);
nor U49935 (N_49935,N_46431,N_45557);
or U49936 (N_49936,N_46724,N_46792);
nand U49937 (N_49937,N_46948,N_46262);
nor U49938 (N_49938,N_46979,N_45732);
xnor U49939 (N_49939,N_45765,N_46490);
nor U49940 (N_49940,N_45981,N_47327);
and U49941 (N_49941,N_46819,N_45674);
and U49942 (N_49942,N_45344,N_47289);
and U49943 (N_49943,N_45302,N_47428);
nand U49944 (N_49944,N_45348,N_47002);
or U49945 (N_49945,N_46044,N_46028);
and U49946 (N_49946,N_47452,N_45495);
nand U49947 (N_49947,N_45553,N_45683);
and U49948 (N_49948,N_45392,N_46769);
xor U49949 (N_49949,N_45906,N_46438);
or U49950 (N_49950,N_47310,N_46182);
nor U49951 (N_49951,N_46892,N_46566);
or U49952 (N_49952,N_45550,N_45835);
nor U49953 (N_49953,N_47034,N_47389);
nand U49954 (N_49954,N_45301,N_47402);
and U49955 (N_49955,N_45048,N_46768);
and U49956 (N_49956,N_46330,N_46379);
nor U49957 (N_49957,N_46521,N_46389);
or U49958 (N_49958,N_46213,N_45579);
and U49959 (N_49959,N_45004,N_46985);
or U49960 (N_49960,N_46128,N_47365);
nor U49961 (N_49961,N_47154,N_46159);
or U49962 (N_49962,N_46958,N_45631);
nor U49963 (N_49963,N_45802,N_46959);
xor U49964 (N_49964,N_46200,N_46113);
nor U49965 (N_49965,N_46112,N_46256);
xor U49966 (N_49966,N_45538,N_47210);
nand U49967 (N_49967,N_46705,N_45489);
nand U49968 (N_49968,N_46289,N_45921);
xor U49969 (N_49969,N_46149,N_45911);
and U49970 (N_49970,N_47414,N_46452);
xnor U49971 (N_49971,N_46470,N_45371);
nor U49972 (N_49972,N_47435,N_46364);
xnor U49973 (N_49973,N_47423,N_45985);
nor U49974 (N_49974,N_47048,N_46720);
and U49975 (N_49975,N_45487,N_45159);
nand U49976 (N_49976,N_45830,N_45315);
nand U49977 (N_49977,N_46444,N_46527);
nor U49978 (N_49978,N_46224,N_46732);
nand U49979 (N_49979,N_46412,N_47256);
or U49980 (N_49980,N_45202,N_45738);
or U49981 (N_49981,N_46808,N_46337);
nor U49982 (N_49982,N_45431,N_46874);
or U49983 (N_49983,N_45369,N_46790);
nor U49984 (N_49984,N_45149,N_47484);
and U49985 (N_49985,N_47275,N_46311);
xnor U49986 (N_49986,N_45901,N_45215);
or U49987 (N_49987,N_45329,N_45323);
xnor U49988 (N_49988,N_45439,N_47208);
and U49989 (N_49989,N_46948,N_46256);
nand U49990 (N_49990,N_45329,N_46564);
nor U49991 (N_49991,N_47152,N_45301);
or U49992 (N_49992,N_46067,N_46045);
nand U49993 (N_49993,N_46027,N_45908);
nor U49994 (N_49994,N_46750,N_46635);
nand U49995 (N_49995,N_47371,N_46926);
or U49996 (N_49996,N_46931,N_46520);
or U49997 (N_49997,N_45128,N_45432);
or U49998 (N_49998,N_46695,N_45165);
xnor U49999 (N_49999,N_45813,N_45640);
nor UO_0 (O_0,N_48361,N_47630);
nand UO_1 (O_1,N_48499,N_47693);
or UO_2 (O_2,N_49230,N_47904);
and UO_3 (O_3,N_48413,N_49574);
and UO_4 (O_4,N_49944,N_48855);
xor UO_5 (O_5,N_48127,N_47856);
or UO_6 (O_6,N_49337,N_47528);
xor UO_7 (O_7,N_49914,N_49778);
and UO_8 (O_8,N_48005,N_47770);
or UO_9 (O_9,N_48387,N_48923);
xor UO_10 (O_10,N_48036,N_49319);
or UO_11 (O_11,N_48489,N_48717);
nand UO_12 (O_12,N_48690,N_49692);
xor UO_13 (O_13,N_48231,N_49322);
and UO_14 (O_14,N_47937,N_48618);
and UO_15 (O_15,N_49225,N_47638);
nor UO_16 (O_16,N_47705,N_47690);
or UO_17 (O_17,N_48630,N_49248);
or UO_18 (O_18,N_49383,N_47820);
nand UO_19 (O_19,N_48471,N_49754);
xor UO_20 (O_20,N_47617,N_47870);
and UO_21 (O_21,N_49338,N_48031);
or UO_22 (O_22,N_49212,N_49279);
or UO_23 (O_23,N_48436,N_49434);
xor UO_24 (O_24,N_48787,N_47780);
or UO_25 (O_25,N_49636,N_48629);
nor UO_26 (O_26,N_48681,N_47939);
xor UO_27 (O_27,N_48383,N_48033);
xor UO_28 (O_28,N_49571,N_48165);
and UO_29 (O_29,N_48175,N_49628);
nor UO_30 (O_30,N_49738,N_49859);
xnor UO_31 (O_31,N_49823,N_49417);
or UO_32 (O_32,N_48002,N_48193);
nand UO_33 (O_33,N_49341,N_49813);
xor UO_34 (O_34,N_49182,N_47711);
xor UO_35 (O_35,N_49824,N_47522);
nor UO_36 (O_36,N_48990,N_47557);
and UO_37 (O_37,N_47980,N_49081);
nor UO_38 (O_38,N_48405,N_49346);
xnor UO_39 (O_39,N_49254,N_49395);
nand UO_40 (O_40,N_48668,N_49489);
or UO_41 (O_41,N_48076,N_49722);
xnor UO_42 (O_42,N_48275,N_47853);
and UO_43 (O_43,N_49334,N_48954);
and UO_44 (O_44,N_49269,N_49374);
nand UO_45 (O_45,N_48983,N_49630);
nor UO_46 (O_46,N_49236,N_49528);
nand UO_47 (O_47,N_48163,N_48708);
and UO_48 (O_48,N_49903,N_48271);
nor UO_49 (O_49,N_49662,N_48652);
nand UO_50 (O_50,N_49093,N_48014);
nor UO_51 (O_51,N_49460,N_47516);
and UO_52 (O_52,N_48173,N_47696);
nor UO_53 (O_53,N_47663,N_49268);
and UO_54 (O_54,N_48540,N_47565);
nor UO_55 (O_55,N_48500,N_48785);
nor UO_56 (O_56,N_47731,N_49157);
or UO_57 (O_57,N_48968,N_49977);
xor UO_58 (O_58,N_49825,N_49991);
xnor UO_59 (O_59,N_48643,N_49314);
and UO_60 (O_60,N_49452,N_48143);
nor UO_61 (O_61,N_48077,N_49062);
and UO_62 (O_62,N_49713,N_49833);
and UO_63 (O_63,N_47725,N_49331);
or UO_64 (O_64,N_49995,N_47763);
nor UO_65 (O_65,N_47969,N_49201);
and UO_66 (O_66,N_48966,N_49919);
nor UO_67 (O_67,N_48010,N_49665);
and UO_68 (O_68,N_47931,N_49476);
nand UO_69 (O_69,N_47584,N_49698);
or UO_70 (O_70,N_48477,N_48117);
xor UO_71 (O_71,N_47607,N_49497);
nor UO_72 (O_72,N_49853,N_48381);
nor UO_73 (O_73,N_47858,N_48376);
nand UO_74 (O_74,N_49088,N_48769);
and UO_75 (O_75,N_49838,N_48441);
xnor UO_76 (O_76,N_49696,N_49987);
nor UO_77 (O_77,N_48311,N_48705);
xnor UO_78 (O_78,N_48693,N_47579);
xnor UO_79 (O_79,N_49339,N_49750);
or UO_80 (O_80,N_49097,N_48307);
nand UO_81 (O_81,N_48921,N_48837);
nand UO_82 (O_82,N_49695,N_49898);
nor UO_83 (O_83,N_49119,N_48216);
xor UO_84 (O_84,N_48816,N_47821);
xor UO_85 (O_85,N_48247,N_49391);
and UO_86 (O_86,N_48277,N_48437);
nand UO_87 (O_87,N_48492,N_48178);
nand UO_88 (O_88,N_48442,N_48498);
or UO_89 (O_89,N_48953,N_48907);
and UO_90 (O_90,N_47677,N_47935);
nor UO_91 (O_91,N_48521,N_47898);
nor UO_92 (O_92,N_49384,N_48246);
xnor UO_93 (O_93,N_48801,N_48885);
and UO_94 (O_94,N_48707,N_48292);
xor UO_95 (O_95,N_48955,N_48223);
nand UO_96 (O_96,N_47542,N_49585);
xnor UO_97 (O_97,N_49701,N_49222);
xnor UO_98 (O_98,N_49749,N_48928);
or UO_99 (O_99,N_49865,N_49207);
xor UO_100 (O_100,N_48034,N_48831);
nand UO_101 (O_101,N_49289,N_48805);
and UO_102 (O_102,N_49109,N_47539);
nor UO_103 (O_103,N_48448,N_49408);
xor UO_104 (O_104,N_47737,N_47768);
nand UO_105 (O_105,N_48653,N_47918);
nand UO_106 (O_106,N_49422,N_49169);
and UO_107 (O_107,N_49507,N_48541);
nand UO_108 (O_108,N_48520,N_49568);
xnor UO_109 (O_109,N_48184,N_48998);
xor UO_110 (O_110,N_47950,N_48768);
or UO_111 (O_111,N_49634,N_48369);
nand UO_112 (O_112,N_49557,N_49603);
nor UO_113 (O_113,N_49085,N_49240);
and UO_114 (O_114,N_48919,N_49753);
or UO_115 (O_115,N_49454,N_49542);
nand UO_116 (O_116,N_48967,N_48762);
nand UO_117 (O_117,N_49617,N_49974);
or UO_118 (O_118,N_49055,N_47752);
xnor UO_119 (O_119,N_48766,N_49581);
and UO_120 (O_120,N_48777,N_48200);
nor UO_121 (O_121,N_49797,N_48651);
xor UO_122 (O_122,N_49027,N_49875);
and UO_123 (O_123,N_48610,N_49465);
nor UO_124 (O_124,N_48323,N_49503);
and UO_125 (O_125,N_49623,N_49608);
or UO_126 (O_126,N_47627,N_49515);
nor UO_127 (O_127,N_48069,N_49596);
and UO_128 (O_128,N_47877,N_48234);
xnor UO_129 (O_129,N_49849,N_49361);
or UO_130 (O_130,N_48543,N_48700);
or UO_131 (O_131,N_49810,N_49801);
xor UO_132 (O_132,N_48462,N_49028);
or UO_133 (O_133,N_48552,N_49734);
nand UO_134 (O_134,N_47642,N_49601);
nand UO_135 (O_135,N_48140,N_49782);
or UO_136 (O_136,N_48289,N_49439);
and UO_137 (O_137,N_48548,N_48470);
nor UO_138 (O_138,N_48112,N_49747);
xnor UO_139 (O_139,N_48506,N_47879);
xnor UO_140 (O_140,N_49659,N_49016);
nand UO_141 (O_141,N_47905,N_47750);
nor UO_142 (O_142,N_48519,N_49049);
and UO_143 (O_143,N_48713,N_49072);
nor UO_144 (O_144,N_49563,N_49845);
nor UO_145 (O_145,N_48438,N_49532);
or UO_146 (O_146,N_48198,N_49057);
or UO_147 (O_147,N_48959,N_49305);
and UO_148 (O_148,N_48624,N_48207);
or UO_149 (O_149,N_49350,N_48974);
and UO_150 (O_150,N_49294,N_49598);
xnor UO_151 (O_151,N_48562,N_49927);
and UO_152 (O_152,N_48429,N_49549);
xnor UO_153 (O_153,N_48722,N_48661);
nor UO_154 (O_154,N_49921,N_49794);
or UO_155 (O_155,N_48759,N_49550);
and UO_156 (O_156,N_48371,N_49008);
and UO_157 (O_157,N_49961,N_48871);
nand UO_158 (O_158,N_49595,N_49590);
or UO_159 (O_159,N_48137,N_48791);
nand UO_160 (O_160,N_47676,N_48633);
and UO_161 (O_161,N_47695,N_49902);
xor UO_162 (O_162,N_48201,N_49803);
or UO_163 (O_163,N_48712,N_47536);
xor UO_164 (O_164,N_48776,N_48620);
and UO_165 (O_165,N_49519,N_47538);
or UO_166 (O_166,N_49631,N_49783);
or UO_167 (O_167,N_49949,N_49150);
nor UO_168 (O_168,N_47922,N_47517);
and UO_169 (O_169,N_49234,N_49473);
xnor UO_170 (O_170,N_49321,N_49398);
nor UO_171 (O_171,N_49437,N_49101);
nand UO_172 (O_172,N_48149,N_49034);
and UO_173 (O_173,N_48674,N_49498);
or UO_174 (O_174,N_48676,N_49180);
nand UO_175 (O_175,N_48314,N_48526);
xnor UO_176 (O_176,N_48586,N_49209);
or UO_177 (O_177,N_48449,N_49655);
nor UO_178 (O_178,N_47976,N_49527);
and UO_179 (O_179,N_47916,N_48751);
nor UO_180 (O_180,N_49788,N_48397);
or UO_181 (O_181,N_47533,N_47609);
nor UO_182 (O_182,N_48073,N_48943);
xnor UO_183 (O_183,N_49671,N_48063);
or UO_184 (O_184,N_49400,N_49872);
nand UO_185 (O_185,N_49160,N_47634);
or UO_186 (O_186,N_48616,N_49271);
nor UO_187 (O_187,N_48293,N_47855);
and UO_188 (O_188,N_48570,N_48932);
xnor UO_189 (O_189,N_48236,N_49638);
and UO_190 (O_190,N_49502,N_48527);
or UO_191 (O_191,N_48428,N_48497);
nor UO_192 (O_192,N_49108,N_49354);
xnor UO_193 (O_193,N_47672,N_49155);
nand UO_194 (O_194,N_49998,N_47691);
xnor UO_195 (O_195,N_47556,N_47745);
nor UO_196 (O_196,N_49270,N_47626);
or UO_197 (O_197,N_48836,N_48186);
xnor UO_198 (O_198,N_48869,N_48822);
xor UO_199 (O_199,N_48233,N_49067);
nor UO_200 (O_200,N_49114,N_48542);
nor UO_201 (O_201,N_48485,N_47515);
nand UO_202 (O_202,N_49310,N_47632);
nor UO_203 (O_203,N_49245,N_49227);
or UO_204 (O_204,N_49570,N_48351);
and UO_205 (O_205,N_48318,N_47830);
and UO_206 (O_206,N_48480,N_49948);
nor UO_207 (O_207,N_49826,N_48695);
or UO_208 (O_208,N_49365,N_48644);
and UO_209 (O_209,N_48905,N_47896);
and UO_210 (O_210,N_48895,N_47839);
nor UO_211 (O_211,N_49247,N_48842);
and UO_212 (O_212,N_49144,N_48995);
or UO_213 (O_213,N_48594,N_47622);
xnor UO_214 (O_214,N_47744,N_48657);
or UO_215 (O_215,N_49128,N_48402);
nand UO_216 (O_216,N_49411,N_48760);
or UO_217 (O_217,N_48414,N_47668);
nor UO_218 (O_218,N_48082,N_49353);
nor UO_219 (O_219,N_49970,N_47551);
nor UO_220 (O_220,N_48299,N_49483);
or UO_221 (O_221,N_48576,N_48993);
and UO_222 (O_222,N_47546,N_49768);
and UO_223 (O_223,N_49781,N_49802);
nand UO_224 (O_224,N_49748,N_47836);
nand UO_225 (O_225,N_48803,N_49369);
and UO_226 (O_226,N_48728,N_49158);
xnor UO_227 (O_227,N_48926,N_48018);
nand UO_228 (O_228,N_48160,N_48450);
or UO_229 (O_229,N_47585,N_48088);
nor UO_230 (O_230,N_49912,N_47851);
nor UO_231 (O_231,N_49074,N_47886);
xor UO_232 (O_232,N_49228,N_49320);
or UO_233 (O_233,N_48194,N_48678);
nand UO_234 (O_234,N_47912,N_48013);
nor UO_235 (O_235,N_49191,N_48296);
xor UO_236 (O_236,N_48560,N_49523);
nand UO_237 (O_237,N_47567,N_48715);
nor UO_238 (O_238,N_47815,N_48403);
nand UO_239 (O_239,N_47955,N_49178);
or UO_240 (O_240,N_49011,N_48040);
or UO_241 (O_241,N_49131,N_49103);
nand UO_242 (O_242,N_49646,N_49772);
nor UO_243 (O_243,N_48172,N_49059);
nor UO_244 (O_244,N_49643,N_47953);
xnor UO_245 (O_245,N_49610,N_48102);
nor UO_246 (O_246,N_48092,N_48346);
xnor UO_247 (O_247,N_47652,N_49421);
or UO_248 (O_248,N_48103,N_49039);
or UO_249 (O_249,N_49640,N_48490);
nor UO_250 (O_250,N_48596,N_49923);
xnor UO_251 (O_251,N_48281,N_48208);
and UO_252 (O_252,N_48495,N_49867);
nand UO_253 (O_253,N_49614,N_47764);
nor UO_254 (O_254,N_48726,N_49500);
and UO_255 (O_255,N_48951,N_48536);
nor UO_256 (O_256,N_47523,N_49834);
xor UO_257 (O_257,N_49141,N_48514);
and UO_258 (O_258,N_47739,N_48870);
and UO_259 (O_259,N_47724,N_49589);
or UO_260 (O_260,N_49934,N_47753);
and UO_261 (O_261,N_47956,N_48673);
and UO_262 (O_262,N_47822,N_49776);
or UO_263 (O_263,N_48790,N_49357);
nand UO_264 (O_264,N_47681,N_49148);
nor UO_265 (O_265,N_48771,N_49540);
and UO_266 (O_266,N_48725,N_48938);
or UO_267 (O_267,N_48187,N_47811);
xnor UO_268 (O_268,N_49467,N_47748);
nand UO_269 (O_269,N_47548,N_48434);
xnor UO_270 (O_270,N_48931,N_49347);
and UO_271 (O_271,N_49830,N_49719);
nor UO_272 (O_272,N_48704,N_48670);
xnor UO_273 (O_273,N_49688,N_49013);
or UO_274 (O_274,N_49984,N_48986);
or UO_275 (O_275,N_48783,N_48058);
xnor UO_276 (O_276,N_48873,N_47894);
nand UO_277 (O_277,N_48125,N_48814);
xor UO_278 (O_278,N_47513,N_49900);
and UO_279 (O_279,N_49962,N_49325);
nand UO_280 (O_280,N_49156,N_49586);
and UO_281 (O_281,N_49204,N_48665);
or UO_282 (O_282,N_47701,N_49746);
or UO_283 (O_283,N_49001,N_48425);
nor UO_284 (O_284,N_49579,N_48961);
or UO_285 (O_285,N_49026,N_47659);
or UO_286 (O_286,N_48081,N_47776);
xor UO_287 (O_287,N_48382,N_49641);
and UO_288 (O_288,N_48411,N_49763);
xnor UO_289 (O_289,N_49683,N_47618);
and UO_290 (O_290,N_49134,N_49704);
nor UO_291 (O_291,N_49443,N_47929);
or UO_292 (O_292,N_49807,N_48363);
nor UO_293 (O_293,N_49186,N_49444);
nor UO_294 (O_294,N_49583,N_47641);
nand UO_295 (O_295,N_48724,N_47646);
nor UO_296 (O_296,N_49355,N_47566);
nand UO_297 (O_297,N_47945,N_49419);
xor UO_298 (O_298,N_49855,N_48048);
or UO_299 (O_299,N_47949,N_49862);
xnor UO_300 (O_300,N_47909,N_49622);
xor UO_301 (O_301,N_49715,N_49602);
and UO_302 (O_302,N_48887,N_47654);
xor UO_303 (O_303,N_47738,N_49396);
and UO_304 (O_304,N_47901,N_47788);
nand UO_305 (O_305,N_48772,N_48879);
nor UO_306 (O_306,N_47583,N_47938);
or UO_307 (O_307,N_48044,N_49371);
and UO_308 (O_308,N_48358,N_48862);
xor UO_309 (O_309,N_48565,N_49584);
xnor UO_310 (O_310,N_49766,N_48511);
nor UO_311 (O_311,N_47616,N_48614);
and UO_312 (O_312,N_47908,N_48893);
or UO_313 (O_313,N_48270,N_49342);
nand UO_314 (O_314,N_48078,N_49442);
nand UO_315 (O_315,N_47686,N_49492);
nand UO_316 (O_316,N_48153,N_48575);
nand UO_317 (O_317,N_49918,N_49508);
nor UO_318 (O_318,N_48973,N_48922);
nor UO_319 (O_319,N_48874,N_47614);
nand UO_320 (O_320,N_49386,N_49745);
and UO_321 (O_321,N_49136,N_49566);
nor UO_322 (O_322,N_48736,N_49423);
or UO_323 (O_323,N_47534,N_47742);
and UO_324 (O_324,N_49769,N_49260);
or UO_325 (O_325,N_48141,N_48891);
nand UO_326 (O_326,N_48020,N_48135);
xnor UO_327 (O_327,N_49135,N_48512);
xnor UO_328 (O_328,N_48667,N_48128);
nor UO_329 (O_329,N_47761,N_47997);
nor UO_330 (O_330,N_48463,N_48316);
xnor UO_331 (O_331,N_48881,N_48568);
nand UO_332 (O_332,N_48601,N_48864);
or UO_333 (O_333,N_49064,N_49928);
nor UO_334 (O_334,N_48537,N_49393);
and UO_335 (O_335,N_47589,N_48792);
nand UO_336 (O_336,N_48045,N_47503);
or UO_337 (O_337,N_48267,N_48743);
nand UO_338 (O_338,N_47511,N_49139);
nor UO_339 (O_339,N_48215,N_47735);
or UO_340 (O_340,N_48256,N_48094);
nand UO_341 (O_341,N_49588,N_49997);
nor UO_342 (O_342,N_48079,N_48640);
nor UO_343 (O_343,N_48431,N_47722);
xnor UO_344 (O_344,N_49068,N_48903);
or UO_345 (O_345,N_49285,N_47595);
and UO_346 (O_346,N_48053,N_48309);
nand UO_347 (O_347,N_48177,N_48445);
nand UO_348 (O_348,N_49162,N_49981);
nand UO_349 (O_349,N_47550,N_49149);
nand UO_350 (O_350,N_48604,N_49477);
nand UO_351 (O_351,N_48003,N_49539);
or UO_352 (O_352,N_48426,N_47925);
xnor UO_353 (O_353,N_48278,N_48074);
nor UO_354 (O_354,N_48529,N_48433);
xor UO_355 (O_355,N_49858,N_48212);
and UO_356 (O_356,N_49387,N_48294);
nor UO_357 (O_357,N_48623,N_49251);
nand UO_358 (O_358,N_48559,N_49448);
nand UO_359 (O_359,N_48213,N_48237);
nand UO_360 (O_360,N_48843,N_49535);
nor UO_361 (O_361,N_49282,N_48828);
or UO_362 (O_362,N_49187,N_49983);
and UO_363 (O_363,N_48494,N_48156);
xnor UO_364 (O_364,N_48016,N_47840);
xnor UO_365 (O_365,N_47610,N_48319);
xnor UO_366 (O_366,N_48528,N_49086);
nor UO_367 (O_367,N_48756,N_49123);
nor UO_368 (O_368,N_49594,N_49717);
nand UO_369 (O_369,N_48295,N_48007);
xor UO_370 (O_370,N_47590,N_49856);
or UO_371 (O_371,N_48355,N_49210);
nand UO_372 (O_372,N_49879,N_49189);
nand UO_373 (O_373,N_48111,N_49516);
or UO_374 (O_374,N_49909,N_48022);
or UO_375 (O_375,N_48284,N_48181);
and UO_376 (O_376,N_47846,N_49551);
nand UO_377 (O_377,N_49891,N_47832);
nand UO_378 (O_378,N_48352,N_49487);
nor UO_379 (O_379,N_48911,N_48254);
nor UO_380 (O_380,N_47620,N_48067);
xnor UO_381 (O_381,N_47795,N_49529);
nor UO_382 (O_382,N_49559,N_49525);
nor UO_383 (O_383,N_48424,N_49220);
xnor UO_384 (O_384,N_48917,N_47869);
or UO_385 (O_385,N_49307,N_49901);
nor UO_386 (O_386,N_48978,N_48846);
or UO_387 (O_387,N_48364,N_49253);
and UO_388 (O_388,N_48444,N_49664);
and UO_389 (O_389,N_48510,N_48844);
nand UO_390 (O_390,N_47773,N_49440);
xnor UO_391 (O_391,N_48386,N_48151);
or UO_392 (O_392,N_49406,N_49988);
nor UO_393 (O_393,N_47604,N_48392);
nand UO_394 (O_394,N_48166,N_49555);
nand UO_395 (O_395,N_49296,N_48268);
xnor UO_396 (O_396,N_49930,N_48116);
nand UO_397 (O_397,N_48976,N_47692);
nor UO_398 (O_398,N_48396,N_49455);
nand UO_399 (O_399,N_48718,N_48041);
nor UO_400 (O_400,N_48287,N_49221);
xor UO_401 (O_401,N_49463,N_47648);
nor UO_402 (O_402,N_48691,N_48159);
nand UO_403 (O_403,N_49561,N_49513);
nor UO_404 (O_404,N_47817,N_48603);
nor UO_405 (O_405,N_49675,N_48343);
nand UO_406 (O_406,N_49061,N_49229);
xnor UO_407 (O_407,N_48349,N_48339);
nor UO_408 (O_408,N_47837,N_49152);
nand UO_409 (O_409,N_48375,N_49416);
nand UO_410 (O_410,N_47719,N_49729);
xor UO_411 (O_411,N_49084,N_48747);
nor UO_412 (O_412,N_48142,N_49179);
nor UO_413 (O_413,N_49790,N_48675);
or UO_414 (O_414,N_47917,N_49520);
nand UO_415 (O_415,N_49197,N_49620);
and UO_416 (O_416,N_49140,N_48336);
or UO_417 (O_417,N_48692,N_47606);
and UO_418 (O_418,N_48035,N_49710);
xor UO_419 (O_419,N_48650,N_47867);
nand UO_420 (O_420,N_47636,N_49739);
or UO_421 (O_421,N_49301,N_49056);
nand UO_422 (O_422,N_49509,N_49107);
xnor UO_423 (O_423,N_48697,N_49318);
xor UO_424 (O_424,N_49741,N_47911);
nor UO_425 (O_425,N_48517,N_49818);
xnor UO_426 (O_426,N_48797,N_47872);
nand UO_427 (O_427,N_49326,N_48694);
or UO_428 (O_428,N_48199,N_49521);
or UO_429 (O_429,N_49814,N_47643);
nand UO_430 (O_430,N_49642,N_48706);
xnor UO_431 (O_431,N_49447,N_47535);
and UO_432 (O_432,N_49380,N_48037);
nand UO_433 (O_433,N_49138,N_49740);
or UO_434 (O_434,N_47504,N_49827);
or UO_435 (O_435,N_49435,N_49940);
nand UO_436 (O_436,N_48466,N_49433);
xor UO_437 (O_437,N_48464,N_48804);
xnor UO_438 (O_438,N_47807,N_49537);
or UO_439 (O_439,N_49171,N_48940);
nand UO_440 (O_440,N_48897,N_48249);
nor UO_441 (O_441,N_49931,N_48326);
nand UO_442 (O_442,N_49118,N_48419);
nand UO_443 (O_443,N_47540,N_49576);
or UO_444 (O_444,N_48407,N_49989);
or UO_445 (O_445,N_48269,N_48344);
xnor UO_446 (O_446,N_49815,N_47678);
and UO_447 (O_447,N_47889,N_48979);
or UO_448 (O_448,N_49226,N_49842);
nor UO_449 (O_449,N_48481,N_48832);
or UO_450 (O_450,N_47860,N_49906);
and UO_451 (O_451,N_47952,N_48461);
nor UO_452 (O_452,N_48120,N_48539);
nor UO_453 (O_453,N_49392,N_48531);
or UO_454 (O_454,N_49684,N_48969);
or UO_455 (O_455,N_49231,N_48291);
xor UO_456 (O_456,N_49445,N_49367);
nor UO_457 (O_457,N_49657,N_48557);
xor UO_458 (O_458,N_47564,N_47895);
nor UO_459 (O_459,N_49257,N_49273);
nand UO_460 (O_460,N_48388,N_49985);
and UO_461 (O_461,N_47749,N_48359);
and UO_462 (O_462,N_48826,N_49420);
nand UO_463 (O_463,N_48068,N_49170);
xnor UO_464 (O_464,N_48158,N_49767);
or UO_465 (O_465,N_49063,N_49724);
and UO_466 (O_466,N_49510,N_47847);
xnor UO_467 (O_467,N_49091,N_49324);
or UO_468 (O_468,N_48915,N_47793);
or UO_469 (O_469,N_48085,N_49647);
nand UO_470 (O_470,N_49894,N_49045);
nor UO_471 (O_471,N_47995,N_49605);
and UO_472 (O_472,N_48852,N_48144);
nor UO_473 (O_473,N_49025,N_47670);
xor UO_474 (O_474,N_48205,N_47628);
xor UO_475 (O_475,N_47802,N_47576);
xnor UO_476 (O_476,N_49565,N_49963);
xor UO_477 (O_477,N_48182,N_48525);
nand UO_478 (O_478,N_49450,N_48948);
and UO_479 (O_479,N_49673,N_49175);
nand UO_480 (O_480,N_47649,N_47828);
and UO_481 (O_481,N_48834,N_47973);
nor UO_482 (O_482,N_48742,N_48865);
or UO_483 (O_483,N_49030,N_48486);
xor UO_484 (O_484,N_49611,N_47657);
and UO_485 (O_485,N_48566,N_48154);
xnor UO_486 (O_486,N_48719,N_49272);
nand UO_487 (O_487,N_47792,N_49362);
or UO_488 (O_488,N_49723,N_48809);
nand UO_489 (O_489,N_47613,N_47891);
nand UO_490 (O_490,N_49569,N_49922);
xnor UO_491 (O_491,N_48427,N_49486);
or UO_492 (O_492,N_49333,N_48171);
nand UO_493 (O_493,N_48658,N_48532);
xor UO_494 (O_494,N_47612,N_49597);
or UO_495 (O_495,N_48059,N_48243);
xor UO_496 (O_496,N_49792,N_48872);
and UO_497 (O_497,N_48645,N_48333);
xor UO_498 (O_498,N_49866,N_47982);
nor UO_499 (O_499,N_47553,N_47924);
nor UO_500 (O_500,N_48342,N_49058);
nor UO_501 (O_501,N_49094,N_48204);
or UO_502 (O_502,N_47702,N_49364);
nor UO_503 (O_503,N_48679,N_49839);
nand UO_504 (O_504,N_47732,N_48518);
nand UO_505 (O_505,N_47530,N_48083);
nand UO_506 (O_506,N_49964,N_47789);
and UO_507 (O_507,N_49399,N_49832);
nor UO_508 (O_508,N_47983,N_49712);
xor UO_509 (O_509,N_48418,N_49945);
and UO_510 (O_510,N_49046,N_49799);
nor UO_511 (O_511,N_49428,N_47527);
or UO_512 (O_512,N_49911,N_47510);
nor UO_513 (O_513,N_47993,N_48752);
nor UO_514 (O_514,N_48929,N_48660);
xor UO_515 (O_515,N_48004,N_47520);
xor UO_516 (O_516,N_49099,N_49313);
and UO_517 (O_517,N_49735,N_49883);
and UO_518 (O_518,N_48356,N_49625);
nand UO_519 (O_519,N_47577,N_49377);
and UO_520 (O_520,N_49146,N_49481);
nand UO_521 (O_521,N_48621,N_47508);
and UO_522 (O_522,N_49404,N_48947);
nand UO_523 (O_523,N_49517,N_48298);
xnor UO_524 (O_524,N_48416,N_49885);
and UO_525 (O_525,N_48026,N_48224);
or UO_526 (O_526,N_48297,N_47717);
and UO_527 (O_527,N_48952,N_48056);
xor UO_528 (O_528,N_47586,N_48446);
xor UO_529 (O_529,N_47600,N_49127);
nor UO_530 (O_530,N_48260,N_49878);
and UO_531 (O_531,N_47706,N_49385);
or UO_532 (O_532,N_48738,N_47833);
and UO_533 (O_533,N_48868,N_49880);
nand UO_534 (O_534,N_47887,N_49764);
nand UO_535 (O_535,N_49065,N_47920);
nand UO_536 (O_536,N_48169,N_48720);
and UO_537 (O_537,N_49658,N_49202);
nand UO_538 (O_538,N_48835,N_47637);
nor UO_539 (O_539,N_49453,N_49779);
nor UO_540 (O_540,N_47665,N_48017);
or UO_541 (O_541,N_48796,N_49896);
xor UO_542 (O_542,N_47653,N_49388);
nor UO_543 (O_543,N_49560,N_48262);
nor UO_544 (O_544,N_47671,N_47741);
or UO_545 (O_545,N_48628,N_48987);
and UO_546 (O_546,N_47906,N_49246);
or UO_547 (O_547,N_47545,N_49777);
nor UO_548 (O_548,N_48909,N_48101);
or UO_549 (O_549,N_48867,N_48334);
and UO_550 (O_550,N_48731,N_49639);
nor UO_551 (O_551,N_49758,N_49685);
and UO_552 (O_552,N_49607,N_48795);
and UO_553 (O_553,N_49265,N_48958);
or UO_554 (O_554,N_49728,N_47876);
and UO_555 (O_555,N_48052,N_48811);
and UO_556 (O_556,N_47915,N_49881);
nor UO_557 (O_557,N_49348,N_48065);
and UO_558 (O_558,N_49714,N_49021);
xnor UO_559 (O_559,N_48936,N_49116);
xor UO_560 (O_560,N_49935,N_49462);
nand UO_561 (O_561,N_48944,N_49785);
or UO_562 (O_562,N_48019,N_48567);
xnor UO_563 (O_563,N_48941,N_47747);
or UO_564 (O_564,N_49087,N_49032);
and UO_565 (O_565,N_48273,N_49441);
or UO_566 (O_566,N_49886,N_48935);
xor UO_567 (O_567,N_49390,N_48251);
nor UO_568 (O_568,N_49295,N_47593);
xor UO_569 (O_569,N_49299,N_49262);
and UO_570 (O_570,N_48075,N_49806);
or UO_571 (O_571,N_48988,N_49887);
xnor UO_572 (O_572,N_47841,N_47838);
nor UO_573 (O_573,N_47720,N_48285);
xor UO_574 (O_574,N_48301,N_49547);
or UO_575 (O_575,N_48686,N_49992);
nand UO_576 (O_576,N_48395,N_49616);
nor UO_577 (O_577,N_48105,N_49471);
xor UO_578 (O_578,N_49208,N_48564);
nand UO_579 (O_579,N_48838,N_49407);
or UO_580 (O_580,N_48977,N_48595);
nand UO_581 (O_581,N_48209,N_48145);
nand UO_582 (O_582,N_48664,N_48245);
nor UO_583 (O_583,N_49041,N_49003);
xor UO_584 (O_584,N_48875,N_49637);
xnor UO_585 (O_585,N_49106,N_49966);
nor UO_586 (O_586,N_49626,N_49177);
and UO_587 (O_587,N_47544,N_48337);
and UO_588 (O_588,N_49426,N_49491);
xnor UO_589 (O_589,N_47884,N_49316);
nand UO_590 (O_590,N_49648,N_49000);
and UO_591 (O_591,N_48098,N_49593);
or UO_592 (O_592,N_48534,N_49402);
or UO_593 (O_593,N_48818,N_47919);
nor UO_594 (O_594,N_49656,N_48920);
or UO_595 (O_595,N_48501,N_47890);
and UO_596 (O_596,N_48839,N_49176);
nor UO_597 (O_597,N_48851,N_49232);
xor UO_598 (O_598,N_48577,N_47987);
nand UO_599 (O_599,N_48721,N_48259);
or UO_600 (O_600,N_47797,N_48242);
nand UO_601 (O_601,N_47984,N_49937);
xor UO_602 (O_602,N_49233,N_48398);
and UO_603 (O_603,N_49691,N_48763);
and UO_604 (O_604,N_49351,N_49938);
nand UO_605 (O_605,N_48677,N_49079);
nor UO_606 (O_606,N_48286,N_47861);
or UO_607 (O_607,N_49939,N_49693);
xnor UO_608 (O_608,N_49405,N_48900);
and UO_609 (O_609,N_48227,N_49494);
nand UO_610 (O_610,N_49242,N_47526);
or UO_611 (O_611,N_48417,N_47581);
xor UO_612 (O_612,N_49791,N_47698);
xor UO_613 (O_613,N_49479,N_49924);
nor UO_614 (O_614,N_48240,N_48906);
or UO_615 (O_615,N_48472,N_47674);
or UO_616 (O_616,N_49415,N_49822);
and UO_617 (O_617,N_48753,N_48191);
and UO_618 (O_618,N_48788,N_48734);
nand UO_619 (O_619,N_48321,N_49165);
nor UO_620 (O_620,N_47818,N_48711);
nor UO_621 (O_621,N_49505,N_49876);
xnor UO_622 (O_622,N_47721,N_47758);
nand UO_623 (O_623,N_47512,N_49744);
and UO_624 (O_624,N_48385,N_48012);
and UO_625 (O_625,N_48432,N_49727);
nor UO_626 (O_626,N_49624,N_49010);
nand UO_627 (O_627,N_49300,N_47900);
nor UO_628 (O_628,N_48469,N_49456);
xor UO_629 (O_629,N_47588,N_47549);
or UO_630 (O_630,N_49050,N_49366);
nor UO_631 (O_631,N_48982,N_48750);
nor UO_632 (O_632,N_49653,N_47796);
nand UO_633 (O_633,N_47843,N_49070);
nand UO_634 (O_634,N_47507,N_49414);
xnor UO_635 (O_635,N_48808,N_48220);
xnor UO_636 (O_636,N_48000,N_47689);
nand UO_637 (O_637,N_47624,N_48138);
nor UO_638 (O_638,N_49373,N_49612);
or UO_639 (O_639,N_47729,N_47771);
and UO_640 (O_640,N_49291,N_48325);
nor UO_641 (O_641,N_47754,N_48524);
or UO_642 (O_642,N_47703,N_49255);
nor UO_643 (O_643,N_49848,N_48550);
nand UO_644 (O_644,N_47597,N_48646);
xor UO_645 (O_645,N_48960,N_49040);
or UO_646 (O_646,N_49192,N_48984);
nand UO_647 (O_647,N_47892,N_49281);
xor UO_648 (O_648,N_48680,N_49147);
xnor UO_649 (O_649,N_47991,N_49143);
xnor UO_650 (O_650,N_48970,N_49737);
and UO_651 (O_651,N_48134,N_48266);
or UO_652 (O_652,N_47733,N_49464);
nor UO_653 (O_653,N_48806,N_49129);
or UO_654 (O_654,N_47778,N_49195);
or UO_655 (O_655,N_49847,N_48773);
and UO_656 (O_656,N_49835,N_48683);
nor UO_657 (O_657,N_47509,N_48710);
or UO_658 (O_658,N_48904,N_49558);
nand UO_659 (O_659,N_47996,N_49345);
nor UO_660 (O_660,N_48228,N_48136);
nor UO_661 (O_661,N_49592,N_49907);
xor UO_662 (O_662,N_48218,N_49293);
or UO_663 (O_663,N_49496,N_47990);
nor UO_664 (O_664,N_49820,N_48331);
xor UO_665 (O_665,N_47714,N_48021);
xnor UO_666 (O_666,N_49812,N_48569);
nor UO_667 (O_667,N_49104,N_48072);
or UO_668 (O_668,N_49112,N_47882);
nor UO_669 (O_669,N_48997,N_47957);
and UO_670 (O_670,N_48183,N_49577);
or UO_671 (O_671,N_47661,N_49436);
nor UO_672 (O_672,N_48043,N_48638);
nor UO_673 (O_673,N_49752,N_47897);
and UO_674 (O_674,N_48884,N_48229);
xnor UO_675 (O_675,N_47781,N_47798);
nor UO_676 (O_676,N_49890,N_49468);
nor UO_677 (O_677,N_47502,N_47740);
or UO_678 (O_678,N_49687,N_48853);
nand UO_679 (O_679,N_49929,N_48100);
nand UO_680 (O_680,N_48584,N_47525);
or UO_681 (O_681,N_49682,N_49022);
nor UO_682 (O_682,N_49286,N_47835);
xor UO_683 (O_683,N_49418,N_48735);
nand UO_684 (O_684,N_49805,N_49275);
nor UO_685 (O_685,N_48636,N_48765);
xnor UO_686 (O_686,N_48152,N_49451);
or UO_687 (O_687,N_48341,N_49976);
or UO_688 (O_688,N_47558,N_49773);
nand UO_689 (O_689,N_47640,N_47831);
xor UO_690 (O_690,N_49604,N_47967);
nand UO_691 (O_691,N_48757,N_49762);
xnor UO_692 (O_692,N_48468,N_48802);
xor UO_693 (O_693,N_47913,N_49315);
nor UO_694 (O_694,N_49854,N_47631);
or UO_695 (O_695,N_49166,N_48108);
and UO_696 (O_696,N_48006,N_49621);
xor UO_697 (O_697,N_49633,N_48157);
and UO_698 (O_698,N_48161,N_48515);
nand UO_699 (O_699,N_48039,N_49668);
nor UO_700 (O_700,N_49298,N_49526);
nand UO_701 (O_701,N_49469,N_49548);
nor UO_702 (O_702,N_49787,N_48367);
xnor UO_703 (O_703,N_49869,N_47709);
or UO_704 (O_704,N_47940,N_48093);
xor UO_705 (O_705,N_48912,N_48114);
or UO_706 (O_706,N_47645,N_48404);
xor UO_707 (O_707,N_48847,N_49667);
or UO_708 (O_708,N_48057,N_48248);
xor UO_709 (O_709,N_49629,N_48423);
or UO_710 (O_710,N_48829,N_48888);
xor UO_711 (O_711,N_48746,N_47941);
nand UO_712 (O_712,N_49007,N_49263);
nand UO_713 (O_713,N_49666,N_49358);
nor UO_714 (O_714,N_47947,N_49522);
or UO_715 (O_715,N_49533,N_48957);
and UO_716 (O_716,N_48168,N_49843);
nor UO_717 (O_717,N_48132,N_49276);
and UO_718 (O_718,N_47932,N_49975);
nand UO_719 (O_719,N_48162,N_49485);
or UO_720 (O_720,N_49283,N_48669);
nand UO_721 (O_721,N_49567,N_48764);
and UO_722 (O_722,N_49863,N_48840);
or UO_723 (O_723,N_49908,N_48880);
nand UO_724 (O_724,N_48613,N_48280);
nand UO_725 (O_725,N_48632,N_47726);
nand UO_726 (O_726,N_49461,N_48588);
nor UO_727 (O_727,N_47878,N_48230);
or UO_728 (O_728,N_49986,N_48551);
nand UO_729 (O_729,N_48555,N_47700);
nor UO_730 (O_730,N_48739,N_49761);
or UO_731 (O_731,N_48197,N_48327);
xnor UO_732 (O_732,N_47907,N_49703);
xor UO_733 (O_733,N_49765,N_48090);
nor UO_734 (O_734,N_47881,N_48579);
nand UO_735 (O_735,N_47962,N_48617);
or UO_736 (O_736,N_48981,N_48589);
and UO_737 (O_737,N_47910,N_49120);
and UO_738 (O_738,N_48605,N_48146);
and UO_739 (O_739,N_49048,N_48399);
or UO_740 (O_740,N_48119,N_49990);
xnor UO_741 (O_741,N_48180,N_48937);
xnor UO_742 (O_742,N_48535,N_49705);
or UO_743 (O_743,N_49036,N_49102);
or UO_744 (O_744,N_48696,N_48748);
and UO_745 (O_745,N_48096,N_47734);
and UO_746 (O_746,N_49680,N_47603);
nor UO_747 (O_747,N_48221,N_49733);
or UO_748 (O_748,N_48538,N_48890);
nor UO_749 (O_749,N_47961,N_49816);
nand UO_750 (O_750,N_48379,N_48647);
nor UO_751 (O_751,N_48479,N_47827);
or UO_752 (O_752,N_49323,N_48025);
xnor UO_753 (O_753,N_49490,N_47888);
nor UO_754 (O_754,N_48338,N_49700);
xor UO_755 (O_755,N_48578,N_48328);
nand UO_756 (O_756,N_49993,N_49852);
nor UO_757 (O_757,N_49105,N_47675);
nand UO_758 (O_758,N_48896,N_47903);
nor UO_759 (O_759,N_48794,N_47829);
nor UO_760 (O_760,N_47660,N_48282);
and UO_761 (O_761,N_48761,N_49368);
or UO_762 (O_762,N_48949,N_49493);
xor UO_763 (O_763,N_48656,N_48820);
nor UO_764 (O_764,N_48698,N_49599);
or UO_765 (O_765,N_49609,N_47757);
nor UO_766 (O_766,N_49330,N_48465);
nor UO_767 (O_767,N_49375,N_48716);
xor UO_768 (O_768,N_49969,N_47809);
or UO_769 (O_769,N_47791,N_49644);
nand UO_770 (O_770,N_49959,N_47769);
xnor UO_771 (O_771,N_48408,N_48590);
nand UO_772 (O_772,N_48467,N_47930);
nand UO_773 (O_773,N_48377,N_49219);
or UO_774 (O_774,N_49870,N_48859);
or UO_775 (O_775,N_49401,N_47800);
nand UO_776 (O_776,N_48741,N_47766);
nand UO_777 (O_777,N_48682,N_49669);
xnor UO_778 (O_778,N_49895,N_48798);
xor UO_779 (O_779,N_49774,N_48689);
or UO_780 (O_780,N_49837,N_49860);
or UO_781 (O_781,N_49352,N_47978);
nor UO_782 (O_782,N_48699,N_48360);
and UO_783 (O_783,N_48129,N_47656);
nand UO_784 (O_784,N_48784,N_49836);
nand UO_785 (O_785,N_49360,N_48264);
and UO_786 (O_786,N_48914,N_48861);
nand UO_787 (O_787,N_49861,N_49654);
xor UO_788 (O_788,N_47893,N_47994);
nand UO_789 (O_789,N_48422,N_49950);
nand UO_790 (O_790,N_49297,N_48807);
xnor UO_791 (O_791,N_49706,N_48622);
nand UO_792 (O_792,N_48410,N_48672);
xor UO_793 (O_793,N_48115,N_48889);
and UO_794 (O_794,N_49804,N_49235);
nor UO_795 (O_795,N_48999,N_49203);
or UO_796 (O_796,N_49038,N_49121);
xor UO_797 (O_797,N_48956,N_49397);
nor UO_798 (O_798,N_49243,N_47767);
and UO_799 (O_799,N_48655,N_49786);
nand UO_800 (O_800,N_48241,N_48824);
nor UO_801 (O_801,N_49999,N_49844);
xor UO_802 (O_802,N_48848,N_47812);
and UO_803 (O_803,N_48516,N_48095);
xnor UO_804 (O_804,N_49478,N_48459);
nor UO_805 (O_805,N_48950,N_48302);
nand UO_806 (O_806,N_49661,N_48439);
nor UO_807 (O_807,N_47934,N_48786);
or UO_808 (O_808,N_47521,N_47951);
and UO_809 (O_809,N_48857,N_48927);
xor UO_810 (O_810,N_49304,N_47923);
nand UO_811 (O_811,N_48609,N_48089);
nor UO_812 (O_812,N_48235,N_48179);
xnor UO_813 (O_813,N_47635,N_49475);
xor UO_814 (O_814,N_49920,N_47799);
xor UO_815 (O_815,N_48345,N_49303);
and UO_816 (O_816,N_48420,N_47902);
nor UO_817 (O_817,N_49514,N_49942);
and UO_818 (O_818,N_48038,N_48239);
nand UO_819 (O_819,N_48097,N_49709);
xnor UO_820 (O_820,N_48458,N_47662);
nand UO_821 (O_821,N_49430,N_48107);
or UO_822 (O_822,N_49954,N_48121);
xor UO_823 (O_823,N_48975,N_49564);
nor UO_824 (O_824,N_47715,N_48930);
nor UO_825 (O_825,N_49488,N_48050);
nand UO_826 (O_826,N_48009,N_47571);
xor UO_827 (O_827,N_49546,N_48819);
xor UO_828 (O_828,N_48167,N_49080);
nor UO_829 (O_829,N_47615,N_48612);
nor UO_830 (O_830,N_49194,N_49256);
and UO_831 (O_831,N_47578,N_48701);
nand UO_832 (O_832,N_49037,N_48203);
or UO_833 (O_833,N_47708,N_48475);
xnor UO_834 (O_834,N_47824,N_47985);
or UO_835 (O_835,N_48400,N_48310);
nand UO_836 (O_836,N_47970,N_48744);
and UO_837 (O_837,N_48780,N_49742);
and UO_838 (O_838,N_48523,N_47806);
and UO_839 (O_839,N_47928,N_47541);
nor UO_840 (O_840,N_49627,N_49237);
or UO_841 (O_841,N_48910,N_49083);
xor UO_842 (O_842,N_47570,N_48250);
nand UO_843 (O_843,N_49943,N_47697);
nand UO_844 (O_844,N_49697,N_49553);
nand UO_845 (O_845,N_48648,N_49308);
nor UO_846 (O_846,N_48390,N_48139);
nand UO_847 (O_847,N_49499,N_47794);
nor UO_848 (O_848,N_47819,N_48723);
and UO_849 (O_849,N_48634,N_48064);
and UO_850 (O_850,N_47813,N_49292);
and UO_851 (O_851,N_47704,N_49552);
xnor UO_852 (O_852,N_47823,N_47899);
nor UO_853 (O_853,N_48597,N_48011);
xnor UO_854 (O_854,N_47506,N_48238);
and UO_855 (O_855,N_49941,N_49725);
nand UO_856 (O_856,N_48211,N_49018);
or UO_857 (O_857,N_48666,N_48572);
nand UO_858 (O_858,N_49874,N_49095);
xor UO_859 (O_859,N_47914,N_49379);
xnor UO_860 (O_860,N_49952,N_47974);
xor UO_861 (O_861,N_49124,N_48164);
or UO_862 (O_862,N_48210,N_49075);
nor UO_863 (O_863,N_48755,N_49800);
or UO_864 (O_864,N_48781,N_49784);
nand UO_865 (O_865,N_47529,N_49394);
nand UO_866 (O_866,N_48599,N_48335);
or UO_867 (O_867,N_49841,N_48394);
xnor UO_868 (O_868,N_48800,N_47682);
nand UO_869 (O_869,N_49932,N_48217);
nor UO_870 (O_870,N_48362,N_49484);
xnor UO_871 (O_871,N_47655,N_47524);
nor UO_872 (O_872,N_48886,N_49910);
nand UO_873 (O_873,N_48150,N_49828);
nor UO_874 (O_874,N_47543,N_48513);
nand UO_875 (O_875,N_48252,N_49261);
and UO_876 (O_876,N_48263,N_47688);
or UO_877 (O_877,N_47814,N_49770);
or UO_878 (O_878,N_49650,N_47568);
or UO_879 (O_879,N_49006,N_49793);
nand UO_880 (O_880,N_49674,N_48898);
nand UO_881 (O_881,N_49751,N_49808);
nand UO_882 (O_882,N_47598,N_48029);
nor UO_883 (O_883,N_48942,N_48963);
nand UO_884 (O_884,N_49743,N_47954);
or UO_885 (O_885,N_48104,N_49916);
nand UO_886 (O_886,N_47639,N_48754);
and UO_887 (O_887,N_48491,N_48866);
xor UO_888 (O_888,N_48313,N_49218);
nor UO_889 (O_889,N_48635,N_47736);
nor UO_890 (O_890,N_48473,N_47633);
nor UO_891 (O_891,N_48729,N_47765);
and UO_892 (O_892,N_49082,N_48625);
and UO_893 (O_893,N_49200,N_48737);
nand UO_894 (O_894,N_48508,N_49720);
xor UO_895 (O_895,N_47537,N_47554);
nor UO_896 (O_896,N_48255,N_47960);
and UO_897 (O_897,N_48587,N_49137);
or UO_898 (O_898,N_49133,N_47927);
nor UO_899 (O_899,N_49370,N_48447);
nand UO_900 (O_900,N_49541,N_47573);
nand UO_901 (O_901,N_49184,N_47713);
or UO_902 (O_902,N_49850,N_48913);
or UO_903 (O_903,N_48106,N_49244);
or UO_904 (O_904,N_49965,N_48195);
or UO_905 (O_905,N_49554,N_49349);
or UO_906 (O_906,N_49306,N_48749);
nand UO_907 (O_907,N_49472,N_47958);
nor UO_908 (O_908,N_48860,N_48188);
xor UO_909 (O_909,N_49239,N_49181);
nor UO_910 (O_910,N_47514,N_48563);
nor UO_911 (O_911,N_49043,N_49652);
nand UO_912 (O_912,N_48830,N_49335);
nor UO_913 (O_913,N_48971,N_48482);
and UO_914 (O_914,N_48354,N_49819);
or UO_915 (O_915,N_49649,N_48435);
nand UO_916 (O_916,N_47518,N_47680);
xnor UO_917 (O_917,N_49012,N_49089);
or UO_918 (O_918,N_49632,N_48190);
xor UO_919 (O_919,N_49676,N_48368);
and UO_920 (O_920,N_47871,N_48366);
nor UO_921 (O_921,N_48124,N_48740);
nand UO_922 (O_922,N_47946,N_49994);
nand UO_923 (O_923,N_48502,N_48047);
or UO_924 (O_924,N_47730,N_48883);
or UO_925 (O_925,N_48133,N_47664);
nor UO_926 (O_926,N_49274,N_49951);
nand UO_927 (O_927,N_49449,N_48054);
and UO_928 (O_928,N_48055,N_47594);
nor UO_929 (O_929,N_49188,N_49796);
and UO_930 (O_930,N_49562,N_49019);
nand UO_931 (O_931,N_48196,N_48027);
nand UO_932 (O_932,N_48393,N_49905);
nor UO_933 (O_933,N_48770,N_49892);
and UO_934 (O_934,N_49780,N_47601);
or UO_935 (O_935,N_49960,N_49511);
and UO_936 (O_936,N_47592,N_49023);
nor UO_937 (O_937,N_49759,N_48357);
nand UO_938 (O_938,N_47679,N_49199);
nor UO_939 (O_939,N_49660,N_47685);
nand UO_940 (O_940,N_48858,N_49775);
and UO_941 (O_941,N_47787,N_48992);
nor UO_942 (O_942,N_47563,N_48598);
xor UO_943 (O_943,N_48946,N_47999);
nor UO_944 (O_944,N_48775,N_48415);
nor UO_945 (O_945,N_48219,N_47619);
xor UO_946 (O_946,N_49249,N_49947);
nor UO_947 (O_947,N_48084,N_48813);
nor UO_948 (O_948,N_49538,N_49044);
xor UO_949 (O_949,N_49020,N_48189);
xor UO_950 (O_950,N_49755,N_48823);
nor UO_951 (O_951,N_49495,N_47505);
xnor UO_952 (O_952,N_48793,N_49372);
or UO_953 (O_953,N_48008,N_49412);
nand UO_954 (O_954,N_48451,N_48639);
nor UO_955 (O_955,N_49917,N_49029);
or UO_956 (O_956,N_47727,N_49967);
xor UO_957 (O_957,N_47555,N_48454);
or UO_958 (O_958,N_49356,N_47669);
and UO_959 (O_959,N_48430,N_48663);
xor UO_960 (O_960,N_48365,N_48779);
xnor UO_961 (O_961,N_48607,N_49726);
nand UO_962 (O_962,N_47666,N_49252);
nand UO_963 (O_963,N_48671,N_48409);
or UO_964 (O_964,N_48899,N_48649);
and UO_965 (O_965,N_49651,N_48080);
nand UO_966 (O_966,N_49732,N_49284);
and UO_967 (O_967,N_49267,N_49317);
nor UO_968 (O_968,N_48496,N_48845);
nand UO_969 (O_969,N_49971,N_49556);
xor UO_970 (O_970,N_47852,N_47964);
nand UO_971 (O_971,N_48258,N_49005);
xor UO_972 (O_972,N_48244,N_48312);
or UO_973 (O_973,N_49789,N_48066);
nand UO_974 (O_974,N_49573,N_49996);
nor UO_975 (O_975,N_47801,N_48642);
or UO_976 (O_976,N_47784,N_48849);
and UO_977 (O_977,N_48626,N_48192);
and UO_978 (O_978,N_47975,N_49877);
xor UO_979 (O_979,N_48878,N_49277);
nand UO_980 (O_980,N_48727,N_48827);
xor UO_981 (O_981,N_49096,N_48989);
or UO_982 (O_982,N_47611,N_47883);
nor UO_983 (O_983,N_48202,N_49957);
or UO_984 (O_984,N_49111,N_49302);
or UO_985 (O_985,N_49047,N_49332);
xnor UO_986 (O_986,N_49699,N_48456);
xor UO_987 (O_987,N_49071,N_47552);
and UO_988 (O_988,N_47921,N_49336);
nor UO_989 (O_989,N_48714,N_48684);
nor UO_990 (O_990,N_47575,N_49287);
and UO_991 (O_991,N_48023,N_48348);
nand UO_992 (O_992,N_49130,N_49359);
or UO_993 (O_993,N_49618,N_48330);
and UO_994 (O_994,N_47972,N_48894);
or UO_995 (O_995,N_48487,N_48374);
nand UO_996 (O_996,N_49871,N_49389);
nor UO_997 (O_997,N_47651,N_47723);
xnor UO_998 (O_998,N_48662,N_49078);
and UO_999 (O_999,N_48733,N_49241);
or UO_1000 (O_1000,N_48585,N_47777);
xnor UO_1001 (O_1001,N_48833,N_48850);
and UO_1002 (O_1002,N_48994,N_48484);
nand UO_1003 (O_1003,N_49238,N_47591);
nor UO_1004 (O_1004,N_49645,N_48505);
xnor UO_1005 (O_1005,N_49363,N_47582);
nand UO_1006 (O_1006,N_49145,N_48991);
and UO_1007 (O_1007,N_47560,N_48730);
nor UO_1008 (O_1008,N_47658,N_49035);
or UO_1009 (O_1009,N_48279,N_49309);
nor UO_1010 (O_1010,N_48745,N_48303);
xnor UO_1011 (O_1011,N_49504,N_49882);
xor UO_1012 (O_1012,N_47673,N_49424);
and UO_1013 (O_1013,N_49288,N_49953);
xor UO_1014 (O_1014,N_47650,N_49459);
or UO_1015 (O_1015,N_48602,N_48812);
or UO_1016 (O_1016,N_48317,N_47880);
nor UO_1017 (O_1017,N_49215,N_49756);
nand UO_1018 (O_1018,N_48608,N_48654);
nand UO_1019 (O_1019,N_48304,N_47760);
nand UO_1020 (O_1020,N_49017,N_49425);
nor UO_1021 (O_1021,N_47559,N_49172);
or UO_1022 (O_1022,N_47868,N_48087);
nor UO_1023 (O_1023,N_48619,N_48476);
nor UO_1024 (O_1024,N_49259,N_48582);
nand UO_1025 (O_1025,N_48483,N_48876);
xor UO_1026 (O_1026,N_47862,N_48687);
nand UO_1027 (O_1027,N_49972,N_49376);
and UO_1028 (O_1028,N_49211,N_47943);
xor UO_1029 (O_1029,N_49409,N_48509);
nor UO_1030 (O_1030,N_47825,N_49857);
nor UO_1031 (O_1031,N_47885,N_49098);
nor UO_1032 (O_1032,N_48685,N_47786);
and UO_1033 (O_1033,N_49198,N_48174);
and UO_1034 (O_1034,N_48148,N_47772);
and UO_1035 (O_1035,N_49343,N_48561);
nand UO_1036 (O_1036,N_47875,N_48453);
nand UO_1037 (O_1037,N_49110,N_48332);
nor UO_1038 (O_1038,N_48109,N_49266);
or UO_1039 (O_1039,N_47808,N_48253);
and UO_1040 (O_1040,N_49760,N_48086);
and UO_1041 (O_1041,N_48350,N_49730);
or UO_1042 (O_1042,N_49042,N_49619);
and UO_1043 (O_1043,N_48370,N_48206);
or UO_1044 (O_1044,N_49458,N_49033);
xor UO_1045 (O_1045,N_47751,N_48123);
or UO_1046 (O_1046,N_48892,N_48962);
or UO_1047 (O_1047,N_48110,N_47500);
and UO_1048 (O_1048,N_47864,N_47587);
and UO_1049 (O_1049,N_49946,N_48815);
nor UO_1050 (O_1050,N_49076,N_49126);
and UO_1051 (O_1051,N_47683,N_49117);
nor UO_1052 (O_1052,N_48789,N_48421);
nand UO_1053 (O_1053,N_47844,N_49708);
nor UO_1054 (O_1054,N_49060,N_47561);
nor UO_1055 (O_1055,N_49069,N_48782);
nand UO_1056 (O_1056,N_49142,N_47779);
nor UO_1057 (O_1057,N_49151,N_48028);
or UO_1058 (O_1058,N_47865,N_47965);
nor UO_1059 (O_1059,N_49980,N_48347);
and UO_1060 (O_1060,N_47531,N_48272);
or UO_1061 (O_1061,N_48627,N_48222);
or UO_1062 (O_1062,N_49873,N_49840);
xnor UO_1063 (O_1063,N_48558,N_49702);
and UO_1064 (O_1064,N_48032,N_49340);
or UO_1065 (O_1065,N_48378,N_48939);
xor UO_1066 (O_1066,N_48778,N_49798);
nand UO_1067 (O_1067,N_48863,N_47712);
nand UO_1068 (O_1068,N_48030,N_48091);
xor UO_1069 (O_1069,N_49015,N_49100);
nor UO_1070 (O_1070,N_48854,N_48071);
or UO_1071 (O_1071,N_47936,N_49587);
xor UO_1072 (O_1072,N_49689,N_48170);
nor UO_1073 (O_1073,N_49161,N_48732);
nor UO_1074 (O_1074,N_49893,N_48046);
and UO_1075 (O_1075,N_48406,N_47532);
nand UO_1076 (O_1076,N_49432,N_47580);
or UO_1077 (O_1077,N_47759,N_48556);
xnor UO_1078 (O_1078,N_47866,N_47684);
nand UO_1079 (O_1079,N_48592,N_48902);
and UO_1080 (O_1080,N_49582,N_48051);
or UO_1081 (O_1081,N_47782,N_47599);
and UO_1082 (O_1082,N_47959,N_49884);
and UO_1083 (O_1083,N_48214,N_48825);
or UO_1084 (O_1084,N_48373,N_48276);
or UO_1085 (O_1085,N_48688,N_48315);
or UO_1086 (O_1086,N_48856,N_47596);
xor UO_1087 (O_1087,N_49206,N_49936);
nor UO_1088 (O_1088,N_48226,N_49470);
or UO_1089 (O_1089,N_47857,N_47775);
nor UO_1090 (O_1090,N_49431,N_49925);
and UO_1091 (O_1091,N_47774,N_49224);
xor UO_1092 (O_1092,N_48580,N_48606);
nor UO_1093 (O_1093,N_48440,N_49092);
and UO_1094 (O_1094,N_48767,N_48443);
and UO_1095 (O_1095,N_49868,N_49915);
nor UO_1096 (O_1096,N_49031,N_49164);
nor UO_1097 (O_1097,N_48641,N_49280);
xor UO_1098 (O_1098,N_49053,N_47979);
nand UO_1099 (O_1099,N_48924,N_47623);
and UO_1100 (O_1100,N_47574,N_49312);
or UO_1101 (O_1101,N_49506,N_48062);
nand UO_1102 (O_1102,N_49205,N_49344);
and UO_1103 (O_1103,N_47718,N_47605);
nor UO_1104 (O_1104,N_49410,N_47743);
nor UO_1105 (O_1105,N_49670,N_48274);
or UO_1106 (O_1106,N_47850,N_49264);
nor UO_1107 (O_1107,N_49536,N_48257);
nor UO_1108 (O_1108,N_49159,N_49004);
or UO_1109 (O_1109,N_49066,N_49672);
or UO_1110 (O_1110,N_47859,N_47989);
nor UO_1111 (O_1111,N_49190,N_48530);
and UO_1112 (O_1112,N_49466,N_49223);
and UO_1113 (O_1113,N_49009,N_47854);
and UO_1114 (O_1114,N_49518,N_48380);
xnor UO_1115 (O_1115,N_49427,N_48972);
and UO_1116 (O_1116,N_48547,N_48070);
xnor UO_1117 (O_1117,N_49531,N_48799);
nor UO_1118 (O_1118,N_49544,N_49196);
nor UO_1119 (O_1119,N_47707,N_48934);
and UO_1120 (O_1120,N_47694,N_49677);
xnor UO_1121 (O_1121,N_48545,N_48901);
nor UO_1122 (O_1122,N_49955,N_48060);
or UO_1123 (O_1123,N_48821,N_49795);
xor UO_1124 (O_1124,N_49051,N_48384);
nor UO_1125 (O_1125,N_49615,N_47998);
nor UO_1126 (O_1126,N_49054,N_48130);
or UO_1127 (O_1127,N_49913,N_49329);
nand UO_1128 (O_1128,N_47687,N_49482);
and UO_1129 (O_1129,N_48024,N_48488);
and UO_1130 (O_1130,N_47716,N_49678);
and UO_1131 (O_1131,N_47986,N_49600);
xor UO_1132 (O_1132,N_48709,N_49718);
nand UO_1133 (O_1133,N_47501,N_48593);
xnor UO_1134 (O_1134,N_49501,N_48810);
nor UO_1135 (O_1135,N_48817,N_47572);
nand UO_1136 (O_1136,N_47981,N_48113);
or UO_1137 (O_1137,N_48554,N_49731);
xor UO_1138 (O_1138,N_49578,N_47625);
nor UO_1139 (O_1139,N_47746,N_47621);
and UO_1140 (O_1140,N_49122,N_48099);
nand UO_1141 (O_1141,N_49580,N_48288);
nand UO_1142 (O_1142,N_49817,N_49829);
nor UO_1143 (O_1143,N_49328,N_48573);
nor UO_1144 (O_1144,N_48147,N_47944);
xnor UO_1145 (O_1145,N_48507,N_48574);
nand UO_1146 (O_1146,N_49958,N_49889);
and UO_1147 (O_1147,N_48544,N_48659);
nand UO_1148 (O_1148,N_47790,N_48155);
xor UO_1149 (O_1149,N_48702,N_49899);
nand UO_1150 (O_1150,N_48965,N_48353);
nand UO_1151 (O_1151,N_47804,N_47988);
nor UO_1152 (O_1152,N_48774,N_48305);
xor UO_1153 (O_1153,N_48615,N_47805);
or UO_1154 (O_1154,N_47874,N_47710);
or UO_1155 (O_1155,N_47926,N_49174);
nand UO_1156 (O_1156,N_49982,N_47755);
nand UO_1157 (O_1157,N_47842,N_47783);
nor UO_1158 (O_1158,N_48455,N_48049);
nor UO_1159 (O_1159,N_48185,N_49757);
or UO_1160 (O_1160,N_49258,N_49413);
or UO_1161 (O_1161,N_49073,N_47873);
nand UO_1162 (O_1162,N_49686,N_49968);
or UO_1163 (O_1163,N_48522,N_48980);
nand UO_1164 (O_1164,N_47699,N_47562);
nand UO_1165 (O_1165,N_48553,N_48001);
xnor UO_1166 (O_1166,N_48015,N_47849);
nand UO_1167 (O_1167,N_49311,N_49904);
nand UO_1168 (O_1168,N_48061,N_49956);
and UO_1169 (O_1169,N_49090,N_48401);
nor UO_1170 (O_1170,N_48758,N_48503);
nor UO_1171 (O_1171,N_49545,N_49635);
xor UO_1172 (O_1172,N_49327,N_48324);
nand UO_1173 (O_1173,N_48600,N_48126);
nor UO_1174 (O_1174,N_48457,N_49534);
xnor UO_1175 (O_1175,N_49183,N_49707);
nand UO_1176 (O_1176,N_48637,N_49771);
or UO_1177 (O_1177,N_47863,N_48591);
xor UO_1178 (O_1178,N_49216,N_47547);
or UO_1179 (O_1179,N_49821,N_48611);
xor UO_1180 (O_1180,N_48306,N_49077);
and UO_1181 (O_1181,N_49002,N_49154);
xor UO_1182 (O_1182,N_47992,N_49052);
or UO_1183 (O_1183,N_48916,N_49694);
and UO_1184 (O_1184,N_48042,N_49530);
nor UO_1185 (O_1185,N_48583,N_49690);
xor UO_1186 (O_1186,N_49113,N_47644);
nor UO_1187 (O_1187,N_49809,N_47762);
or UO_1188 (O_1188,N_47602,N_48118);
or UO_1189 (O_1189,N_48985,N_47647);
nand UO_1190 (O_1190,N_48581,N_48340);
nor UO_1191 (O_1191,N_47816,N_48474);
or UO_1192 (O_1192,N_47963,N_48122);
and UO_1193 (O_1193,N_49446,N_49591);
nand UO_1194 (O_1194,N_48322,N_48908);
nand UO_1195 (O_1195,N_48964,N_49512);
nand UO_1196 (O_1196,N_47826,N_49438);
nand UO_1197 (O_1197,N_48533,N_48372);
and UO_1198 (O_1198,N_47933,N_47667);
or UO_1199 (O_1199,N_48391,N_48389);
xnor UO_1200 (O_1200,N_47971,N_48918);
nand UO_1201 (O_1201,N_49811,N_49846);
and UO_1202 (O_1202,N_49606,N_49378);
or UO_1203 (O_1203,N_48933,N_49524);
nor UO_1204 (O_1204,N_49543,N_48329);
nor UO_1205 (O_1205,N_49480,N_49429);
and UO_1206 (O_1206,N_47803,N_49173);
xnor UO_1207 (O_1207,N_49933,N_47756);
or UO_1208 (O_1208,N_47629,N_49115);
and UO_1209 (O_1209,N_47519,N_48703);
and UO_1210 (O_1210,N_49864,N_48283);
nand UO_1211 (O_1211,N_48504,N_48452);
nor UO_1212 (O_1212,N_49721,N_47834);
nor UO_1213 (O_1213,N_48300,N_48631);
nand UO_1214 (O_1214,N_47966,N_48925);
nand UO_1215 (O_1215,N_48261,N_48996);
nor UO_1216 (O_1216,N_49024,N_49851);
xor UO_1217 (O_1217,N_48320,N_49250);
nor UO_1218 (O_1218,N_49217,N_47848);
or UO_1219 (O_1219,N_49185,N_49290);
xor UO_1220 (O_1220,N_49278,N_49926);
xnor UO_1221 (O_1221,N_49572,N_49214);
nor UO_1222 (O_1222,N_49163,N_47845);
nand UO_1223 (O_1223,N_49474,N_48232);
nor UO_1224 (O_1224,N_47968,N_48546);
or UO_1225 (O_1225,N_47948,N_49457);
xnor UO_1226 (O_1226,N_48225,N_49575);
nand UO_1227 (O_1227,N_48460,N_48478);
xnor UO_1228 (O_1228,N_48290,N_48412);
nor UO_1229 (O_1229,N_49168,N_47785);
or UO_1230 (O_1230,N_48265,N_47569);
nand UO_1231 (O_1231,N_49681,N_49736);
and UO_1232 (O_1232,N_49973,N_48882);
nor UO_1233 (O_1233,N_48945,N_49979);
and UO_1234 (O_1234,N_49213,N_49711);
or UO_1235 (O_1235,N_49978,N_49382);
or UO_1236 (O_1236,N_49613,N_47608);
and UO_1237 (O_1237,N_49167,N_47810);
nand UO_1238 (O_1238,N_47942,N_49125);
nor UO_1239 (O_1239,N_48308,N_49381);
nor UO_1240 (O_1240,N_48176,N_48841);
xnor UO_1241 (O_1241,N_49679,N_49831);
nand UO_1242 (O_1242,N_49897,N_49132);
xnor UO_1243 (O_1243,N_49153,N_48877);
or UO_1244 (O_1244,N_47728,N_49716);
nor UO_1245 (O_1245,N_49403,N_48571);
or UO_1246 (O_1246,N_49888,N_48549);
xor UO_1247 (O_1247,N_49193,N_49014);
xnor UO_1248 (O_1248,N_47977,N_49663);
nor UO_1249 (O_1249,N_48493,N_48131);
or UO_1250 (O_1250,N_47518,N_49468);
nand UO_1251 (O_1251,N_49413,N_48426);
or UO_1252 (O_1252,N_48252,N_49941);
and UO_1253 (O_1253,N_48575,N_47795);
or UO_1254 (O_1254,N_47745,N_48572);
nor UO_1255 (O_1255,N_49103,N_49426);
xor UO_1256 (O_1256,N_48632,N_48622);
xnor UO_1257 (O_1257,N_47507,N_49612);
and UO_1258 (O_1258,N_48300,N_48362);
or UO_1259 (O_1259,N_48259,N_47954);
and UO_1260 (O_1260,N_49446,N_49824);
or UO_1261 (O_1261,N_47598,N_47501);
or UO_1262 (O_1262,N_48447,N_49798);
or UO_1263 (O_1263,N_49854,N_48897);
nor UO_1264 (O_1264,N_47939,N_48676);
or UO_1265 (O_1265,N_49377,N_49199);
nand UO_1266 (O_1266,N_47681,N_49358);
nor UO_1267 (O_1267,N_47883,N_48453);
nor UO_1268 (O_1268,N_48623,N_49882);
nor UO_1269 (O_1269,N_48651,N_49335);
or UO_1270 (O_1270,N_49901,N_48901);
and UO_1271 (O_1271,N_47687,N_47806);
nand UO_1272 (O_1272,N_49090,N_48861);
nand UO_1273 (O_1273,N_49125,N_49789);
and UO_1274 (O_1274,N_49024,N_48150);
and UO_1275 (O_1275,N_48680,N_49843);
nor UO_1276 (O_1276,N_49371,N_48635);
and UO_1277 (O_1277,N_47677,N_48969);
or UO_1278 (O_1278,N_48889,N_49430);
nand UO_1279 (O_1279,N_49576,N_47633);
or UO_1280 (O_1280,N_49349,N_48711);
or UO_1281 (O_1281,N_48356,N_49421);
nand UO_1282 (O_1282,N_47675,N_47622);
nand UO_1283 (O_1283,N_49872,N_49398);
nand UO_1284 (O_1284,N_48963,N_49980);
nand UO_1285 (O_1285,N_49884,N_48768);
xnor UO_1286 (O_1286,N_49432,N_48967);
and UO_1287 (O_1287,N_47951,N_48681);
xor UO_1288 (O_1288,N_47864,N_48610);
nand UO_1289 (O_1289,N_49201,N_47832);
xnor UO_1290 (O_1290,N_48263,N_47757);
or UO_1291 (O_1291,N_49037,N_48932);
and UO_1292 (O_1292,N_48764,N_49004);
nand UO_1293 (O_1293,N_48332,N_49555);
and UO_1294 (O_1294,N_48662,N_49782);
xnor UO_1295 (O_1295,N_48708,N_48374);
nand UO_1296 (O_1296,N_48945,N_49234);
and UO_1297 (O_1297,N_48305,N_49253);
or UO_1298 (O_1298,N_47811,N_49398);
nor UO_1299 (O_1299,N_48391,N_48899);
or UO_1300 (O_1300,N_49473,N_49761);
and UO_1301 (O_1301,N_49384,N_48301);
and UO_1302 (O_1302,N_49620,N_48567);
and UO_1303 (O_1303,N_49305,N_48742);
and UO_1304 (O_1304,N_47535,N_49636);
nor UO_1305 (O_1305,N_49962,N_47894);
nor UO_1306 (O_1306,N_48014,N_48900);
and UO_1307 (O_1307,N_49134,N_48035);
or UO_1308 (O_1308,N_48612,N_49461);
or UO_1309 (O_1309,N_48528,N_48608);
and UO_1310 (O_1310,N_47821,N_48425);
nor UO_1311 (O_1311,N_49341,N_49136);
and UO_1312 (O_1312,N_49733,N_48189);
nor UO_1313 (O_1313,N_49502,N_48359);
and UO_1314 (O_1314,N_49690,N_49532);
or UO_1315 (O_1315,N_48874,N_49667);
xnor UO_1316 (O_1316,N_47811,N_49093);
and UO_1317 (O_1317,N_47865,N_49446);
and UO_1318 (O_1318,N_48788,N_47917);
xnor UO_1319 (O_1319,N_48101,N_48020);
nor UO_1320 (O_1320,N_49413,N_49475);
xnor UO_1321 (O_1321,N_49100,N_49469);
nor UO_1322 (O_1322,N_49142,N_47595);
or UO_1323 (O_1323,N_49494,N_49733);
or UO_1324 (O_1324,N_49784,N_48162);
nand UO_1325 (O_1325,N_49888,N_48080);
nand UO_1326 (O_1326,N_49585,N_49073);
xnor UO_1327 (O_1327,N_47699,N_49094);
and UO_1328 (O_1328,N_48816,N_49699);
and UO_1329 (O_1329,N_49669,N_49812);
nand UO_1330 (O_1330,N_47635,N_48120);
or UO_1331 (O_1331,N_48728,N_47637);
xnor UO_1332 (O_1332,N_47739,N_49733);
xnor UO_1333 (O_1333,N_48900,N_49307);
or UO_1334 (O_1334,N_48392,N_49606);
nand UO_1335 (O_1335,N_48814,N_48315);
nand UO_1336 (O_1336,N_47862,N_49725);
and UO_1337 (O_1337,N_47570,N_48571);
nand UO_1338 (O_1338,N_47645,N_49320);
and UO_1339 (O_1339,N_49977,N_49217);
nor UO_1340 (O_1340,N_49121,N_49670);
or UO_1341 (O_1341,N_48488,N_48896);
nand UO_1342 (O_1342,N_48085,N_48020);
and UO_1343 (O_1343,N_48526,N_49565);
xor UO_1344 (O_1344,N_48526,N_49246);
xnor UO_1345 (O_1345,N_49341,N_49914);
nand UO_1346 (O_1346,N_48518,N_48875);
and UO_1347 (O_1347,N_49211,N_48154);
and UO_1348 (O_1348,N_49758,N_48282);
xor UO_1349 (O_1349,N_48801,N_48935);
nor UO_1350 (O_1350,N_47985,N_48421);
nand UO_1351 (O_1351,N_49894,N_48723);
xnor UO_1352 (O_1352,N_48729,N_49192);
nor UO_1353 (O_1353,N_48097,N_47669);
and UO_1354 (O_1354,N_49756,N_49924);
and UO_1355 (O_1355,N_49289,N_48219);
and UO_1356 (O_1356,N_48850,N_48101);
or UO_1357 (O_1357,N_47990,N_47982);
nor UO_1358 (O_1358,N_49267,N_49385);
xnor UO_1359 (O_1359,N_47819,N_49085);
xnor UO_1360 (O_1360,N_48732,N_48760);
and UO_1361 (O_1361,N_48416,N_47726);
xnor UO_1362 (O_1362,N_48920,N_47808);
or UO_1363 (O_1363,N_49881,N_49747);
or UO_1364 (O_1364,N_47678,N_47911);
nor UO_1365 (O_1365,N_48848,N_49059);
or UO_1366 (O_1366,N_49584,N_49187);
xnor UO_1367 (O_1367,N_49835,N_49076);
and UO_1368 (O_1368,N_49210,N_48063);
nor UO_1369 (O_1369,N_49640,N_48683);
nor UO_1370 (O_1370,N_49775,N_48423);
nor UO_1371 (O_1371,N_49534,N_48957);
and UO_1372 (O_1372,N_48036,N_48912);
and UO_1373 (O_1373,N_47750,N_49950);
and UO_1374 (O_1374,N_49382,N_48546);
xor UO_1375 (O_1375,N_48224,N_48722);
xor UO_1376 (O_1376,N_47561,N_48255);
and UO_1377 (O_1377,N_47514,N_48511);
xor UO_1378 (O_1378,N_49303,N_48962);
or UO_1379 (O_1379,N_48154,N_48551);
and UO_1380 (O_1380,N_49253,N_49491);
or UO_1381 (O_1381,N_49433,N_49652);
nand UO_1382 (O_1382,N_47791,N_49310);
xnor UO_1383 (O_1383,N_49460,N_48353);
xnor UO_1384 (O_1384,N_47605,N_47678);
and UO_1385 (O_1385,N_49172,N_49508);
nor UO_1386 (O_1386,N_49594,N_49940);
or UO_1387 (O_1387,N_48216,N_47794);
nor UO_1388 (O_1388,N_48789,N_47760);
nand UO_1389 (O_1389,N_49370,N_49810);
or UO_1390 (O_1390,N_48575,N_47586);
xnor UO_1391 (O_1391,N_49979,N_47528);
and UO_1392 (O_1392,N_47530,N_47825);
or UO_1393 (O_1393,N_49193,N_47540);
nand UO_1394 (O_1394,N_48055,N_48658);
xnor UO_1395 (O_1395,N_47956,N_48786);
or UO_1396 (O_1396,N_47519,N_47903);
or UO_1397 (O_1397,N_49829,N_49588);
xnor UO_1398 (O_1398,N_48975,N_49816);
or UO_1399 (O_1399,N_48166,N_48969);
and UO_1400 (O_1400,N_47979,N_48687);
xnor UO_1401 (O_1401,N_49310,N_49366);
and UO_1402 (O_1402,N_49322,N_49642);
nor UO_1403 (O_1403,N_49655,N_49487);
nand UO_1404 (O_1404,N_47566,N_49788);
or UO_1405 (O_1405,N_48692,N_47961);
xnor UO_1406 (O_1406,N_48452,N_48050);
or UO_1407 (O_1407,N_47948,N_47751);
nand UO_1408 (O_1408,N_48094,N_48842);
xor UO_1409 (O_1409,N_48673,N_47803);
nand UO_1410 (O_1410,N_47807,N_48971);
or UO_1411 (O_1411,N_48259,N_49869);
xor UO_1412 (O_1412,N_48068,N_49754);
nor UO_1413 (O_1413,N_48704,N_48002);
nand UO_1414 (O_1414,N_48432,N_49344);
and UO_1415 (O_1415,N_48169,N_48441);
and UO_1416 (O_1416,N_49158,N_49996);
xor UO_1417 (O_1417,N_49589,N_49316);
xnor UO_1418 (O_1418,N_49415,N_49007);
or UO_1419 (O_1419,N_49324,N_47679);
nand UO_1420 (O_1420,N_49341,N_49435);
nor UO_1421 (O_1421,N_49382,N_48014);
nand UO_1422 (O_1422,N_48181,N_48936);
nand UO_1423 (O_1423,N_48897,N_49091);
xor UO_1424 (O_1424,N_47765,N_49203);
nand UO_1425 (O_1425,N_49676,N_48945);
xnor UO_1426 (O_1426,N_48837,N_47713);
nor UO_1427 (O_1427,N_49439,N_48328);
nand UO_1428 (O_1428,N_48888,N_49935);
and UO_1429 (O_1429,N_48761,N_49091);
nand UO_1430 (O_1430,N_49976,N_48823);
nand UO_1431 (O_1431,N_47582,N_48041);
nor UO_1432 (O_1432,N_49882,N_49148);
xor UO_1433 (O_1433,N_49727,N_48765);
or UO_1434 (O_1434,N_48309,N_48574);
and UO_1435 (O_1435,N_49066,N_49663);
or UO_1436 (O_1436,N_48051,N_48583);
and UO_1437 (O_1437,N_48684,N_48091);
nor UO_1438 (O_1438,N_48605,N_48925);
and UO_1439 (O_1439,N_49244,N_48883);
nand UO_1440 (O_1440,N_49390,N_47914);
nor UO_1441 (O_1441,N_49698,N_47812);
xnor UO_1442 (O_1442,N_48096,N_47518);
xnor UO_1443 (O_1443,N_49278,N_48740);
or UO_1444 (O_1444,N_48062,N_47972);
xnor UO_1445 (O_1445,N_48317,N_49479);
nor UO_1446 (O_1446,N_48609,N_48093);
xnor UO_1447 (O_1447,N_47966,N_47949);
or UO_1448 (O_1448,N_49109,N_48298);
nor UO_1449 (O_1449,N_47769,N_48459);
xnor UO_1450 (O_1450,N_49262,N_48195);
or UO_1451 (O_1451,N_48470,N_48748);
or UO_1452 (O_1452,N_49240,N_49476);
xnor UO_1453 (O_1453,N_48113,N_49486);
nor UO_1454 (O_1454,N_49880,N_49636);
or UO_1455 (O_1455,N_47604,N_49137);
and UO_1456 (O_1456,N_48793,N_48588);
or UO_1457 (O_1457,N_49176,N_49076);
or UO_1458 (O_1458,N_47522,N_48697);
or UO_1459 (O_1459,N_49943,N_49799);
and UO_1460 (O_1460,N_49385,N_49817);
nand UO_1461 (O_1461,N_48014,N_47906);
xor UO_1462 (O_1462,N_49481,N_48373);
and UO_1463 (O_1463,N_47736,N_49427);
or UO_1464 (O_1464,N_48870,N_48108);
and UO_1465 (O_1465,N_49158,N_47773);
and UO_1466 (O_1466,N_47905,N_48485);
and UO_1467 (O_1467,N_47615,N_47519);
nor UO_1468 (O_1468,N_48882,N_49645);
and UO_1469 (O_1469,N_49021,N_47948);
and UO_1470 (O_1470,N_48623,N_47898);
or UO_1471 (O_1471,N_49193,N_49191);
and UO_1472 (O_1472,N_48724,N_47586);
nor UO_1473 (O_1473,N_49731,N_47539);
and UO_1474 (O_1474,N_49970,N_48351);
xor UO_1475 (O_1475,N_48835,N_48589);
or UO_1476 (O_1476,N_47522,N_49986);
xnor UO_1477 (O_1477,N_48992,N_49246);
or UO_1478 (O_1478,N_48056,N_49090);
and UO_1479 (O_1479,N_47640,N_49867);
nor UO_1480 (O_1480,N_48383,N_48390);
xnor UO_1481 (O_1481,N_49622,N_49551);
nor UO_1482 (O_1482,N_47691,N_49308);
and UO_1483 (O_1483,N_49657,N_49156);
xnor UO_1484 (O_1484,N_48733,N_48888);
xor UO_1485 (O_1485,N_48256,N_49351);
or UO_1486 (O_1486,N_48979,N_48356);
and UO_1487 (O_1487,N_49885,N_47917);
xor UO_1488 (O_1488,N_47755,N_48544);
nor UO_1489 (O_1489,N_48549,N_48303);
xnor UO_1490 (O_1490,N_48316,N_49916);
nand UO_1491 (O_1491,N_49057,N_47542);
and UO_1492 (O_1492,N_48172,N_49595);
or UO_1493 (O_1493,N_48537,N_48203);
and UO_1494 (O_1494,N_48219,N_49753);
and UO_1495 (O_1495,N_49437,N_48951);
nand UO_1496 (O_1496,N_48845,N_48435);
or UO_1497 (O_1497,N_48608,N_49578);
xnor UO_1498 (O_1498,N_48640,N_49408);
nand UO_1499 (O_1499,N_49525,N_48374);
or UO_1500 (O_1500,N_47502,N_49777);
or UO_1501 (O_1501,N_48653,N_47719);
nand UO_1502 (O_1502,N_49589,N_47635);
nor UO_1503 (O_1503,N_49092,N_47801);
nor UO_1504 (O_1504,N_48222,N_48753);
nand UO_1505 (O_1505,N_48411,N_48999);
nor UO_1506 (O_1506,N_49844,N_47590);
and UO_1507 (O_1507,N_48723,N_48936);
or UO_1508 (O_1508,N_49449,N_49689);
and UO_1509 (O_1509,N_49938,N_49658);
nand UO_1510 (O_1510,N_48451,N_48083);
and UO_1511 (O_1511,N_49578,N_49445);
nand UO_1512 (O_1512,N_47715,N_49797);
nand UO_1513 (O_1513,N_49867,N_48008);
nand UO_1514 (O_1514,N_47889,N_47718);
nor UO_1515 (O_1515,N_49255,N_47796);
nor UO_1516 (O_1516,N_49795,N_48687);
or UO_1517 (O_1517,N_48114,N_48202);
nand UO_1518 (O_1518,N_48256,N_48597);
nand UO_1519 (O_1519,N_47976,N_47790);
nor UO_1520 (O_1520,N_48283,N_48446);
xnor UO_1521 (O_1521,N_47988,N_47726);
and UO_1522 (O_1522,N_49036,N_48891);
xor UO_1523 (O_1523,N_47939,N_48506);
nand UO_1524 (O_1524,N_47717,N_48108);
or UO_1525 (O_1525,N_49252,N_47779);
and UO_1526 (O_1526,N_49783,N_48742);
nand UO_1527 (O_1527,N_48721,N_49583);
nand UO_1528 (O_1528,N_49633,N_49302);
nand UO_1529 (O_1529,N_48438,N_48478);
and UO_1530 (O_1530,N_48555,N_48450);
xor UO_1531 (O_1531,N_47824,N_48159);
and UO_1532 (O_1532,N_47540,N_48734);
and UO_1533 (O_1533,N_48211,N_47804);
xor UO_1534 (O_1534,N_47726,N_49448);
and UO_1535 (O_1535,N_47655,N_47554);
and UO_1536 (O_1536,N_49900,N_49845);
nor UO_1537 (O_1537,N_49555,N_49081);
nor UO_1538 (O_1538,N_48354,N_49776);
and UO_1539 (O_1539,N_47838,N_48746);
nand UO_1540 (O_1540,N_49554,N_48862);
xnor UO_1541 (O_1541,N_49158,N_48924);
and UO_1542 (O_1542,N_49878,N_49678);
nand UO_1543 (O_1543,N_47504,N_49120);
nor UO_1544 (O_1544,N_49417,N_47516);
nor UO_1545 (O_1545,N_48475,N_48276);
nor UO_1546 (O_1546,N_47677,N_49531);
xnor UO_1547 (O_1547,N_49145,N_49285);
nand UO_1548 (O_1548,N_48302,N_48000);
nand UO_1549 (O_1549,N_48229,N_48177);
xnor UO_1550 (O_1550,N_48354,N_48470);
or UO_1551 (O_1551,N_48378,N_49418);
nor UO_1552 (O_1552,N_49905,N_49940);
xor UO_1553 (O_1553,N_47937,N_48471);
or UO_1554 (O_1554,N_48652,N_49779);
nand UO_1555 (O_1555,N_49300,N_49813);
xor UO_1556 (O_1556,N_49279,N_47554);
and UO_1557 (O_1557,N_48161,N_49114);
or UO_1558 (O_1558,N_48176,N_48239);
nand UO_1559 (O_1559,N_47538,N_48607);
nor UO_1560 (O_1560,N_48607,N_49253);
or UO_1561 (O_1561,N_49476,N_49971);
and UO_1562 (O_1562,N_48749,N_47714);
nor UO_1563 (O_1563,N_48119,N_47893);
and UO_1564 (O_1564,N_48913,N_48073);
nor UO_1565 (O_1565,N_48775,N_49247);
nor UO_1566 (O_1566,N_49279,N_48207);
xnor UO_1567 (O_1567,N_49391,N_49868);
nand UO_1568 (O_1568,N_49217,N_47663);
or UO_1569 (O_1569,N_48507,N_48008);
nor UO_1570 (O_1570,N_49529,N_48533);
xnor UO_1571 (O_1571,N_49245,N_49344);
and UO_1572 (O_1572,N_48843,N_47897);
nor UO_1573 (O_1573,N_48676,N_49973);
nand UO_1574 (O_1574,N_49652,N_49072);
nor UO_1575 (O_1575,N_49510,N_49570);
nand UO_1576 (O_1576,N_48580,N_47766);
nor UO_1577 (O_1577,N_47531,N_48503);
xor UO_1578 (O_1578,N_49150,N_49684);
nor UO_1579 (O_1579,N_49351,N_49296);
nand UO_1580 (O_1580,N_47950,N_47846);
or UO_1581 (O_1581,N_49989,N_48114);
xnor UO_1582 (O_1582,N_48999,N_47698);
and UO_1583 (O_1583,N_48601,N_48792);
nor UO_1584 (O_1584,N_49171,N_49302);
and UO_1585 (O_1585,N_49728,N_48591);
or UO_1586 (O_1586,N_49244,N_49159);
xor UO_1587 (O_1587,N_49097,N_47975);
nand UO_1588 (O_1588,N_47556,N_48207);
and UO_1589 (O_1589,N_49142,N_47966);
xor UO_1590 (O_1590,N_48922,N_48971);
and UO_1591 (O_1591,N_47932,N_47750);
and UO_1592 (O_1592,N_48428,N_49038);
and UO_1593 (O_1593,N_49378,N_48992);
or UO_1594 (O_1594,N_47817,N_48489);
and UO_1595 (O_1595,N_49321,N_49775);
and UO_1596 (O_1596,N_47820,N_49005);
nand UO_1597 (O_1597,N_48223,N_48809);
xnor UO_1598 (O_1598,N_49916,N_47696);
nor UO_1599 (O_1599,N_49650,N_48971);
nor UO_1600 (O_1600,N_48732,N_47798);
nor UO_1601 (O_1601,N_48125,N_49829);
nor UO_1602 (O_1602,N_49999,N_49066);
xor UO_1603 (O_1603,N_48343,N_48374);
or UO_1604 (O_1604,N_48314,N_49081);
nor UO_1605 (O_1605,N_49628,N_48354);
or UO_1606 (O_1606,N_49779,N_48972);
nor UO_1607 (O_1607,N_48012,N_49348);
or UO_1608 (O_1608,N_49119,N_48258);
or UO_1609 (O_1609,N_48403,N_49905);
xor UO_1610 (O_1610,N_48896,N_49439);
and UO_1611 (O_1611,N_47800,N_47541);
nor UO_1612 (O_1612,N_47509,N_48720);
and UO_1613 (O_1613,N_47617,N_48003);
and UO_1614 (O_1614,N_49031,N_49969);
xor UO_1615 (O_1615,N_47530,N_47523);
xor UO_1616 (O_1616,N_48534,N_48969);
or UO_1617 (O_1617,N_48680,N_47597);
xnor UO_1618 (O_1618,N_48687,N_48291);
or UO_1619 (O_1619,N_49193,N_49217);
xor UO_1620 (O_1620,N_48005,N_48192);
nor UO_1621 (O_1621,N_49399,N_48464);
and UO_1622 (O_1622,N_49607,N_49212);
and UO_1623 (O_1623,N_48806,N_48540);
nand UO_1624 (O_1624,N_48942,N_48880);
nand UO_1625 (O_1625,N_48258,N_48584);
nor UO_1626 (O_1626,N_48179,N_47776);
xnor UO_1627 (O_1627,N_48976,N_48154);
nand UO_1628 (O_1628,N_49669,N_49557);
nor UO_1629 (O_1629,N_49219,N_49411);
or UO_1630 (O_1630,N_49507,N_49321);
xnor UO_1631 (O_1631,N_48278,N_49517);
and UO_1632 (O_1632,N_49043,N_49475);
nand UO_1633 (O_1633,N_48515,N_48222);
nand UO_1634 (O_1634,N_48670,N_49952);
nand UO_1635 (O_1635,N_49708,N_48725);
nand UO_1636 (O_1636,N_47723,N_49294);
nand UO_1637 (O_1637,N_49835,N_47936);
nand UO_1638 (O_1638,N_49569,N_49658);
nand UO_1639 (O_1639,N_49141,N_48964);
xor UO_1640 (O_1640,N_47616,N_49691);
and UO_1641 (O_1641,N_48122,N_49894);
nand UO_1642 (O_1642,N_47657,N_48574);
nand UO_1643 (O_1643,N_48279,N_49942);
nand UO_1644 (O_1644,N_49845,N_48572);
and UO_1645 (O_1645,N_49789,N_48177);
xor UO_1646 (O_1646,N_47677,N_49288);
nor UO_1647 (O_1647,N_47511,N_49498);
nor UO_1648 (O_1648,N_48127,N_49927);
and UO_1649 (O_1649,N_47659,N_49276);
or UO_1650 (O_1650,N_49171,N_48419);
nor UO_1651 (O_1651,N_49984,N_47797);
nor UO_1652 (O_1652,N_47850,N_47781);
nand UO_1653 (O_1653,N_48238,N_47561);
nor UO_1654 (O_1654,N_48357,N_49548);
nor UO_1655 (O_1655,N_48857,N_49854);
or UO_1656 (O_1656,N_49847,N_48629);
nor UO_1657 (O_1657,N_49513,N_48481);
or UO_1658 (O_1658,N_49758,N_47944);
and UO_1659 (O_1659,N_47949,N_49177);
xor UO_1660 (O_1660,N_48201,N_48987);
or UO_1661 (O_1661,N_47993,N_48088);
or UO_1662 (O_1662,N_48146,N_48914);
and UO_1663 (O_1663,N_49992,N_48086);
nor UO_1664 (O_1664,N_48772,N_48567);
nand UO_1665 (O_1665,N_49820,N_48965);
xnor UO_1666 (O_1666,N_47684,N_49725);
and UO_1667 (O_1667,N_48623,N_47982);
and UO_1668 (O_1668,N_49413,N_47768);
or UO_1669 (O_1669,N_48462,N_48293);
nor UO_1670 (O_1670,N_47798,N_49804);
nand UO_1671 (O_1671,N_49324,N_48188);
or UO_1672 (O_1672,N_47687,N_47880);
nor UO_1673 (O_1673,N_49825,N_49417);
and UO_1674 (O_1674,N_49169,N_49248);
nor UO_1675 (O_1675,N_49277,N_48141);
or UO_1676 (O_1676,N_48983,N_49450);
nor UO_1677 (O_1677,N_49125,N_47717);
or UO_1678 (O_1678,N_48710,N_48980);
and UO_1679 (O_1679,N_48764,N_49480);
nor UO_1680 (O_1680,N_49204,N_48003);
and UO_1681 (O_1681,N_47616,N_48932);
or UO_1682 (O_1682,N_47519,N_49479);
xnor UO_1683 (O_1683,N_47975,N_47904);
and UO_1684 (O_1684,N_49719,N_49498);
xnor UO_1685 (O_1685,N_48984,N_49845);
or UO_1686 (O_1686,N_48932,N_49167);
nand UO_1687 (O_1687,N_47971,N_49943);
and UO_1688 (O_1688,N_48018,N_49234);
nand UO_1689 (O_1689,N_48878,N_49283);
or UO_1690 (O_1690,N_48157,N_49381);
nand UO_1691 (O_1691,N_49977,N_48502);
or UO_1692 (O_1692,N_48982,N_49891);
xor UO_1693 (O_1693,N_48708,N_47939);
nor UO_1694 (O_1694,N_47657,N_48972);
nand UO_1695 (O_1695,N_49018,N_48546);
nor UO_1696 (O_1696,N_49129,N_48387);
or UO_1697 (O_1697,N_48159,N_49976);
xnor UO_1698 (O_1698,N_49839,N_48806);
xor UO_1699 (O_1699,N_49039,N_49989);
or UO_1700 (O_1700,N_48099,N_49259);
nand UO_1701 (O_1701,N_49310,N_48156);
nor UO_1702 (O_1702,N_49689,N_48856);
or UO_1703 (O_1703,N_48045,N_47786);
xor UO_1704 (O_1704,N_49287,N_48069);
nor UO_1705 (O_1705,N_48862,N_47941);
nor UO_1706 (O_1706,N_49263,N_48756);
nand UO_1707 (O_1707,N_48644,N_48808);
and UO_1708 (O_1708,N_49911,N_48721);
or UO_1709 (O_1709,N_47540,N_47838);
xnor UO_1710 (O_1710,N_49553,N_48401);
xor UO_1711 (O_1711,N_48907,N_47531);
or UO_1712 (O_1712,N_48726,N_47791);
and UO_1713 (O_1713,N_49568,N_47667);
nor UO_1714 (O_1714,N_49369,N_48337);
and UO_1715 (O_1715,N_49648,N_49478);
xor UO_1716 (O_1716,N_48723,N_49571);
or UO_1717 (O_1717,N_48769,N_49942);
and UO_1718 (O_1718,N_47803,N_49037);
or UO_1719 (O_1719,N_47821,N_49676);
or UO_1720 (O_1720,N_47886,N_49547);
nor UO_1721 (O_1721,N_48732,N_47513);
nor UO_1722 (O_1722,N_48170,N_48076);
and UO_1723 (O_1723,N_47570,N_48014);
nand UO_1724 (O_1724,N_49178,N_49091);
and UO_1725 (O_1725,N_49312,N_48733);
xnor UO_1726 (O_1726,N_48336,N_49225);
or UO_1727 (O_1727,N_48156,N_48587);
or UO_1728 (O_1728,N_48622,N_48794);
nor UO_1729 (O_1729,N_48570,N_48739);
and UO_1730 (O_1730,N_49761,N_48560);
xor UO_1731 (O_1731,N_48354,N_47809);
nor UO_1732 (O_1732,N_49086,N_49027);
xnor UO_1733 (O_1733,N_48021,N_49826);
nor UO_1734 (O_1734,N_49262,N_48200);
xnor UO_1735 (O_1735,N_49874,N_48148);
nor UO_1736 (O_1736,N_48735,N_49507);
or UO_1737 (O_1737,N_49756,N_47973);
nor UO_1738 (O_1738,N_49471,N_47920);
nor UO_1739 (O_1739,N_47508,N_49150);
or UO_1740 (O_1740,N_48702,N_48748);
xnor UO_1741 (O_1741,N_48841,N_48469);
or UO_1742 (O_1742,N_49934,N_49219);
and UO_1743 (O_1743,N_49897,N_47513);
nor UO_1744 (O_1744,N_48448,N_47836);
or UO_1745 (O_1745,N_48363,N_48760);
nor UO_1746 (O_1746,N_49375,N_49813);
and UO_1747 (O_1747,N_49111,N_49865);
nor UO_1748 (O_1748,N_49927,N_49487);
and UO_1749 (O_1749,N_48941,N_48326);
nor UO_1750 (O_1750,N_49924,N_48100);
and UO_1751 (O_1751,N_49241,N_49629);
and UO_1752 (O_1752,N_47743,N_47522);
nand UO_1753 (O_1753,N_48988,N_49308);
nor UO_1754 (O_1754,N_48491,N_47914);
nor UO_1755 (O_1755,N_48447,N_49469);
or UO_1756 (O_1756,N_49269,N_48156);
nor UO_1757 (O_1757,N_49742,N_47589);
nor UO_1758 (O_1758,N_47901,N_48518);
nand UO_1759 (O_1759,N_48966,N_48838);
and UO_1760 (O_1760,N_48496,N_48936);
xor UO_1761 (O_1761,N_47833,N_49054);
xor UO_1762 (O_1762,N_48943,N_48277);
xnor UO_1763 (O_1763,N_49091,N_48660);
nand UO_1764 (O_1764,N_49707,N_48409);
and UO_1765 (O_1765,N_49996,N_49609);
nor UO_1766 (O_1766,N_49915,N_48039);
nor UO_1767 (O_1767,N_47997,N_48203);
nor UO_1768 (O_1768,N_49347,N_49533);
xnor UO_1769 (O_1769,N_47734,N_49044);
nor UO_1770 (O_1770,N_47558,N_47529);
xor UO_1771 (O_1771,N_49199,N_48149);
or UO_1772 (O_1772,N_48554,N_48784);
nor UO_1773 (O_1773,N_48290,N_49197);
and UO_1774 (O_1774,N_48961,N_49157);
and UO_1775 (O_1775,N_49615,N_49483);
xor UO_1776 (O_1776,N_48864,N_49442);
or UO_1777 (O_1777,N_48375,N_49753);
nand UO_1778 (O_1778,N_49519,N_47767);
and UO_1779 (O_1779,N_49680,N_49381);
nor UO_1780 (O_1780,N_48299,N_49107);
xnor UO_1781 (O_1781,N_48943,N_48620);
or UO_1782 (O_1782,N_49363,N_47763);
nor UO_1783 (O_1783,N_48059,N_48483);
nand UO_1784 (O_1784,N_47615,N_48843);
xor UO_1785 (O_1785,N_49188,N_47957);
or UO_1786 (O_1786,N_49885,N_47754);
or UO_1787 (O_1787,N_47669,N_47527);
xnor UO_1788 (O_1788,N_47783,N_49565);
xor UO_1789 (O_1789,N_48048,N_49139);
xor UO_1790 (O_1790,N_47798,N_49505);
nand UO_1791 (O_1791,N_47639,N_48300);
nand UO_1792 (O_1792,N_49514,N_48731);
or UO_1793 (O_1793,N_47614,N_48388);
xnor UO_1794 (O_1794,N_48385,N_48325);
and UO_1795 (O_1795,N_48107,N_47934);
or UO_1796 (O_1796,N_49455,N_48493);
and UO_1797 (O_1797,N_49187,N_48227);
and UO_1798 (O_1798,N_49998,N_49828);
nand UO_1799 (O_1799,N_49504,N_49151);
or UO_1800 (O_1800,N_49910,N_49159);
nand UO_1801 (O_1801,N_48102,N_49170);
xnor UO_1802 (O_1802,N_48835,N_48950);
nor UO_1803 (O_1803,N_48136,N_48699);
xnor UO_1804 (O_1804,N_48158,N_49339);
or UO_1805 (O_1805,N_47679,N_49675);
or UO_1806 (O_1806,N_48125,N_48284);
and UO_1807 (O_1807,N_48323,N_49781);
nor UO_1808 (O_1808,N_48612,N_47586);
nand UO_1809 (O_1809,N_48975,N_47628);
or UO_1810 (O_1810,N_49424,N_49472);
and UO_1811 (O_1811,N_48534,N_49284);
or UO_1812 (O_1812,N_47842,N_48557);
nor UO_1813 (O_1813,N_48934,N_47686);
nand UO_1814 (O_1814,N_49645,N_48831);
or UO_1815 (O_1815,N_48803,N_49440);
nor UO_1816 (O_1816,N_47682,N_49949);
xnor UO_1817 (O_1817,N_48884,N_47918);
and UO_1818 (O_1818,N_47736,N_49415);
xnor UO_1819 (O_1819,N_48572,N_47827);
or UO_1820 (O_1820,N_48103,N_49216);
or UO_1821 (O_1821,N_48650,N_48068);
nand UO_1822 (O_1822,N_49849,N_49759);
xnor UO_1823 (O_1823,N_49409,N_49282);
and UO_1824 (O_1824,N_47568,N_49502);
xor UO_1825 (O_1825,N_49412,N_49878);
xor UO_1826 (O_1826,N_49314,N_49450);
and UO_1827 (O_1827,N_48332,N_49348);
or UO_1828 (O_1828,N_47977,N_48533);
nand UO_1829 (O_1829,N_48272,N_49993);
xor UO_1830 (O_1830,N_49281,N_49585);
nor UO_1831 (O_1831,N_49473,N_47570);
and UO_1832 (O_1832,N_48356,N_49777);
and UO_1833 (O_1833,N_49464,N_49800);
xor UO_1834 (O_1834,N_48738,N_47900);
nand UO_1835 (O_1835,N_49497,N_49591);
and UO_1836 (O_1836,N_48033,N_48264);
nor UO_1837 (O_1837,N_48762,N_47846);
or UO_1838 (O_1838,N_47607,N_49973);
or UO_1839 (O_1839,N_47829,N_49331);
nand UO_1840 (O_1840,N_49258,N_47562);
nor UO_1841 (O_1841,N_49934,N_49163);
and UO_1842 (O_1842,N_47973,N_48538);
nor UO_1843 (O_1843,N_48440,N_48629);
nand UO_1844 (O_1844,N_48965,N_47789);
and UO_1845 (O_1845,N_47699,N_47528);
or UO_1846 (O_1846,N_49672,N_47930);
xnor UO_1847 (O_1847,N_49992,N_47698);
nand UO_1848 (O_1848,N_48759,N_49728);
or UO_1849 (O_1849,N_48277,N_49212);
nor UO_1850 (O_1850,N_48394,N_48230);
xor UO_1851 (O_1851,N_48394,N_48243);
and UO_1852 (O_1852,N_49556,N_47679);
nor UO_1853 (O_1853,N_47532,N_47681);
nand UO_1854 (O_1854,N_48111,N_48734);
xor UO_1855 (O_1855,N_47991,N_47665);
xnor UO_1856 (O_1856,N_48364,N_48844);
nand UO_1857 (O_1857,N_48842,N_48262);
nand UO_1858 (O_1858,N_49546,N_49831);
or UO_1859 (O_1859,N_48211,N_47882);
and UO_1860 (O_1860,N_49678,N_48385);
nor UO_1861 (O_1861,N_49199,N_47568);
nand UO_1862 (O_1862,N_49055,N_49367);
xnor UO_1863 (O_1863,N_47759,N_49727);
nand UO_1864 (O_1864,N_49306,N_47539);
nand UO_1865 (O_1865,N_47772,N_49639);
and UO_1866 (O_1866,N_49531,N_49173);
nor UO_1867 (O_1867,N_49674,N_49204);
or UO_1868 (O_1868,N_47518,N_48501);
xor UO_1869 (O_1869,N_48561,N_49834);
and UO_1870 (O_1870,N_48022,N_48261);
xnor UO_1871 (O_1871,N_48967,N_47655);
xnor UO_1872 (O_1872,N_49858,N_47532);
nand UO_1873 (O_1873,N_49272,N_47760);
and UO_1874 (O_1874,N_47774,N_49353);
and UO_1875 (O_1875,N_48812,N_47596);
xnor UO_1876 (O_1876,N_49580,N_47542);
xor UO_1877 (O_1877,N_49233,N_48963);
xnor UO_1878 (O_1878,N_47565,N_49275);
xor UO_1879 (O_1879,N_49085,N_47714);
nor UO_1880 (O_1880,N_49505,N_49531);
xor UO_1881 (O_1881,N_49893,N_49522);
and UO_1882 (O_1882,N_49814,N_47874);
and UO_1883 (O_1883,N_49621,N_49653);
and UO_1884 (O_1884,N_47818,N_49138);
xnor UO_1885 (O_1885,N_48123,N_49084);
and UO_1886 (O_1886,N_48195,N_49028);
nand UO_1887 (O_1887,N_47665,N_49605);
and UO_1888 (O_1888,N_49294,N_47877);
xor UO_1889 (O_1889,N_48916,N_48148);
and UO_1890 (O_1890,N_47819,N_49096);
nor UO_1891 (O_1891,N_49440,N_47894);
and UO_1892 (O_1892,N_49099,N_48558);
and UO_1893 (O_1893,N_48548,N_49644);
and UO_1894 (O_1894,N_48099,N_49661);
and UO_1895 (O_1895,N_47629,N_49945);
or UO_1896 (O_1896,N_48059,N_47672);
nand UO_1897 (O_1897,N_48621,N_48705);
and UO_1898 (O_1898,N_48246,N_48733);
nand UO_1899 (O_1899,N_47650,N_47833);
nor UO_1900 (O_1900,N_47568,N_48551);
nand UO_1901 (O_1901,N_48609,N_49804);
and UO_1902 (O_1902,N_48254,N_49313);
or UO_1903 (O_1903,N_48119,N_48285);
or UO_1904 (O_1904,N_47704,N_47915);
nand UO_1905 (O_1905,N_49075,N_48136);
nand UO_1906 (O_1906,N_49103,N_48572);
and UO_1907 (O_1907,N_48139,N_48218);
or UO_1908 (O_1908,N_47741,N_49848);
nand UO_1909 (O_1909,N_48964,N_49041);
or UO_1910 (O_1910,N_48417,N_49675);
nand UO_1911 (O_1911,N_49275,N_48764);
nand UO_1912 (O_1912,N_49617,N_48023);
xnor UO_1913 (O_1913,N_48043,N_49355);
nor UO_1914 (O_1914,N_49104,N_48205);
nand UO_1915 (O_1915,N_49025,N_47927);
xor UO_1916 (O_1916,N_49475,N_48196);
nand UO_1917 (O_1917,N_49145,N_47715);
or UO_1918 (O_1918,N_49177,N_47887);
and UO_1919 (O_1919,N_47876,N_48942);
xnor UO_1920 (O_1920,N_49958,N_49227);
nor UO_1921 (O_1921,N_47935,N_49097);
nor UO_1922 (O_1922,N_49768,N_49657);
and UO_1923 (O_1923,N_48478,N_48525);
nor UO_1924 (O_1924,N_49860,N_48809);
nor UO_1925 (O_1925,N_48993,N_49442);
nand UO_1926 (O_1926,N_48676,N_48961);
or UO_1927 (O_1927,N_48268,N_48183);
and UO_1928 (O_1928,N_49021,N_48365);
nand UO_1929 (O_1929,N_49725,N_47636);
nand UO_1930 (O_1930,N_48203,N_48282);
xor UO_1931 (O_1931,N_49881,N_48840);
nand UO_1932 (O_1932,N_48581,N_49935);
or UO_1933 (O_1933,N_49106,N_47734);
nor UO_1934 (O_1934,N_48112,N_49534);
xnor UO_1935 (O_1935,N_49623,N_48292);
nor UO_1936 (O_1936,N_47558,N_49584);
and UO_1937 (O_1937,N_47997,N_48803);
or UO_1938 (O_1938,N_48941,N_47839);
nand UO_1939 (O_1939,N_49158,N_48901);
nand UO_1940 (O_1940,N_49317,N_48617);
nand UO_1941 (O_1941,N_49098,N_48457);
and UO_1942 (O_1942,N_47858,N_49961);
and UO_1943 (O_1943,N_48285,N_47820);
and UO_1944 (O_1944,N_49060,N_48452);
xor UO_1945 (O_1945,N_49331,N_48259);
and UO_1946 (O_1946,N_48046,N_48314);
nand UO_1947 (O_1947,N_49394,N_48435);
xnor UO_1948 (O_1948,N_48629,N_49315);
nand UO_1949 (O_1949,N_47715,N_48403);
xor UO_1950 (O_1950,N_47667,N_49454);
nand UO_1951 (O_1951,N_49116,N_48032);
and UO_1952 (O_1952,N_49128,N_49263);
and UO_1953 (O_1953,N_47637,N_47751);
or UO_1954 (O_1954,N_47502,N_49253);
nor UO_1955 (O_1955,N_49848,N_48315);
xnor UO_1956 (O_1956,N_49148,N_48120);
and UO_1957 (O_1957,N_49215,N_48627);
xnor UO_1958 (O_1958,N_49381,N_49251);
or UO_1959 (O_1959,N_49941,N_48763);
nor UO_1960 (O_1960,N_48890,N_49221);
xnor UO_1961 (O_1961,N_49637,N_48783);
and UO_1962 (O_1962,N_47964,N_48459);
or UO_1963 (O_1963,N_48863,N_49130);
xnor UO_1964 (O_1964,N_47637,N_48851);
or UO_1965 (O_1965,N_47776,N_49779);
nand UO_1966 (O_1966,N_49402,N_48768);
and UO_1967 (O_1967,N_48263,N_48413);
xnor UO_1968 (O_1968,N_47674,N_48512);
and UO_1969 (O_1969,N_48774,N_47671);
or UO_1970 (O_1970,N_49930,N_48479);
nand UO_1971 (O_1971,N_48305,N_48569);
xnor UO_1972 (O_1972,N_48477,N_47806);
or UO_1973 (O_1973,N_49217,N_48028);
nand UO_1974 (O_1974,N_49663,N_48139);
and UO_1975 (O_1975,N_48925,N_48992);
or UO_1976 (O_1976,N_47854,N_49147);
or UO_1977 (O_1977,N_49908,N_48056);
and UO_1978 (O_1978,N_47774,N_47991);
nor UO_1979 (O_1979,N_48705,N_49791);
and UO_1980 (O_1980,N_49861,N_49155);
or UO_1981 (O_1981,N_49923,N_49527);
xor UO_1982 (O_1982,N_47913,N_49128);
nand UO_1983 (O_1983,N_49695,N_47898);
and UO_1984 (O_1984,N_48508,N_48221);
or UO_1985 (O_1985,N_48741,N_49725);
nor UO_1986 (O_1986,N_48113,N_47937);
and UO_1987 (O_1987,N_48616,N_49186);
xor UO_1988 (O_1988,N_48017,N_48592);
xnor UO_1989 (O_1989,N_47779,N_49999);
xnor UO_1990 (O_1990,N_48380,N_49875);
nand UO_1991 (O_1991,N_48444,N_48025);
xor UO_1992 (O_1992,N_48994,N_49806);
nor UO_1993 (O_1993,N_48083,N_47623);
and UO_1994 (O_1994,N_48580,N_47528);
or UO_1995 (O_1995,N_49552,N_48423);
xnor UO_1996 (O_1996,N_49978,N_48669);
nand UO_1997 (O_1997,N_49505,N_48229);
xnor UO_1998 (O_1998,N_49118,N_48191);
or UO_1999 (O_1999,N_47915,N_48447);
xnor UO_2000 (O_2000,N_47818,N_49938);
nor UO_2001 (O_2001,N_47880,N_49313);
or UO_2002 (O_2002,N_48787,N_48726);
and UO_2003 (O_2003,N_48923,N_49295);
nor UO_2004 (O_2004,N_49219,N_48986);
and UO_2005 (O_2005,N_47599,N_48109);
nand UO_2006 (O_2006,N_49514,N_47830);
nand UO_2007 (O_2007,N_48554,N_48677);
xnor UO_2008 (O_2008,N_48665,N_47956);
nor UO_2009 (O_2009,N_48958,N_48487);
and UO_2010 (O_2010,N_48331,N_48541);
or UO_2011 (O_2011,N_48482,N_48426);
nand UO_2012 (O_2012,N_48666,N_49907);
nand UO_2013 (O_2013,N_49152,N_49491);
or UO_2014 (O_2014,N_48431,N_49225);
or UO_2015 (O_2015,N_47885,N_49529);
nand UO_2016 (O_2016,N_49466,N_48037);
xnor UO_2017 (O_2017,N_47913,N_48033);
xor UO_2018 (O_2018,N_49386,N_48187);
or UO_2019 (O_2019,N_49144,N_49275);
and UO_2020 (O_2020,N_49680,N_48667);
xor UO_2021 (O_2021,N_49421,N_48575);
or UO_2022 (O_2022,N_49830,N_47806);
or UO_2023 (O_2023,N_49184,N_47589);
nor UO_2024 (O_2024,N_47750,N_48027);
nor UO_2025 (O_2025,N_48182,N_48318);
and UO_2026 (O_2026,N_47780,N_48449);
and UO_2027 (O_2027,N_48200,N_49632);
xor UO_2028 (O_2028,N_49230,N_47986);
nor UO_2029 (O_2029,N_47940,N_48145);
nor UO_2030 (O_2030,N_47833,N_48776);
or UO_2031 (O_2031,N_48711,N_49640);
or UO_2032 (O_2032,N_47522,N_49134);
or UO_2033 (O_2033,N_48419,N_47912);
or UO_2034 (O_2034,N_48165,N_48024);
and UO_2035 (O_2035,N_47861,N_48799);
nor UO_2036 (O_2036,N_48487,N_49761);
nand UO_2037 (O_2037,N_47987,N_48095);
or UO_2038 (O_2038,N_47634,N_49941);
nor UO_2039 (O_2039,N_48987,N_48892);
or UO_2040 (O_2040,N_48262,N_48220);
xor UO_2041 (O_2041,N_48752,N_48182);
or UO_2042 (O_2042,N_47611,N_48362);
and UO_2043 (O_2043,N_49915,N_47551);
nand UO_2044 (O_2044,N_47764,N_48500);
xor UO_2045 (O_2045,N_48758,N_48274);
or UO_2046 (O_2046,N_47612,N_48471);
or UO_2047 (O_2047,N_47546,N_49292);
and UO_2048 (O_2048,N_49157,N_47723);
and UO_2049 (O_2049,N_49785,N_47800);
nand UO_2050 (O_2050,N_49487,N_48814);
or UO_2051 (O_2051,N_48267,N_48421);
xnor UO_2052 (O_2052,N_49439,N_47805);
or UO_2053 (O_2053,N_49384,N_48627);
nor UO_2054 (O_2054,N_49241,N_49595);
nor UO_2055 (O_2055,N_49280,N_47860);
nand UO_2056 (O_2056,N_48395,N_49144);
or UO_2057 (O_2057,N_48998,N_48934);
or UO_2058 (O_2058,N_48580,N_49928);
xnor UO_2059 (O_2059,N_49732,N_47627);
or UO_2060 (O_2060,N_49510,N_49870);
and UO_2061 (O_2061,N_49487,N_48990);
nor UO_2062 (O_2062,N_49454,N_49371);
nor UO_2063 (O_2063,N_48918,N_48728);
nand UO_2064 (O_2064,N_49648,N_48403);
nand UO_2065 (O_2065,N_49617,N_47806);
nor UO_2066 (O_2066,N_48235,N_49874);
or UO_2067 (O_2067,N_49239,N_48377);
and UO_2068 (O_2068,N_49071,N_48841);
or UO_2069 (O_2069,N_48877,N_48408);
xnor UO_2070 (O_2070,N_48770,N_48651);
xnor UO_2071 (O_2071,N_48824,N_47818);
xor UO_2072 (O_2072,N_49418,N_49332);
nand UO_2073 (O_2073,N_48601,N_48423);
and UO_2074 (O_2074,N_49144,N_48280);
nor UO_2075 (O_2075,N_49861,N_47647);
nor UO_2076 (O_2076,N_48736,N_48758);
or UO_2077 (O_2077,N_47653,N_48931);
and UO_2078 (O_2078,N_47885,N_47930);
xor UO_2079 (O_2079,N_49817,N_47892);
xnor UO_2080 (O_2080,N_48659,N_49234);
xnor UO_2081 (O_2081,N_48574,N_47879);
xnor UO_2082 (O_2082,N_49029,N_48139);
nor UO_2083 (O_2083,N_49440,N_47578);
nor UO_2084 (O_2084,N_47671,N_47807);
xor UO_2085 (O_2085,N_48115,N_49906);
or UO_2086 (O_2086,N_48660,N_49880);
or UO_2087 (O_2087,N_48777,N_47738);
nand UO_2088 (O_2088,N_48918,N_49794);
and UO_2089 (O_2089,N_48222,N_49905);
xnor UO_2090 (O_2090,N_47856,N_49380);
xnor UO_2091 (O_2091,N_48319,N_49655);
nand UO_2092 (O_2092,N_48153,N_47507);
and UO_2093 (O_2093,N_49703,N_49049);
or UO_2094 (O_2094,N_48925,N_48151);
nand UO_2095 (O_2095,N_47969,N_47844);
xor UO_2096 (O_2096,N_49897,N_47550);
and UO_2097 (O_2097,N_48159,N_49119);
xor UO_2098 (O_2098,N_49582,N_48513);
nand UO_2099 (O_2099,N_49929,N_49117);
and UO_2100 (O_2100,N_47912,N_49008);
nand UO_2101 (O_2101,N_47639,N_49406);
xnor UO_2102 (O_2102,N_48959,N_48275);
nor UO_2103 (O_2103,N_48243,N_49658);
xnor UO_2104 (O_2104,N_49610,N_47873);
and UO_2105 (O_2105,N_49426,N_48507);
and UO_2106 (O_2106,N_49890,N_48017);
xor UO_2107 (O_2107,N_48194,N_49888);
xnor UO_2108 (O_2108,N_48829,N_48070);
and UO_2109 (O_2109,N_48534,N_48912);
and UO_2110 (O_2110,N_48955,N_47737);
and UO_2111 (O_2111,N_48617,N_48156);
or UO_2112 (O_2112,N_47759,N_48100);
xnor UO_2113 (O_2113,N_48785,N_49049);
or UO_2114 (O_2114,N_49101,N_48521);
nand UO_2115 (O_2115,N_49423,N_49330);
nor UO_2116 (O_2116,N_47678,N_49228);
nand UO_2117 (O_2117,N_49727,N_48556);
nand UO_2118 (O_2118,N_47756,N_48557);
xor UO_2119 (O_2119,N_48529,N_47672);
nor UO_2120 (O_2120,N_48053,N_49355);
nor UO_2121 (O_2121,N_49457,N_48602);
xor UO_2122 (O_2122,N_47564,N_49095);
nor UO_2123 (O_2123,N_48780,N_48152);
xnor UO_2124 (O_2124,N_48209,N_48951);
nand UO_2125 (O_2125,N_49630,N_49557);
or UO_2126 (O_2126,N_49766,N_47659);
and UO_2127 (O_2127,N_48927,N_47822);
nand UO_2128 (O_2128,N_49282,N_49751);
xnor UO_2129 (O_2129,N_49380,N_49384);
xnor UO_2130 (O_2130,N_49650,N_49169);
xor UO_2131 (O_2131,N_49183,N_47669);
xnor UO_2132 (O_2132,N_48416,N_49702);
or UO_2133 (O_2133,N_48353,N_48523);
xor UO_2134 (O_2134,N_47784,N_47888);
and UO_2135 (O_2135,N_49243,N_48898);
or UO_2136 (O_2136,N_48252,N_48234);
xnor UO_2137 (O_2137,N_49513,N_49227);
and UO_2138 (O_2138,N_47737,N_49272);
nand UO_2139 (O_2139,N_49867,N_49027);
and UO_2140 (O_2140,N_48640,N_49015);
nand UO_2141 (O_2141,N_49264,N_48153);
and UO_2142 (O_2142,N_48366,N_49957);
nand UO_2143 (O_2143,N_48376,N_49861);
nor UO_2144 (O_2144,N_47958,N_47773);
nand UO_2145 (O_2145,N_47881,N_48148);
nor UO_2146 (O_2146,N_49164,N_48002);
and UO_2147 (O_2147,N_49724,N_49339);
or UO_2148 (O_2148,N_48145,N_48510);
xor UO_2149 (O_2149,N_47612,N_49720);
and UO_2150 (O_2150,N_47700,N_48104);
nand UO_2151 (O_2151,N_48210,N_47946);
or UO_2152 (O_2152,N_47755,N_47610);
and UO_2153 (O_2153,N_48155,N_48654);
and UO_2154 (O_2154,N_47740,N_47837);
nor UO_2155 (O_2155,N_47821,N_47681);
nand UO_2156 (O_2156,N_49434,N_48026);
and UO_2157 (O_2157,N_48982,N_48918);
nor UO_2158 (O_2158,N_48477,N_48145);
or UO_2159 (O_2159,N_48500,N_49562);
xor UO_2160 (O_2160,N_48706,N_49143);
nand UO_2161 (O_2161,N_49615,N_48442);
xor UO_2162 (O_2162,N_49960,N_47510);
nand UO_2163 (O_2163,N_48583,N_48345);
or UO_2164 (O_2164,N_47875,N_48281);
nand UO_2165 (O_2165,N_48939,N_48925);
nand UO_2166 (O_2166,N_48070,N_48184);
xnor UO_2167 (O_2167,N_49912,N_48486);
xor UO_2168 (O_2168,N_49643,N_49383);
nand UO_2169 (O_2169,N_47562,N_48763);
and UO_2170 (O_2170,N_49947,N_48135);
or UO_2171 (O_2171,N_49682,N_49928);
and UO_2172 (O_2172,N_47708,N_49621);
or UO_2173 (O_2173,N_47844,N_47733);
xor UO_2174 (O_2174,N_47907,N_48109);
nor UO_2175 (O_2175,N_48996,N_49914);
and UO_2176 (O_2176,N_49122,N_48828);
and UO_2177 (O_2177,N_47559,N_47787);
or UO_2178 (O_2178,N_48814,N_49775);
or UO_2179 (O_2179,N_48987,N_47693);
xnor UO_2180 (O_2180,N_48458,N_49724);
and UO_2181 (O_2181,N_49998,N_48533);
nor UO_2182 (O_2182,N_48423,N_49953);
and UO_2183 (O_2183,N_49507,N_48296);
xor UO_2184 (O_2184,N_48514,N_47780);
nand UO_2185 (O_2185,N_48823,N_48940);
nor UO_2186 (O_2186,N_49149,N_49637);
xnor UO_2187 (O_2187,N_48147,N_49183);
and UO_2188 (O_2188,N_47558,N_48741);
nand UO_2189 (O_2189,N_48552,N_48427);
nand UO_2190 (O_2190,N_48805,N_48004);
nand UO_2191 (O_2191,N_48733,N_47629);
nand UO_2192 (O_2192,N_48456,N_49522);
nand UO_2193 (O_2193,N_48024,N_48518);
or UO_2194 (O_2194,N_47734,N_47556);
nand UO_2195 (O_2195,N_48083,N_47617);
xor UO_2196 (O_2196,N_48482,N_49229);
xor UO_2197 (O_2197,N_49773,N_47890);
nor UO_2198 (O_2198,N_47590,N_48488);
nand UO_2199 (O_2199,N_49560,N_48225);
and UO_2200 (O_2200,N_47907,N_49298);
nor UO_2201 (O_2201,N_49696,N_48761);
nor UO_2202 (O_2202,N_48887,N_48900);
xor UO_2203 (O_2203,N_48212,N_49806);
nor UO_2204 (O_2204,N_47905,N_48056);
and UO_2205 (O_2205,N_49757,N_47837);
or UO_2206 (O_2206,N_49453,N_47814);
nand UO_2207 (O_2207,N_47604,N_48397);
or UO_2208 (O_2208,N_47705,N_47932);
nor UO_2209 (O_2209,N_48688,N_47518);
or UO_2210 (O_2210,N_47748,N_48057);
xor UO_2211 (O_2211,N_47741,N_49458);
nand UO_2212 (O_2212,N_49718,N_49868);
nor UO_2213 (O_2213,N_48389,N_48013);
nand UO_2214 (O_2214,N_48342,N_48198);
and UO_2215 (O_2215,N_48812,N_48369);
nor UO_2216 (O_2216,N_49105,N_48468);
nand UO_2217 (O_2217,N_48153,N_48232);
or UO_2218 (O_2218,N_47571,N_49409);
nor UO_2219 (O_2219,N_49082,N_48381);
nand UO_2220 (O_2220,N_47520,N_48632);
nand UO_2221 (O_2221,N_48251,N_47598);
and UO_2222 (O_2222,N_48643,N_49820);
or UO_2223 (O_2223,N_49018,N_47953);
xnor UO_2224 (O_2224,N_49094,N_49514);
or UO_2225 (O_2225,N_48764,N_49762);
nand UO_2226 (O_2226,N_49109,N_48727);
nor UO_2227 (O_2227,N_47628,N_48103);
and UO_2228 (O_2228,N_48536,N_49562);
nor UO_2229 (O_2229,N_49743,N_48161);
nand UO_2230 (O_2230,N_48336,N_48246);
and UO_2231 (O_2231,N_49205,N_49352);
and UO_2232 (O_2232,N_48340,N_49505);
or UO_2233 (O_2233,N_48165,N_49760);
nor UO_2234 (O_2234,N_48642,N_48482);
xor UO_2235 (O_2235,N_49338,N_49396);
nand UO_2236 (O_2236,N_49994,N_48131);
and UO_2237 (O_2237,N_49490,N_47663);
and UO_2238 (O_2238,N_49312,N_49963);
xnor UO_2239 (O_2239,N_49969,N_48342);
and UO_2240 (O_2240,N_47783,N_48172);
xnor UO_2241 (O_2241,N_48109,N_48484);
nand UO_2242 (O_2242,N_49083,N_49081);
or UO_2243 (O_2243,N_48864,N_47923);
or UO_2244 (O_2244,N_48308,N_48049);
or UO_2245 (O_2245,N_48974,N_48191);
or UO_2246 (O_2246,N_49884,N_49232);
or UO_2247 (O_2247,N_47798,N_49563);
nor UO_2248 (O_2248,N_49178,N_49045);
nand UO_2249 (O_2249,N_49456,N_48295);
or UO_2250 (O_2250,N_48115,N_48492);
or UO_2251 (O_2251,N_49807,N_49421);
xor UO_2252 (O_2252,N_47888,N_48499);
nor UO_2253 (O_2253,N_47544,N_49973);
xnor UO_2254 (O_2254,N_47655,N_47598);
nor UO_2255 (O_2255,N_48641,N_48823);
xor UO_2256 (O_2256,N_49086,N_49555);
xor UO_2257 (O_2257,N_48545,N_49913);
and UO_2258 (O_2258,N_49414,N_47696);
xnor UO_2259 (O_2259,N_47695,N_47666);
nand UO_2260 (O_2260,N_49071,N_49669);
xor UO_2261 (O_2261,N_48689,N_49054);
and UO_2262 (O_2262,N_47968,N_49707);
nor UO_2263 (O_2263,N_47520,N_48775);
and UO_2264 (O_2264,N_49753,N_47814);
nor UO_2265 (O_2265,N_47582,N_48307);
nand UO_2266 (O_2266,N_47976,N_48534);
and UO_2267 (O_2267,N_48228,N_47884);
and UO_2268 (O_2268,N_47620,N_49177);
or UO_2269 (O_2269,N_47506,N_48219);
xnor UO_2270 (O_2270,N_49980,N_47967);
nand UO_2271 (O_2271,N_48918,N_48765);
nor UO_2272 (O_2272,N_48698,N_47513);
nor UO_2273 (O_2273,N_49084,N_49767);
nand UO_2274 (O_2274,N_48972,N_47921);
xor UO_2275 (O_2275,N_49742,N_49576);
and UO_2276 (O_2276,N_49032,N_49179);
nand UO_2277 (O_2277,N_49719,N_48953);
and UO_2278 (O_2278,N_49296,N_49219);
nand UO_2279 (O_2279,N_49607,N_49947);
xnor UO_2280 (O_2280,N_48364,N_48193);
nor UO_2281 (O_2281,N_49322,N_47581);
nor UO_2282 (O_2282,N_47606,N_47716);
and UO_2283 (O_2283,N_49285,N_49769);
or UO_2284 (O_2284,N_49280,N_49425);
xor UO_2285 (O_2285,N_48076,N_47882);
and UO_2286 (O_2286,N_49753,N_49946);
and UO_2287 (O_2287,N_49003,N_47711);
xor UO_2288 (O_2288,N_49280,N_49037);
and UO_2289 (O_2289,N_47703,N_49170);
and UO_2290 (O_2290,N_49058,N_48509);
nand UO_2291 (O_2291,N_48296,N_47542);
or UO_2292 (O_2292,N_47736,N_47825);
nand UO_2293 (O_2293,N_49954,N_48881);
nand UO_2294 (O_2294,N_49866,N_48115);
nor UO_2295 (O_2295,N_49457,N_48053);
and UO_2296 (O_2296,N_47684,N_48663);
or UO_2297 (O_2297,N_48313,N_49888);
or UO_2298 (O_2298,N_48253,N_49539);
xnor UO_2299 (O_2299,N_49713,N_48335);
xnor UO_2300 (O_2300,N_49887,N_49541);
nor UO_2301 (O_2301,N_47501,N_48296);
and UO_2302 (O_2302,N_49097,N_48532);
or UO_2303 (O_2303,N_47597,N_48652);
xor UO_2304 (O_2304,N_47648,N_49981);
nand UO_2305 (O_2305,N_49541,N_48992);
or UO_2306 (O_2306,N_49945,N_48182);
nand UO_2307 (O_2307,N_49849,N_49511);
nor UO_2308 (O_2308,N_48290,N_48410);
nand UO_2309 (O_2309,N_48902,N_49204);
nand UO_2310 (O_2310,N_49639,N_47884);
and UO_2311 (O_2311,N_48444,N_48467);
nor UO_2312 (O_2312,N_49588,N_48998);
or UO_2313 (O_2313,N_48324,N_47588);
nor UO_2314 (O_2314,N_47834,N_49513);
and UO_2315 (O_2315,N_48355,N_48927);
or UO_2316 (O_2316,N_49947,N_49986);
xor UO_2317 (O_2317,N_48338,N_48964);
nand UO_2318 (O_2318,N_48599,N_47966);
or UO_2319 (O_2319,N_47754,N_49850);
and UO_2320 (O_2320,N_49200,N_48325);
nor UO_2321 (O_2321,N_48540,N_49838);
or UO_2322 (O_2322,N_49040,N_48547);
and UO_2323 (O_2323,N_48085,N_49527);
xnor UO_2324 (O_2324,N_49298,N_49852);
or UO_2325 (O_2325,N_48340,N_48047);
nor UO_2326 (O_2326,N_49208,N_48321);
nand UO_2327 (O_2327,N_49809,N_47552);
nor UO_2328 (O_2328,N_49605,N_48047);
and UO_2329 (O_2329,N_49541,N_48096);
nor UO_2330 (O_2330,N_48137,N_48149);
or UO_2331 (O_2331,N_47541,N_47944);
nand UO_2332 (O_2332,N_48237,N_47887);
nor UO_2333 (O_2333,N_49272,N_48640);
and UO_2334 (O_2334,N_48631,N_48438);
or UO_2335 (O_2335,N_48739,N_47835);
xor UO_2336 (O_2336,N_49121,N_49406);
and UO_2337 (O_2337,N_48639,N_48031);
nor UO_2338 (O_2338,N_49858,N_47525);
or UO_2339 (O_2339,N_48021,N_47671);
or UO_2340 (O_2340,N_47872,N_48793);
xnor UO_2341 (O_2341,N_49508,N_47568);
xor UO_2342 (O_2342,N_48198,N_48497);
or UO_2343 (O_2343,N_48579,N_49118);
nand UO_2344 (O_2344,N_48316,N_49673);
nand UO_2345 (O_2345,N_48705,N_48168);
and UO_2346 (O_2346,N_48733,N_49995);
nand UO_2347 (O_2347,N_47703,N_48476);
xnor UO_2348 (O_2348,N_49745,N_47687);
xor UO_2349 (O_2349,N_49173,N_48984);
and UO_2350 (O_2350,N_47701,N_47533);
and UO_2351 (O_2351,N_48941,N_47619);
and UO_2352 (O_2352,N_49842,N_49031);
nor UO_2353 (O_2353,N_49762,N_49945);
xor UO_2354 (O_2354,N_48399,N_49744);
xnor UO_2355 (O_2355,N_48935,N_48516);
or UO_2356 (O_2356,N_48026,N_48779);
xor UO_2357 (O_2357,N_48635,N_49916);
or UO_2358 (O_2358,N_47634,N_49607);
or UO_2359 (O_2359,N_48750,N_49616);
and UO_2360 (O_2360,N_49833,N_48054);
nand UO_2361 (O_2361,N_49998,N_49204);
xnor UO_2362 (O_2362,N_48876,N_48264);
or UO_2363 (O_2363,N_49095,N_49744);
or UO_2364 (O_2364,N_48969,N_47536);
nand UO_2365 (O_2365,N_49521,N_49074);
xor UO_2366 (O_2366,N_49668,N_49759);
xnor UO_2367 (O_2367,N_49605,N_49457);
nor UO_2368 (O_2368,N_49728,N_47733);
xor UO_2369 (O_2369,N_47733,N_49128);
xnor UO_2370 (O_2370,N_47712,N_48014);
nand UO_2371 (O_2371,N_48891,N_49437);
or UO_2372 (O_2372,N_48516,N_48442);
nand UO_2373 (O_2373,N_49065,N_48257);
xor UO_2374 (O_2374,N_47718,N_49205);
nand UO_2375 (O_2375,N_47671,N_48985);
nor UO_2376 (O_2376,N_47546,N_49212);
or UO_2377 (O_2377,N_48618,N_49667);
nand UO_2378 (O_2378,N_47569,N_49415);
and UO_2379 (O_2379,N_47969,N_49939);
nor UO_2380 (O_2380,N_48758,N_48475);
xor UO_2381 (O_2381,N_48946,N_48402);
xor UO_2382 (O_2382,N_48499,N_49545);
nand UO_2383 (O_2383,N_48717,N_48496);
nor UO_2384 (O_2384,N_49034,N_49100);
nand UO_2385 (O_2385,N_49759,N_49676);
xor UO_2386 (O_2386,N_49609,N_49276);
nand UO_2387 (O_2387,N_49457,N_49717);
nand UO_2388 (O_2388,N_49289,N_49038);
or UO_2389 (O_2389,N_48864,N_49167);
and UO_2390 (O_2390,N_49079,N_48430);
and UO_2391 (O_2391,N_47582,N_47726);
nor UO_2392 (O_2392,N_48728,N_47616);
nand UO_2393 (O_2393,N_48306,N_49471);
and UO_2394 (O_2394,N_49658,N_47544);
nor UO_2395 (O_2395,N_49292,N_47758);
nand UO_2396 (O_2396,N_49407,N_49393);
xnor UO_2397 (O_2397,N_49511,N_48861);
nand UO_2398 (O_2398,N_49762,N_49416);
and UO_2399 (O_2399,N_49118,N_47675);
or UO_2400 (O_2400,N_49732,N_47743);
xor UO_2401 (O_2401,N_48886,N_47966);
xnor UO_2402 (O_2402,N_47891,N_48787);
xor UO_2403 (O_2403,N_49977,N_49199);
nand UO_2404 (O_2404,N_47853,N_48416);
or UO_2405 (O_2405,N_48668,N_49910);
nand UO_2406 (O_2406,N_48641,N_48042);
xor UO_2407 (O_2407,N_49609,N_49004);
nand UO_2408 (O_2408,N_49881,N_49793);
xnor UO_2409 (O_2409,N_48156,N_48582);
or UO_2410 (O_2410,N_48192,N_49922);
or UO_2411 (O_2411,N_49901,N_49000);
xor UO_2412 (O_2412,N_47902,N_47516);
and UO_2413 (O_2413,N_49577,N_48754);
xnor UO_2414 (O_2414,N_49418,N_47822);
or UO_2415 (O_2415,N_48876,N_49142);
nand UO_2416 (O_2416,N_48747,N_47663);
and UO_2417 (O_2417,N_49924,N_49445);
and UO_2418 (O_2418,N_49077,N_47724);
xnor UO_2419 (O_2419,N_48670,N_48095);
and UO_2420 (O_2420,N_48450,N_48223);
or UO_2421 (O_2421,N_49097,N_48564);
xnor UO_2422 (O_2422,N_48919,N_48371);
nor UO_2423 (O_2423,N_48567,N_49771);
nor UO_2424 (O_2424,N_47735,N_49540);
nor UO_2425 (O_2425,N_48621,N_47641);
nand UO_2426 (O_2426,N_49286,N_48506);
and UO_2427 (O_2427,N_47539,N_49559);
nand UO_2428 (O_2428,N_49265,N_49520);
and UO_2429 (O_2429,N_49327,N_48573);
or UO_2430 (O_2430,N_48892,N_47703);
nand UO_2431 (O_2431,N_47861,N_49413);
xor UO_2432 (O_2432,N_47549,N_48110);
xnor UO_2433 (O_2433,N_48845,N_48640);
or UO_2434 (O_2434,N_48876,N_49544);
xnor UO_2435 (O_2435,N_48778,N_49159);
or UO_2436 (O_2436,N_49608,N_47650);
or UO_2437 (O_2437,N_49125,N_49581);
and UO_2438 (O_2438,N_49309,N_49079);
or UO_2439 (O_2439,N_47580,N_48645);
and UO_2440 (O_2440,N_48977,N_49177);
xnor UO_2441 (O_2441,N_49360,N_47609);
nand UO_2442 (O_2442,N_48681,N_48013);
nand UO_2443 (O_2443,N_48581,N_49356);
and UO_2444 (O_2444,N_48763,N_48455);
and UO_2445 (O_2445,N_49294,N_47622);
nor UO_2446 (O_2446,N_47685,N_47562);
nor UO_2447 (O_2447,N_48600,N_48234);
or UO_2448 (O_2448,N_49261,N_47550);
xor UO_2449 (O_2449,N_48776,N_47613);
nor UO_2450 (O_2450,N_49736,N_48822);
nor UO_2451 (O_2451,N_48327,N_48927);
and UO_2452 (O_2452,N_49415,N_48080);
and UO_2453 (O_2453,N_47655,N_48045);
xnor UO_2454 (O_2454,N_49865,N_48350);
xor UO_2455 (O_2455,N_48115,N_48777);
nor UO_2456 (O_2456,N_48716,N_49658);
or UO_2457 (O_2457,N_49881,N_49516);
nor UO_2458 (O_2458,N_49225,N_49538);
xor UO_2459 (O_2459,N_48971,N_49553);
xnor UO_2460 (O_2460,N_47837,N_49349);
or UO_2461 (O_2461,N_48593,N_48935);
xor UO_2462 (O_2462,N_48489,N_49626);
nand UO_2463 (O_2463,N_48323,N_47692);
xnor UO_2464 (O_2464,N_49453,N_49550);
nor UO_2465 (O_2465,N_48013,N_49500);
or UO_2466 (O_2466,N_48285,N_49453);
nor UO_2467 (O_2467,N_47576,N_48385);
and UO_2468 (O_2468,N_49504,N_48468);
and UO_2469 (O_2469,N_47816,N_49143);
and UO_2470 (O_2470,N_48424,N_48501);
and UO_2471 (O_2471,N_48757,N_49947);
xnor UO_2472 (O_2472,N_47747,N_48877);
nand UO_2473 (O_2473,N_48705,N_49813);
xor UO_2474 (O_2474,N_47827,N_49093);
xnor UO_2475 (O_2475,N_48990,N_48500);
nor UO_2476 (O_2476,N_48237,N_49980);
nor UO_2477 (O_2477,N_48183,N_49270);
xnor UO_2478 (O_2478,N_49933,N_48644);
nand UO_2479 (O_2479,N_49947,N_48451);
nand UO_2480 (O_2480,N_49277,N_47585);
xor UO_2481 (O_2481,N_49101,N_49717);
and UO_2482 (O_2482,N_49512,N_49205);
or UO_2483 (O_2483,N_49338,N_48103);
or UO_2484 (O_2484,N_49402,N_49849);
xnor UO_2485 (O_2485,N_49844,N_49256);
xnor UO_2486 (O_2486,N_48006,N_48223);
and UO_2487 (O_2487,N_49122,N_48186);
or UO_2488 (O_2488,N_48944,N_49424);
nand UO_2489 (O_2489,N_48903,N_49924);
nor UO_2490 (O_2490,N_47518,N_49794);
or UO_2491 (O_2491,N_49352,N_49506);
nand UO_2492 (O_2492,N_47982,N_48913);
nand UO_2493 (O_2493,N_49007,N_49354);
and UO_2494 (O_2494,N_48287,N_49753);
or UO_2495 (O_2495,N_49165,N_47779);
and UO_2496 (O_2496,N_49360,N_48867);
nor UO_2497 (O_2497,N_49862,N_49476);
nand UO_2498 (O_2498,N_49697,N_48288);
nand UO_2499 (O_2499,N_48477,N_49450);
xor UO_2500 (O_2500,N_48676,N_47946);
and UO_2501 (O_2501,N_48693,N_49369);
or UO_2502 (O_2502,N_49266,N_48675);
nand UO_2503 (O_2503,N_49743,N_47583);
nor UO_2504 (O_2504,N_49258,N_47633);
nand UO_2505 (O_2505,N_48583,N_47743);
nand UO_2506 (O_2506,N_48469,N_48449);
xnor UO_2507 (O_2507,N_49466,N_49781);
nand UO_2508 (O_2508,N_49055,N_49439);
xnor UO_2509 (O_2509,N_49433,N_49696);
or UO_2510 (O_2510,N_47935,N_48149);
or UO_2511 (O_2511,N_48439,N_47551);
nor UO_2512 (O_2512,N_48780,N_48702);
or UO_2513 (O_2513,N_48797,N_49312);
nor UO_2514 (O_2514,N_48424,N_48514);
nor UO_2515 (O_2515,N_48170,N_48939);
or UO_2516 (O_2516,N_47904,N_49923);
nor UO_2517 (O_2517,N_49430,N_48017);
nand UO_2518 (O_2518,N_49912,N_48697);
and UO_2519 (O_2519,N_47856,N_49094);
or UO_2520 (O_2520,N_48833,N_49659);
and UO_2521 (O_2521,N_48747,N_49142);
nor UO_2522 (O_2522,N_47591,N_48102);
nor UO_2523 (O_2523,N_48143,N_48533);
nor UO_2524 (O_2524,N_49370,N_48232);
or UO_2525 (O_2525,N_48936,N_49110);
xor UO_2526 (O_2526,N_48489,N_49830);
and UO_2527 (O_2527,N_48954,N_47758);
or UO_2528 (O_2528,N_49521,N_47643);
nand UO_2529 (O_2529,N_49166,N_47750);
nand UO_2530 (O_2530,N_48818,N_47584);
nand UO_2531 (O_2531,N_49921,N_49337);
nand UO_2532 (O_2532,N_49352,N_49816);
xnor UO_2533 (O_2533,N_48156,N_47824);
or UO_2534 (O_2534,N_49057,N_49577);
or UO_2535 (O_2535,N_49120,N_49665);
and UO_2536 (O_2536,N_49115,N_49370);
nand UO_2537 (O_2537,N_49775,N_48136);
xnor UO_2538 (O_2538,N_48090,N_48504);
or UO_2539 (O_2539,N_49494,N_49862);
nand UO_2540 (O_2540,N_48739,N_48716);
and UO_2541 (O_2541,N_49635,N_48125);
nor UO_2542 (O_2542,N_49817,N_49602);
xor UO_2543 (O_2543,N_47948,N_48678);
xor UO_2544 (O_2544,N_49728,N_49691);
and UO_2545 (O_2545,N_48990,N_49071);
nand UO_2546 (O_2546,N_47664,N_48383);
nand UO_2547 (O_2547,N_47587,N_49851);
nor UO_2548 (O_2548,N_47631,N_48237);
and UO_2549 (O_2549,N_48803,N_47599);
xnor UO_2550 (O_2550,N_49995,N_47621);
nor UO_2551 (O_2551,N_49222,N_49450);
xor UO_2552 (O_2552,N_49513,N_49747);
xor UO_2553 (O_2553,N_49692,N_48263);
and UO_2554 (O_2554,N_48934,N_49448);
or UO_2555 (O_2555,N_47890,N_48554);
or UO_2556 (O_2556,N_48952,N_49603);
nand UO_2557 (O_2557,N_49798,N_49015);
or UO_2558 (O_2558,N_49463,N_48874);
nor UO_2559 (O_2559,N_49301,N_48499);
or UO_2560 (O_2560,N_49003,N_48489);
or UO_2561 (O_2561,N_49260,N_47653);
nor UO_2562 (O_2562,N_47804,N_47817);
or UO_2563 (O_2563,N_48040,N_49924);
or UO_2564 (O_2564,N_49464,N_48727);
or UO_2565 (O_2565,N_48180,N_48666);
nand UO_2566 (O_2566,N_49404,N_47684);
and UO_2567 (O_2567,N_48151,N_49869);
nand UO_2568 (O_2568,N_49372,N_48990);
nand UO_2569 (O_2569,N_49244,N_49458);
nand UO_2570 (O_2570,N_47879,N_47626);
xnor UO_2571 (O_2571,N_47577,N_49453);
and UO_2572 (O_2572,N_48593,N_47992);
nand UO_2573 (O_2573,N_48370,N_49098);
and UO_2574 (O_2574,N_49895,N_49426);
xnor UO_2575 (O_2575,N_47857,N_48668);
and UO_2576 (O_2576,N_47669,N_49806);
and UO_2577 (O_2577,N_48222,N_49448);
nor UO_2578 (O_2578,N_49641,N_49964);
nor UO_2579 (O_2579,N_47831,N_48463);
nor UO_2580 (O_2580,N_48633,N_47532);
or UO_2581 (O_2581,N_47981,N_48748);
and UO_2582 (O_2582,N_48988,N_48634);
nor UO_2583 (O_2583,N_47778,N_49179);
xor UO_2584 (O_2584,N_47757,N_49878);
and UO_2585 (O_2585,N_48066,N_48211);
and UO_2586 (O_2586,N_49355,N_49017);
xor UO_2587 (O_2587,N_48053,N_47789);
xor UO_2588 (O_2588,N_49056,N_47502);
and UO_2589 (O_2589,N_49756,N_49931);
nor UO_2590 (O_2590,N_48169,N_49638);
nor UO_2591 (O_2591,N_48515,N_47836);
xnor UO_2592 (O_2592,N_48073,N_49159);
nand UO_2593 (O_2593,N_47976,N_48912);
and UO_2594 (O_2594,N_48071,N_48934);
or UO_2595 (O_2595,N_48063,N_47662);
xnor UO_2596 (O_2596,N_49799,N_49212);
nand UO_2597 (O_2597,N_47738,N_48893);
xnor UO_2598 (O_2598,N_48371,N_48216);
nor UO_2599 (O_2599,N_49480,N_48943);
nand UO_2600 (O_2600,N_48444,N_49083);
xor UO_2601 (O_2601,N_48007,N_47696);
nor UO_2602 (O_2602,N_49457,N_48338);
nor UO_2603 (O_2603,N_48199,N_48284);
nor UO_2604 (O_2604,N_49950,N_49033);
nand UO_2605 (O_2605,N_48430,N_48256);
xnor UO_2606 (O_2606,N_48783,N_48797);
xor UO_2607 (O_2607,N_48878,N_47932);
and UO_2608 (O_2608,N_48898,N_47773);
and UO_2609 (O_2609,N_47829,N_49560);
nand UO_2610 (O_2610,N_47539,N_49274);
nand UO_2611 (O_2611,N_49158,N_48105);
xor UO_2612 (O_2612,N_48414,N_48813);
xnor UO_2613 (O_2613,N_49671,N_49927);
or UO_2614 (O_2614,N_49698,N_48501);
nor UO_2615 (O_2615,N_48414,N_49439);
xnor UO_2616 (O_2616,N_48123,N_47938);
nor UO_2617 (O_2617,N_49556,N_48909);
and UO_2618 (O_2618,N_48378,N_48546);
xnor UO_2619 (O_2619,N_49370,N_48937);
nand UO_2620 (O_2620,N_48406,N_49833);
xor UO_2621 (O_2621,N_48239,N_49121);
and UO_2622 (O_2622,N_48466,N_48288);
nor UO_2623 (O_2623,N_48555,N_48522);
xnor UO_2624 (O_2624,N_47768,N_49740);
or UO_2625 (O_2625,N_48913,N_48967);
nand UO_2626 (O_2626,N_48820,N_49501);
nand UO_2627 (O_2627,N_48037,N_49667);
xnor UO_2628 (O_2628,N_48654,N_49193);
or UO_2629 (O_2629,N_48879,N_48243);
xnor UO_2630 (O_2630,N_47666,N_48726);
and UO_2631 (O_2631,N_49680,N_47594);
and UO_2632 (O_2632,N_47932,N_47996);
nor UO_2633 (O_2633,N_48861,N_49317);
and UO_2634 (O_2634,N_49293,N_49763);
xnor UO_2635 (O_2635,N_47720,N_48033);
and UO_2636 (O_2636,N_49511,N_49067);
and UO_2637 (O_2637,N_47989,N_48079);
and UO_2638 (O_2638,N_49333,N_47711);
nor UO_2639 (O_2639,N_48426,N_48166);
or UO_2640 (O_2640,N_49343,N_48346);
or UO_2641 (O_2641,N_49763,N_48508);
or UO_2642 (O_2642,N_48473,N_48186);
nor UO_2643 (O_2643,N_47546,N_47737);
and UO_2644 (O_2644,N_48958,N_48240);
nand UO_2645 (O_2645,N_48971,N_47867);
or UO_2646 (O_2646,N_48658,N_48775);
xor UO_2647 (O_2647,N_48818,N_48828);
nor UO_2648 (O_2648,N_49388,N_48975);
xor UO_2649 (O_2649,N_49843,N_48601);
xnor UO_2650 (O_2650,N_48967,N_48253);
nand UO_2651 (O_2651,N_47528,N_49537);
or UO_2652 (O_2652,N_48230,N_49529);
nand UO_2653 (O_2653,N_48127,N_47807);
xnor UO_2654 (O_2654,N_49650,N_47783);
or UO_2655 (O_2655,N_47943,N_48645);
nor UO_2656 (O_2656,N_49176,N_48339);
nor UO_2657 (O_2657,N_47585,N_49962);
or UO_2658 (O_2658,N_48261,N_48290);
or UO_2659 (O_2659,N_48433,N_49383);
and UO_2660 (O_2660,N_49084,N_49749);
and UO_2661 (O_2661,N_49745,N_48525);
xnor UO_2662 (O_2662,N_48709,N_49127);
and UO_2663 (O_2663,N_48841,N_49926);
nand UO_2664 (O_2664,N_49854,N_48935);
xor UO_2665 (O_2665,N_48659,N_49251);
or UO_2666 (O_2666,N_49777,N_49335);
nand UO_2667 (O_2667,N_47627,N_48123);
or UO_2668 (O_2668,N_49641,N_47629);
xor UO_2669 (O_2669,N_48456,N_48820);
or UO_2670 (O_2670,N_47994,N_48412);
xnor UO_2671 (O_2671,N_48721,N_48083);
nor UO_2672 (O_2672,N_49362,N_48983);
nor UO_2673 (O_2673,N_49782,N_49500);
xor UO_2674 (O_2674,N_49743,N_47958);
or UO_2675 (O_2675,N_48525,N_47969);
and UO_2676 (O_2676,N_48329,N_49648);
or UO_2677 (O_2677,N_49503,N_48335);
and UO_2678 (O_2678,N_49742,N_49499);
nand UO_2679 (O_2679,N_49589,N_48929);
nand UO_2680 (O_2680,N_48821,N_49184);
and UO_2681 (O_2681,N_48410,N_49766);
nor UO_2682 (O_2682,N_47934,N_49717);
and UO_2683 (O_2683,N_48994,N_49714);
or UO_2684 (O_2684,N_49910,N_49106);
and UO_2685 (O_2685,N_47790,N_49163);
nand UO_2686 (O_2686,N_48079,N_48082);
or UO_2687 (O_2687,N_47726,N_48278);
and UO_2688 (O_2688,N_49199,N_49629);
nand UO_2689 (O_2689,N_49197,N_48324);
and UO_2690 (O_2690,N_49270,N_48349);
nor UO_2691 (O_2691,N_48796,N_49758);
nand UO_2692 (O_2692,N_49633,N_47685);
or UO_2693 (O_2693,N_49734,N_48600);
nor UO_2694 (O_2694,N_49890,N_48022);
and UO_2695 (O_2695,N_49612,N_47851);
or UO_2696 (O_2696,N_49779,N_48008);
nand UO_2697 (O_2697,N_48266,N_47708);
and UO_2698 (O_2698,N_47650,N_47636);
nor UO_2699 (O_2699,N_49115,N_49488);
or UO_2700 (O_2700,N_49524,N_48525);
or UO_2701 (O_2701,N_49803,N_48133);
nor UO_2702 (O_2702,N_48972,N_47798);
nor UO_2703 (O_2703,N_48550,N_49453);
nor UO_2704 (O_2704,N_48285,N_47948);
or UO_2705 (O_2705,N_48700,N_49890);
and UO_2706 (O_2706,N_49134,N_48232);
xor UO_2707 (O_2707,N_49570,N_47834);
or UO_2708 (O_2708,N_49681,N_48267);
and UO_2709 (O_2709,N_49129,N_48627);
nor UO_2710 (O_2710,N_48727,N_48951);
nor UO_2711 (O_2711,N_48880,N_49241);
nor UO_2712 (O_2712,N_49881,N_49406);
nor UO_2713 (O_2713,N_49663,N_47959);
or UO_2714 (O_2714,N_47736,N_47667);
xor UO_2715 (O_2715,N_49677,N_48876);
and UO_2716 (O_2716,N_49529,N_48766);
and UO_2717 (O_2717,N_48438,N_49470);
and UO_2718 (O_2718,N_49900,N_49614);
nand UO_2719 (O_2719,N_49455,N_49111);
and UO_2720 (O_2720,N_48576,N_48307);
nand UO_2721 (O_2721,N_49716,N_49147);
xnor UO_2722 (O_2722,N_48276,N_48000);
or UO_2723 (O_2723,N_47662,N_48759);
nand UO_2724 (O_2724,N_47856,N_48214);
nor UO_2725 (O_2725,N_48183,N_48327);
nor UO_2726 (O_2726,N_47834,N_49642);
nand UO_2727 (O_2727,N_48892,N_49003);
xnor UO_2728 (O_2728,N_49953,N_48741);
nor UO_2729 (O_2729,N_48739,N_49731);
and UO_2730 (O_2730,N_49296,N_49798);
nand UO_2731 (O_2731,N_48581,N_49172);
and UO_2732 (O_2732,N_48319,N_47631);
or UO_2733 (O_2733,N_48230,N_48448);
and UO_2734 (O_2734,N_47537,N_48699);
or UO_2735 (O_2735,N_49436,N_49533);
nand UO_2736 (O_2736,N_48846,N_48121);
nor UO_2737 (O_2737,N_49401,N_48667);
and UO_2738 (O_2738,N_47628,N_48848);
xor UO_2739 (O_2739,N_47713,N_49217);
nor UO_2740 (O_2740,N_48779,N_47632);
nand UO_2741 (O_2741,N_49910,N_48688);
or UO_2742 (O_2742,N_48314,N_47578);
nor UO_2743 (O_2743,N_48810,N_48940);
and UO_2744 (O_2744,N_48548,N_48384);
and UO_2745 (O_2745,N_49066,N_48430);
nor UO_2746 (O_2746,N_48339,N_49772);
or UO_2747 (O_2747,N_47892,N_49607);
xor UO_2748 (O_2748,N_49457,N_47601);
nor UO_2749 (O_2749,N_48795,N_49233);
nand UO_2750 (O_2750,N_47765,N_48244);
nand UO_2751 (O_2751,N_49332,N_48914);
xor UO_2752 (O_2752,N_47773,N_49244);
or UO_2753 (O_2753,N_49595,N_47590);
xnor UO_2754 (O_2754,N_47505,N_48370);
or UO_2755 (O_2755,N_48752,N_49859);
xor UO_2756 (O_2756,N_49677,N_49988);
and UO_2757 (O_2757,N_49054,N_49161);
or UO_2758 (O_2758,N_47936,N_48611);
or UO_2759 (O_2759,N_48708,N_48493);
nand UO_2760 (O_2760,N_49085,N_49355);
and UO_2761 (O_2761,N_47964,N_48923);
or UO_2762 (O_2762,N_49816,N_48052);
nor UO_2763 (O_2763,N_48127,N_49843);
or UO_2764 (O_2764,N_47667,N_49688);
nand UO_2765 (O_2765,N_49652,N_49038);
or UO_2766 (O_2766,N_48970,N_48299);
nor UO_2767 (O_2767,N_48283,N_47550);
or UO_2768 (O_2768,N_48091,N_49372);
and UO_2769 (O_2769,N_48058,N_49494);
and UO_2770 (O_2770,N_49670,N_48320);
nand UO_2771 (O_2771,N_47795,N_49274);
nand UO_2772 (O_2772,N_48174,N_49310);
xnor UO_2773 (O_2773,N_48477,N_48175);
nand UO_2774 (O_2774,N_48930,N_49121);
and UO_2775 (O_2775,N_48005,N_47972);
or UO_2776 (O_2776,N_48466,N_49852);
or UO_2777 (O_2777,N_48503,N_47892);
nor UO_2778 (O_2778,N_49667,N_48943);
and UO_2779 (O_2779,N_48289,N_48017);
nor UO_2780 (O_2780,N_49753,N_49866);
nor UO_2781 (O_2781,N_48141,N_48478);
xnor UO_2782 (O_2782,N_49664,N_48604);
and UO_2783 (O_2783,N_49868,N_48585);
xnor UO_2784 (O_2784,N_48912,N_49910);
nand UO_2785 (O_2785,N_48119,N_47997);
nor UO_2786 (O_2786,N_49050,N_48798);
xnor UO_2787 (O_2787,N_47816,N_49217);
xnor UO_2788 (O_2788,N_48173,N_49650);
nand UO_2789 (O_2789,N_47949,N_48215);
xor UO_2790 (O_2790,N_47922,N_47674);
xor UO_2791 (O_2791,N_49425,N_48497);
or UO_2792 (O_2792,N_48730,N_48380);
nand UO_2793 (O_2793,N_47658,N_49367);
nand UO_2794 (O_2794,N_49905,N_47905);
xor UO_2795 (O_2795,N_48006,N_48812);
nand UO_2796 (O_2796,N_48182,N_48734);
nand UO_2797 (O_2797,N_48801,N_47682);
xor UO_2798 (O_2798,N_48836,N_48615);
nor UO_2799 (O_2799,N_49364,N_49822);
and UO_2800 (O_2800,N_49398,N_47719);
xor UO_2801 (O_2801,N_49572,N_48172);
or UO_2802 (O_2802,N_48889,N_49685);
nor UO_2803 (O_2803,N_49977,N_49975);
nor UO_2804 (O_2804,N_48145,N_48518);
nor UO_2805 (O_2805,N_48367,N_49828);
or UO_2806 (O_2806,N_48867,N_49503);
and UO_2807 (O_2807,N_49261,N_49701);
nand UO_2808 (O_2808,N_48636,N_49404);
nand UO_2809 (O_2809,N_49825,N_49369);
xor UO_2810 (O_2810,N_48795,N_48818);
and UO_2811 (O_2811,N_49531,N_48238);
nand UO_2812 (O_2812,N_49610,N_49555);
nor UO_2813 (O_2813,N_48802,N_49964);
or UO_2814 (O_2814,N_48791,N_47811);
nand UO_2815 (O_2815,N_49424,N_47819);
nor UO_2816 (O_2816,N_48945,N_49230);
or UO_2817 (O_2817,N_48857,N_47695);
or UO_2818 (O_2818,N_49160,N_47932);
or UO_2819 (O_2819,N_49351,N_47829);
nand UO_2820 (O_2820,N_48296,N_48940);
xor UO_2821 (O_2821,N_49204,N_49133);
xnor UO_2822 (O_2822,N_49052,N_49393);
nand UO_2823 (O_2823,N_49613,N_48414);
nor UO_2824 (O_2824,N_49162,N_48841);
or UO_2825 (O_2825,N_48176,N_49696);
xor UO_2826 (O_2826,N_48364,N_48287);
and UO_2827 (O_2827,N_49691,N_47821);
nand UO_2828 (O_2828,N_49849,N_48797);
or UO_2829 (O_2829,N_48343,N_47777);
xnor UO_2830 (O_2830,N_48529,N_48620);
or UO_2831 (O_2831,N_48738,N_48140);
nand UO_2832 (O_2832,N_48560,N_49016);
or UO_2833 (O_2833,N_47669,N_49789);
or UO_2834 (O_2834,N_47666,N_48195);
nand UO_2835 (O_2835,N_47736,N_48978);
and UO_2836 (O_2836,N_49932,N_48962);
nor UO_2837 (O_2837,N_48084,N_48119);
and UO_2838 (O_2838,N_49349,N_48681);
and UO_2839 (O_2839,N_49960,N_47673);
and UO_2840 (O_2840,N_49399,N_49313);
nand UO_2841 (O_2841,N_47682,N_49712);
or UO_2842 (O_2842,N_49139,N_48679);
nand UO_2843 (O_2843,N_49592,N_49311);
and UO_2844 (O_2844,N_48675,N_49392);
nor UO_2845 (O_2845,N_49839,N_48541);
or UO_2846 (O_2846,N_49930,N_49029);
nand UO_2847 (O_2847,N_48707,N_47689);
or UO_2848 (O_2848,N_47706,N_48491);
nor UO_2849 (O_2849,N_49676,N_47830);
xor UO_2850 (O_2850,N_49171,N_47780);
nor UO_2851 (O_2851,N_49375,N_47822);
or UO_2852 (O_2852,N_49414,N_49270);
xor UO_2853 (O_2853,N_48768,N_48564);
xnor UO_2854 (O_2854,N_48584,N_47932);
or UO_2855 (O_2855,N_48214,N_47524);
xnor UO_2856 (O_2856,N_49105,N_48783);
or UO_2857 (O_2857,N_49444,N_48452);
xor UO_2858 (O_2858,N_48419,N_48434);
or UO_2859 (O_2859,N_48188,N_49700);
nand UO_2860 (O_2860,N_49243,N_48481);
or UO_2861 (O_2861,N_49230,N_49458);
nand UO_2862 (O_2862,N_49802,N_49660);
or UO_2863 (O_2863,N_49996,N_47947);
nand UO_2864 (O_2864,N_48694,N_47741);
and UO_2865 (O_2865,N_49134,N_48936);
or UO_2866 (O_2866,N_49580,N_49108);
xnor UO_2867 (O_2867,N_49884,N_49560);
nand UO_2868 (O_2868,N_49408,N_49680);
and UO_2869 (O_2869,N_47592,N_48172);
nand UO_2870 (O_2870,N_49877,N_48583);
or UO_2871 (O_2871,N_47841,N_47794);
and UO_2872 (O_2872,N_47803,N_49961);
or UO_2873 (O_2873,N_49844,N_49466);
and UO_2874 (O_2874,N_49704,N_47605);
xor UO_2875 (O_2875,N_49836,N_47578);
nor UO_2876 (O_2876,N_48697,N_48653);
or UO_2877 (O_2877,N_49260,N_49379);
xnor UO_2878 (O_2878,N_48960,N_49440);
nand UO_2879 (O_2879,N_49628,N_48467);
or UO_2880 (O_2880,N_48047,N_48521);
nand UO_2881 (O_2881,N_49121,N_49282);
xnor UO_2882 (O_2882,N_49281,N_49851);
and UO_2883 (O_2883,N_48161,N_48301);
or UO_2884 (O_2884,N_48945,N_47804);
nand UO_2885 (O_2885,N_48382,N_48515);
nand UO_2886 (O_2886,N_48028,N_49960);
nand UO_2887 (O_2887,N_49620,N_49333);
nor UO_2888 (O_2888,N_47522,N_47656);
and UO_2889 (O_2889,N_48487,N_47549);
xor UO_2890 (O_2890,N_49103,N_48130);
nor UO_2891 (O_2891,N_47943,N_47859);
and UO_2892 (O_2892,N_49348,N_48394);
or UO_2893 (O_2893,N_48073,N_48909);
and UO_2894 (O_2894,N_49450,N_49889);
and UO_2895 (O_2895,N_49933,N_49895);
and UO_2896 (O_2896,N_49923,N_49162);
xor UO_2897 (O_2897,N_47679,N_49096);
nor UO_2898 (O_2898,N_49333,N_49104);
nor UO_2899 (O_2899,N_48956,N_49679);
or UO_2900 (O_2900,N_49789,N_47753);
nor UO_2901 (O_2901,N_48996,N_48329);
and UO_2902 (O_2902,N_49528,N_47566);
nand UO_2903 (O_2903,N_48212,N_48255);
xnor UO_2904 (O_2904,N_49570,N_48274);
and UO_2905 (O_2905,N_49275,N_49491);
and UO_2906 (O_2906,N_48182,N_48794);
xor UO_2907 (O_2907,N_48799,N_48384);
or UO_2908 (O_2908,N_49676,N_49851);
nor UO_2909 (O_2909,N_47725,N_49629);
and UO_2910 (O_2910,N_48581,N_48385);
and UO_2911 (O_2911,N_48492,N_49707);
nor UO_2912 (O_2912,N_47911,N_48926);
nand UO_2913 (O_2913,N_48639,N_48564);
and UO_2914 (O_2914,N_48133,N_48408);
xor UO_2915 (O_2915,N_48383,N_47850);
xnor UO_2916 (O_2916,N_49494,N_48701);
and UO_2917 (O_2917,N_48001,N_48221);
or UO_2918 (O_2918,N_49519,N_48637);
or UO_2919 (O_2919,N_49190,N_48641);
nor UO_2920 (O_2920,N_48338,N_49444);
or UO_2921 (O_2921,N_48913,N_49073);
and UO_2922 (O_2922,N_48574,N_49266);
nand UO_2923 (O_2923,N_48688,N_49118);
xnor UO_2924 (O_2924,N_48330,N_47726);
nor UO_2925 (O_2925,N_48847,N_48383);
nand UO_2926 (O_2926,N_48470,N_49539);
nand UO_2927 (O_2927,N_48202,N_48197);
xnor UO_2928 (O_2928,N_48460,N_48801);
nor UO_2929 (O_2929,N_48078,N_48418);
or UO_2930 (O_2930,N_47547,N_49149);
nor UO_2931 (O_2931,N_48419,N_48263);
nor UO_2932 (O_2932,N_49794,N_48192);
xor UO_2933 (O_2933,N_49701,N_47698);
xnor UO_2934 (O_2934,N_48777,N_49964);
nand UO_2935 (O_2935,N_49810,N_49942);
xor UO_2936 (O_2936,N_49920,N_49007);
nor UO_2937 (O_2937,N_48748,N_49341);
and UO_2938 (O_2938,N_49281,N_49717);
or UO_2939 (O_2939,N_48808,N_49418);
or UO_2940 (O_2940,N_49643,N_48345);
or UO_2941 (O_2941,N_47618,N_47661);
nand UO_2942 (O_2942,N_49207,N_48472);
nor UO_2943 (O_2943,N_49598,N_49788);
or UO_2944 (O_2944,N_47588,N_49427);
nor UO_2945 (O_2945,N_48912,N_48254);
nand UO_2946 (O_2946,N_47770,N_48033);
xnor UO_2947 (O_2947,N_49160,N_48247);
or UO_2948 (O_2948,N_49398,N_47809);
nand UO_2949 (O_2949,N_49513,N_48519);
and UO_2950 (O_2950,N_49212,N_49843);
or UO_2951 (O_2951,N_48049,N_48172);
nor UO_2952 (O_2952,N_48496,N_48304);
nor UO_2953 (O_2953,N_48426,N_48671);
and UO_2954 (O_2954,N_48597,N_49805);
and UO_2955 (O_2955,N_48144,N_49753);
nand UO_2956 (O_2956,N_48658,N_49959);
or UO_2957 (O_2957,N_49652,N_48597);
nor UO_2958 (O_2958,N_49567,N_49449);
nor UO_2959 (O_2959,N_49790,N_48269);
or UO_2960 (O_2960,N_49375,N_47884);
or UO_2961 (O_2961,N_49758,N_49268);
or UO_2962 (O_2962,N_48124,N_48263);
or UO_2963 (O_2963,N_47556,N_49121);
xnor UO_2964 (O_2964,N_48684,N_48619);
and UO_2965 (O_2965,N_49524,N_47712);
nor UO_2966 (O_2966,N_47934,N_47930);
xor UO_2967 (O_2967,N_48508,N_47676);
xnor UO_2968 (O_2968,N_48718,N_47788);
xor UO_2969 (O_2969,N_48939,N_48412);
xor UO_2970 (O_2970,N_49072,N_47977);
xnor UO_2971 (O_2971,N_49848,N_48106);
or UO_2972 (O_2972,N_48933,N_49047);
or UO_2973 (O_2973,N_47771,N_47511);
nor UO_2974 (O_2974,N_47825,N_47574);
xor UO_2975 (O_2975,N_49905,N_48966);
xor UO_2976 (O_2976,N_48326,N_48868);
or UO_2977 (O_2977,N_47511,N_48176);
nor UO_2978 (O_2978,N_49867,N_47868);
or UO_2979 (O_2979,N_49829,N_48262);
and UO_2980 (O_2980,N_48927,N_48816);
xnor UO_2981 (O_2981,N_49965,N_49266);
or UO_2982 (O_2982,N_48486,N_47789);
nand UO_2983 (O_2983,N_49121,N_49224);
xor UO_2984 (O_2984,N_49304,N_49761);
nand UO_2985 (O_2985,N_48017,N_48970);
xnor UO_2986 (O_2986,N_49436,N_48331);
and UO_2987 (O_2987,N_49302,N_49460);
xnor UO_2988 (O_2988,N_48048,N_47523);
xnor UO_2989 (O_2989,N_47543,N_48802);
xor UO_2990 (O_2990,N_47817,N_47699);
and UO_2991 (O_2991,N_47741,N_48320);
or UO_2992 (O_2992,N_47574,N_49408);
xnor UO_2993 (O_2993,N_49137,N_47616);
nor UO_2994 (O_2994,N_48254,N_48647);
nor UO_2995 (O_2995,N_47732,N_49930);
and UO_2996 (O_2996,N_48945,N_47850);
nand UO_2997 (O_2997,N_47874,N_48833);
nor UO_2998 (O_2998,N_49905,N_48994);
nand UO_2999 (O_2999,N_48027,N_48940);
or UO_3000 (O_3000,N_48102,N_48577);
and UO_3001 (O_3001,N_49414,N_49929);
xnor UO_3002 (O_3002,N_49670,N_47528);
nor UO_3003 (O_3003,N_49062,N_48477);
or UO_3004 (O_3004,N_49188,N_48171);
nand UO_3005 (O_3005,N_48263,N_49362);
xor UO_3006 (O_3006,N_47586,N_48033);
xnor UO_3007 (O_3007,N_49787,N_47765);
and UO_3008 (O_3008,N_48210,N_47738);
nand UO_3009 (O_3009,N_49462,N_49400);
and UO_3010 (O_3010,N_48834,N_49541);
nand UO_3011 (O_3011,N_49103,N_49879);
nor UO_3012 (O_3012,N_47853,N_47764);
nor UO_3013 (O_3013,N_47569,N_48498);
xnor UO_3014 (O_3014,N_47857,N_48000);
or UO_3015 (O_3015,N_48494,N_48913);
and UO_3016 (O_3016,N_49916,N_48022);
xor UO_3017 (O_3017,N_48896,N_49384);
and UO_3018 (O_3018,N_49699,N_49038);
nand UO_3019 (O_3019,N_47590,N_49408);
or UO_3020 (O_3020,N_49903,N_49166);
nand UO_3021 (O_3021,N_47756,N_48699);
nand UO_3022 (O_3022,N_48806,N_47728);
or UO_3023 (O_3023,N_48520,N_49988);
nor UO_3024 (O_3024,N_49861,N_47936);
or UO_3025 (O_3025,N_48189,N_48903);
xnor UO_3026 (O_3026,N_49428,N_48155);
xor UO_3027 (O_3027,N_48714,N_48643);
xor UO_3028 (O_3028,N_48642,N_48916);
xor UO_3029 (O_3029,N_48456,N_48202);
nand UO_3030 (O_3030,N_49049,N_47659);
nor UO_3031 (O_3031,N_49675,N_47865);
or UO_3032 (O_3032,N_49551,N_48169);
nand UO_3033 (O_3033,N_49136,N_48318);
or UO_3034 (O_3034,N_48741,N_48496);
and UO_3035 (O_3035,N_48702,N_49495);
nor UO_3036 (O_3036,N_48899,N_49014);
and UO_3037 (O_3037,N_49382,N_47716);
and UO_3038 (O_3038,N_49760,N_48932);
nor UO_3039 (O_3039,N_49723,N_49899);
xor UO_3040 (O_3040,N_49593,N_48410);
nand UO_3041 (O_3041,N_48901,N_47789);
nor UO_3042 (O_3042,N_47553,N_48961);
and UO_3043 (O_3043,N_47845,N_47582);
nor UO_3044 (O_3044,N_49283,N_48286);
or UO_3045 (O_3045,N_49690,N_47717);
xnor UO_3046 (O_3046,N_49912,N_49893);
nor UO_3047 (O_3047,N_47917,N_47877);
xor UO_3048 (O_3048,N_48710,N_47992);
nor UO_3049 (O_3049,N_48978,N_49569);
nor UO_3050 (O_3050,N_47680,N_47899);
nand UO_3051 (O_3051,N_49956,N_48837);
xor UO_3052 (O_3052,N_47725,N_49294);
or UO_3053 (O_3053,N_49584,N_47834);
nor UO_3054 (O_3054,N_48960,N_47831);
xor UO_3055 (O_3055,N_47618,N_49104);
nand UO_3056 (O_3056,N_49315,N_49366);
and UO_3057 (O_3057,N_49411,N_48894);
or UO_3058 (O_3058,N_49997,N_49033);
xor UO_3059 (O_3059,N_47572,N_49151);
nor UO_3060 (O_3060,N_47722,N_48778);
or UO_3061 (O_3061,N_48313,N_47750);
and UO_3062 (O_3062,N_47521,N_49680);
nor UO_3063 (O_3063,N_49435,N_49813);
or UO_3064 (O_3064,N_48137,N_49488);
xor UO_3065 (O_3065,N_48169,N_47932);
nor UO_3066 (O_3066,N_49507,N_48523);
nor UO_3067 (O_3067,N_49574,N_49986);
and UO_3068 (O_3068,N_49997,N_49581);
xor UO_3069 (O_3069,N_49804,N_48172);
nor UO_3070 (O_3070,N_49013,N_47640);
nand UO_3071 (O_3071,N_49964,N_47737);
nand UO_3072 (O_3072,N_48032,N_47963);
nor UO_3073 (O_3073,N_49300,N_48315);
or UO_3074 (O_3074,N_49042,N_47660);
nor UO_3075 (O_3075,N_48735,N_48621);
or UO_3076 (O_3076,N_48605,N_49928);
xnor UO_3077 (O_3077,N_48984,N_48127);
nand UO_3078 (O_3078,N_49236,N_49376);
and UO_3079 (O_3079,N_48953,N_48063);
xor UO_3080 (O_3080,N_49394,N_47803);
and UO_3081 (O_3081,N_48316,N_48093);
and UO_3082 (O_3082,N_49632,N_49581);
xor UO_3083 (O_3083,N_47957,N_48375);
and UO_3084 (O_3084,N_48868,N_48250);
nand UO_3085 (O_3085,N_49323,N_49589);
or UO_3086 (O_3086,N_48716,N_48361);
xor UO_3087 (O_3087,N_48024,N_49751);
or UO_3088 (O_3088,N_47930,N_47538);
nand UO_3089 (O_3089,N_47676,N_48838);
nor UO_3090 (O_3090,N_49788,N_49754);
or UO_3091 (O_3091,N_49383,N_49617);
or UO_3092 (O_3092,N_48829,N_48387);
or UO_3093 (O_3093,N_49171,N_48204);
and UO_3094 (O_3094,N_48509,N_47874);
xor UO_3095 (O_3095,N_47520,N_48065);
nor UO_3096 (O_3096,N_49150,N_49999);
xnor UO_3097 (O_3097,N_49538,N_49166);
xnor UO_3098 (O_3098,N_49383,N_47594);
nor UO_3099 (O_3099,N_48715,N_49047);
nor UO_3100 (O_3100,N_48503,N_48296);
or UO_3101 (O_3101,N_47850,N_49912);
nand UO_3102 (O_3102,N_49578,N_49333);
nor UO_3103 (O_3103,N_47916,N_48080);
or UO_3104 (O_3104,N_47633,N_48973);
nor UO_3105 (O_3105,N_49701,N_49558);
and UO_3106 (O_3106,N_49668,N_47874);
nor UO_3107 (O_3107,N_48539,N_48542);
or UO_3108 (O_3108,N_47914,N_49891);
nand UO_3109 (O_3109,N_48004,N_48888);
or UO_3110 (O_3110,N_48893,N_48343);
or UO_3111 (O_3111,N_49673,N_47662);
nand UO_3112 (O_3112,N_49440,N_47810);
and UO_3113 (O_3113,N_49209,N_48644);
nor UO_3114 (O_3114,N_49893,N_47747);
or UO_3115 (O_3115,N_47606,N_48400);
nand UO_3116 (O_3116,N_49337,N_47612);
nand UO_3117 (O_3117,N_48727,N_47866);
and UO_3118 (O_3118,N_49253,N_47583);
xor UO_3119 (O_3119,N_49034,N_48977);
nor UO_3120 (O_3120,N_48457,N_48797);
nor UO_3121 (O_3121,N_47818,N_47616);
xor UO_3122 (O_3122,N_49425,N_49781);
nor UO_3123 (O_3123,N_49644,N_49398);
and UO_3124 (O_3124,N_48911,N_48211);
xor UO_3125 (O_3125,N_48595,N_49641);
or UO_3126 (O_3126,N_47607,N_49269);
or UO_3127 (O_3127,N_48790,N_47824);
or UO_3128 (O_3128,N_49931,N_49375);
or UO_3129 (O_3129,N_48562,N_49756);
or UO_3130 (O_3130,N_49929,N_48450);
and UO_3131 (O_3131,N_49636,N_49002);
or UO_3132 (O_3132,N_48681,N_48133);
and UO_3133 (O_3133,N_47504,N_48600);
nor UO_3134 (O_3134,N_49034,N_48971);
xnor UO_3135 (O_3135,N_47950,N_48253);
xor UO_3136 (O_3136,N_49787,N_47862);
or UO_3137 (O_3137,N_48435,N_47910);
nand UO_3138 (O_3138,N_48556,N_47959);
nor UO_3139 (O_3139,N_47749,N_47887);
xor UO_3140 (O_3140,N_49463,N_49467);
xnor UO_3141 (O_3141,N_48931,N_48377);
nor UO_3142 (O_3142,N_48861,N_48630);
nand UO_3143 (O_3143,N_49633,N_48933);
and UO_3144 (O_3144,N_48555,N_48447);
and UO_3145 (O_3145,N_47816,N_48397);
or UO_3146 (O_3146,N_49801,N_48507);
nor UO_3147 (O_3147,N_48818,N_47789);
nand UO_3148 (O_3148,N_48845,N_49349);
nor UO_3149 (O_3149,N_49962,N_48300);
nand UO_3150 (O_3150,N_48125,N_48456);
nand UO_3151 (O_3151,N_49964,N_47740);
nand UO_3152 (O_3152,N_48881,N_49654);
nor UO_3153 (O_3153,N_47549,N_48262);
nand UO_3154 (O_3154,N_47561,N_48595);
or UO_3155 (O_3155,N_48366,N_49565);
nor UO_3156 (O_3156,N_49966,N_49370);
xnor UO_3157 (O_3157,N_49037,N_48331);
and UO_3158 (O_3158,N_48703,N_48033);
xor UO_3159 (O_3159,N_48622,N_47541);
nand UO_3160 (O_3160,N_49832,N_48203);
xor UO_3161 (O_3161,N_49487,N_49283);
nor UO_3162 (O_3162,N_47587,N_47989);
or UO_3163 (O_3163,N_47702,N_48430);
nand UO_3164 (O_3164,N_47644,N_49946);
or UO_3165 (O_3165,N_48390,N_47987);
and UO_3166 (O_3166,N_49128,N_48953);
xnor UO_3167 (O_3167,N_49297,N_48654);
or UO_3168 (O_3168,N_48326,N_48095);
nand UO_3169 (O_3169,N_49996,N_49093);
xor UO_3170 (O_3170,N_49022,N_48480);
and UO_3171 (O_3171,N_49835,N_48190);
or UO_3172 (O_3172,N_48137,N_47983);
or UO_3173 (O_3173,N_48964,N_48664);
or UO_3174 (O_3174,N_49290,N_47975);
nand UO_3175 (O_3175,N_48603,N_48430);
xnor UO_3176 (O_3176,N_49603,N_49248);
and UO_3177 (O_3177,N_48453,N_49491);
xnor UO_3178 (O_3178,N_48534,N_48401);
or UO_3179 (O_3179,N_48273,N_48397);
xor UO_3180 (O_3180,N_49393,N_49085);
xnor UO_3181 (O_3181,N_48588,N_47966);
xor UO_3182 (O_3182,N_47726,N_48988);
nand UO_3183 (O_3183,N_49530,N_47992);
or UO_3184 (O_3184,N_48298,N_48307);
nor UO_3185 (O_3185,N_48391,N_47917);
nor UO_3186 (O_3186,N_48526,N_48975);
and UO_3187 (O_3187,N_49049,N_47947);
nand UO_3188 (O_3188,N_49685,N_48735);
nand UO_3189 (O_3189,N_47594,N_47597);
or UO_3190 (O_3190,N_49103,N_48290);
nor UO_3191 (O_3191,N_49382,N_48222);
and UO_3192 (O_3192,N_48658,N_49776);
and UO_3193 (O_3193,N_49074,N_49753);
and UO_3194 (O_3194,N_47728,N_47906);
xor UO_3195 (O_3195,N_47639,N_48707);
nand UO_3196 (O_3196,N_48718,N_48695);
nor UO_3197 (O_3197,N_48686,N_48605);
nor UO_3198 (O_3198,N_47866,N_49607);
or UO_3199 (O_3199,N_48638,N_48761);
nand UO_3200 (O_3200,N_48156,N_48713);
nor UO_3201 (O_3201,N_49655,N_47828);
or UO_3202 (O_3202,N_48362,N_47839);
or UO_3203 (O_3203,N_49176,N_48719);
xor UO_3204 (O_3204,N_48468,N_48367);
and UO_3205 (O_3205,N_49866,N_49002);
and UO_3206 (O_3206,N_48074,N_48082);
or UO_3207 (O_3207,N_48011,N_49561);
and UO_3208 (O_3208,N_49897,N_49299);
or UO_3209 (O_3209,N_47616,N_47793);
xor UO_3210 (O_3210,N_47507,N_49495);
and UO_3211 (O_3211,N_49336,N_48366);
xor UO_3212 (O_3212,N_48117,N_49959);
nand UO_3213 (O_3213,N_47978,N_49817);
nand UO_3214 (O_3214,N_48237,N_47958);
nand UO_3215 (O_3215,N_49257,N_49521);
nor UO_3216 (O_3216,N_48219,N_48550);
or UO_3217 (O_3217,N_49597,N_48640);
and UO_3218 (O_3218,N_48191,N_48300);
nor UO_3219 (O_3219,N_48715,N_49429);
nor UO_3220 (O_3220,N_48865,N_47976);
nand UO_3221 (O_3221,N_48002,N_49510);
or UO_3222 (O_3222,N_47644,N_49254);
or UO_3223 (O_3223,N_48279,N_47502);
or UO_3224 (O_3224,N_48435,N_49370);
or UO_3225 (O_3225,N_49704,N_49015);
or UO_3226 (O_3226,N_47509,N_49628);
xor UO_3227 (O_3227,N_48094,N_47936);
and UO_3228 (O_3228,N_48831,N_48628);
xor UO_3229 (O_3229,N_48224,N_48049);
xnor UO_3230 (O_3230,N_48482,N_48275);
or UO_3231 (O_3231,N_49406,N_48903);
nor UO_3232 (O_3232,N_49052,N_48695);
xnor UO_3233 (O_3233,N_49217,N_47806);
or UO_3234 (O_3234,N_48261,N_49312);
nand UO_3235 (O_3235,N_48917,N_48961);
xnor UO_3236 (O_3236,N_48828,N_47784);
or UO_3237 (O_3237,N_48597,N_48526);
or UO_3238 (O_3238,N_47532,N_47686);
and UO_3239 (O_3239,N_48334,N_47694);
and UO_3240 (O_3240,N_49603,N_48366);
nand UO_3241 (O_3241,N_48324,N_49451);
and UO_3242 (O_3242,N_48533,N_48740);
xor UO_3243 (O_3243,N_47607,N_49869);
xor UO_3244 (O_3244,N_48313,N_49986);
nor UO_3245 (O_3245,N_49455,N_48191);
xor UO_3246 (O_3246,N_48117,N_47915);
xnor UO_3247 (O_3247,N_47591,N_49440);
or UO_3248 (O_3248,N_47574,N_48941);
nand UO_3249 (O_3249,N_47901,N_48376);
nor UO_3250 (O_3250,N_48170,N_49446);
or UO_3251 (O_3251,N_49132,N_48978);
and UO_3252 (O_3252,N_49729,N_48937);
nand UO_3253 (O_3253,N_49262,N_48246);
or UO_3254 (O_3254,N_47648,N_49649);
xnor UO_3255 (O_3255,N_49132,N_48204);
nand UO_3256 (O_3256,N_47895,N_49991);
or UO_3257 (O_3257,N_49987,N_48012);
and UO_3258 (O_3258,N_48039,N_48746);
or UO_3259 (O_3259,N_49272,N_48252);
and UO_3260 (O_3260,N_49266,N_47572);
or UO_3261 (O_3261,N_48606,N_49817);
and UO_3262 (O_3262,N_47921,N_48218);
xnor UO_3263 (O_3263,N_48758,N_47721);
nor UO_3264 (O_3264,N_48767,N_49433);
nand UO_3265 (O_3265,N_47616,N_48516);
or UO_3266 (O_3266,N_48774,N_47886);
xnor UO_3267 (O_3267,N_48280,N_47962);
or UO_3268 (O_3268,N_48028,N_47740);
and UO_3269 (O_3269,N_48609,N_49465);
nand UO_3270 (O_3270,N_47825,N_49464);
xnor UO_3271 (O_3271,N_49834,N_47982);
nor UO_3272 (O_3272,N_49209,N_47979);
or UO_3273 (O_3273,N_48130,N_49907);
nor UO_3274 (O_3274,N_49158,N_49204);
xnor UO_3275 (O_3275,N_47752,N_48525);
nand UO_3276 (O_3276,N_47983,N_49420);
xnor UO_3277 (O_3277,N_48856,N_49897);
and UO_3278 (O_3278,N_47873,N_48384);
xor UO_3279 (O_3279,N_48446,N_49135);
nor UO_3280 (O_3280,N_49546,N_47709);
nand UO_3281 (O_3281,N_49471,N_49507);
nor UO_3282 (O_3282,N_49726,N_49587);
and UO_3283 (O_3283,N_47629,N_48034);
nor UO_3284 (O_3284,N_49251,N_48990);
or UO_3285 (O_3285,N_49737,N_49405);
and UO_3286 (O_3286,N_49954,N_47607);
nand UO_3287 (O_3287,N_47781,N_48055);
or UO_3288 (O_3288,N_49579,N_47765);
or UO_3289 (O_3289,N_47770,N_49374);
and UO_3290 (O_3290,N_49546,N_47855);
nor UO_3291 (O_3291,N_47740,N_48323);
and UO_3292 (O_3292,N_47929,N_49556);
or UO_3293 (O_3293,N_49280,N_49788);
and UO_3294 (O_3294,N_48107,N_47524);
and UO_3295 (O_3295,N_48378,N_49410);
nand UO_3296 (O_3296,N_47886,N_48398);
xnor UO_3297 (O_3297,N_49753,N_48536);
nor UO_3298 (O_3298,N_48530,N_48660);
xnor UO_3299 (O_3299,N_47834,N_48600);
and UO_3300 (O_3300,N_49536,N_48830);
xnor UO_3301 (O_3301,N_48240,N_48740);
xnor UO_3302 (O_3302,N_49311,N_49730);
or UO_3303 (O_3303,N_49644,N_48365);
or UO_3304 (O_3304,N_48024,N_48862);
xnor UO_3305 (O_3305,N_47657,N_48030);
xor UO_3306 (O_3306,N_49299,N_49138);
xor UO_3307 (O_3307,N_49698,N_48833);
and UO_3308 (O_3308,N_48631,N_47779);
nor UO_3309 (O_3309,N_48053,N_47835);
xnor UO_3310 (O_3310,N_49952,N_49494);
nor UO_3311 (O_3311,N_49673,N_49387);
or UO_3312 (O_3312,N_49911,N_48493);
and UO_3313 (O_3313,N_49150,N_49446);
and UO_3314 (O_3314,N_49022,N_49855);
or UO_3315 (O_3315,N_48726,N_49169);
xor UO_3316 (O_3316,N_49692,N_49105);
xnor UO_3317 (O_3317,N_49838,N_48308);
nand UO_3318 (O_3318,N_48769,N_49910);
nor UO_3319 (O_3319,N_48852,N_48792);
xnor UO_3320 (O_3320,N_48646,N_48513);
and UO_3321 (O_3321,N_48975,N_49175);
xnor UO_3322 (O_3322,N_49901,N_49870);
nor UO_3323 (O_3323,N_49110,N_49258);
or UO_3324 (O_3324,N_48346,N_49080);
or UO_3325 (O_3325,N_47876,N_49131);
or UO_3326 (O_3326,N_47965,N_49798);
or UO_3327 (O_3327,N_48089,N_47719);
nand UO_3328 (O_3328,N_49649,N_48138);
and UO_3329 (O_3329,N_48209,N_48846);
xnor UO_3330 (O_3330,N_48190,N_48818);
nor UO_3331 (O_3331,N_47607,N_49024);
and UO_3332 (O_3332,N_48288,N_48011);
xnor UO_3333 (O_3333,N_49741,N_47733);
or UO_3334 (O_3334,N_49422,N_49423);
nand UO_3335 (O_3335,N_49246,N_47545);
and UO_3336 (O_3336,N_49225,N_49309);
nor UO_3337 (O_3337,N_49390,N_49983);
or UO_3338 (O_3338,N_49500,N_49089);
and UO_3339 (O_3339,N_49689,N_49302);
or UO_3340 (O_3340,N_49369,N_49957);
or UO_3341 (O_3341,N_49090,N_48270);
nand UO_3342 (O_3342,N_49801,N_47852);
nor UO_3343 (O_3343,N_48389,N_47993);
nor UO_3344 (O_3344,N_48571,N_48950);
nand UO_3345 (O_3345,N_47995,N_48339);
nand UO_3346 (O_3346,N_49539,N_49175);
or UO_3347 (O_3347,N_48125,N_49875);
xnor UO_3348 (O_3348,N_48777,N_47842);
and UO_3349 (O_3349,N_48554,N_47863);
and UO_3350 (O_3350,N_47666,N_49070);
or UO_3351 (O_3351,N_48247,N_49351);
nand UO_3352 (O_3352,N_49349,N_49779);
or UO_3353 (O_3353,N_49252,N_48500);
or UO_3354 (O_3354,N_48077,N_48480);
or UO_3355 (O_3355,N_48629,N_49590);
nor UO_3356 (O_3356,N_48008,N_49112);
and UO_3357 (O_3357,N_48269,N_48831);
or UO_3358 (O_3358,N_49149,N_47895);
nand UO_3359 (O_3359,N_47533,N_49824);
xnor UO_3360 (O_3360,N_47720,N_48464);
xnor UO_3361 (O_3361,N_49503,N_49666);
nand UO_3362 (O_3362,N_47655,N_48867);
or UO_3363 (O_3363,N_49704,N_48394);
or UO_3364 (O_3364,N_48452,N_49109);
or UO_3365 (O_3365,N_49063,N_49577);
or UO_3366 (O_3366,N_49101,N_48126);
and UO_3367 (O_3367,N_48483,N_48050);
or UO_3368 (O_3368,N_48476,N_49368);
nor UO_3369 (O_3369,N_48778,N_47614);
nor UO_3370 (O_3370,N_49737,N_49862);
nor UO_3371 (O_3371,N_47630,N_49803);
and UO_3372 (O_3372,N_49527,N_47510);
or UO_3373 (O_3373,N_48116,N_48560);
and UO_3374 (O_3374,N_47522,N_49633);
nand UO_3375 (O_3375,N_48011,N_48603);
nand UO_3376 (O_3376,N_48327,N_49778);
or UO_3377 (O_3377,N_48593,N_49611);
nand UO_3378 (O_3378,N_47725,N_47753);
or UO_3379 (O_3379,N_48714,N_48982);
and UO_3380 (O_3380,N_49202,N_49987);
nor UO_3381 (O_3381,N_48764,N_47629);
nand UO_3382 (O_3382,N_49961,N_48606);
or UO_3383 (O_3383,N_49066,N_49123);
or UO_3384 (O_3384,N_48355,N_47942);
xor UO_3385 (O_3385,N_49605,N_48281);
or UO_3386 (O_3386,N_48974,N_47813);
nand UO_3387 (O_3387,N_48246,N_48863);
nand UO_3388 (O_3388,N_49480,N_48278);
and UO_3389 (O_3389,N_49464,N_47731);
and UO_3390 (O_3390,N_48626,N_47574);
xor UO_3391 (O_3391,N_49654,N_47576);
or UO_3392 (O_3392,N_47628,N_49289);
and UO_3393 (O_3393,N_48741,N_48710);
nand UO_3394 (O_3394,N_49662,N_49593);
or UO_3395 (O_3395,N_49491,N_49211);
and UO_3396 (O_3396,N_49342,N_49537);
xnor UO_3397 (O_3397,N_49464,N_49227);
nand UO_3398 (O_3398,N_49686,N_49629);
nand UO_3399 (O_3399,N_48741,N_48621);
nor UO_3400 (O_3400,N_48558,N_47986);
xnor UO_3401 (O_3401,N_48529,N_48066);
and UO_3402 (O_3402,N_47553,N_49293);
nand UO_3403 (O_3403,N_48900,N_48175);
xor UO_3404 (O_3404,N_47654,N_49864);
or UO_3405 (O_3405,N_47843,N_48956);
and UO_3406 (O_3406,N_49230,N_48690);
xnor UO_3407 (O_3407,N_49969,N_48358);
xor UO_3408 (O_3408,N_48140,N_49265);
and UO_3409 (O_3409,N_48536,N_48206);
xor UO_3410 (O_3410,N_48350,N_47727);
nand UO_3411 (O_3411,N_47614,N_49825);
or UO_3412 (O_3412,N_47976,N_47920);
xor UO_3413 (O_3413,N_48483,N_49338);
xor UO_3414 (O_3414,N_48208,N_48222);
or UO_3415 (O_3415,N_48050,N_49041);
or UO_3416 (O_3416,N_49796,N_48068);
nor UO_3417 (O_3417,N_48106,N_47832);
nor UO_3418 (O_3418,N_48763,N_49682);
or UO_3419 (O_3419,N_48093,N_49677);
and UO_3420 (O_3420,N_48701,N_47640);
and UO_3421 (O_3421,N_49933,N_48810);
xor UO_3422 (O_3422,N_48568,N_48551);
xnor UO_3423 (O_3423,N_47845,N_47819);
nand UO_3424 (O_3424,N_48672,N_48643);
or UO_3425 (O_3425,N_48802,N_49591);
or UO_3426 (O_3426,N_48597,N_48398);
or UO_3427 (O_3427,N_47547,N_47549);
nor UO_3428 (O_3428,N_49420,N_49853);
nor UO_3429 (O_3429,N_49621,N_48432);
xor UO_3430 (O_3430,N_48682,N_47737);
xor UO_3431 (O_3431,N_49784,N_48499);
nor UO_3432 (O_3432,N_48339,N_48916);
xnor UO_3433 (O_3433,N_48342,N_49336);
xor UO_3434 (O_3434,N_49121,N_48644);
or UO_3435 (O_3435,N_49265,N_48266);
xnor UO_3436 (O_3436,N_49675,N_47907);
nand UO_3437 (O_3437,N_48241,N_47762);
xnor UO_3438 (O_3438,N_49075,N_47845);
and UO_3439 (O_3439,N_49193,N_47549);
xor UO_3440 (O_3440,N_47665,N_49895);
or UO_3441 (O_3441,N_49863,N_48972);
or UO_3442 (O_3442,N_49766,N_48168);
and UO_3443 (O_3443,N_47524,N_48331);
or UO_3444 (O_3444,N_47688,N_47626);
nand UO_3445 (O_3445,N_47681,N_49117);
nand UO_3446 (O_3446,N_47920,N_49123);
or UO_3447 (O_3447,N_48683,N_49883);
or UO_3448 (O_3448,N_49703,N_49707);
xnor UO_3449 (O_3449,N_49619,N_49151);
and UO_3450 (O_3450,N_48123,N_48883);
or UO_3451 (O_3451,N_48699,N_48832);
or UO_3452 (O_3452,N_48803,N_47680);
xor UO_3453 (O_3453,N_48450,N_48665);
nand UO_3454 (O_3454,N_49392,N_49623);
or UO_3455 (O_3455,N_48483,N_49320);
nor UO_3456 (O_3456,N_49056,N_47617);
nor UO_3457 (O_3457,N_48651,N_48847);
or UO_3458 (O_3458,N_49680,N_49251);
nor UO_3459 (O_3459,N_48158,N_49645);
or UO_3460 (O_3460,N_49696,N_48690);
or UO_3461 (O_3461,N_48062,N_47597);
xnor UO_3462 (O_3462,N_49177,N_49881);
nor UO_3463 (O_3463,N_48803,N_47620);
and UO_3464 (O_3464,N_49855,N_47882);
or UO_3465 (O_3465,N_48375,N_49816);
nand UO_3466 (O_3466,N_47562,N_47561);
and UO_3467 (O_3467,N_47506,N_49800);
or UO_3468 (O_3468,N_49227,N_47605);
and UO_3469 (O_3469,N_48328,N_47554);
or UO_3470 (O_3470,N_47575,N_48309);
or UO_3471 (O_3471,N_48723,N_48575);
xor UO_3472 (O_3472,N_47886,N_49833);
nor UO_3473 (O_3473,N_47978,N_47654);
nor UO_3474 (O_3474,N_49936,N_48996);
or UO_3475 (O_3475,N_49004,N_48976);
and UO_3476 (O_3476,N_49686,N_47980);
nand UO_3477 (O_3477,N_48746,N_48639);
nand UO_3478 (O_3478,N_47678,N_47790);
and UO_3479 (O_3479,N_47606,N_47898);
xor UO_3480 (O_3480,N_47682,N_48446);
and UO_3481 (O_3481,N_47808,N_48291);
nand UO_3482 (O_3482,N_48063,N_49746);
and UO_3483 (O_3483,N_49607,N_48721);
nor UO_3484 (O_3484,N_48196,N_49365);
xor UO_3485 (O_3485,N_49702,N_49764);
or UO_3486 (O_3486,N_49662,N_48608);
and UO_3487 (O_3487,N_49842,N_49565);
nor UO_3488 (O_3488,N_48798,N_48408);
and UO_3489 (O_3489,N_48426,N_49628);
and UO_3490 (O_3490,N_49077,N_48916);
xnor UO_3491 (O_3491,N_47878,N_49022);
nor UO_3492 (O_3492,N_47862,N_49834);
nand UO_3493 (O_3493,N_49231,N_48822);
nand UO_3494 (O_3494,N_49871,N_49142);
nor UO_3495 (O_3495,N_48418,N_47987);
or UO_3496 (O_3496,N_48502,N_48421);
nand UO_3497 (O_3497,N_47564,N_47646);
nor UO_3498 (O_3498,N_48263,N_48671);
or UO_3499 (O_3499,N_49856,N_48888);
or UO_3500 (O_3500,N_49506,N_48626);
and UO_3501 (O_3501,N_49944,N_47998);
nor UO_3502 (O_3502,N_49895,N_49791);
and UO_3503 (O_3503,N_47656,N_48566);
nand UO_3504 (O_3504,N_48499,N_48151);
nand UO_3505 (O_3505,N_49641,N_49284);
and UO_3506 (O_3506,N_47673,N_48456);
nor UO_3507 (O_3507,N_49209,N_47742);
nor UO_3508 (O_3508,N_47584,N_47723);
or UO_3509 (O_3509,N_49256,N_47946);
xnor UO_3510 (O_3510,N_49048,N_48766);
xnor UO_3511 (O_3511,N_47937,N_49693);
or UO_3512 (O_3512,N_48067,N_49259);
or UO_3513 (O_3513,N_48730,N_48902);
and UO_3514 (O_3514,N_49331,N_49245);
xnor UO_3515 (O_3515,N_48240,N_49155);
nor UO_3516 (O_3516,N_48176,N_49052);
nor UO_3517 (O_3517,N_49356,N_49924);
nand UO_3518 (O_3518,N_49087,N_49049);
xnor UO_3519 (O_3519,N_49263,N_48968);
nor UO_3520 (O_3520,N_49056,N_47959);
and UO_3521 (O_3521,N_47973,N_48233);
xor UO_3522 (O_3522,N_48207,N_48886);
nor UO_3523 (O_3523,N_48769,N_48535);
xor UO_3524 (O_3524,N_48943,N_48831);
nand UO_3525 (O_3525,N_48782,N_47516);
nor UO_3526 (O_3526,N_49192,N_48980);
nand UO_3527 (O_3527,N_48406,N_47896);
and UO_3528 (O_3528,N_48728,N_48563);
nor UO_3529 (O_3529,N_49357,N_48495);
nand UO_3530 (O_3530,N_49642,N_48967);
nor UO_3531 (O_3531,N_47546,N_47826);
and UO_3532 (O_3532,N_49164,N_49751);
or UO_3533 (O_3533,N_49836,N_47750);
nand UO_3534 (O_3534,N_49050,N_48820);
nand UO_3535 (O_3535,N_49035,N_49540);
nand UO_3536 (O_3536,N_48196,N_49180);
nand UO_3537 (O_3537,N_48395,N_47935);
or UO_3538 (O_3538,N_49667,N_49708);
or UO_3539 (O_3539,N_47953,N_49259);
and UO_3540 (O_3540,N_48114,N_47681);
or UO_3541 (O_3541,N_49079,N_48050);
or UO_3542 (O_3542,N_49882,N_49767);
nor UO_3543 (O_3543,N_49248,N_48908);
nor UO_3544 (O_3544,N_48337,N_49520);
xor UO_3545 (O_3545,N_49773,N_48845);
xnor UO_3546 (O_3546,N_48244,N_47858);
xnor UO_3547 (O_3547,N_49823,N_49396);
and UO_3548 (O_3548,N_48518,N_48557);
xnor UO_3549 (O_3549,N_48728,N_48171);
and UO_3550 (O_3550,N_48423,N_48766);
and UO_3551 (O_3551,N_48263,N_47946);
and UO_3552 (O_3552,N_49652,N_49870);
or UO_3553 (O_3553,N_48754,N_49149);
xor UO_3554 (O_3554,N_48066,N_49224);
nand UO_3555 (O_3555,N_49846,N_48355);
xnor UO_3556 (O_3556,N_48507,N_49798);
nand UO_3557 (O_3557,N_49259,N_49002);
xnor UO_3558 (O_3558,N_49011,N_47636);
or UO_3559 (O_3559,N_49416,N_48662);
nand UO_3560 (O_3560,N_48238,N_49617);
nor UO_3561 (O_3561,N_47725,N_47880);
or UO_3562 (O_3562,N_48789,N_49183);
and UO_3563 (O_3563,N_48540,N_48608);
nor UO_3564 (O_3564,N_49738,N_49316);
xnor UO_3565 (O_3565,N_49954,N_48044);
xnor UO_3566 (O_3566,N_49543,N_49127);
and UO_3567 (O_3567,N_49320,N_49459);
xnor UO_3568 (O_3568,N_49485,N_49547);
and UO_3569 (O_3569,N_48604,N_47591);
xnor UO_3570 (O_3570,N_48352,N_49250);
nor UO_3571 (O_3571,N_49194,N_49609);
and UO_3572 (O_3572,N_48440,N_48616);
or UO_3573 (O_3573,N_47920,N_49693);
or UO_3574 (O_3574,N_47584,N_49586);
xnor UO_3575 (O_3575,N_48159,N_48270);
or UO_3576 (O_3576,N_47885,N_48060);
nor UO_3577 (O_3577,N_48168,N_49913);
xnor UO_3578 (O_3578,N_48729,N_48887);
and UO_3579 (O_3579,N_49015,N_49148);
and UO_3580 (O_3580,N_48700,N_47730);
and UO_3581 (O_3581,N_48042,N_48245);
or UO_3582 (O_3582,N_49248,N_48509);
nor UO_3583 (O_3583,N_47898,N_47748);
nand UO_3584 (O_3584,N_49780,N_48384);
and UO_3585 (O_3585,N_49788,N_48452);
or UO_3586 (O_3586,N_48767,N_48327);
nand UO_3587 (O_3587,N_47578,N_47570);
nand UO_3588 (O_3588,N_49227,N_49677);
and UO_3589 (O_3589,N_47571,N_47963);
and UO_3590 (O_3590,N_49600,N_48267);
nand UO_3591 (O_3591,N_48380,N_48096);
or UO_3592 (O_3592,N_49446,N_47795);
nand UO_3593 (O_3593,N_47644,N_49613);
or UO_3594 (O_3594,N_49951,N_49099);
nor UO_3595 (O_3595,N_47628,N_47602);
nand UO_3596 (O_3596,N_48396,N_47869);
and UO_3597 (O_3597,N_49993,N_48093);
nor UO_3598 (O_3598,N_47587,N_47933);
xor UO_3599 (O_3599,N_48972,N_48976);
or UO_3600 (O_3600,N_47894,N_49847);
and UO_3601 (O_3601,N_48680,N_48177);
xor UO_3602 (O_3602,N_49661,N_48566);
xnor UO_3603 (O_3603,N_49532,N_48711);
nor UO_3604 (O_3604,N_48893,N_47652);
and UO_3605 (O_3605,N_48506,N_47597);
or UO_3606 (O_3606,N_48713,N_49741);
or UO_3607 (O_3607,N_48792,N_48761);
nor UO_3608 (O_3608,N_48863,N_48158);
or UO_3609 (O_3609,N_48314,N_48572);
nand UO_3610 (O_3610,N_48452,N_49018);
nand UO_3611 (O_3611,N_47937,N_48821);
nor UO_3612 (O_3612,N_47932,N_49229);
nor UO_3613 (O_3613,N_49813,N_49420);
or UO_3614 (O_3614,N_49813,N_49671);
nor UO_3615 (O_3615,N_47692,N_49575);
and UO_3616 (O_3616,N_48240,N_48777);
nand UO_3617 (O_3617,N_48615,N_49743);
and UO_3618 (O_3618,N_48356,N_49850);
and UO_3619 (O_3619,N_48620,N_49196);
nor UO_3620 (O_3620,N_47970,N_48731);
nor UO_3621 (O_3621,N_49036,N_49023);
or UO_3622 (O_3622,N_48734,N_49630);
nor UO_3623 (O_3623,N_49453,N_49936);
nor UO_3624 (O_3624,N_48236,N_49766);
nor UO_3625 (O_3625,N_47866,N_48175);
xnor UO_3626 (O_3626,N_48401,N_47762);
and UO_3627 (O_3627,N_48005,N_49536);
nand UO_3628 (O_3628,N_49190,N_48453);
xnor UO_3629 (O_3629,N_49663,N_49467);
and UO_3630 (O_3630,N_49644,N_49427);
nand UO_3631 (O_3631,N_49373,N_49488);
or UO_3632 (O_3632,N_49782,N_49567);
or UO_3633 (O_3633,N_48539,N_48357);
and UO_3634 (O_3634,N_49793,N_49444);
and UO_3635 (O_3635,N_48819,N_47881);
or UO_3636 (O_3636,N_48939,N_48100);
and UO_3637 (O_3637,N_49128,N_48431);
xnor UO_3638 (O_3638,N_49570,N_47515);
and UO_3639 (O_3639,N_48509,N_49867);
xor UO_3640 (O_3640,N_47655,N_49841);
nor UO_3641 (O_3641,N_47942,N_48456);
xnor UO_3642 (O_3642,N_48136,N_49061);
and UO_3643 (O_3643,N_49179,N_47908);
and UO_3644 (O_3644,N_47753,N_49886);
nor UO_3645 (O_3645,N_48886,N_48999);
xnor UO_3646 (O_3646,N_49911,N_47978);
and UO_3647 (O_3647,N_49006,N_49432);
nor UO_3648 (O_3648,N_48743,N_47753);
and UO_3649 (O_3649,N_48719,N_48627);
and UO_3650 (O_3650,N_49155,N_49022);
nand UO_3651 (O_3651,N_48710,N_49902);
or UO_3652 (O_3652,N_48308,N_48141);
nand UO_3653 (O_3653,N_48846,N_48277);
nand UO_3654 (O_3654,N_47835,N_48349);
or UO_3655 (O_3655,N_49721,N_49513);
or UO_3656 (O_3656,N_47505,N_49351);
xor UO_3657 (O_3657,N_48360,N_49677);
and UO_3658 (O_3658,N_48555,N_48469);
xor UO_3659 (O_3659,N_49861,N_48524);
nor UO_3660 (O_3660,N_49979,N_49152);
xor UO_3661 (O_3661,N_49078,N_49636);
nor UO_3662 (O_3662,N_48745,N_47680);
and UO_3663 (O_3663,N_49141,N_48941);
nand UO_3664 (O_3664,N_49559,N_47993);
nor UO_3665 (O_3665,N_49237,N_49260);
xnor UO_3666 (O_3666,N_48604,N_48744);
nor UO_3667 (O_3667,N_48633,N_48435);
and UO_3668 (O_3668,N_49419,N_49718);
or UO_3669 (O_3669,N_48305,N_48339);
nor UO_3670 (O_3670,N_47981,N_49388);
nand UO_3671 (O_3671,N_49454,N_48580);
xnor UO_3672 (O_3672,N_48406,N_49823);
or UO_3673 (O_3673,N_49973,N_48932);
xnor UO_3674 (O_3674,N_48377,N_48343);
nor UO_3675 (O_3675,N_48302,N_48866);
nand UO_3676 (O_3676,N_48614,N_49861);
nor UO_3677 (O_3677,N_49419,N_48764);
and UO_3678 (O_3678,N_49585,N_48659);
nand UO_3679 (O_3679,N_47963,N_48642);
xor UO_3680 (O_3680,N_49589,N_49903);
xor UO_3681 (O_3681,N_48445,N_48408);
nand UO_3682 (O_3682,N_48334,N_48230);
or UO_3683 (O_3683,N_48204,N_49406);
or UO_3684 (O_3684,N_47924,N_49231);
or UO_3685 (O_3685,N_49110,N_48181);
and UO_3686 (O_3686,N_48460,N_48463);
xnor UO_3687 (O_3687,N_49354,N_48951);
nor UO_3688 (O_3688,N_48196,N_47768);
nor UO_3689 (O_3689,N_48775,N_49760);
nor UO_3690 (O_3690,N_48702,N_49194);
nand UO_3691 (O_3691,N_48988,N_47563);
and UO_3692 (O_3692,N_47756,N_49766);
and UO_3693 (O_3693,N_48855,N_48858);
or UO_3694 (O_3694,N_47513,N_47711);
xnor UO_3695 (O_3695,N_48061,N_48593);
nand UO_3696 (O_3696,N_48605,N_49192);
or UO_3697 (O_3697,N_48007,N_49859);
nor UO_3698 (O_3698,N_49638,N_48266);
or UO_3699 (O_3699,N_48307,N_49195);
or UO_3700 (O_3700,N_48255,N_49213);
or UO_3701 (O_3701,N_47534,N_48923);
nor UO_3702 (O_3702,N_49133,N_48943);
xor UO_3703 (O_3703,N_49747,N_49527);
nand UO_3704 (O_3704,N_48142,N_47636);
or UO_3705 (O_3705,N_48607,N_49897);
nand UO_3706 (O_3706,N_49358,N_48831);
nor UO_3707 (O_3707,N_47782,N_49929);
xnor UO_3708 (O_3708,N_48751,N_48517);
xnor UO_3709 (O_3709,N_49475,N_48526);
nor UO_3710 (O_3710,N_49996,N_47612);
nor UO_3711 (O_3711,N_49337,N_49751);
nor UO_3712 (O_3712,N_49672,N_48891);
nand UO_3713 (O_3713,N_48575,N_47739);
or UO_3714 (O_3714,N_49226,N_48164);
xnor UO_3715 (O_3715,N_47678,N_49528);
and UO_3716 (O_3716,N_48745,N_48976);
nand UO_3717 (O_3717,N_48440,N_47838);
xnor UO_3718 (O_3718,N_49018,N_47966);
or UO_3719 (O_3719,N_48015,N_49204);
nor UO_3720 (O_3720,N_47635,N_48600);
and UO_3721 (O_3721,N_49349,N_47657);
xnor UO_3722 (O_3722,N_48664,N_47717);
nand UO_3723 (O_3723,N_48180,N_48254);
or UO_3724 (O_3724,N_48033,N_47589);
xor UO_3725 (O_3725,N_48122,N_48915);
xor UO_3726 (O_3726,N_47577,N_49499);
nand UO_3727 (O_3727,N_48870,N_49465);
xnor UO_3728 (O_3728,N_49073,N_47852);
nand UO_3729 (O_3729,N_48367,N_47822);
xnor UO_3730 (O_3730,N_48524,N_49519);
nor UO_3731 (O_3731,N_48117,N_48709);
xor UO_3732 (O_3732,N_48217,N_48441);
or UO_3733 (O_3733,N_49585,N_47915);
nand UO_3734 (O_3734,N_48655,N_48393);
nand UO_3735 (O_3735,N_49283,N_48880);
xnor UO_3736 (O_3736,N_48268,N_48326);
xnor UO_3737 (O_3737,N_48326,N_48654);
xnor UO_3738 (O_3738,N_47593,N_49136);
nand UO_3739 (O_3739,N_49025,N_49239);
or UO_3740 (O_3740,N_49254,N_49774);
or UO_3741 (O_3741,N_49295,N_49480);
or UO_3742 (O_3742,N_49691,N_47804);
nor UO_3743 (O_3743,N_48884,N_48524);
nor UO_3744 (O_3744,N_47619,N_47539);
nand UO_3745 (O_3745,N_49494,N_48699);
nor UO_3746 (O_3746,N_48699,N_48282);
and UO_3747 (O_3747,N_47557,N_48684);
nor UO_3748 (O_3748,N_48158,N_48761);
nor UO_3749 (O_3749,N_47505,N_49846);
nor UO_3750 (O_3750,N_48999,N_48345);
nand UO_3751 (O_3751,N_48457,N_48283);
nand UO_3752 (O_3752,N_48925,N_49734);
and UO_3753 (O_3753,N_48288,N_49985);
nand UO_3754 (O_3754,N_49478,N_49320);
xnor UO_3755 (O_3755,N_48327,N_47854);
nand UO_3756 (O_3756,N_48263,N_48332);
nand UO_3757 (O_3757,N_49477,N_48179);
and UO_3758 (O_3758,N_49802,N_49830);
or UO_3759 (O_3759,N_48317,N_48500);
and UO_3760 (O_3760,N_49542,N_48033);
or UO_3761 (O_3761,N_48004,N_49233);
and UO_3762 (O_3762,N_47997,N_48060);
nor UO_3763 (O_3763,N_48362,N_49979);
nor UO_3764 (O_3764,N_47841,N_48166);
xor UO_3765 (O_3765,N_48237,N_49217);
and UO_3766 (O_3766,N_48261,N_49196);
or UO_3767 (O_3767,N_48381,N_49758);
and UO_3768 (O_3768,N_47500,N_48314);
or UO_3769 (O_3769,N_48115,N_49430);
and UO_3770 (O_3770,N_49799,N_48862);
xor UO_3771 (O_3771,N_49699,N_47853);
xor UO_3772 (O_3772,N_49164,N_49677);
xor UO_3773 (O_3773,N_48088,N_48863);
nand UO_3774 (O_3774,N_49362,N_48336);
nor UO_3775 (O_3775,N_48239,N_48188);
nand UO_3776 (O_3776,N_49782,N_48706);
nor UO_3777 (O_3777,N_47745,N_48586);
or UO_3778 (O_3778,N_47879,N_48580);
and UO_3779 (O_3779,N_48403,N_48894);
xor UO_3780 (O_3780,N_48824,N_49847);
or UO_3781 (O_3781,N_49191,N_48936);
nor UO_3782 (O_3782,N_47790,N_47514);
or UO_3783 (O_3783,N_49847,N_48020);
and UO_3784 (O_3784,N_48497,N_48384);
xor UO_3785 (O_3785,N_48857,N_47518);
and UO_3786 (O_3786,N_49082,N_49138);
nand UO_3787 (O_3787,N_49806,N_48113);
xor UO_3788 (O_3788,N_49041,N_49721);
nand UO_3789 (O_3789,N_48281,N_49496);
xor UO_3790 (O_3790,N_47806,N_48258);
nand UO_3791 (O_3791,N_47945,N_47867);
nor UO_3792 (O_3792,N_47755,N_47772);
nand UO_3793 (O_3793,N_48436,N_47866);
nand UO_3794 (O_3794,N_48414,N_49760);
or UO_3795 (O_3795,N_48195,N_49843);
xor UO_3796 (O_3796,N_49432,N_49251);
and UO_3797 (O_3797,N_49324,N_48891);
and UO_3798 (O_3798,N_49241,N_48258);
and UO_3799 (O_3799,N_49065,N_49995);
nor UO_3800 (O_3800,N_49352,N_48539);
nor UO_3801 (O_3801,N_48393,N_49822);
nor UO_3802 (O_3802,N_47651,N_49397);
nor UO_3803 (O_3803,N_47547,N_48701);
and UO_3804 (O_3804,N_47865,N_47565);
or UO_3805 (O_3805,N_47570,N_49817);
xnor UO_3806 (O_3806,N_48410,N_48235);
xnor UO_3807 (O_3807,N_47657,N_48957);
nor UO_3808 (O_3808,N_49861,N_47565);
or UO_3809 (O_3809,N_49692,N_47578);
nor UO_3810 (O_3810,N_49041,N_49987);
xor UO_3811 (O_3811,N_48453,N_48983);
or UO_3812 (O_3812,N_47992,N_47707);
nand UO_3813 (O_3813,N_48004,N_49121);
nand UO_3814 (O_3814,N_47876,N_47631);
and UO_3815 (O_3815,N_48131,N_49602);
or UO_3816 (O_3816,N_48156,N_48698);
and UO_3817 (O_3817,N_48012,N_48579);
or UO_3818 (O_3818,N_49319,N_47955);
or UO_3819 (O_3819,N_48513,N_47800);
nor UO_3820 (O_3820,N_48468,N_49821);
or UO_3821 (O_3821,N_47993,N_48998);
nor UO_3822 (O_3822,N_48034,N_48444);
nor UO_3823 (O_3823,N_48283,N_49552);
nor UO_3824 (O_3824,N_48044,N_47917);
and UO_3825 (O_3825,N_49497,N_47921);
xor UO_3826 (O_3826,N_49144,N_48444);
and UO_3827 (O_3827,N_48403,N_49352);
xor UO_3828 (O_3828,N_49145,N_47626);
xor UO_3829 (O_3829,N_49960,N_48370);
nand UO_3830 (O_3830,N_49696,N_47681);
nand UO_3831 (O_3831,N_49473,N_49248);
and UO_3832 (O_3832,N_47676,N_49418);
xnor UO_3833 (O_3833,N_48156,N_47583);
nand UO_3834 (O_3834,N_49365,N_49005);
or UO_3835 (O_3835,N_49630,N_48231);
or UO_3836 (O_3836,N_49653,N_47723);
and UO_3837 (O_3837,N_49328,N_48835);
nand UO_3838 (O_3838,N_48035,N_49153);
xnor UO_3839 (O_3839,N_49004,N_49980);
and UO_3840 (O_3840,N_48037,N_49980);
and UO_3841 (O_3841,N_48443,N_49874);
or UO_3842 (O_3842,N_48898,N_48890);
xor UO_3843 (O_3843,N_49269,N_47968);
and UO_3844 (O_3844,N_48837,N_49470);
nor UO_3845 (O_3845,N_48053,N_47939);
xor UO_3846 (O_3846,N_49405,N_48768);
nand UO_3847 (O_3847,N_48708,N_48402);
nor UO_3848 (O_3848,N_48984,N_47594);
xnor UO_3849 (O_3849,N_48957,N_49120);
or UO_3850 (O_3850,N_48520,N_49905);
xor UO_3851 (O_3851,N_47530,N_47549);
and UO_3852 (O_3852,N_49985,N_48151);
nor UO_3853 (O_3853,N_48535,N_49324);
or UO_3854 (O_3854,N_48641,N_49747);
xor UO_3855 (O_3855,N_48578,N_48126);
and UO_3856 (O_3856,N_48552,N_49740);
and UO_3857 (O_3857,N_48842,N_49150);
nand UO_3858 (O_3858,N_48220,N_49047);
xor UO_3859 (O_3859,N_47936,N_47846);
nand UO_3860 (O_3860,N_49574,N_47964);
xor UO_3861 (O_3861,N_48554,N_48466);
and UO_3862 (O_3862,N_49138,N_48295);
or UO_3863 (O_3863,N_49300,N_48230);
xnor UO_3864 (O_3864,N_48650,N_48206);
nand UO_3865 (O_3865,N_48564,N_47802);
and UO_3866 (O_3866,N_47706,N_48920);
and UO_3867 (O_3867,N_49372,N_48645);
nor UO_3868 (O_3868,N_48491,N_48410);
xnor UO_3869 (O_3869,N_47899,N_48943);
xnor UO_3870 (O_3870,N_47540,N_49251);
or UO_3871 (O_3871,N_47835,N_48694);
nand UO_3872 (O_3872,N_48083,N_49926);
or UO_3873 (O_3873,N_49251,N_48105);
or UO_3874 (O_3874,N_49529,N_47916);
xnor UO_3875 (O_3875,N_49697,N_48799);
or UO_3876 (O_3876,N_49111,N_47513);
or UO_3877 (O_3877,N_48123,N_48763);
or UO_3878 (O_3878,N_49672,N_48020);
nor UO_3879 (O_3879,N_49960,N_49934);
xnor UO_3880 (O_3880,N_49268,N_48640);
and UO_3881 (O_3881,N_48911,N_48842);
nand UO_3882 (O_3882,N_48290,N_47812);
and UO_3883 (O_3883,N_48541,N_48244);
xor UO_3884 (O_3884,N_47933,N_49839);
and UO_3885 (O_3885,N_49314,N_48575);
or UO_3886 (O_3886,N_49351,N_47916);
nand UO_3887 (O_3887,N_48329,N_48093);
xor UO_3888 (O_3888,N_49176,N_47801);
nand UO_3889 (O_3889,N_49012,N_48652);
nor UO_3890 (O_3890,N_49045,N_49722);
and UO_3891 (O_3891,N_48434,N_47538);
xnor UO_3892 (O_3892,N_49150,N_47796);
or UO_3893 (O_3893,N_49103,N_48384);
xor UO_3894 (O_3894,N_49799,N_49220);
and UO_3895 (O_3895,N_48194,N_47637);
or UO_3896 (O_3896,N_48266,N_49536);
or UO_3897 (O_3897,N_49127,N_48677);
or UO_3898 (O_3898,N_47587,N_47927);
xnor UO_3899 (O_3899,N_49516,N_49163);
or UO_3900 (O_3900,N_48849,N_49854);
xor UO_3901 (O_3901,N_47939,N_48406);
and UO_3902 (O_3902,N_47884,N_48610);
nand UO_3903 (O_3903,N_49916,N_48214);
or UO_3904 (O_3904,N_49542,N_48977);
nor UO_3905 (O_3905,N_49059,N_49333);
and UO_3906 (O_3906,N_49942,N_49035);
nand UO_3907 (O_3907,N_47856,N_49193);
nor UO_3908 (O_3908,N_48033,N_47686);
or UO_3909 (O_3909,N_47617,N_49917);
or UO_3910 (O_3910,N_49040,N_49861);
xnor UO_3911 (O_3911,N_49760,N_48248);
nor UO_3912 (O_3912,N_48129,N_48251);
xnor UO_3913 (O_3913,N_48346,N_49497);
and UO_3914 (O_3914,N_49028,N_49171);
nand UO_3915 (O_3915,N_49119,N_49683);
or UO_3916 (O_3916,N_49100,N_47607);
xnor UO_3917 (O_3917,N_49619,N_48661);
xor UO_3918 (O_3918,N_48295,N_49394);
and UO_3919 (O_3919,N_49299,N_47970);
or UO_3920 (O_3920,N_49391,N_49894);
nor UO_3921 (O_3921,N_48325,N_49957);
and UO_3922 (O_3922,N_49349,N_49363);
nor UO_3923 (O_3923,N_47881,N_47804);
nor UO_3924 (O_3924,N_48750,N_48569);
xnor UO_3925 (O_3925,N_48190,N_48183);
or UO_3926 (O_3926,N_47527,N_48905);
nand UO_3927 (O_3927,N_49340,N_48694);
or UO_3928 (O_3928,N_48637,N_49533);
or UO_3929 (O_3929,N_49733,N_48491);
or UO_3930 (O_3930,N_49481,N_48366);
xnor UO_3931 (O_3931,N_49743,N_49519);
xor UO_3932 (O_3932,N_49154,N_49211);
nand UO_3933 (O_3933,N_48891,N_48024);
nor UO_3934 (O_3934,N_49319,N_49860);
nor UO_3935 (O_3935,N_48186,N_47695);
nand UO_3936 (O_3936,N_48281,N_48342);
nor UO_3937 (O_3937,N_47580,N_49920);
xnor UO_3938 (O_3938,N_47517,N_48046);
nor UO_3939 (O_3939,N_49027,N_48507);
or UO_3940 (O_3940,N_48673,N_48333);
xnor UO_3941 (O_3941,N_49306,N_49152);
or UO_3942 (O_3942,N_47966,N_48012);
xnor UO_3943 (O_3943,N_49290,N_48777);
nand UO_3944 (O_3944,N_47577,N_49598);
or UO_3945 (O_3945,N_47504,N_47848);
nor UO_3946 (O_3946,N_49488,N_47941);
xor UO_3947 (O_3947,N_49320,N_47995);
and UO_3948 (O_3948,N_49614,N_48658);
or UO_3949 (O_3949,N_47502,N_49249);
or UO_3950 (O_3950,N_49592,N_48196);
or UO_3951 (O_3951,N_49653,N_48731);
or UO_3952 (O_3952,N_49904,N_49059);
and UO_3953 (O_3953,N_49917,N_48429);
nand UO_3954 (O_3954,N_49932,N_48101);
nor UO_3955 (O_3955,N_49755,N_47928);
or UO_3956 (O_3956,N_49196,N_48785);
and UO_3957 (O_3957,N_49402,N_48734);
or UO_3958 (O_3958,N_48443,N_49460);
and UO_3959 (O_3959,N_49411,N_49481);
and UO_3960 (O_3960,N_48234,N_47535);
or UO_3961 (O_3961,N_48997,N_49007);
or UO_3962 (O_3962,N_48788,N_49970);
nor UO_3963 (O_3963,N_48228,N_49037);
xor UO_3964 (O_3964,N_48519,N_49065);
or UO_3965 (O_3965,N_49590,N_49653);
and UO_3966 (O_3966,N_49685,N_48072);
xor UO_3967 (O_3967,N_47663,N_48732);
xnor UO_3968 (O_3968,N_48718,N_49702);
nand UO_3969 (O_3969,N_48578,N_49027);
nor UO_3970 (O_3970,N_49238,N_49934);
or UO_3971 (O_3971,N_49784,N_48667);
xor UO_3972 (O_3972,N_47825,N_48416);
or UO_3973 (O_3973,N_49250,N_48062);
nand UO_3974 (O_3974,N_48043,N_49698);
or UO_3975 (O_3975,N_49200,N_49893);
xor UO_3976 (O_3976,N_49448,N_49351);
nand UO_3977 (O_3977,N_48910,N_47580);
xnor UO_3978 (O_3978,N_47543,N_49238);
nand UO_3979 (O_3979,N_48626,N_48379);
and UO_3980 (O_3980,N_48393,N_48140);
and UO_3981 (O_3981,N_48439,N_49931);
xor UO_3982 (O_3982,N_48863,N_47999);
or UO_3983 (O_3983,N_48536,N_49979);
xnor UO_3984 (O_3984,N_49154,N_47865);
xnor UO_3985 (O_3985,N_49112,N_49363);
nor UO_3986 (O_3986,N_48821,N_48156);
nor UO_3987 (O_3987,N_49970,N_49186);
nand UO_3988 (O_3988,N_48770,N_49608);
nor UO_3989 (O_3989,N_48442,N_48133);
nor UO_3990 (O_3990,N_49601,N_47951);
xor UO_3991 (O_3991,N_49071,N_49457);
and UO_3992 (O_3992,N_49100,N_48091);
xnor UO_3993 (O_3993,N_48360,N_47688);
and UO_3994 (O_3994,N_47520,N_47851);
and UO_3995 (O_3995,N_48714,N_48400);
nand UO_3996 (O_3996,N_47946,N_49047);
xor UO_3997 (O_3997,N_49751,N_48431);
or UO_3998 (O_3998,N_49190,N_49132);
nor UO_3999 (O_3999,N_49982,N_49226);
xnor UO_4000 (O_4000,N_49738,N_49762);
xor UO_4001 (O_4001,N_47768,N_49313);
and UO_4002 (O_4002,N_48273,N_48734);
nor UO_4003 (O_4003,N_48002,N_49450);
and UO_4004 (O_4004,N_47631,N_47619);
and UO_4005 (O_4005,N_48984,N_48090);
nand UO_4006 (O_4006,N_49074,N_48191);
nand UO_4007 (O_4007,N_49662,N_49999);
or UO_4008 (O_4008,N_48083,N_49632);
nor UO_4009 (O_4009,N_48587,N_47622);
nor UO_4010 (O_4010,N_48109,N_48604);
and UO_4011 (O_4011,N_48625,N_48245);
and UO_4012 (O_4012,N_47843,N_48884);
xor UO_4013 (O_4013,N_49118,N_47580);
or UO_4014 (O_4014,N_48363,N_49894);
or UO_4015 (O_4015,N_48277,N_48740);
or UO_4016 (O_4016,N_49509,N_49262);
nor UO_4017 (O_4017,N_49901,N_47637);
xor UO_4018 (O_4018,N_49849,N_48510);
or UO_4019 (O_4019,N_48251,N_47557);
nor UO_4020 (O_4020,N_48411,N_48654);
nor UO_4021 (O_4021,N_49198,N_48752);
nor UO_4022 (O_4022,N_47919,N_49355);
xor UO_4023 (O_4023,N_49517,N_49725);
or UO_4024 (O_4024,N_49829,N_49281);
nand UO_4025 (O_4025,N_47652,N_49078);
nor UO_4026 (O_4026,N_49911,N_48141);
nand UO_4027 (O_4027,N_47616,N_49805);
nand UO_4028 (O_4028,N_49304,N_49826);
or UO_4029 (O_4029,N_48442,N_48196);
nand UO_4030 (O_4030,N_47857,N_49529);
nor UO_4031 (O_4031,N_49847,N_48982);
nor UO_4032 (O_4032,N_49872,N_49843);
nor UO_4033 (O_4033,N_47587,N_48960);
and UO_4034 (O_4034,N_47705,N_48273);
or UO_4035 (O_4035,N_49604,N_49480);
nand UO_4036 (O_4036,N_47933,N_49645);
nor UO_4037 (O_4037,N_47635,N_49858);
and UO_4038 (O_4038,N_48995,N_48696);
nor UO_4039 (O_4039,N_48915,N_47852);
or UO_4040 (O_4040,N_49439,N_47616);
or UO_4041 (O_4041,N_48591,N_49837);
and UO_4042 (O_4042,N_48584,N_49268);
and UO_4043 (O_4043,N_49385,N_48449);
xor UO_4044 (O_4044,N_48027,N_49322);
nand UO_4045 (O_4045,N_48899,N_48767);
or UO_4046 (O_4046,N_48970,N_48513);
nand UO_4047 (O_4047,N_48461,N_49727);
nor UO_4048 (O_4048,N_48914,N_49084);
nor UO_4049 (O_4049,N_49277,N_48565);
and UO_4050 (O_4050,N_49407,N_49626);
nand UO_4051 (O_4051,N_49764,N_48012);
nor UO_4052 (O_4052,N_48464,N_49794);
nand UO_4053 (O_4053,N_49159,N_47609);
nor UO_4054 (O_4054,N_49111,N_49835);
and UO_4055 (O_4055,N_48908,N_47593);
or UO_4056 (O_4056,N_48491,N_49696);
or UO_4057 (O_4057,N_48954,N_48631);
nand UO_4058 (O_4058,N_48164,N_47698);
nand UO_4059 (O_4059,N_48346,N_47943);
and UO_4060 (O_4060,N_49631,N_47877);
or UO_4061 (O_4061,N_49608,N_49666);
nor UO_4062 (O_4062,N_47582,N_49526);
or UO_4063 (O_4063,N_48339,N_48917);
xnor UO_4064 (O_4064,N_49995,N_48916);
nor UO_4065 (O_4065,N_49342,N_48166);
or UO_4066 (O_4066,N_48803,N_49047);
xnor UO_4067 (O_4067,N_48275,N_48992);
nor UO_4068 (O_4068,N_47917,N_48446);
nor UO_4069 (O_4069,N_48284,N_49718);
xor UO_4070 (O_4070,N_48622,N_49003);
or UO_4071 (O_4071,N_48740,N_48951);
nor UO_4072 (O_4072,N_49339,N_48170);
nor UO_4073 (O_4073,N_49273,N_47806);
xor UO_4074 (O_4074,N_48930,N_49965);
and UO_4075 (O_4075,N_49241,N_49795);
and UO_4076 (O_4076,N_49523,N_49576);
nor UO_4077 (O_4077,N_48787,N_48100);
nand UO_4078 (O_4078,N_47975,N_47872);
and UO_4079 (O_4079,N_49382,N_49069);
and UO_4080 (O_4080,N_48316,N_48029);
or UO_4081 (O_4081,N_47840,N_48929);
or UO_4082 (O_4082,N_48386,N_49703);
xnor UO_4083 (O_4083,N_49898,N_49663);
xnor UO_4084 (O_4084,N_49506,N_47541);
or UO_4085 (O_4085,N_48194,N_47909);
xor UO_4086 (O_4086,N_49727,N_47827);
nand UO_4087 (O_4087,N_48288,N_49790);
nor UO_4088 (O_4088,N_49320,N_48299);
xor UO_4089 (O_4089,N_48742,N_48470);
or UO_4090 (O_4090,N_48339,N_49361);
and UO_4091 (O_4091,N_48458,N_48201);
or UO_4092 (O_4092,N_49042,N_48587);
nand UO_4093 (O_4093,N_49618,N_48966);
and UO_4094 (O_4094,N_48524,N_48862);
nor UO_4095 (O_4095,N_49290,N_49194);
nand UO_4096 (O_4096,N_47636,N_48461);
nor UO_4097 (O_4097,N_48695,N_48379);
or UO_4098 (O_4098,N_49119,N_48111);
or UO_4099 (O_4099,N_49502,N_47996);
xor UO_4100 (O_4100,N_48481,N_48542);
nor UO_4101 (O_4101,N_47699,N_49691);
and UO_4102 (O_4102,N_48416,N_49945);
nor UO_4103 (O_4103,N_49291,N_49079);
nand UO_4104 (O_4104,N_48771,N_47755);
nand UO_4105 (O_4105,N_49453,N_47630);
or UO_4106 (O_4106,N_49241,N_49097);
nor UO_4107 (O_4107,N_47505,N_48003);
and UO_4108 (O_4108,N_48402,N_49749);
nor UO_4109 (O_4109,N_49763,N_48982);
nand UO_4110 (O_4110,N_48929,N_48442);
or UO_4111 (O_4111,N_49831,N_48631);
and UO_4112 (O_4112,N_48403,N_48842);
nor UO_4113 (O_4113,N_49410,N_49910);
nor UO_4114 (O_4114,N_48162,N_47552);
xnor UO_4115 (O_4115,N_49891,N_47518);
and UO_4116 (O_4116,N_49503,N_48674);
or UO_4117 (O_4117,N_49156,N_47694);
or UO_4118 (O_4118,N_48790,N_48153);
or UO_4119 (O_4119,N_48565,N_48582);
nor UO_4120 (O_4120,N_49451,N_49135);
nand UO_4121 (O_4121,N_48098,N_49922);
nand UO_4122 (O_4122,N_49457,N_48835);
nand UO_4123 (O_4123,N_48835,N_49848);
and UO_4124 (O_4124,N_48417,N_48760);
and UO_4125 (O_4125,N_48252,N_49185);
xor UO_4126 (O_4126,N_48386,N_48986);
nand UO_4127 (O_4127,N_48887,N_49299);
xnor UO_4128 (O_4128,N_47822,N_48672);
or UO_4129 (O_4129,N_47789,N_48001);
xnor UO_4130 (O_4130,N_49305,N_47763);
nor UO_4131 (O_4131,N_47724,N_49536);
and UO_4132 (O_4132,N_48490,N_47651);
or UO_4133 (O_4133,N_48058,N_49945);
nor UO_4134 (O_4134,N_47797,N_49332);
nand UO_4135 (O_4135,N_48629,N_48789);
xnor UO_4136 (O_4136,N_49009,N_48769);
and UO_4137 (O_4137,N_49303,N_49602);
nand UO_4138 (O_4138,N_49152,N_47603);
and UO_4139 (O_4139,N_48516,N_48338);
xnor UO_4140 (O_4140,N_47895,N_49926);
nor UO_4141 (O_4141,N_47627,N_49314);
and UO_4142 (O_4142,N_48452,N_48722);
nor UO_4143 (O_4143,N_48238,N_48414);
xnor UO_4144 (O_4144,N_49774,N_47850);
and UO_4145 (O_4145,N_48821,N_47574);
nor UO_4146 (O_4146,N_47513,N_49738);
xnor UO_4147 (O_4147,N_49064,N_48318);
or UO_4148 (O_4148,N_48718,N_47597);
or UO_4149 (O_4149,N_47635,N_48530);
and UO_4150 (O_4150,N_48646,N_48320);
nor UO_4151 (O_4151,N_48948,N_47842);
xnor UO_4152 (O_4152,N_48962,N_48303);
or UO_4153 (O_4153,N_47550,N_49064);
xnor UO_4154 (O_4154,N_49879,N_49258);
xor UO_4155 (O_4155,N_49214,N_48814);
xor UO_4156 (O_4156,N_48409,N_48707);
nand UO_4157 (O_4157,N_48205,N_48432);
nand UO_4158 (O_4158,N_48408,N_49615);
nor UO_4159 (O_4159,N_49300,N_48201);
and UO_4160 (O_4160,N_47981,N_49622);
xor UO_4161 (O_4161,N_48412,N_48042);
xnor UO_4162 (O_4162,N_48297,N_47582);
nor UO_4163 (O_4163,N_49974,N_47630);
or UO_4164 (O_4164,N_47856,N_48345);
nand UO_4165 (O_4165,N_49381,N_47993);
and UO_4166 (O_4166,N_48051,N_49170);
or UO_4167 (O_4167,N_49363,N_47727);
nor UO_4168 (O_4168,N_48175,N_49663);
nand UO_4169 (O_4169,N_48189,N_49586);
and UO_4170 (O_4170,N_48426,N_49742);
xnor UO_4171 (O_4171,N_48329,N_49510);
or UO_4172 (O_4172,N_49908,N_47617);
xnor UO_4173 (O_4173,N_47944,N_49399);
xor UO_4174 (O_4174,N_47811,N_47799);
nor UO_4175 (O_4175,N_47553,N_49664);
nand UO_4176 (O_4176,N_49103,N_49466);
and UO_4177 (O_4177,N_48035,N_48121);
and UO_4178 (O_4178,N_49759,N_48414);
or UO_4179 (O_4179,N_48555,N_49508);
nor UO_4180 (O_4180,N_49665,N_48832);
or UO_4181 (O_4181,N_49926,N_48946);
or UO_4182 (O_4182,N_47613,N_49363);
or UO_4183 (O_4183,N_49960,N_47803);
and UO_4184 (O_4184,N_49962,N_49762);
or UO_4185 (O_4185,N_47704,N_48967);
nand UO_4186 (O_4186,N_49822,N_48337);
nor UO_4187 (O_4187,N_49375,N_47798);
nor UO_4188 (O_4188,N_49687,N_48027);
xor UO_4189 (O_4189,N_49816,N_49530);
nor UO_4190 (O_4190,N_47991,N_47751);
or UO_4191 (O_4191,N_48141,N_47520);
nand UO_4192 (O_4192,N_49330,N_47577);
and UO_4193 (O_4193,N_49225,N_49567);
or UO_4194 (O_4194,N_49285,N_47768);
xnor UO_4195 (O_4195,N_48850,N_47948);
nor UO_4196 (O_4196,N_48764,N_49764);
and UO_4197 (O_4197,N_47701,N_49301);
xnor UO_4198 (O_4198,N_47786,N_48969);
or UO_4199 (O_4199,N_47904,N_47587);
xnor UO_4200 (O_4200,N_47614,N_48564);
xor UO_4201 (O_4201,N_49384,N_47590);
nor UO_4202 (O_4202,N_47903,N_49621);
nor UO_4203 (O_4203,N_49990,N_48096);
or UO_4204 (O_4204,N_48111,N_48061);
nor UO_4205 (O_4205,N_48213,N_48106);
nand UO_4206 (O_4206,N_47958,N_48442);
or UO_4207 (O_4207,N_48010,N_49208);
nor UO_4208 (O_4208,N_48144,N_49239);
xor UO_4209 (O_4209,N_48820,N_49388);
xnor UO_4210 (O_4210,N_48928,N_49600);
nand UO_4211 (O_4211,N_47975,N_49158);
xnor UO_4212 (O_4212,N_48215,N_49970);
and UO_4213 (O_4213,N_49588,N_47854);
nand UO_4214 (O_4214,N_47770,N_48816);
xnor UO_4215 (O_4215,N_47741,N_49669);
nand UO_4216 (O_4216,N_48344,N_48014);
xnor UO_4217 (O_4217,N_49267,N_48403);
xnor UO_4218 (O_4218,N_49624,N_48742);
nand UO_4219 (O_4219,N_47607,N_49183);
nor UO_4220 (O_4220,N_49872,N_47581);
and UO_4221 (O_4221,N_47678,N_47824);
or UO_4222 (O_4222,N_49282,N_47649);
nor UO_4223 (O_4223,N_49478,N_49749);
nand UO_4224 (O_4224,N_49846,N_49441);
and UO_4225 (O_4225,N_48756,N_49324);
nor UO_4226 (O_4226,N_49306,N_49585);
nor UO_4227 (O_4227,N_49772,N_49509);
and UO_4228 (O_4228,N_49920,N_49586);
nand UO_4229 (O_4229,N_48987,N_48753);
nor UO_4230 (O_4230,N_48674,N_48188);
and UO_4231 (O_4231,N_48787,N_48723);
nand UO_4232 (O_4232,N_49954,N_49667);
nand UO_4233 (O_4233,N_47756,N_48436);
or UO_4234 (O_4234,N_48831,N_47608);
or UO_4235 (O_4235,N_49881,N_49954);
nand UO_4236 (O_4236,N_48221,N_49209);
or UO_4237 (O_4237,N_48929,N_48150);
and UO_4238 (O_4238,N_47694,N_47606);
nand UO_4239 (O_4239,N_48497,N_49371);
nand UO_4240 (O_4240,N_48102,N_49747);
and UO_4241 (O_4241,N_49394,N_49269);
and UO_4242 (O_4242,N_49277,N_49762);
nor UO_4243 (O_4243,N_49609,N_49604);
or UO_4244 (O_4244,N_49389,N_49092);
or UO_4245 (O_4245,N_49832,N_47567);
nand UO_4246 (O_4246,N_48124,N_48423);
nor UO_4247 (O_4247,N_49005,N_49382);
nand UO_4248 (O_4248,N_47851,N_49979);
or UO_4249 (O_4249,N_48449,N_48557);
nand UO_4250 (O_4250,N_49492,N_49339);
xor UO_4251 (O_4251,N_49119,N_48497);
and UO_4252 (O_4252,N_47869,N_47925);
xnor UO_4253 (O_4253,N_47688,N_48747);
nor UO_4254 (O_4254,N_48907,N_47617);
and UO_4255 (O_4255,N_48484,N_47678);
and UO_4256 (O_4256,N_49893,N_47808);
nand UO_4257 (O_4257,N_48143,N_49647);
xor UO_4258 (O_4258,N_49771,N_48348);
nand UO_4259 (O_4259,N_49222,N_49135);
nor UO_4260 (O_4260,N_47632,N_49093);
nor UO_4261 (O_4261,N_48755,N_47651);
and UO_4262 (O_4262,N_49007,N_48474);
or UO_4263 (O_4263,N_49282,N_47909);
xor UO_4264 (O_4264,N_49306,N_47740);
and UO_4265 (O_4265,N_49011,N_47751);
nand UO_4266 (O_4266,N_48367,N_48864);
nand UO_4267 (O_4267,N_49653,N_48354);
and UO_4268 (O_4268,N_49942,N_49187);
or UO_4269 (O_4269,N_47625,N_49579);
nor UO_4270 (O_4270,N_49980,N_48829);
xnor UO_4271 (O_4271,N_49991,N_47729);
nand UO_4272 (O_4272,N_47674,N_47743);
nand UO_4273 (O_4273,N_49577,N_47524);
nand UO_4274 (O_4274,N_47550,N_48162);
and UO_4275 (O_4275,N_47748,N_48560);
xor UO_4276 (O_4276,N_49381,N_48429);
and UO_4277 (O_4277,N_48182,N_48371);
nand UO_4278 (O_4278,N_47610,N_49899);
xnor UO_4279 (O_4279,N_49046,N_47716);
or UO_4280 (O_4280,N_49513,N_48111);
nand UO_4281 (O_4281,N_47645,N_48716);
xor UO_4282 (O_4282,N_47975,N_49680);
or UO_4283 (O_4283,N_49239,N_49106);
xor UO_4284 (O_4284,N_48206,N_48979);
nor UO_4285 (O_4285,N_49171,N_48608);
and UO_4286 (O_4286,N_47699,N_47685);
nor UO_4287 (O_4287,N_47630,N_48432);
or UO_4288 (O_4288,N_49996,N_47627);
nand UO_4289 (O_4289,N_48107,N_48337);
nor UO_4290 (O_4290,N_48004,N_48065);
nand UO_4291 (O_4291,N_48566,N_49662);
nor UO_4292 (O_4292,N_48620,N_49622);
xnor UO_4293 (O_4293,N_48323,N_48723);
nand UO_4294 (O_4294,N_48771,N_49351);
or UO_4295 (O_4295,N_48128,N_49516);
xnor UO_4296 (O_4296,N_48937,N_49665);
xnor UO_4297 (O_4297,N_47738,N_47890);
nand UO_4298 (O_4298,N_49772,N_48244);
and UO_4299 (O_4299,N_48548,N_48206);
xnor UO_4300 (O_4300,N_49347,N_48340);
nand UO_4301 (O_4301,N_48672,N_48843);
or UO_4302 (O_4302,N_49951,N_48860);
and UO_4303 (O_4303,N_47554,N_48832);
and UO_4304 (O_4304,N_49812,N_48757);
nand UO_4305 (O_4305,N_49362,N_48416);
nor UO_4306 (O_4306,N_48207,N_49703);
or UO_4307 (O_4307,N_47655,N_49542);
xnor UO_4308 (O_4308,N_47861,N_49285);
nor UO_4309 (O_4309,N_47630,N_49876);
nor UO_4310 (O_4310,N_49919,N_49304);
nand UO_4311 (O_4311,N_49750,N_49568);
nand UO_4312 (O_4312,N_48610,N_47819);
or UO_4313 (O_4313,N_48070,N_47894);
xor UO_4314 (O_4314,N_49134,N_49422);
and UO_4315 (O_4315,N_49765,N_47982);
xnor UO_4316 (O_4316,N_48275,N_48395);
nor UO_4317 (O_4317,N_48863,N_48375);
and UO_4318 (O_4318,N_47653,N_48719);
xor UO_4319 (O_4319,N_47902,N_47586);
nand UO_4320 (O_4320,N_48657,N_47566);
xnor UO_4321 (O_4321,N_49961,N_47573);
nor UO_4322 (O_4322,N_49924,N_47954);
nand UO_4323 (O_4323,N_47838,N_48706);
and UO_4324 (O_4324,N_48776,N_48070);
xnor UO_4325 (O_4325,N_49322,N_48316);
or UO_4326 (O_4326,N_48519,N_48238);
nand UO_4327 (O_4327,N_48999,N_47665);
nand UO_4328 (O_4328,N_48786,N_49146);
nand UO_4329 (O_4329,N_48783,N_48342);
or UO_4330 (O_4330,N_48782,N_49945);
and UO_4331 (O_4331,N_48978,N_48886);
nor UO_4332 (O_4332,N_49572,N_49843);
nor UO_4333 (O_4333,N_49845,N_47951);
and UO_4334 (O_4334,N_49301,N_49629);
and UO_4335 (O_4335,N_49737,N_49656);
xor UO_4336 (O_4336,N_49890,N_48274);
or UO_4337 (O_4337,N_49030,N_47628);
nor UO_4338 (O_4338,N_48982,N_49648);
or UO_4339 (O_4339,N_47702,N_49608);
or UO_4340 (O_4340,N_47715,N_49107);
xnor UO_4341 (O_4341,N_48591,N_49305);
nor UO_4342 (O_4342,N_49284,N_47837);
nor UO_4343 (O_4343,N_48370,N_49679);
nand UO_4344 (O_4344,N_48877,N_48975);
nor UO_4345 (O_4345,N_48982,N_49857);
xnor UO_4346 (O_4346,N_48152,N_49040);
nand UO_4347 (O_4347,N_48660,N_48405);
nand UO_4348 (O_4348,N_48958,N_49878);
nand UO_4349 (O_4349,N_48925,N_49222);
or UO_4350 (O_4350,N_47727,N_48038);
xor UO_4351 (O_4351,N_48017,N_47624);
or UO_4352 (O_4352,N_49341,N_49195);
xnor UO_4353 (O_4353,N_48115,N_49580);
nor UO_4354 (O_4354,N_47957,N_48222);
or UO_4355 (O_4355,N_49266,N_47711);
or UO_4356 (O_4356,N_49339,N_48957);
nor UO_4357 (O_4357,N_48101,N_49069);
or UO_4358 (O_4358,N_47560,N_48427);
or UO_4359 (O_4359,N_48803,N_49326);
xor UO_4360 (O_4360,N_49495,N_49271);
nand UO_4361 (O_4361,N_48438,N_49396);
xnor UO_4362 (O_4362,N_49719,N_49627);
nor UO_4363 (O_4363,N_49803,N_49783);
nor UO_4364 (O_4364,N_48603,N_48234);
or UO_4365 (O_4365,N_48757,N_47668);
nand UO_4366 (O_4366,N_48778,N_49779);
or UO_4367 (O_4367,N_49986,N_48330);
or UO_4368 (O_4368,N_48018,N_47902);
and UO_4369 (O_4369,N_49828,N_48611);
or UO_4370 (O_4370,N_48110,N_49754);
or UO_4371 (O_4371,N_48422,N_49175);
nor UO_4372 (O_4372,N_47820,N_47577);
and UO_4373 (O_4373,N_47536,N_47620);
or UO_4374 (O_4374,N_48391,N_48588);
nor UO_4375 (O_4375,N_49252,N_48395);
and UO_4376 (O_4376,N_48331,N_49057);
nor UO_4377 (O_4377,N_48372,N_48819);
nand UO_4378 (O_4378,N_48490,N_48743);
nor UO_4379 (O_4379,N_48490,N_48822);
xnor UO_4380 (O_4380,N_48694,N_47588);
and UO_4381 (O_4381,N_49605,N_49641);
xor UO_4382 (O_4382,N_48523,N_47719);
or UO_4383 (O_4383,N_49424,N_47802);
nand UO_4384 (O_4384,N_49530,N_49329);
and UO_4385 (O_4385,N_48092,N_48219);
xor UO_4386 (O_4386,N_48508,N_48352);
xnor UO_4387 (O_4387,N_48089,N_49552);
xnor UO_4388 (O_4388,N_48465,N_47658);
xnor UO_4389 (O_4389,N_49115,N_49562);
nor UO_4390 (O_4390,N_49404,N_48037);
xor UO_4391 (O_4391,N_49141,N_48831);
or UO_4392 (O_4392,N_48120,N_48582);
nor UO_4393 (O_4393,N_48817,N_47749);
nor UO_4394 (O_4394,N_49384,N_47617);
xor UO_4395 (O_4395,N_48527,N_49015);
or UO_4396 (O_4396,N_47928,N_49812);
or UO_4397 (O_4397,N_49952,N_48358);
xnor UO_4398 (O_4398,N_48340,N_48738);
xor UO_4399 (O_4399,N_49019,N_47957);
nor UO_4400 (O_4400,N_47861,N_48222);
and UO_4401 (O_4401,N_49789,N_49732);
or UO_4402 (O_4402,N_48672,N_48287);
and UO_4403 (O_4403,N_49799,N_48103);
nor UO_4404 (O_4404,N_49942,N_49401);
or UO_4405 (O_4405,N_48211,N_48758);
and UO_4406 (O_4406,N_48912,N_48374);
nor UO_4407 (O_4407,N_48736,N_49951);
nand UO_4408 (O_4408,N_47805,N_48890);
nor UO_4409 (O_4409,N_47608,N_47500);
or UO_4410 (O_4410,N_48724,N_49774);
nand UO_4411 (O_4411,N_49752,N_49295);
and UO_4412 (O_4412,N_48624,N_49653);
nor UO_4413 (O_4413,N_48281,N_48622);
or UO_4414 (O_4414,N_47758,N_47549);
nand UO_4415 (O_4415,N_49558,N_48231);
nor UO_4416 (O_4416,N_48080,N_48045);
nor UO_4417 (O_4417,N_47603,N_48474);
xnor UO_4418 (O_4418,N_48176,N_49367);
nor UO_4419 (O_4419,N_49553,N_49421);
xor UO_4420 (O_4420,N_48717,N_49770);
xnor UO_4421 (O_4421,N_49290,N_48832);
nor UO_4422 (O_4422,N_49521,N_48152);
nor UO_4423 (O_4423,N_48558,N_47640);
nand UO_4424 (O_4424,N_48161,N_48919);
xnor UO_4425 (O_4425,N_48281,N_48242);
and UO_4426 (O_4426,N_47695,N_48571);
xor UO_4427 (O_4427,N_49828,N_49147);
nand UO_4428 (O_4428,N_47930,N_48116);
or UO_4429 (O_4429,N_49996,N_49424);
or UO_4430 (O_4430,N_49717,N_48322);
xor UO_4431 (O_4431,N_48271,N_47581);
xnor UO_4432 (O_4432,N_47949,N_48926);
nand UO_4433 (O_4433,N_49143,N_47854);
nor UO_4434 (O_4434,N_47784,N_48984);
xor UO_4435 (O_4435,N_47516,N_48970);
and UO_4436 (O_4436,N_47882,N_48861);
nor UO_4437 (O_4437,N_48154,N_49275);
nor UO_4438 (O_4438,N_48887,N_48694);
nand UO_4439 (O_4439,N_48913,N_49570);
xnor UO_4440 (O_4440,N_47567,N_49858);
or UO_4441 (O_4441,N_48093,N_49452);
nand UO_4442 (O_4442,N_49540,N_47649);
and UO_4443 (O_4443,N_48860,N_49827);
and UO_4444 (O_4444,N_48476,N_48899);
nand UO_4445 (O_4445,N_48331,N_47916);
nor UO_4446 (O_4446,N_47937,N_48851);
nand UO_4447 (O_4447,N_48796,N_48223);
nand UO_4448 (O_4448,N_47605,N_48765);
or UO_4449 (O_4449,N_48059,N_49287);
nor UO_4450 (O_4450,N_49130,N_48499);
nor UO_4451 (O_4451,N_47732,N_48175);
nor UO_4452 (O_4452,N_49002,N_49928);
xnor UO_4453 (O_4453,N_49478,N_49517);
nor UO_4454 (O_4454,N_48755,N_49861);
and UO_4455 (O_4455,N_48620,N_49910);
nand UO_4456 (O_4456,N_47542,N_47651);
nand UO_4457 (O_4457,N_48006,N_48159);
and UO_4458 (O_4458,N_47994,N_48898);
and UO_4459 (O_4459,N_49341,N_48250);
nand UO_4460 (O_4460,N_48488,N_47847);
xnor UO_4461 (O_4461,N_48362,N_47828);
and UO_4462 (O_4462,N_47902,N_48398);
and UO_4463 (O_4463,N_47628,N_49354);
and UO_4464 (O_4464,N_49960,N_48644);
xor UO_4465 (O_4465,N_49641,N_49299);
xor UO_4466 (O_4466,N_49290,N_49030);
and UO_4467 (O_4467,N_48652,N_48743);
or UO_4468 (O_4468,N_48210,N_49839);
xor UO_4469 (O_4469,N_49874,N_47701);
nor UO_4470 (O_4470,N_48518,N_49862);
nor UO_4471 (O_4471,N_49829,N_49351);
nor UO_4472 (O_4472,N_49321,N_48169);
or UO_4473 (O_4473,N_47578,N_48203);
and UO_4474 (O_4474,N_48752,N_48105);
nand UO_4475 (O_4475,N_49701,N_48195);
xnor UO_4476 (O_4476,N_48301,N_48072);
xor UO_4477 (O_4477,N_48144,N_48505);
xor UO_4478 (O_4478,N_47639,N_49904);
nand UO_4479 (O_4479,N_48883,N_49975);
and UO_4480 (O_4480,N_48812,N_47789);
and UO_4481 (O_4481,N_49565,N_49745);
nor UO_4482 (O_4482,N_49108,N_48649);
xnor UO_4483 (O_4483,N_47660,N_49939);
xor UO_4484 (O_4484,N_48275,N_48403);
nand UO_4485 (O_4485,N_48645,N_48658);
xor UO_4486 (O_4486,N_47782,N_49936);
nor UO_4487 (O_4487,N_48755,N_47602);
and UO_4488 (O_4488,N_47739,N_48758);
and UO_4489 (O_4489,N_48276,N_48478);
xor UO_4490 (O_4490,N_47955,N_47548);
nand UO_4491 (O_4491,N_48394,N_49598);
nor UO_4492 (O_4492,N_49940,N_49371);
and UO_4493 (O_4493,N_48897,N_49792);
or UO_4494 (O_4494,N_48317,N_47755);
nor UO_4495 (O_4495,N_49111,N_48279);
nor UO_4496 (O_4496,N_47768,N_48389);
or UO_4497 (O_4497,N_48111,N_48855);
and UO_4498 (O_4498,N_47569,N_49304);
and UO_4499 (O_4499,N_48879,N_49808);
nor UO_4500 (O_4500,N_49433,N_48217);
nand UO_4501 (O_4501,N_48303,N_48472);
nor UO_4502 (O_4502,N_47903,N_49595);
or UO_4503 (O_4503,N_47912,N_47619);
nor UO_4504 (O_4504,N_49939,N_49072);
xor UO_4505 (O_4505,N_48195,N_47545);
nand UO_4506 (O_4506,N_47913,N_49977);
or UO_4507 (O_4507,N_47990,N_49692);
or UO_4508 (O_4508,N_47610,N_48808);
nand UO_4509 (O_4509,N_48681,N_49666);
xor UO_4510 (O_4510,N_49679,N_49530);
or UO_4511 (O_4511,N_48638,N_48267);
and UO_4512 (O_4512,N_48227,N_47897);
nor UO_4513 (O_4513,N_48003,N_49936);
or UO_4514 (O_4514,N_48550,N_49608);
and UO_4515 (O_4515,N_47698,N_48592);
nor UO_4516 (O_4516,N_49708,N_47941);
or UO_4517 (O_4517,N_48746,N_49917);
nor UO_4518 (O_4518,N_48893,N_48714);
or UO_4519 (O_4519,N_49155,N_49172);
xor UO_4520 (O_4520,N_47755,N_49585);
nand UO_4521 (O_4521,N_48252,N_48044);
nand UO_4522 (O_4522,N_47594,N_49044);
nor UO_4523 (O_4523,N_48559,N_49760);
xor UO_4524 (O_4524,N_48854,N_49876);
xor UO_4525 (O_4525,N_48282,N_48632);
nor UO_4526 (O_4526,N_48862,N_49610);
nand UO_4527 (O_4527,N_49824,N_49140);
nor UO_4528 (O_4528,N_48068,N_49195);
xnor UO_4529 (O_4529,N_49512,N_47605);
nand UO_4530 (O_4530,N_47934,N_49908);
and UO_4531 (O_4531,N_47556,N_48122);
nor UO_4532 (O_4532,N_48085,N_48515);
xor UO_4533 (O_4533,N_49228,N_49599);
nor UO_4534 (O_4534,N_49992,N_49944);
and UO_4535 (O_4535,N_48048,N_48752);
xor UO_4536 (O_4536,N_49836,N_48263);
xnor UO_4537 (O_4537,N_49530,N_48470);
and UO_4538 (O_4538,N_48495,N_48777);
nand UO_4539 (O_4539,N_48266,N_49329);
or UO_4540 (O_4540,N_49264,N_49045);
nor UO_4541 (O_4541,N_48616,N_49700);
or UO_4542 (O_4542,N_48412,N_48223);
nand UO_4543 (O_4543,N_49579,N_48748);
nand UO_4544 (O_4544,N_49010,N_47827);
and UO_4545 (O_4545,N_48904,N_47918);
or UO_4546 (O_4546,N_47684,N_48642);
xnor UO_4547 (O_4547,N_49046,N_49164);
and UO_4548 (O_4548,N_49730,N_47789);
or UO_4549 (O_4549,N_49345,N_47982);
and UO_4550 (O_4550,N_48707,N_48032);
nand UO_4551 (O_4551,N_48404,N_48996);
nor UO_4552 (O_4552,N_48472,N_48261);
nor UO_4553 (O_4553,N_49872,N_49255);
xor UO_4554 (O_4554,N_48189,N_49490);
xor UO_4555 (O_4555,N_48185,N_48222);
xnor UO_4556 (O_4556,N_49553,N_49623);
nor UO_4557 (O_4557,N_49815,N_49045);
nand UO_4558 (O_4558,N_48153,N_47642);
nand UO_4559 (O_4559,N_49901,N_48766);
and UO_4560 (O_4560,N_49798,N_47665);
or UO_4561 (O_4561,N_49095,N_48802);
or UO_4562 (O_4562,N_49304,N_49374);
xnor UO_4563 (O_4563,N_49802,N_49040);
nand UO_4564 (O_4564,N_49866,N_49935);
nor UO_4565 (O_4565,N_48747,N_48777);
or UO_4566 (O_4566,N_49254,N_48205);
and UO_4567 (O_4567,N_48237,N_48670);
nand UO_4568 (O_4568,N_48435,N_49323);
and UO_4569 (O_4569,N_48835,N_49379);
and UO_4570 (O_4570,N_48834,N_47771);
or UO_4571 (O_4571,N_47878,N_48981);
and UO_4572 (O_4572,N_49967,N_49527);
or UO_4573 (O_4573,N_48284,N_48329);
and UO_4574 (O_4574,N_49801,N_48842);
xor UO_4575 (O_4575,N_48442,N_48345);
xnor UO_4576 (O_4576,N_49034,N_47657);
and UO_4577 (O_4577,N_48049,N_48200);
or UO_4578 (O_4578,N_47754,N_47983);
or UO_4579 (O_4579,N_48771,N_49111);
nor UO_4580 (O_4580,N_49034,N_49127);
and UO_4581 (O_4581,N_49011,N_49454);
xnor UO_4582 (O_4582,N_49815,N_49226);
nor UO_4583 (O_4583,N_48847,N_49893);
xor UO_4584 (O_4584,N_49658,N_47847);
and UO_4585 (O_4585,N_47633,N_48396);
or UO_4586 (O_4586,N_49783,N_48672);
or UO_4587 (O_4587,N_48934,N_49917);
xnor UO_4588 (O_4588,N_48501,N_48446);
and UO_4589 (O_4589,N_48875,N_49147);
and UO_4590 (O_4590,N_48971,N_48710);
xnor UO_4591 (O_4591,N_49016,N_48779);
or UO_4592 (O_4592,N_49393,N_48975);
nor UO_4593 (O_4593,N_49449,N_49406);
and UO_4594 (O_4594,N_48905,N_49384);
and UO_4595 (O_4595,N_49057,N_49224);
and UO_4596 (O_4596,N_48900,N_48865);
xor UO_4597 (O_4597,N_49147,N_48654);
or UO_4598 (O_4598,N_47605,N_49230);
and UO_4599 (O_4599,N_48375,N_48188);
xnor UO_4600 (O_4600,N_49618,N_47675);
nor UO_4601 (O_4601,N_47803,N_48211);
and UO_4602 (O_4602,N_48535,N_49922);
or UO_4603 (O_4603,N_48755,N_48191);
or UO_4604 (O_4604,N_49852,N_47595);
or UO_4605 (O_4605,N_48829,N_49121);
or UO_4606 (O_4606,N_49410,N_48615);
nand UO_4607 (O_4607,N_49208,N_49025);
nor UO_4608 (O_4608,N_48998,N_49707);
nand UO_4609 (O_4609,N_48856,N_49508);
or UO_4610 (O_4610,N_49989,N_49572);
nand UO_4611 (O_4611,N_48823,N_47535);
nor UO_4612 (O_4612,N_49797,N_48119);
or UO_4613 (O_4613,N_49608,N_49891);
and UO_4614 (O_4614,N_48821,N_49101);
nor UO_4615 (O_4615,N_49031,N_48993);
xor UO_4616 (O_4616,N_48249,N_49271);
xor UO_4617 (O_4617,N_48703,N_48330);
xor UO_4618 (O_4618,N_48932,N_48039);
nor UO_4619 (O_4619,N_49731,N_47757);
nor UO_4620 (O_4620,N_47813,N_47658);
and UO_4621 (O_4621,N_49466,N_49559);
or UO_4622 (O_4622,N_48060,N_48274);
and UO_4623 (O_4623,N_47860,N_48657);
xor UO_4624 (O_4624,N_48451,N_49841);
xor UO_4625 (O_4625,N_49565,N_49234);
or UO_4626 (O_4626,N_49464,N_48927);
xnor UO_4627 (O_4627,N_48789,N_47848);
and UO_4628 (O_4628,N_49445,N_48127);
xnor UO_4629 (O_4629,N_49926,N_48553);
or UO_4630 (O_4630,N_49143,N_48227);
xnor UO_4631 (O_4631,N_49518,N_47531);
nor UO_4632 (O_4632,N_47691,N_49590);
xnor UO_4633 (O_4633,N_49881,N_49598);
or UO_4634 (O_4634,N_48010,N_49879);
xor UO_4635 (O_4635,N_49026,N_47787);
or UO_4636 (O_4636,N_48324,N_48753);
nand UO_4637 (O_4637,N_48659,N_49321);
and UO_4638 (O_4638,N_47768,N_48614);
or UO_4639 (O_4639,N_48541,N_49662);
and UO_4640 (O_4640,N_47886,N_47977);
nand UO_4641 (O_4641,N_48209,N_47528);
and UO_4642 (O_4642,N_49553,N_47593);
or UO_4643 (O_4643,N_48247,N_48230);
xnor UO_4644 (O_4644,N_48955,N_47736);
nand UO_4645 (O_4645,N_49423,N_49611);
nand UO_4646 (O_4646,N_49462,N_49465);
and UO_4647 (O_4647,N_48742,N_48069);
nand UO_4648 (O_4648,N_48125,N_48344);
or UO_4649 (O_4649,N_49462,N_48644);
and UO_4650 (O_4650,N_48130,N_48390);
or UO_4651 (O_4651,N_49515,N_48938);
or UO_4652 (O_4652,N_47670,N_48488);
xnor UO_4653 (O_4653,N_48941,N_49889);
nand UO_4654 (O_4654,N_49156,N_48274);
nand UO_4655 (O_4655,N_49856,N_49199);
xnor UO_4656 (O_4656,N_49759,N_47691);
or UO_4657 (O_4657,N_49033,N_47731);
and UO_4658 (O_4658,N_49862,N_47617);
nor UO_4659 (O_4659,N_47537,N_48558);
or UO_4660 (O_4660,N_49415,N_48525);
xnor UO_4661 (O_4661,N_48191,N_49020);
nor UO_4662 (O_4662,N_47557,N_48288);
nor UO_4663 (O_4663,N_47963,N_48980);
or UO_4664 (O_4664,N_48155,N_47840);
nor UO_4665 (O_4665,N_48631,N_49140);
or UO_4666 (O_4666,N_48053,N_47959);
xor UO_4667 (O_4667,N_49560,N_47954);
xor UO_4668 (O_4668,N_49375,N_49122);
nand UO_4669 (O_4669,N_49791,N_48600);
nor UO_4670 (O_4670,N_47707,N_47615);
nor UO_4671 (O_4671,N_49161,N_49239);
xnor UO_4672 (O_4672,N_49401,N_49563);
xnor UO_4673 (O_4673,N_49640,N_49878);
xor UO_4674 (O_4674,N_49092,N_49274);
nand UO_4675 (O_4675,N_47800,N_49885);
nand UO_4676 (O_4676,N_48528,N_49716);
nor UO_4677 (O_4677,N_48219,N_47664);
or UO_4678 (O_4678,N_48058,N_49166);
and UO_4679 (O_4679,N_49587,N_47700);
nand UO_4680 (O_4680,N_48064,N_47688);
nor UO_4681 (O_4681,N_49702,N_49708);
and UO_4682 (O_4682,N_48211,N_47575);
nand UO_4683 (O_4683,N_49886,N_49548);
nand UO_4684 (O_4684,N_47561,N_48540);
nor UO_4685 (O_4685,N_49570,N_49778);
and UO_4686 (O_4686,N_48089,N_48736);
nand UO_4687 (O_4687,N_47794,N_48333);
xnor UO_4688 (O_4688,N_49207,N_47757);
or UO_4689 (O_4689,N_48700,N_48770);
nand UO_4690 (O_4690,N_48631,N_49639);
or UO_4691 (O_4691,N_47547,N_47695);
and UO_4692 (O_4692,N_49044,N_49831);
xnor UO_4693 (O_4693,N_48569,N_48598);
nand UO_4694 (O_4694,N_47793,N_48886);
xnor UO_4695 (O_4695,N_47785,N_49643);
nand UO_4696 (O_4696,N_47876,N_49615);
or UO_4697 (O_4697,N_49045,N_47996);
and UO_4698 (O_4698,N_47984,N_49362);
and UO_4699 (O_4699,N_48473,N_47614);
and UO_4700 (O_4700,N_49794,N_47718);
nand UO_4701 (O_4701,N_48710,N_49299);
or UO_4702 (O_4702,N_49967,N_49155);
or UO_4703 (O_4703,N_49537,N_48779);
nor UO_4704 (O_4704,N_47921,N_48055);
xor UO_4705 (O_4705,N_49913,N_48069);
nand UO_4706 (O_4706,N_48900,N_48724);
xor UO_4707 (O_4707,N_49599,N_49363);
xnor UO_4708 (O_4708,N_48272,N_49363);
and UO_4709 (O_4709,N_49229,N_47561);
xnor UO_4710 (O_4710,N_48129,N_48525);
or UO_4711 (O_4711,N_48882,N_49741);
nor UO_4712 (O_4712,N_49324,N_47591);
nand UO_4713 (O_4713,N_48676,N_47588);
nor UO_4714 (O_4714,N_49905,N_49928);
or UO_4715 (O_4715,N_48304,N_47699);
or UO_4716 (O_4716,N_48772,N_49945);
nor UO_4717 (O_4717,N_49004,N_47655);
xnor UO_4718 (O_4718,N_49004,N_48061);
and UO_4719 (O_4719,N_49274,N_47665);
or UO_4720 (O_4720,N_47514,N_49880);
nand UO_4721 (O_4721,N_48305,N_49655);
and UO_4722 (O_4722,N_48181,N_47942);
or UO_4723 (O_4723,N_48852,N_48534);
and UO_4724 (O_4724,N_47674,N_49656);
or UO_4725 (O_4725,N_49325,N_48204);
nor UO_4726 (O_4726,N_47982,N_48946);
nand UO_4727 (O_4727,N_48211,N_48728);
or UO_4728 (O_4728,N_49205,N_48481);
or UO_4729 (O_4729,N_48349,N_47718);
and UO_4730 (O_4730,N_49698,N_48100);
xor UO_4731 (O_4731,N_48091,N_49668);
nand UO_4732 (O_4732,N_48369,N_48288);
and UO_4733 (O_4733,N_49928,N_49848);
nor UO_4734 (O_4734,N_49426,N_48097);
and UO_4735 (O_4735,N_49621,N_48384);
or UO_4736 (O_4736,N_47636,N_47694);
nand UO_4737 (O_4737,N_48778,N_49379);
nor UO_4738 (O_4738,N_49821,N_48912);
nor UO_4739 (O_4739,N_49913,N_49909);
or UO_4740 (O_4740,N_49510,N_49639);
or UO_4741 (O_4741,N_49888,N_48626);
nor UO_4742 (O_4742,N_49638,N_49677);
nor UO_4743 (O_4743,N_47835,N_48166);
nand UO_4744 (O_4744,N_48072,N_49368);
and UO_4745 (O_4745,N_48979,N_48625);
nor UO_4746 (O_4746,N_49965,N_47890);
or UO_4747 (O_4747,N_49910,N_48106);
and UO_4748 (O_4748,N_48088,N_49783);
nand UO_4749 (O_4749,N_47766,N_49901);
and UO_4750 (O_4750,N_48943,N_49214);
xnor UO_4751 (O_4751,N_49442,N_49506);
or UO_4752 (O_4752,N_48645,N_48043);
or UO_4753 (O_4753,N_47956,N_48010);
xor UO_4754 (O_4754,N_47640,N_48537);
nor UO_4755 (O_4755,N_48585,N_49852);
nand UO_4756 (O_4756,N_49224,N_48834);
xor UO_4757 (O_4757,N_48285,N_49215);
nor UO_4758 (O_4758,N_49727,N_49378);
or UO_4759 (O_4759,N_48518,N_47610);
nand UO_4760 (O_4760,N_49769,N_49241);
nand UO_4761 (O_4761,N_48217,N_49233);
or UO_4762 (O_4762,N_48300,N_49230);
nor UO_4763 (O_4763,N_49206,N_49340);
or UO_4764 (O_4764,N_49643,N_49540);
and UO_4765 (O_4765,N_48572,N_47829);
nor UO_4766 (O_4766,N_48725,N_48399);
xnor UO_4767 (O_4767,N_49023,N_49524);
and UO_4768 (O_4768,N_48971,N_47826);
xor UO_4769 (O_4769,N_49238,N_47851);
or UO_4770 (O_4770,N_49060,N_48946);
xor UO_4771 (O_4771,N_48306,N_47580);
nor UO_4772 (O_4772,N_49035,N_49983);
xor UO_4773 (O_4773,N_48512,N_48195);
and UO_4774 (O_4774,N_48269,N_48008);
or UO_4775 (O_4775,N_49368,N_47737);
or UO_4776 (O_4776,N_48505,N_48635);
nor UO_4777 (O_4777,N_49998,N_47670);
nand UO_4778 (O_4778,N_48601,N_48595);
xor UO_4779 (O_4779,N_48447,N_49605);
nand UO_4780 (O_4780,N_48214,N_49452);
and UO_4781 (O_4781,N_49893,N_48556);
nor UO_4782 (O_4782,N_49858,N_47665);
xor UO_4783 (O_4783,N_48248,N_48212);
nand UO_4784 (O_4784,N_47886,N_48215);
and UO_4785 (O_4785,N_48584,N_48695);
and UO_4786 (O_4786,N_49440,N_48993);
xor UO_4787 (O_4787,N_47882,N_49562);
nand UO_4788 (O_4788,N_49329,N_49220);
or UO_4789 (O_4789,N_48096,N_49677);
xor UO_4790 (O_4790,N_48189,N_47817);
nand UO_4791 (O_4791,N_48264,N_47949);
nor UO_4792 (O_4792,N_49526,N_48564);
or UO_4793 (O_4793,N_48707,N_49020);
or UO_4794 (O_4794,N_49763,N_47640);
nand UO_4795 (O_4795,N_49507,N_48572);
or UO_4796 (O_4796,N_48843,N_48215);
and UO_4797 (O_4797,N_49031,N_48802);
nor UO_4798 (O_4798,N_49304,N_48330);
nand UO_4799 (O_4799,N_49472,N_48842);
nor UO_4800 (O_4800,N_48460,N_49862);
nor UO_4801 (O_4801,N_47642,N_49206);
or UO_4802 (O_4802,N_48276,N_48620);
and UO_4803 (O_4803,N_48035,N_49529);
nor UO_4804 (O_4804,N_48455,N_48277);
and UO_4805 (O_4805,N_48768,N_49104);
nor UO_4806 (O_4806,N_48410,N_48896);
nand UO_4807 (O_4807,N_47903,N_47933);
or UO_4808 (O_4808,N_48772,N_47663);
xor UO_4809 (O_4809,N_48806,N_47538);
or UO_4810 (O_4810,N_48999,N_48018);
xnor UO_4811 (O_4811,N_49561,N_49376);
and UO_4812 (O_4812,N_49699,N_49973);
and UO_4813 (O_4813,N_49993,N_49064);
nand UO_4814 (O_4814,N_49793,N_49299);
or UO_4815 (O_4815,N_48715,N_48081);
and UO_4816 (O_4816,N_47650,N_48176);
and UO_4817 (O_4817,N_49289,N_49233);
xnor UO_4818 (O_4818,N_48522,N_49072);
xnor UO_4819 (O_4819,N_47902,N_48787);
nor UO_4820 (O_4820,N_47736,N_48456);
nor UO_4821 (O_4821,N_48005,N_49180);
nand UO_4822 (O_4822,N_49023,N_48328);
and UO_4823 (O_4823,N_47874,N_48125);
and UO_4824 (O_4824,N_48986,N_48842);
xor UO_4825 (O_4825,N_48365,N_48740);
and UO_4826 (O_4826,N_48543,N_49287);
or UO_4827 (O_4827,N_49529,N_48857);
nand UO_4828 (O_4828,N_47737,N_49887);
nor UO_4829 (O_4829,N_47793,N_48840);
nand UO_4830 (O_4830,N_49944,N_47877);
or UO_4831 (O_4831,N_48689,N_49393);
or UO_4832 (O_4832,N_48801,N_47886);
xnor UO_4833 (O_4833,N_47531,N_47825);
or UO_4834 (O_4834,N_49842,N_48725);
or UO_4835 (O_4835,N_47556,N_49027);
nor UO_4836 (O_4836,N_48616,N_48629);
xnor UO_4837 (O_4837,N_48038,N_47884);
or UO_4838 (O_4838,N_49203,N_48205);
xor UO_4839 (O_4839,N_48141,N_48601);
and UO_4840 (O_4840,N_49936,N_49610);
nor UO_4841 (O_4841,N_47912,N_48563);
xnor UO_4842 (O_4842,N_47760,N_48581);
nand UO_4843 (O_4843,N_49026,N_48587);
nor UO_4844 (O_4844,N_49731,N_49361);
nor UO_4845 (O_4845,N_48582,N_49055);
nor UO_4846 (O_4846,N_48727,N_49533);
xor UO_4847 (O_4847,N_48091,N_47527);
nand UO_4848 (O_4848,N_48491,N_47771);
nor UO_4849 (O_4849,N_48204,N_48394);
nand UO_4850 (O_4850,N_48477,N_48958);
nor UO_4851 (O_4851,N_49470,N_49244);
or UO_4852 (O_4852,N_48445,N_49962);
nor UO_4853 (O_4853,N_48822,N_49774);
nand UO_4854 (O_4854,N_49126,N_49484);
or UO_4855 (O_4855,N_48838,N_48826);
or UO_4856 (O_4856,N_48044,N_48810);
or UO_4857 (O_4857,N_48433,N_49602);
or UO_4858 (O_4858,N_48860,N_48167);
nor UO_4859 (O_4859,N_48046,N_49411);
nand UO_4860 (O_4860,N_49076,N_49743);
or UO_4861 (O_4861,N_49545,N_49409);
xor UO_4862 (O_4862,N_49280,N_48773);
nor UO_4863 (O_4863,N_49451,N_48414);
or UO_4864 (O_4864,N_48674,N_49637);
or UO_4865 (O_4865,N_48155,N_49789);
and UO_4866 (O_4866,N_49478,N_48926);
nand UO_4867 (O_4867,N_49625,N_48017);
xnor UO_4868 (O_4868,N_47742,N_48231);
nand UO_4869 (O_4869,N_48523,N_48140);
or UO_4870 (O_4870,N_47962,N_47746);
nor UO_4871 (O_4871,N_48908,N_48997);
nand UO_4872 (O_4872,N_49501,N_47824);
nand UO_4873 (O_4873,N_48928,N_49668);
nor UO_4874 (O_4874,N_48226,N_49577);
xor UO_4875 (O_4875,N_48207,N_48975);
nand UO_4876 (O_4876,N_47687,N_49018);
nand UO_4877 (O_4877,N_48325,N_49371);
nand UO_4878 (O_4878,N_49574,N_49877);
nor UO_4879 (O_4879,N_49193,N_48750);
nand UO_4880 (O_4880,N_47711,N_48123);
nand UO_4881 (O_4881,N_49185,N_48355);
nor UO_4882 (O_4882,N_49305,N_49080);
nor UO_4883 (O_4883,N_47762,N_48468);
xor UO_4884 (O_4884,N_49893,N_48521);
xor UO_4885 (O_4885,N_48581,N_47673);
nand UO_4886 (O_4886,N_48466,N_49454);
or UO_4887 (O_4887,N_49433,N_48933);
nor UO_4888 (O_4888,N_47545,N_48441);
nand UO_4889 (O_4889,N_47665,N_48908);
nor UO_4890 (O_4890,N_47759,N_47734);
or UO_4891 (O_4891,N_47750,N_49901);
or UO_4892 (O_4892,N_48330,N_47548);
and UO_4893 (O_4893,N_49252,N_47736);
nand UO_4894 (O_4894,N_49803,N_49429);
nor UO_4895 (O_4895,N_49202,N_49788);
nor UO_4896 (O_4896,N_48632,N_47735);
nand UO_4897 (O_4897,N_49938,N_48583);
xor UO_4898 (O_4898,N_48483,N_49894);
or UO_4899 (O_4899,N_48547,N_49152);
nor UO_4900 (O_4900,N_48520,N_49806);
and UO_4901 (O_4901,N_48801,N_47526);
or UO_4902 (O_4902,N_49420,N_47552);
nor UO_4903 (O_4903,N_48782,N_49006);
or UO_4904 (O_4904,N_48937,N_47778);
xnor UO_4905 (O_4905,N_47585,N_49190);
xnor UO_4906 (O_4906,N_48600,N_47690);
nor UO_4907 (O_4907,N_49205,N_48097);
xnor UO_4908 (O_4908,N_49592,N_49048);
or UO_4909 (O_4909,N_48259,N_48776);
nand UO_4910 (O_4910,N_48359,N_47837);
or UO_4911 (O_4911,N_48618,N_48660);
xnor UO_4912 (O_4912,N_49365,N_49659);
or UO_4913 (O_4913,N_48983,N_47620);
or UO_4914 (O_4914,N_47533,N_48823);
nor UO_4915 (O_4915,N_49148,N_48091);
xnor UO_4916 (O_4916,N_49774,N_47954);
nor UO_4917 (O_4917,N_48772,N_47695);
and UO_4918 (O_4918,N_48561,N_48842);
xor UO_4919 (O_4919,N_48871,N_49223);
or UO_4920 (O_4920,N_49512,N_48425);
and UO_4921 (O_4921,N_49810,N_48661);
xor UO_4922 (O_4922,N_48871,N_49850);
nor UO_4923 (O_4923,N_48712,N_48603);
nand UO_4924 (O_4924,N_49023,N_47788);
and UO_4925 (O_4925,N_47620,N_49824);
nand UO_4926 (O_4926,N_48107,N_49113);
xor UO_4927 (O_4927,N_48276,N_48496);
and UO_4928 (O_4928,N_48914,N_49847);
xnor UO_4929 (O_4929,N_48856,N_49405);
and UO_4930 (O_4930,N_48202,N_48379);
nand UO_4931 (O_4931,N_47673,N_49160);
or UO_4932 (O_4932,N_48284,N_48349);
nand UO_4933 (O_4933,N_47757,N_49871);
or UO_4934 (O_4934,N_47613,N_47967);
and UO_4935 (O_4935,N_47873,N_49622);
xor UO_4936 (O_4936,N_49003,N_48246);
and UO_4937 (O_4937,N_49239,N_48940);
xnor UO_4938 (O_4938,N_48383,N_47640);
or UO_4939 (O_4939,N_48295,N_49085);
nand UO_4940 (O_4940,N_49041,N_48801);
nor UO_4941 (O_4941,N_49036,N_48486);
nor UO_4942 (O_4942,N_49089,N_48629);
and UO_4943 (O_4943,N_48609,N_49798);
nand UO_4944 (O_4944,N_48668,N_49405);
or UO_4945 (O_4945,N_49533,N_49574);
nand UO_4946 (O_4946,N_48250,N_49778);
nor UO_4947 (O_4947,N_49783,N_49854);
and UO_4948 (O_4948,N_49409,N_47528);
and UO_4949 (O_4949,N_47702,N_48465);
nor UO_4950 (O_4950,N_48814,N_49076);
or UO_4951 (O_4951,N_49875,N_48713);
or UO_4952 (O_4952,N_48675,N_49979);
xor UO_4953 (O_4953,N_48491,N_48977);
or UO_4954 (O_4954,N_48084,N_47642);
xor UO_4955 (O_4955,N_49670,N_49325);
xor UO_4956 (O_4956,N_49132,N_47851);
nor UO_4957 (O_4957,N_49970,N_48758);
xor UO_4958 (O_4958,N_48495,N_48908);
xnor UO_4959 (O_4959,N_48565,N_48797);
and UO_4960 (O_4960,N_49375,N_47776);
or UO_4961 (O_4961,N_49421,N_48362);
nor UO_4962 (O_4962,N_49856,N_49015);
or UO_4963 (O_4963,N_48057,N_49156);
or UO_4964 (O_4964,N_49644,N_49926);
and UO_4965 (O_4965,N_47614,N_48700);
and UO_4966 (O_4966,N_49144,N_47503);
nand UO_4967 (O_4967,N_47735,N_48001);
and UO_4968 (O_4968,N_47887,N_49514);
xnor UO_4969 (O_4969,N_49227,N_49876);
xor UO_4970 (O_4970,N_49086,N_48608);
nand UO_4971 (O_4971,N_48232,N_48795);
nand UO_4972 (O_4972,N_48018,N_48213);
or UO_4973 (O_4973,N_48380,N_48912);
and UO_4974 (O_4974,N_47752,N_49750);
and UO_4975 (O_4975,N_48995,N_48602);
nand UO_4976 (O_4976,N_48690,N_49772);
xnor UO_4977 (O_4977,N_48655,N_49240);
nor UO_4978 (O_4978,N_48330,N_48962);
nand UO_4979 (O_4979,N_49438,N_49156);
xnor UO_4980 (O_4980,N_49973,N_48644);
nand UO_4981 (O_4981,N_49842,N_49413);
nor UO_4982 (O_4982,N_49833,N_48689);
nand UO_4983 (O_4983,N_48677,N_49896);
nand UO_4984 (O_4984,N_49382,N_47737);
or UO_4985 (O_4985,N_49649,N_49947);
and UO_4986 (O_4986,N_48026,N_48123);
and UO_4987 (O_4987,N_48967,N_48500);
xnor UO_4988 (O_4988,N_49168,N_49797);
nor UO_4989 (O_4989,N_48320,N_49400);
nand UO_4990 (O_4990,N_49910,N_49331);
or UO_4991 (O_4991,N_49503,N_49325);
xnor UO_4992 (O_4992,N_49629,N_49461);
and UO_4993 (O_4993,N_48206,N_49820);
nor UO_4994 (O_4994,N_49945,N_49281);
and UO_4995 (O_4995,N_47601,N_49704);
xor UO_4996 (O_4996,N_47810,N_49883);
nor UO_4997 (O_4997,N_47537,N_48886);
nor UO_4998 (O_4998,N_49034,N_49176);
nor UO_4999 (O_4999,N_49396,N_49885);
endmodule